--------------------------------------------------------- 
-- Ce programme a ete developpe a CENTRALESUPELEC
-- Merci de conserver ce cartouche
-- Copyright  (c) 2021  CENTRALESUPELEC   
-- Dpartement Systmes lectroniques
-- ------------------------------------------------------
--
-- fichier : testbench_e.vhd
-- auteur  : P.BENABES   
-- Copyright (c) 2021 CENTRALE-SUPELEC
-- Revision: 1.0  Date: 04/01/2021
--
---------------------------------------------------------
---------------------------------------------------------
--
-- DESCRIPTION DU CODE :
-- ce module est le plus haut niveau du testbench de la pll 
--
----------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.all;
use IEEE.numeric_std.ALL;
use work.coeff.all ;


ENTITY testbench IS
END testbench;
