-------------------------------------------------------
-- Ce programme a été développé à CENTRALE-SUPELEC
-- Merci de conserver ce cartouche
-- Copyright  (c) 2022  CENTRALE-SUPELEC   
-- Département Systèmes électroniques
-- ---------------------------------------------------
--
-- fichier : testbench_Cpresynth_0.vhd
-- auteur  : P.BENABES   
-- Copyright (c) 2022 CENTRALE-SUPELEC
-- Revision: 4.1  Date: 22/02/2022
--
-- ---------------------------------------------------
-- ---------------------------------------------------
--
-- DESCRIPTION DU SCRIPT :
-- Configuration pour la simulation initiale avant synthèse 
-- route_io=0 lowpower=0 multialim=0
--
--------------------------------------------------------

configuration Cpresynth of testbench is 
  for A1
  end for;
end Cpresynth ;

