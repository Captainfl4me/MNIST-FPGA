LIBRARY ieee,work;
USE ieee.std_logic_1164.all;
use IEEE.numeric_std.ALL;
use std.textio.all;
use ieee.fixed_pkg.all;
use ieee.fixed_float_types.all;

package coeff is
 
    constant lngimag : integer := 784 ; 
    constant lngfilt : integer := 680 ; 
    constant nbneuron : integer := 70 ; 
    constant nbsymbol : integer := 10 ; 
    constant nbitq : integer := 8 ; 

type typtabup is array(0 to lngimag-1) of std_logic ;								-- tableau indiquant les pixels effectivement utilisés lors des calculs
type typtabcst is array(natural range <>) of sfixed(1 downto -nbitq) ;				-- tableau des constantes du premier étage de neurones
type typtabaccu is array(0 to nbneuron-1) of sfixed(5 downto -2*nbitq) ;
type typtabaccu2 is array(0 to nbsymbol-1) of sfixed(5 downto -2*nbitq) ;
subtype usng4 is unsigned(3 downto 0) ;
type typlabel is array(0 to 4) of usng4 ;


constant ccf : integer := 4 ; 
constant ccf2 : integer := 4 ; 
constant cct : integer := 16 ; 
constant cct2 : integer := 1 ; 

constant usedpix : typtabup := ( '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0'  ) ; 

constant allcoef1 : typtabcst := ( to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(63.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(62.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-61.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-58.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(62.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-61.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-63.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(62.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-62.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(63.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-71.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-73.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-93.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(62.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-56.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-68.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-73.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-62.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-81.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-62.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-70.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(63.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(74.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(81.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-103.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-63.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(65.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-72.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(64.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(62.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-62.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-56.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(75.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-64.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-87.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(79.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(139.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-97.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(93.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-64.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(62.0/256.0,1,-nbitq), 
to_sfixed(-61.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-66.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-63.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-67.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-60.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-61.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(66.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(63.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(62.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(74.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-74.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-71.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(72.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-63.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(77.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-69.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(83.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(72.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(70.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(62.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-74.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(62.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-68.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(125.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(89.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(70.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(63.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-60.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(-56.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(75.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(76.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(67.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-66.0/256.0,1,-nbitq), 
to_sfixed(78.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-59.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(79.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(62.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(63.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(81.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-61.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-58.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-73.0/256.0,1,-nbitq), 
to_sfixed(-67.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(77.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(64.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-72.0/256.0,1,-nbitq), 
to_sfixed(-67.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-69.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(64.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-73.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(72.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(78.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-56.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-61.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-59.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(62.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(98.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(66.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-56.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-73.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-72.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(76.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(63.0/256.0,1,-nbitq), 
to_sfixed(87.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(64.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(69.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(78.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-58.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(96.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(70.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-77.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-95.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-59.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(69.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-72.0/256.0,1,-nbitq), 
to_sfixed(-76.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(63.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-69.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-63.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(63.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(64.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(65.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-67.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-56.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-63.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(64.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(62.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(71.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-86.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(67.0/256.0,1,-nbitq), 
to_sfixed(71.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-59.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(66.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-60.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(81.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-75.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(71.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(80.0/256.0,1,-nbitq), 
to_sfixed(65.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-90.0/256.0,1,-nbitq), 
to_sfixed(-63.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(83.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(81.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(95.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-77.0/256.0,1,-nbitq), 
to_sfixed(-71.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-62.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(71.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-63.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-56.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-103.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(72.0/256.0,1,-nbitq), 
to_sfixed(70.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(63.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-105.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(70.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(76.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-61.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-56.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-58.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(65.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(-58.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(80.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-58.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-67.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(68.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-68.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(62.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-62.0/256.0,1,-nbitq), 
to_sfixed(-69.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(65.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(75.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(86.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-71.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(62.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(87.0/256.0,1,-nbitq), 
to_sfixed(84.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(80.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(-72.0/256.0,1,-nbitq), 
to_sfixed(-116.0/256.0,1,-nbitq), 
to_sfixed(-84.0/256.0,1,-nbitq), 
to_sfixed(-61.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(74.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-67.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-59.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(83.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(-107.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(62.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-90.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-60.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(68.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-67.0/256.0,1,-nbitq), 
to_sfixed(-70.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-59.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-83.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(73.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-56.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(86.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(68.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-56.0/256.0,1,-nbitq), 
to_sfixed(70.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-56.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(79.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(64.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-60.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-66.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-60.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-59.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(89.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-61.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(83.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-64.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(75.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(81.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(77.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(92.0/256.0,1,-nbitq), 
to_sfixed(67.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(109.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-66.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-59.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(64.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(70.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-71.0/256.0,1,-nbitq), 
to_sfixed(-67.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-76.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-64.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-81.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-72.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-56.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(63.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-59.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(68.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-63.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-79.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-67.0/256.0,1,-nbitq), 
to_sfixed(69.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-58.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-58.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(69.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(-79.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-60.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(65.0/256.0,1,-nbitq), 
to_sfixed(70.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-58.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(68.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(69.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-63.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(-66.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-84.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-80.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-70.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-59.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(72.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-61.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(68.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-68.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(63.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-59.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-62.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-66.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq) ) ; 

constant allcoef2 : typtabcst := ( to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(67.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(62.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-60.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-70.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-61.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-59.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(63.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(75.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(63.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(86.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(75.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-63.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-67.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(68.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(70.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(64.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(65.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(74.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-60.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(76.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(78.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(67.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(80.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(83.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(78.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(70.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-64.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(66.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(78.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(87.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(67.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(83.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-29.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(-10.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-215.0/256.0,1,-nbitq), 
to_sfixed(74.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-110.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(96.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-59.0/256.0,1,-nbitq), 
to_sfixed(79.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(67.0/256.0,1,-nbitq), 
to_sfixed(-69.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(97.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(120.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-56.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(98.0/256.0,1,-nbitq), 
to_sfixed(-2.0/256.0,1,-nbitq), 
to_sfixed(-138.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(75.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(-61.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(73.0/256.0,1,-nbitq), 
to_sfixed(-63.0/256.0,1,-nbitq), 
to_sfixed(-56.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(75.0/256.0,1,-nbitq), 
to_sfixed(-100.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(66.0/256.0,1,-nbitq), 
to_sfixed(97.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-88.0/256.0,1,-nbitq), 
to_sfixed(-115.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(-70.0/256.0,1,-nbitq), 
to_sfixed(-85.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-82.0/256.0,1,-nbitq), 
to_sfixed(72.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(75.0/256.0,1,-nbitq), 
to_sfixed(84.0/256.0,1,-nbitq), 
to_sfixed(-140.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(66.0/256.0,1,-nbitq), 
to_sfixed(78.0/256.0,1,-nbitq), 
to_sfixed(57.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(-82.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(86.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-71.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-123.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(-64.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(82.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-96.0/256.0,1,-nbitq), 
to_sfixed(-55.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-90.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(76.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(-99.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-79.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-60.0/256.0,1,-nbitq), 
to_sfixed(-62.0/256.0,1,-nbitq), 
to_sfixed(71.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-95.0/256.0,1,-nbitq), 
to_sfixed(108.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-99.0/256.0,1,-nbitq), 
to_sfixed(77.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(94.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(85.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-23.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-64.0/256.0,1,-nbitq), 
to_sfixed(84.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-87.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(69.0/256.0,1,-nbitq), 
to_sfixed(-105.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(-90.0/256.0,1,-nbitq), 
to_sfixed(-131.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(133.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(96.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(107.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-69.0/256.0,1,-nbitq), 
to_sfixed(-62.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(34.0/256.0,1,-nbitq), 
to_sfixed(66.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(80.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-40.0/256.0,1,-nbitq), 
to_sfixed(-63.0/256.0,1,-nbitq), 
to_sfixed(-110.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(153.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(69.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-117.0/256.0,1,-nbitq), 
to_sfixed(87.0/256.0,1,-nbitq), 
to_sfixed(68.0/256.0,1,-nbitq), 
to_sfixed(110.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(-69.0/256.0,1,-nbitq), 
to_sfixed(76.0/256.0,1,-nbitq), 
to_sfixed(-101.0/256.0,1,-nbitq), 
to_sfixed(92.0/256.0,1,-nbitq), 
to_sfixed(-96.0/256.0,1,-nbitq), 
to_sfixed(-85.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(66.0/256.0,1,-nbitq), 
to_sfixed(-85.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(-69.0/256.0,1,-nbitq), 
to_sfixed(69.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-78.0/256.0,1,-nbitq), 
to_sfixed(78.0/256.0,1,-nbitq), 
to_sfixed(-91.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-35.0/256.0,1,-nbitq), 
to_sfixed(99.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-60.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(-57.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-93.0/256.0,1,-nbitq), 
to_sfixed(-84.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(87.0/256.0,1,-nbitq), 
to_sfixed(-92.0/256.0,1,-nbitq), 
to_sfixed(118.0/256.0,1,-nbitq), 
to_sfixed(143.0/256.0,1,-nbitq), 
to_sfixed(94.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(-43.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-103.0/256.0,1,-nbitq), 
to_sfixed(-58.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(-83.0/256.0,1,-nbitq), 
to_sfixed(-119.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(96.0/256.0,1,-nbitq), 
to_sfixed(28.0/256.0,1,-nbitq), 
to_sfixed(143.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-70.0/256.0,1,-nbitq), 
to_sfixed(85.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(-81.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(94.0/256.0,1,-nbitq), 
to_sfixed(-48.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(63.0/256.0,1,-nbitq), 
to_sfixed(83.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(82.0/256.0,1,-nbitq), 
to_sfixed(-137.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(-115.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(-84.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(65.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(89.0/256.0,1,-nbitq), 
to_sfixed(-89.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(101.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(-86.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(-61.0/256.0,1,-nbitq), 
to_sfixed(100.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-62.0/256.0,1,-nbitq), 
to_sfixed(8.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(72.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(115.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(13.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(-6.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-80.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(9.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(1.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(-58.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(91.0/256.0,1,-nbitq), 
to_sfixed(101.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-19.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(85.0/256.0,1,-nbitq), 
to_sfixed(55.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(-102.0/256.0,1,-nbitq), 
to_sfixed(-17.0/256.0,1,-nbitq), 
to_sfixed(49.0/256.0,1,-nbitq), 
to_sfixed(76.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(122.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(128.0/256.0,1,-nbitq), 
to_sfixed(120.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-88.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(-94.0/256.0,1,-nbitq), 
to_sfixed(-87.0/256.0,1,-nbitq), 
to_sfixed(-32.0/256.0,1,-nbitq), 
to_sfixed(-99.0/256.0,1,-nbitq), 
to_sfixed(-44.0/256.0,1,-nbitq), 
to_sfixed(80.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(64.0/256.0,1,-nbitq), 
to_sfixed(10.0/256.0,1,-nbitq), 
to_sfixed(97.0/256.0,1,-nbitq), 
to_sfixed(-77.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(135.0/256.0,1,-nbitq), 
to_sfixed(12.0/256.0,1,-nbitq), 
to_sfixed(-117.0/256.0,1,-nbitq), 
to_sfixed(-61.0/256.0,1,-nbitq), 
to_sfixed(-92.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(93.0/256.0,1,-nbitq), 
to_sfixed(81.0/256.0,1,-nbitq), 
to_sfixed(-51.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(68.0/256.0,1,-nbitq), 
to_sfixed(-36.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(-58.0/256.0,1,-nbitq), 
to_sfixed(-82.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-103.0/256.0,1,-nbitq), 
to_sfixed(114.0/256.0,1,-nbitq), 
to_sfixed(-105.0/256.0,1,-nbitq), 
to_sfixed(100.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(44.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(25.0/256.0,1,-nbitq), 
to_sfixed(29.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(73.0/256.0,1,-nbitq), 
to_sfixed(30.0/256.0,1,-nbitq), 
to_sfixed(65.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(-4.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-58.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-11.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(7.0/256.0,1,-nbitq), 
to_sfixed(-28.0/256.0,1,-nbitq), 
to_sfixed(-75.0/256.0,1,-nbitq), 
to_sfixed(70.0/256.0,1,-nbitq), 
to_sfixed(-71.0/256.0,1,-nbitq), 
to_sfixed(39.0/256.0,1,-nbitq), 
to_sfixed(93.0/256.0,1,-nbitq), 
to_sfixed(-76.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(64.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(-67.0/256.0,1,-nbitq), 
to_sfixed(66.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-66.0/256.0,1,-nbitq), 
to_sfixed(-62.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(73.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(-47.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(16.0/256.0,1,-nbitq), 
to_sfixed(-60.0/256.0,1,-nbitq), 
to_sfixed(-30.0/256.0,1,-nbitq), 
to_sfixed(74.0/256.0,1,-nbitq), 
to_sfixed(-65.0/256.0,1,-nbitq), 
to_sfixed(66.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-77.0/256.0,1,-nbitq), 
to_sfixed(-72.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(58.0/256.0,1,-nbitq), 
to_sfixed(5.0/256.0,1,-nbitq), 
to_sfixed(69.0/256.0,1,-nbitq), 
to_sfixed(76.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(-90.0/256.0,1,-nbitq), 
to_sfixed(54.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(51.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(65.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(48.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(66.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(18.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(-15.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(-49.0/256.0,1,-nbitq), 
to_sfixed(-41.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-56.0/256.0,1,-nbitq), 
to_sfixed(74.0/256.0,1,-nbitq), 
to_sfixed(56.0/256.0,1,-nbitq), 
to_sfixed(-112.0/256.0,1,-nbitq), 
to_sfixed(-42.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(69.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-53.0/256.0,1,-nbitq), 
to_sfixed(-27.0/256.0,1,-nbitq), 
to_sfixed(45.0/256.0,1,-nbitq), 
to_sfixed(-68.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(42.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(60.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(33.0/256.0,1,-nbitq), 
to_sfixed(-64.0/256.0,1,-nbitq), 
to_sfixed(-39.0/256.0,1,-nbitq), 
to_sfixed(-12.0/256.0,1,-nbitq), 
to_sfixed(15.0/256.0,1,-nbitq), 
to_sfixed(0.0/256.0,1,-nbitq), 
to_sfixed(-64.0/256.0,1,-nbitq), 
to_sfixed(-33.0/256.0,1,-nbitq), 
to_sfixed(-20.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(36.0/256.0,1,-nbitq), 
to_sfixed(144.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(95.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(-58.0/256.0,1,-nbitq), 
to_sfixed(-91.0/256.0,1,-nbitq), 
to_sfixed(-38.0/256.0,1,-nbitq), 
to_sfixed(-78.0/256.0,1,-nbitq), 
to_sfixed(-83.0/256.0,1,-nbitq), 
to_sfixed(-73.0/256.0,1,-nbitq), 
to_sfixed(-31.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-67.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-67.0/256.0,1,-nbitq), 
to_sfixed(-25.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(23.0/256.0,1,-nbitq), 
to_sfixed(22.0/256.0,1,-nbitq), 
to_sfixed(26.0/256.0,1,-nbitq), 
to_sfixed(-8.0/256.0,1,-nbitq), 
to_sfixed(31.0/256.0,1,-nbitq), 
to_sfixed(-7.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(-60.0/256.0,1,-nbitq), 
to_sfixed(-56.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(-13.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(24.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(74.0/256.0,1,-nbitq), 
to_sfixed(59.0/256.0,1,-nbitq), 
to_sfixed(-105.0/256.0,1,-nbitq), 
to_sfixed(-9.0/256.0,1,-nbitq), 
to_sfixed(21.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(11.0/256.0,1,-nbitq), 
to_sfixed(96.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-1.0/256.0,1,-nbitq), 
to_sfixed(40.0/256.0,1,-nbitq), 
to_sfixed(41.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(69.0/256.0,1,-nbitq), 
to_sfixed(17.0/256.0,1,-nbitq), 
to_sfixed(-52.0/256.0,1,-nbitq), 
to_sfixed(35.0/256.0,1,-nbitq), 
to_sfixed(-72.0/256.0,1,-nbitq), 
to_sfixed(65.0/256.0,1,-nbitq), 
to_sfixed(4.0/256.0,1,-nbitq), 
to_sfixed(2.0/256.0,1,-nbitq), 
to_sfixed(-3.0/256.0,1,-nbitq), 
to_sfixed(-91.0/256.0,1,-nbitq), 
to_sfixed(14.0/256.0,1,-nbitq), 
to_sfixed(-68.0/256.0,1,-nbitq), 
to_sfixed(46.0/256.0,1,-nbitq), 
to_sfixed(-129.0/256.0,1,-nbitq), 
to_sfixed(90.0/256.0,1,-nbitq), 
to_sfixed(74.0/256.0,1,-nbitq), 
to_sfixed(-5.0/256.0,1,-nbitq), 
to_sfixed(43.0/256.0,1,-nbitq), 
to_sfixed(47.0/256.0,1,-nbitq), 
to_sfixed(-82.0/256.0,1,-nbitq), 
to_sfixed(52.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-50.0/256.0,1,-nbitq), 
to_sfixed(53.0/256.0,1,-nbitq), 
to_sfixed(-14.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(27.0/256.0,1,-nbitq), 
to_sfixed(-54.0/256.0,1,-nbitq), 
to_sfixed(-68.0/256.0,1,-nbitq), 
to_sfixed(50.0/256.0,1,-nbitq), 
to_sfixed(-85.0/256.0,1,-nbitq), 
to_sfixed(20.0/256.0,1,-nbitq), 
to_sfixed(88.0/256.0,1,-nbitq), 
to_sfixed(-24.0/256.0,1,-nbitq), 
to_sfixed(-89.0/256.0,1,-nbitq), 
to_sfixed(-34.0/256.0,1,-nbitq), 
to_sfixed(-46.0/256.0,1,-nbitq), 
to_sfixed(63.0/256.0,1,-nbitq), 
to_sfixed(67.0/256.0,1,-nbitq), 
to_sfixed(3.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(32.0/256.0,1,-nbitq), 
to_sfixed(-45.0/256.0,1,-nbitq), 
to_sfixed(19.0/256.0,1,-nbitq), 
to_sfixed(-64.0/256.0,1,-nbitq), 
to_sfixed(66.0/256.0,1,-nbitq), 
to_sfixed(-37.0/256.0,1,-nbitq), 
to_sfixed(-18.0/256.0,1,-nbitq), 
to_sfixed(37.0/256.0,1,-nbitq), 
to_sfixed(6.0/256.0,1,-nbitq), 
to_sfixed(90.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(71.0/256.0,1,-nbitq), 
to_sfixed(38.0/256.0,1,-nbitq), 
to_sfixed(-21.0/256.0,1,-nbitq), 
to_sfixed(-84.0/256.0,1,-nbitq), 
to_sfixed(82.0/256.0,1,-nbitq), 
to_sfixed(-22.0/256.0,1,-nbitq), 
to_sfixed(67.0/256.0,1,-nbitq), 
to_sfixed(-16.0/256.0,1,-nbitq), 
to_sfixed(72.0/256.0,1,-nbitq), 
to_sfixed(-86.0/256.0,1,-nbitq), 
to_sfixed(186.0/256.0,1,-nbitq), 
to_sfixed(61.0/256.0,1,-nbitq), 
to_sfixed(-209.0/256.0,1,-nbitq), 
to_sfixed(202.0/256.0,1,-nbitq), 
to_sfixed(95.0/256.0,1,-nbitq), 
to_sfixed(88.0/256.0,1,-nbitq), 
to_sfixed(-221.0/256.0,1,-nbitq), 
to_sfixed(-135.0/256.0,1,-nbitq), 
to_sfixed(-196.0/256.0,1,-nbitq), 
to_sfixed(-26.0/256.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq), 
to_sfixed(0.0,1,-nbitq) 
 ) ;

 end package coeff;