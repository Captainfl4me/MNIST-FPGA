LIBRARY ieee,work;
USE ieee.std_logic_1164.all;
use IEEE.numeric_std.ALL;
use std.textio.all;
use ieee.fixed_pkg.all;
use ieee.fixed_float_types.all;

package coeff is
 
constant lngimag : integer := 784 ; 
constant lngfilt : integer := 784 ; 
constant nbneuron : integer := 80 ; 
constant nbsymbol : integer := 10 ; 
constant nbitq : integer := 16 ; 


constant ccf : integer := 4 ; 
constant ccf2 : integer := 4 ; 
constant cct : integer := 32 ; 
constant cct2 : integer := 1 ; 

type typtabup is array(0 to lngimag-1) of std_logic ;								-- tableau indiquant les pixels effectivement utilisés lors des calculs
type typtabmul is array(natural range <>) of sfixed(3 downto -nbitq);
type typtabcst is array(natural range <>) of sfixed(1 downto -nbitq);
type typtabcnf1 is array(0 to lngimag-1, 0 to nbneuron-1) of sfixed(1 downto -nbitq);
type typtabcnf2 is array(0 to nbneuron-1, 0 to nbsymbol-1) of sfixed(1 downto -nbitq);
type typtabaccu is array(0 to nbneuron-1) of sfixed(8 downto -2*nbitq) ;
type typtabaccu2 is array(0 to nbsymbol-1) of sfixed(8 downto -2*nbitq) ;
subtype usng4 is unsigned(3 downto 0) ;
type typlabel is array(0 to 4) of usng4 ;

constant usedpix : typtabup := ( '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1'  ) ; 

constant cst1 : typtabcst := ( to_sfixed(-3824.0/65536.0,1,-nbitq), to_sfixed(-1411.0/65536.0,1,-nbitq), to_sfixed(512.0/65536.0,1,-nbitq), to_sfixed(3511.0/65536.0,1,-nbitq), to_sfixed(3803.0/65536.0,1,-nbitq), to_sfixed(-1067.0/65536.0,1,-nbitq), to_sfixed(8672.0/65536.0,1,-nbitq), to_sfixed(-6464.0/65536.0,1,-nbitq), to_sfixed(802.0/65536.0,1,-nbitq), to_sfixed(-9087.0/65536.0,1,-nbitq), to_sfixed(-20425.0/65536.0,1,-nbitq), to_sfixed(-6127.0/65536.0,1,-nbitq), to_sfixed(-12375.0/65536.0,1,-nbitq), to_sfixed(7300.0/65536.0,1,-nbitq), to_sfixed(-868.0/65536.0,1,-nbitq), to_sfixed(-6519.0/65536.0,1,-nbitq), to_sfixed(7937.0/65536.0,1,-nbitq), to_sfixed(-1420.0/65536.0,1,-nbitq), to_sfixed(-5481.0/65536.0,1,-nbitq), to_sfixed(-13506.0/65536.0,1,-nbitq), to_sfixed(3556.0/65536.0,1,-nbitq), to_sfixed(8978.0/65536.0,1,-nbitq), to_sfixed(3851.0/65536.0,1,-nbitq), to_sfixed(-669.0/65536.0,1,-nbitq), to_sfixed(-4365.0/65536.0,1,-nbitq), to_sfixed(295.0/65536.0,1,-nbitq), to_sfixed(-1979.0/65536.0,1,-nbitq), to_sfixed(3466.0/65536.0,1,-nbitq), to_sfixed(-1071.0/65536.0,1,-nbitq), to_sfixed(2099.0/65536.0,1,-nbitq), to_sfixed(8684.0/65536.0,1,-nbitq), to_sfixed(-1952.0/65536.0,1,-nbitq), to_sfixed(8709.0/65536.0,1,-nbitq), to_sfixed(3305.0/65536.0,1,-nbitq), to_sfixed(16628.0/65536.0,1,-nbitq), to_sfixed(1895.0/65536.0,1,-nbitq), to_sfixed(5726.0/65536.0,1,-nbitq), to_sfixed(2644.0/65536.0,1,-nbitq), to_sfixed(3194.0/65536.0,1,-nbitq), to_sfixed(12063.0/65536.0,1,-nbitq), to_sfixed(-536.0/65536.0,1,-nbitq), to_sfixed(13148.0/65536.0,1,-nbitq), to_sfixed(3137.0/65536.0,1,-nbitq), to_sfixed(-807.0/65536.0,1,-nbitq), to_sfixed(-12406.0/65536.0,1,-nbitq), to_sfixed(-1280.0/65536.0,1,-nbitq), to_sfixed(11770.0/65536.0,1,-nbitq), to_sfixed(999.0/65536.0,1,-nbitq), to_sfixed(-26517.0/65536.0,1,-nbitq), to_sfixed(-52994.0/65536.0,1,-nbitq), to_sfixed(-11455.0/65536.0,1,-nbitq), to_sfixed(3127.0/65536.0,1,-nbitq), to_sfixed(-4367.0/65536.0,1,-nbitq), to_sfixed(-2077.0/65536.0,1,-nbitq), to_sfixed(-8691.0/65536.0,1,-nbitq), to_sfixed(7857.0/65536.0,1,-nbitq), to_sfixed(-8925.0/65536.0,1,-nbitq), to_sfixed(-1211.0/65536.0,1,-nbitq), to_sfixed(-2849.0/65536.0,1,-nbitq), to_sfixed(-9242.0/65536.0,1,-nbitq), to_sfixed(3912.0/65536.0,1,-nbitq), to_sfixed(10044.0/65536.0,1,-nbitq), to_sfixed(-10465.0/65536.0,1,-nbitq), to_sfixed(12922.0/65536.0,1,-nbitq), to_sfixed(2233.0/65536.0,1,-nbitq), to_sfixed(2987.0/65536.0,1,-nbitq), to_sfixed(21110.0/65536.0,1,-nbitq), to_sfixed(4299.0/65536.0,1,-nbitq), to_sfixed(2850.0/65536.0,1,-nbitq), to_sfixed(-4575.0/65536.0,1,-nbitq), to_sfixed(-2977.0/65536.0,1,-nbitq), to_sfixed(1618.0/65536.0,1,-nbitq), to_sfixed(-3692.0/65536.0,1,-nbitq), to_sfixed(14018.0/65536.0,1,-nbitq), to_sfixed(9485.0/65536.0,1,-nbitq), to_sfixed(2307.0/65536.0,1,-nbitq), to_sfixed(6002.0/65536.0,1,-nbitq), to_sfixed(-499.0/65536.0,1,-nbitq), to_sfixed(9093.0/65536.0,1,-nbitq), to_sfixed(-6588.0/65536.0,1,-nbitq)  ) ;

constant cst2 : typtabcst := ( to_sfixed(-51014.0/65536.0,1,-nbitq), to_sfixed(-51918.0/65536.0,1,-nbitq), to_sfixed(35896.0/65536.0,1,-nbitq), to_sfixed(-56605.0/65536.0,1,-nbitq), to_sfixed(-52934.0/65536.0,1,-nbitq), to_sfixed(-63534.0/65536.0,1,-nbitq), to_sfixed(-11642.0/65536.0,1,-nbitq), to_sfixed(-58542.0/65536.0,1,-nbitq), to_sfixed(-64144.0/65536.0,1,-nbitq), to_sfixed(11664.0/65536.0,1,-nbitq)  ) ;

constant coef1 : typtabcnf1 := ( ( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1211.0/65536.0,1,-nbitq), 
to_sfixed(2176.0/65536.0,1,-nbitq), 
to_sfixed(-226.0/65536.0,1,-nbitq), 
to_sfixed(-713.0/65536.0,1,-nbitq), 
to_sfixed(-2434.0/65536.0,1,-nbitq), 
to_sfixed(-824.0/65536.0,1,-nbitq), 
to_sfixed(873.0/65536.0,1,-nbitq), 
to_sfixed(1506.0/65536.0,1,-nbitq), 
to_sfixed(-2036.0/65536.0,1,-nbitq), 
to_sfixed(1165.0/65536.0,1,-nbitq), 
to_sfixed(-86.0/65536.0,1,-nbitq), 
to_sfixed(-3795.0/65536.0,1,-nbitq), 
to_sfixed(-2379.0/65536.0,1,-nbitq), 
to_sfixed(-1445.0/65536.0,1,-nbitq), 
to_sfixed(3283.0/65536.0,1,-nbitq), 
to_sfixed(-779.0/65536.0,1,-nbitq), 
to_sfixed(415.0/65536.0,1,-nbitq), 
to_sfixed(-746.0/65536.0,1,-nbitq), 
to_sfixed(2805.0/65536.0,1,-nbitq), 
to_sfixed(-1004.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(1322.0/65536.0,1,-nbitq), 
to_sfixed(2225.0/65536.0,1,-nbitq), 
to_sfixed(4308.0/65536.0,1,-nbitq), 
to_sfixed(469.0/65536.0,1,-nbitq), 
to_sfixed(-1599.0/65536.0,1,-nbitq), 
to_sfixed(-3273.0/65536.0,1,-nbitq), 
to_sfixed(-2058.0/65536.0,1,-nbitq), 
to_sfixed(1282.0/65536.0,1,-nbitq), 
to_sfixed(-2387.0/65536.0,1,-nbitq), 
to_sfixed(1839.0/65536.0,1,-nbitq), 
to_sfixed(-1683.0/65536.0,1,-nbitq), 
to_sfixed(-219.0/65536.0,1,-nbitq), 
to_sfixed(-3498.0/65536.0,1,-nbitq), 
to_sfixed(-1791.0/65536.0,1,-nbitq), 
to_sfixed(-1752.0/65536.0,1,-nbitq), 
to_sfixed(206.0/65536.0,1,-nbitq), 
to_sfixed(-1274.0/65536.0,1,-nbitq), 
to_sfixed(-1702.0/65536.0,1,-nbitq), 
to_sfixed(2182.0/65536.0,1,-nbitq), 
to_sfixed(253.0/65536.0,1,-nbitq), 
to_sfixed(12.0/65536.0,1,-nbitq), 
to_sfixed(550.0/65536.0,1,-nbitq), 
to_sfixed(-353.0/65536.0,1,-nbitq), 
to_sfixed(1891.0/65536.0,1,-nbitq), 
to_sfixed(4334.0/65536.0,1,-nbitq), 
to_sfixed(-657.0/65536.0,1,-nbitq), 
to_sfixed(19.0/65536.0,1,-nbitq), 
to_sfixed(-1964.0/65536.0,1,-nbitq), 
to_sfixed(-955.0/65536.0,1,-nbitq), 
to_sfixed(587.0/65536.0,1,-nbitq), 
to_sfixed(2146.0/65536.0,1,-nbitq), 
to_sfixed(3212.0/65536.0,1,-nbitq), 
to_sfixed(-3024.0/65536.0,1,-nbitq), 
to_sfixed(1556.0/65536.0,1,-nbitq), 
to_sfixed(78.0/65536.0,1,-nbitq), 
to_sfixed(-2754.0/65536.0,1,-nbitq), 
to_sfixed(-648.0/65536.0,1,-nbitq), 
to_sfixed(-2218.0/65536.0,1,-nbitq), 
to_sfixed(4526.0/65536.0,1,-nbitq), 
to_sfixed(-2094.0/65536.0,1,-nbitq), 
to_sfixed(-61.0/65536.0,1,-nbitq), 
to_sfixed(-1857.0/65536.0,1,-nbitq), 
to_sfixed(221.0/65536.0,1,-nbitq), 
to_sfixed(-558.0/65536.0,1,-nbitq), 
to_sfixed(651.0/65536.0,1,-nbitq), 
to_sfixed(1577.0/65536.0,1,-nbitq), 
to_sfixed(-142.0/65536.0,1,-nbitq), 
to_sfixed(1003.0/65536.0,1,-nbitq), 
to_sfixed(-2253.0/65536.0,1,-nbitq), 
to_sfixed(-1369.0/65536.0,1,-nbitq), 
to_sfixed(2820.0/65536.0,1,-nbitq), 
to_sfixed(-802.0/65536.0,1,-nbitq), 
to_sfixed(1634.0/65536.0,1,-nbitq), 
to_sfixed(31.0/65536.0,1,-nbitq), 
to_sfixed(4187.0/65536.0,1,-nbitq), 
to_sfixed(-3579.0/65536.0,1,-nbitq), 
to_sfixed(2254.0/65536.0,1,-nbitq), 
to_sfixed(-2548.0/65536.0,1,-nbitq), 
to_sfixed(5317.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3455.0/65536.0,1,-nbitq), 
to_sfixed(2174.0/65536.0,1,-nbitq), 
to_sfixed(4484.0/65536.0,1,-nbitq), 
to_sfixed(1557.0/65536.0,1,-nbitq), 
to_sfixed(-4793.0/65536.0,1,-nbitq), 
to_sfixed(-2716.0/65536.0,1,-nbitq), 
to_sfixed(-1759.0/65536.0,1,-nbitq), 
to_sfixed(1309.0/65536.0,1,-nbitq), 
to_sfixed(-1114.0/65536.0,1,-nbitq), 
to_sfixed(2527.0/65536.0,1,-nbitq), 
to_sfixed(-2905.0/65536.0,1,-nbitq), 
to_sfixed(-3537.0/65536.0,1,-nbitq), 
to_sfixed(-2222.0/65536.0,1,-nbitq), 
to_sfixed(-4126.0/65536.0,1,-nbitq), 
to_sfixed(2766.0/65536.0,1,-nbitq), 
to_sfixed(683.0/65536.0,1,-nbitq), 
to_sfixed(191.0/65536.0,1,-nbitq), 
to_sfixed(-2022.0/65536.0,1,-nbitq), 
to_sfixed(3396.0/65536.0,1,-nbitq), 
to_sfixed(1211.0/65536.0,1,-nbitq), 
to_sfixed(-1815.0/65536.0,1,-nbitq), 
to_sfixed(958.0/65536.0,1,-nbitq), 
to_sfixed(-688.0/65536.0,1,-nbitq), 
to_sfixed(-1261.0/65536.0,1,-nbitq), 
to_sfixed(-1419.0/65536.0,1,-nbitq), 
to_sfixed(-2069.0/65536.0,1,-nbitq), 
to_sfixed(-3087.0/65536.0,1,-nbitq), 
to_sfixed(-2512.0/65536.0,1,-nbitq), 
to_sfixed(-1262.0/65536.0,1,-nbitq), 
to_sfixed(-3566.0/65536.0,1,-nbitq), 
to_sfixed(2489.0/65536.0,1,-nbitq), 
to_sfixed(2628.0/65536.0,1,-nbitq), 
to_sfixed(-2879.0/65536.0,1,-nbitq), 
to_sfixed(-2686.0/65536.0,1,-nbitq), 
to_sfixed(-923.0/65536.0,1,-nbitq), 
to_sfixed(2045.0/65536.0,1,-nbitq), 
to_sfixed(-1151.0/65536.0,1,-nbitq), 
to_sfixed(-3575.0/65536.0,1,-nbitq), 
to_sfixed(1203.0/65536.0,1,-nbitq), 
to_sfixed(-545.0/65536.0,1,-nbitq), 
to_sfixed(-1243.0/65536.0,1,-nbitq), 
to_sfixed(-875.0/65536.0,1,-nbitq), 
to_sfixed(-4251.0/65536.0,1,-nbitq), 
to_sfixed(-1522.0/65536.0,1,-nbitq), 
to_sfixed(2984.0/65536.0,1,-nbitq), 
to_sfixed(5583.0/65536.0,1,-nbitq), 
to_sfixed(528.0/65536.0,1,-nbitq), 
to_sfixed(-3326.0/65536.0,1,-nbitq), 
to_sfixed(-1013.0/65536.0,1,-nbitq), 
to_sfixed(815.0/65536.0,1,-nbitq), 
to_sfixed(2310.0/65536.0,1,-nbitq), 
to_sfixed(-2481.0/65536.0,1,-nbitq), 
to_sfixed(-2156.0/65536.0,1,-nbitq), 
to_sfixed(-2809.0/65536.0,1,-nbitq), 
to_sfixed(2040.0/65536.0,1,-nbitq), 
to_sfixed(1586.0/65536.0,1,-nbitq), 
to_sfixed(1031.0/65536.0,1,-nbitq), 
to_sfixed(18.0/65536.0,1,-nbitq), 
to_sfixed(121.0/65536.0,1,-nbitq), 
to_sfixed(1536.0/65536.0,1,-nbitq), 
to_sfixed(732.0/65536.0,1,-nbitq), 
to_sfixed(-2043.0/65536.0,1,-nbitq), 
to_sfixed(1296.0/65536.0,1,-nbitq), 
to_sfixed(-2322.0/65536.0,1,-nbitq), 
to_sfixed(813.0/65536.0,1,-nbitq), 
to_sfixed(515.0/65536.0,1,-nbitq), 
to_sfixed(2130.0/65536.0,1,-nbitq), 
to_sfixed(-4680.0/65536.0,1,-nbitq), 
to_sfixed(4127.0/65536.0,1,-nbitq), 
to_sfixed(1876.0/65536.0,1,-nbitq), 
to_sfixed(157.0/65536.0,1,-nbitq), 
to_sfixed(-49.0/65536.0,1,-nbitq), 
to_sfixed(1015.0/65536.0,1,-nbitq), 
to_sfixed(-1455.0/65536.0,1,-nbitq), 
to_sfixed(-158.0/65536.0,1,-nbitq), 
to_sfixed(1164.0/65536.0,1,-nbitq), 
to_sfixed(976.0/65536.0,1,-nbitq), 
to_sfixed(4430.0/65536.0,1,-nbitq), 
to_sfixed(687.0/65536.0,1,-nbitq), 
to_sfixed(2028.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1489.0/65536.0,1,-nbitq), 
to_sfixed(337.0/65536.0,1,-nbitq), 
to_sfixed(1583.0/65536.0,1,-nbitq), 
to_sfixed(1983.0/65536.0,1,-nbitq), 
to_sfixed(616.0/65536.0,1,-nbitq), 
to_sfixed(-1761.0/65536.0,1,-nbitq), 
to_sfixed(154.0/65536.0,1,-nbitq), 
to_sfixed(54.0/65536.0,1,-nbitq), 
to_sfixed(-2256.0/65536.0,1,-nbitq), 
to_sfixed(-1067.0/65536.0,1,-nbitq), 
to_sfixed(-1156.0/65536.0,1,-nbitq), 
to_sfixed(-3434.0/65536.0,1,-nbitq), 
to_sfixed(1889.0/65536.0,1,-nbitq), 
to_sfixed(-3572.0/65536.0,1,-nbitq), 
to_sfixed(-1206.0/65536.0,1,-nbitq), 
to_sfixed(-1813.0/65536.0,1,-nbitq), 
to_sfixed(-1808.0/65536.0,1,-nbitq), 
to_sfixed(-252.0/65536.0,1,-nbitq), 
to_sfixed(-144.0/65536.0,1,-nbitq), 
to_sfixed(3018.0/65536.0,1,-nbitq), 
to_sfixed(-1341.0/65536.0,1,-nbitq), 
to_sfixed(-1312.0/65536.0,1,-nbitq), 
to_sfixed(2209.0/65536.0,1,-nbitq), 
to_sfixed(4104.0/65536.0,1,-nbitq), 
to_sfixed(-315.0/65536.0,1,-nbitq), 
to_sfixed(-2007.0/65536.0,1,-nbitq), 
to_sfixed(-2604.0/65536.0,1,-nbitq), 
to_sfixed(-1102.0/65536.0,1,-nbitq), 
to_sfixed(-396.0/65536.0,1,-nbitq), 
to_sfixed(-2275.0/65536.0,1,-nbitq), 
to_sfixed(686.0/65536.0,1,-nbitq), 
to_sfixed(1246.0/65536.0,1,-nbitq), 
to_sfixed(-4462.0/65536.0,1,-nbitq), 
to_sfixed(-4867.0/65536.0,1,-nbitq), 
to_sfixed(-1172.0/65536.0,1,-nbitq), 
to_sfixed(-1362.0/65536.0,1,-nbitq), 
to_sfixed(-866.0/65536.0,1,-nbitq), 
to_sfixed(-1210.0/65536.0,1,-nbitq), 
to_sfixed(-3384.0/65536.0,1,-nbitq), 
to_sfixed(-1428.0/65536.0,1,-nbitq), 
to_sfixed(1883.0/65536.0,1,-nbitq), 
to_sfixed(-3153.0/65536.0,1,-nbitq), 
to_sfixed(827.0/65536.0,1,-nbitq), 
to_sfixed(2643.0/65536.0,1,-nbitq), 
to_sfixed(268.0/65536.0,1,-nbitq), 
to_sfixed(3298.0/65536.0,1,-nbitq), 
to_sfixed(-1403.0/65536.0,1,-nbitq), 
to_sfixed(-685.0/65536.0,1,-nbitq), 
to_sfixed(3322.0/65536.0,1,-nbitq), 
to_sfixed(1701.0/65536.0,1,-nbitq), 
to_sfixed(533.0/65536.0,1,-nbitq), 
to_sfixed(-1155.0/65536.0,1,-nbitq), 
to_sfixed(472.0/65536.0,1,-nbitq), 
to_sfixed(-145.0/65536.0,1,-nbitq), 
to_sfixed(2222.0/65536.0,1,-nbitq), 
to_sfixed(-356.0/65536.0,1,-nbitq), 
to_sfixed(-640.0/65536.0,1,-nbitq), 
to_sfixed(3284.0/65536.0,1,-nbitq), 
to_sfixed(-2984.0/65536.0,1,-nbitq), 
to_sfixed(5233.0/65536.0,1,-nbitq), 
to_sfixed(1728.0/65536.0,1,-nbitq), 
to_sfixed(1517.0/65536.0,1,-nbitq), 
to_sfixed(-2264.0/65536.0,1,-nbitq), 
to_sfixed(-1851.0/65536.0,1,-nbitq), 
to_sfixed(542.0/65536.0,1,-nbitq), 
to_sfixed(1342.0/65536.0,1,-nbitq), 
to_sfixed(-1715.0/65536.0,1,-nbitq), 
to_sfixed(-714.0/65536.0,1,-nbitq), 
to_sfixed(-1010.0/65536.0,1,-nbitq), 
to_sfixed(1154.0/65536.0,1,-nbitq), 
to_sfixed(256.0/65536.0,1,-nbitq), 
to_sfixed(1784.0/65536.0,1,-nbitq), 
to_sfixed(2646.0/65536.0,1,-nbitq), 
to_sfixed(2097.0/65536.0,1,-nbitq), 
to_sfixed(2137.0/65536.0,1,-nbitq), 
to_sfixed(64.0/65536.0,1,-nbitq), 
to_sfixed(502.0/65536.0,1,-nbitq), 
to_sfixed(562.0/65536.0,1,-nbitq), 
to_sfixed(-3015.0/65536.0,1,-nbitq), 
to_sfixed(4261.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-420.0/65536.0,1,-nbitq), 
to_sfixed(-338.0/65536.0,1,-nbitq), 
to_sfixed(4298.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(-278.0/65536.0,1,-nbitq), 
to_sfixed(357.0/65536.0,1,-nbitq), 
to_sfixed(1030.0/65536.0,1,-nbitq), 
to_sfixed(399.0/65536.0,1,-nbitq), 
to_sfixed(-2308.0/65536.0,1,-nbitq), 
to_sfixed(-1429.0/65536.0,1,-nbitq), 
to_sfixed(1329.0/65536.0,1,-nbitq), 
to_sfixed(-4404.0/65536.0,1,-nbitq), 
to_sfixed(-197.0/65536.0,1,-nbitq), 
to_sfixed(-3383.0/65536.0,1,-nbitq), 
to_sfixed(3404.0/65536.0,1,-nbitq), 
to_sfixed(1497.0/65536.0,1,-nbitq), 
to_sfixed(-121.0/65536.0,1,-nbitq), 
to_sfixed(646.0/65536.0,1,-nbitq), 
to_sfixed(-1793.0/65536.0,1,-nbitq), 
to_sfixed(1552.0/65536.0,1,-nbitq), 
to_sfixed(-3713.0/65536.0,1,-nbitq), 
to_sfixed(-2564.0/65536.0,1,-nbitq), 
to_sfixed(-119.0/65536.0,1,-nbitq), 
to_sfixed(-1135.0/65536.0,1,-nbitq), 
to_sfixed(1948.0/65536.0,1,-nbitq), 
to_sfixed(2560.0/65536.0,1,-nbitq), 
to_sfixed(184.0/65536.0,1,-nbitq), 
to_sfixed(-2064.0/65536.0,1,-nbitq), 
to_sfixed(-177.0/65536.0,1,-nbitq), 
to_sfixed(-762.0/65536.0,1,-nbitq), 
to_sfixed(2816.0/65536.0,1,-nbitq), 
to_sfixed(897.0/65536.0,1,-nbitq), 
to_sfixed(-1000.0/65536.0,1,-nbitq), 
to_sfixed(-2891.0/65536.0,1,-nbitq), 
to_sfixed(-366.0/65536.0,1,-nbitq), 
to_sfixed(1604.0/65536.0,1,-nbitq), 
to_sfixed(-3069.0/65536.0,1,-nbitq), 
to_sfixed(-3343.0/65536.0,1,-nbitq), 
to_sfixed(-3181.0/65536.0,1,-nbitq), 
to_sfixed(-697.0/65536.0,1,-nbitq), 
to_sfixed(1484.0/65536.0,1,-nbitq), 
to_sfixed(1558.0/65536.0,1,-nbitq), 
to_sfixed(-4403.0/65536.0,1,-nbitq), 
to_sfixed(1213.0/65536.0,1,-nbitq), 
to_sfixed(510.0/65536.0,1,-nbitq), 
to_sfixed(2341.0/65536.0,1,-nbitq), 
to_sfixed(1165.0/65536.0,1,-nbitq), 
to_sfixed(489.0/65536.0,1,-nbitq), 
to_sfixed(-669.0/65536.0,1,-nbitq), 
to_sfixed(861.0/65536.0,1,-nbitq), 
to_sfixed(-2464.0/65536.0,1,-nbitq), 
to_sfixed(3405.0/65536.0,1,-nbitq), 
to_sfixed(-1423.0/65536.0,1,-nbitq), 
to_sfixed(-3264.0/65536.0,1,-nbitq), 
to_sfixed(306.0/65536.0,1,-nbitq), 
to_sfixed(-1474.0/65536.0,1,-nbitq), 
to_sfixed(88.0/65536.0,1,-nbitq), 
to_sfixed(-801.0/65536.0,1,-nbitq), 
to_sfixed(2575.0/65536.0,1,-nbitq), 
to_sfixed(5582.0/65536.0,1,-nbitq), 
to_sfixed(-3456.0/65536.0,1,-nbitq), 
to_sfixed(1171.0/65536.0,1,-nbitq), 
to_sfixed(-1233.0/65536.0,1,-nbitq), 
to_sfixed(-876.0/65536.0,1,-nbitq), 
to_sfixed(1386.0/65536.0,1,-nbitq), 
to_sfixed(3343.0/65536.0,1,-nbitq), 
to_sfixed(-147.0/65536.0,1,-nbitq), 
to_sfixed(1378.0/65536.0,1,-nbitq), 
to_sfixed(-141.0/65536.0,1,-nbitq), 
to_sfixed(1434.0/65536.0,1,-nbitq), 
to_sfixed(1342.0/65536.0,1,-nbitq), 
to_sfixed(312.0/65536.0,1,-nbitq), 
to_sfixed(2517.0/65536.0,1,-nbitq), 
to_sfixed(685.0/65536.0,1,-nbitq), 
to_sfixed(-2122.0/65536.0,1,-nbitq), 
to_sfixed(-1216.0/65536.0,1,-nbitq), 
to_sfixed(2173.0/65536.0,1,-nbitq), 
to_sfixed(281.0/65536.0,1,-nbitq), 
to_sfixed(-3007.0/65536.0,1,-nbitq), 
to_sfixed(2849.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1916.0/65536.0,1,-nbitq), 
to_sfixed(721.0/65536.0,1,-nbitq), 
to_sfixed(-298.0/65536.0,1,-nbitq), 
to_sfixed(-1402.0/65536.0,1,-nbitq), 
to_sfixed(-1114.0/65536.0,1,-nbitq), 
to_sfixed(1165.0/65536.0,1,-nbitq), 
to_sfixed(-2996.0/65536.0,1,-nbitq), 
to_sfixed(2144.0/65536.0,1,-nbitq), 
to_sfixed(525.0/65536.0,1,-nbitq), 
to_sfixed(-626.0/65536.0,1,-nbitq), 
to_sfixed(-2805.0/65536.0,1,-nbitq), 
to_sfixed(-1716.0/65536.0,1,-nbitq), 
to_sfixed(-241.0/65536.0,1,-nbitq), 
to_sfixed(-3541.0/65536.0,1,-nbitq), 
to_sfixed(941.0/65536.0,1,-nbitq), 
to_sfixed(-1474.0/65536.0,1,-nbitq), 
to_sfixed(-834.0/65536.0,1,-nbitq), 
to_sfixed(1423.0/65536.0,1,-nbitq), 
to_sfixed(-799.0/65536.0,1,-nbitq), 
to_sfixed(-823.0/65536.0,1,-nbitq), 
to_sfixed(-290.0/65536.0,1,-nbitq), 
to_sfixed(-1664.0/65536.0,1,-nbitq), 
to_sfixed(1610.0/65536.0,1,-nbitq), 
to_sfixed(4182.0/65536.0,1,-nbitq), 
to_sfixed(1460.0/65536.0,1,-nbitq), 
to_sfixed(-243.0/65536.0,1,-nbitq), 
to_sfixed(-614.0/65536.0,1,-nbitq), 
to_sfixed(-2154.0/65536.0,1,-nbitq), 
to_sfixed(1130.0/65536.0,1,-nbitq), 
to_sfixed(1339.0/65536.0,1,-nbitq), 
to_sfixed(1835.0/65536.0,1,-nbitq), 
to_sfixed(-1464.0/65536.0,1,-nbitq), 
to_sfixed(-2167.0/65536.0,1,-nbitq), 
to_sfixed(-5174.0/65536.0,1,-nbitq), 
to_sfixed(-407.0/65536.0,1,-nbitq), 
to_sfixed(-1383.0/65536.0,1,-nbitq), 
to_sfixed(-2661.0/65536.0,1,-nbitq), 
to_sfixed(-3054.0/65536.0,1,-nbitq), 
to_sfixed(-1774.0/65536.0,1,-nbitq), 
to_sfixed(-2621.0/65536.0,1,-nbitq), 
to_sfixed(-89.0/65536.0,1,-nbitq), 
to_sfixed(-465.0/65536.0,1,-nbitq), 
to_sfixed(-530.0/65536.0,1,-nbitq), 
to_sfixed(3362.0/65536.0,1,-nbitq), 
to_sfixed(1181.0/65536.0,1,-nbitq), 
to_sfixed(15.0/65536.0,1,-nbitq), 
to_sfixed(-2338.0/65536.0,1,-nbitq), 
to_sfixed(-1447.0/65536.0,1,-nbitq), 
to_sfixed(746.0/65536.0,1,-nbitq), 
to_sfixed(2078.0/65536.0,1,-nbitq), 
to_sfixed(-143.0/65536.0,1,-nbitq), 
to_sfixed(2360.0/65536.0,1,-nbitq), 
to_sfixed(1954.0/65536.0,1,-nbitq), 
to_sfixed(1836.0/65536.0,1,-nbitq), 
to_sfixed(1360.0/65536.0,1,-nbitq), 
to_sfixed(-728.0/65536.0,1,-nbitq), 
to_sfixed(-2199.0/65536.0,1,-nbitq), 
to_sfixed(849.0/65536.0,1,-nbitq), 
to_sfixed(1525.0/65536.0,1,-nbitq), 
to_sfixed(2687.0/65536.0,1,-nbitq), 
to_sfixed(-3266.0/65536.0,1,-nbitq), 
to_sfixed(-1593.0/65536.0,1,-nbitq), 
to_sfixed(-1930.0/65536.0,1,-nbitq), 
to_sfixed(-1741.0/65536.0,1,-nbitq), 
to_sfixed(613.0/65536.0,1,-nbitq), 
to_sfixed(892.0/65536.0,1,-nbitq), 
to_sfixed(44.0/65536.0,1,-nbitq), 
to_sfixed(853.0/65536.0,1,-nbitq), 
to_sfixed(1036.0/65536.0,1,-nbitq), 
to_sfixed(2759.0/65536.0,1,-nbitq), 
to_sfixed(1198.0/65536.0,1,-nbitq), 
to_sfixed(2802.0/65536.0,1,-nbitq), 
to_sfixed(-321.0/65536.0,1,-nbitq), 
to_sfixed(742.0/65536.0,1,-nbitq), 
to_sfixed(-1456.0/65536.0,1,-nbitq), 
to_sfixed(2049.0/65536.0,1,-nbitq), 
to_sfixed(375.0/65536.0,1,-nbitq), 
to_sfixed(-509.0/65536.0,1,-nbitq), 
to_sfixed(-1674.0/65536.0,1,-nbitq), 
to_sfixed(628.0/65536.0,1,-nbitq)  ), 
( to_sfixed(512.0/65536.0,1,-nbitq), 
to_sfixed(1867.0/65536.0,1,-nbitq), 
to_sfixed(-31.0/65536.0,1,-nbitq), 
to_sfixed(1210.0/65536.0,1,-nbitq), 
to_sfixed(42.0/65536.0,1,-nbitq), 
to_sfixed(-4542.0/65536.0,1,-nbitq), 
to_sfixed(-471.0/65536.0,1,-nbitq), 
to_sfixed(-651.0/65536.0,1,-nbitq), 
to_sfixed(2218.0/65536.0,1,-nbitq), 
to_sfixed(-2838.0/65536.0,1,-nbitq), 
to_sfixed(-1100.0/65536.0,1,-nbitq), 
to_sfixed(-1419.0/65536.0,1,-nbitq), 
to_sfixed(-355.0/65536.0,1,-nbitq), 
to_sfixed(446.0/65536.0,1,-nbitq), 
to_sfixed(-856.0/65536.0,1,-nbitq), 
to_sfixed(1917.0/65536.0,1,-nbitq), 
to_sfixed(-304.0/65536.0,1,-nbitq), 
to_sfixed(-1672.0/65536.0,1,-nbitq), 
to_sfixed(-1551.0/65536.0,1,-nbitq), 
to_sfixed(1788.0/65536.0,1,-nbitq), 
to_sfixed(-1312.0/65536.0,1,-nbitq), 
to_sfixed(-2470.0/65536.0,1,-nbitq), 
to_sfixed(-1565.0/65536.0,1,-nbitq), 
to_sfixed(2026.0/65536.0,1,-nbitq), 
to_sfixed(-1689.0/65536.0,1,-nbitq), 
to_sfixed(2242.0/65536.0,1,-nbitq), 
to_sfixed(-2515.0/65536.0,1,-nbitq), 
to_sfixed(2777.0/65536.0,1,-nbitq), 
to_sfixed(-2928.0/65536.0,1,-nbitq), 
to_sfixed(672.0/65536.0,1,-nbitq), 
to_sfixed(-2166.0/65536.0,1,-nbitq), 
to_sfixed(-1336.0/65536.0,1,-nbitq), 
to_sfixed(-4636.0/65536.0,1,-nbitq), 
to_sfixed(-951.0/65536.0,1,-nbitq), 
to_sfixed(1142.0/65536.0,1,-nbitq), 
to_sfixed(46.0/65536.0,1,-nbitq), 
to_sfixed(-1173.0/65536.0,1,-nbitq), 
to_sfixed(-270.0/65536.0,1,-nbitq), 
to_sfixed(-370.0/65536.0,1,-nbitq), 
to_sfixed(917.0/65536.0,1,-nbitq), 
to_sfixed(-3.0/65536.0,1,-nbitq), 
to_sfixed(2421.0/65536.0,1,-nbitq), 
to_sfixed(-3512.0/65536.0,1,-nbitq), 
to_sfixed(3349.0/65536.0,1,-nbitq), 
to_sfixed(-1227.0/65536.0,1,-nbitq), 
to_sfixed(473.0/65536.0,1,-nbitq), 
to_sfixed(821.0/65536.0,1,-nbitq), 
to_sfixed(-576.0/65536.0,1,-nbitq), 
to_sfixed(314.0/65536.0,1,-nbitq), 
to_sfixed(2245.0/65536.0,1,-nbitq), 
to_sfixed(2005.0/65536.0,1,-nbitq), 
to_sfixed(-654.0/65536.0,1,-nbitq), 
to_sfixed(1657.0/65536.0,1,-nbitq), 
to_sfixed(-1531.0/65536.0,1,-nbitq), 
to_sfixed(3808.0/65536.0,1,-nbitq), 
to_sfixed(1865.0/65536.0,1,-nbitq), 
to_sfixed(-1296.0/65536.0,1,-nbitq), 
to_sfixed(859.0/65536.0,1,-nbitq), 
to_sfixed(340.0/65536.0,1,-nbitq), 
to_sfixed(3295.0/65536.0,1,-nbitq), 
to_sfixed(1230.0/65536.0,1,-nbitq), 
to_sfixed(-1599.0/65536.0,1,-nbitq), 
to_sfixed(-932.0/65536.0,1,-nbitq), 
to_sfixed(-2735.0/65536.0,1,-nbitq), 
to_sfixed(3389.0/65536.0,1,-nbitq), 
to_sfixed(1779.0/65536.0,1,-nbitq), 
to_sfixed(154.0/65536.0,1,-nbitq), 
to_sfixed(-403.0/65536.0,1,-nbitq), 
to_sfixed(919.0/65536.0,1,-nbitq), 
to_sfixed(568.0/65536.0,1,-nbitq), 
to_sfixed(589.0/65536.0,1,-nbitq), 
to_sfixed(1463.0/65536.0,1,-nbitq), 
to_sfixed(1353.0/65536.0,1,-nbitq), 
to_sfixed(2632.0/65536.0,1,-nbitq), 
to_sfixed(-1874.0/65536.0,1,-nbitq), 
to_sfixed(-1457.0/65536.0,1,-nbitq), 
to_sfixed(-3123.0/65536.0,1,-nbitq), 
to_sfixed(-755.0/65536.0,1,-nbitq), 
to_sfixed(-771.0/65536.0,1,-nbitq), 
to_sfixed(1788.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1515.0/65536.0,1,-nbitq), 
to_sfixed(1448.0/65536.0,1,-nbitq), 
to_sfixed(1168.0/65536.0,1,-nbitq), 
to_sfixed(1144.0/65536.0,1,-nbitq), 
to_sfixed(1811.0/65536.0,1,-nbitq), 
to_sfixed(1375.0/65536.0,1,-nbitq), 
to_sfixed(-2924.0/65536.0,1,-nbitq), 
to_sfixed(-2269.0/65536.0,1,-nbitq), 
to_sfixed(1327.0/65536.0,1,-nbitq), 
to_sfixed(-2291.0/65536.0,1,-nbitq), 
to_sfixed(-1265.0/65536.0,1,-nbitq), 
to_sfixed(-656.0/65536.0,1,-nbitq), 
to_sfixed(2014.0/65536.0,1,-nbitq), 
to_sfixed(-1495.0/65536.0,1,-nbitq), 
to_sfixed(52.0/65536.0,1,-nbitq), 
to_sfixed(1264.0/65536.0,1,-nbitq), 
to_sfixed(1375.0/65536.0,1,-nbitq), 
to_sfixed(1199.0/65536.0,1,-nbitq), 
to_sfixed(-900.0/65536.0,1,-nbitq), 
to_sfixed(-1667.0/65536.0,1,-nbitq), 
to_sfixed(-582.0/65536.0,1,-nbitq), 
to_sfixed(-1572.0/65536.0,1,-nbitq), 
to_sfixed(-3443.0/65536.0,1,-nbitq), 
to_sfixed(2732.0/65536.0,1,-nbitq), 
to_sfixed(-1384.0/65536.0,1,-nbitq), 
to_sfixed(676.0/65536.0,1,-nbitq), 
to_sfixed(-229.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(-978.0/65536.0,1,-nbitq), 
to_sfixed(-1374.0/65536.0,1,-nbitq), 
to_sfixed(1164.0/65536.0,1,-nbitq), 
to_sfixed(1527.0/65536.0,1,-nbitq), 
to_sfixed(-1901.0/65536.0,1,-nbitq), 
to_sfixed(-3563.0/65536.0,1,-nbitq), 
to_sfixed(-946.0/65536.0,1,-nbitq), 
to_sfixed(-575.0/65536.0,1,-nbitq), 
to_sfixed(-2187.0/65536.0,1,-nbitq), 
to_sfixed(-2866.0/65536.0,1,-nbitq), 
to_sfixed(1198.0/65536.0,1,-nbitq), 
to_sfixed(-651.0/65536.0,1,-nbitq), 
to_sfixed(1832.0/65536.0,1,-nbitq), 
to_sfixed(-957.0/65536.0,1,-nbitq), 
to_sfixed(-38.0/65536.0,1,-nbitq), 
to_sfixed(1581.0/65536.0,1,-nbitq), 
to_sfixed(2207.0/65536.0,1,-nbitq), 
to_sfixed(4170.0/65536.0,1,-nbitq), 
to_sfixed(-131.0/65536.0,1,-nbitq), 
to_sfixed(-2105.0/65536.0,1,-nbitq), 
to_sfixed(2301.0/65536.0,1,-nbitq), 
to_sfixed(3902.0/65536.0,1,-nbitq), 
to_sfixed(-615.0/65536.0,1,-nbitq), 
to_sfixed(1237.0/65536.0,1,-nbitq), 
to_sfixed(552.0/65536.0,1,-nbitq), 
to_sfixed(-296.0/65536.0,1,-nbitq), 
to_sfixed(4110.0/65536.0,1,-nbitq), 
to_sfixed(-2787.0/65536.0,1,-nbitq), 
to_sfixed(2246.0/65536.0,1,-nbitq), 
to_sfixed(3171.0/65536.0,1,-nbitq), 
to_sfixed(-106.0/65536.0,1,-nbitq), 
to_sfixed(6338.0/65536.0,1,-nbitq), 
to_sfixed(-497.0/65536.0,1,-nbitq), 
to_sfixed(-2236.0/65536.0,1,-nbitq), 
to_sfixed(-1639.0/65536.0,1,-nbitq), 
to_sfixed(-1014.0/65536.0,1,-nbitq), 
to_sfixed(2472.0/65536.0,1,-nbitq), 
to_sfixed(3024.0/65536.0,1,-nbitq), 
to_sfixed(1999.0/65536.0,1,-nbitq), 
to_sfixed(-2297.0/65536.0,1,-nbitq), 
to_sfixed(593.0/65536.0,1,-nbitq), 
to_sfixed(-3048.0/65536.0,1,-nbitq), 
to_sfixed(-1671.0/65536.0,1,-nbitq), 
to_sfixed(-2475.0/65536.0,1,-nbitq), 
to_sfixed(1672.0/65536.0,1,-nbitq), 
to_sfixed(-332.0/65536.0,1,-nbitq), 
to_sfixed(-2051.0/65536.0,1,-nbitq), 
to_sfixed(841.0/65536.0,1,-nbitq), 
to_sfixed(-3399.0/65536.0,1,-nbitq), 
to_sfixed(-957.0/65536.0,1,-nbitq), 
to_sfixed(1915.0/65536.0,1,-nbitq), 
to_sfixed(2469.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1936.0/65536.0,1,-nbitq), 
to_sfixed(1085.0/65536.0,1,-nbitq), 
to_sfixed(830.0/65536.0,1,-nbitq), 
to_sfixed(1552.0/65536.0,1,-nbitq), 
to_sfixed(1771.0/65536.0,1,-nbitq), 
to_sfixed(1537.0/65536.0,1,-nbitq), 
to_sfixed(-3799.0/65536.0,1,-nbitq), 
to_sfixed(1940.0/65536.0,1,-nbitq), 
to_sfixed(1185.0/65536.0,1,-nbitq), 
to_sfixed(2996.0/65536.0,1,-nbitq), 
to_sfixed(-1106.0/65536.0,1,-nbitq), 
to_sfixed(-835.0/65536.0,1,-nbitq), 
to_sfixed(1674.0/65536.0,1,-nbitq), 
to_sfixed(-2991.0/65536.0,1,-nbitq), 
to_sfixed(1130.0/65536.0,1,-nbitq), 
to_sfixed(2733.0/65536.0,1,-nbitq), 
to_sfixed(356.0/65536.0,1,-nbitq), 
to_sfixed(3068.0/65536.0,1,-nbitq), 
to_sfixed(1310.0/65536.0,1,-nbitq), 
to_sfixed(969.0/65536.0,1,-nbitq), 
to_sfixed(-2551.0/65536.0,1,-nbitq), 
to_sfixed(1176.0/65536.0,1,-nbitq), 
to_sfixed(-3449.0/65536.0,1,-nbitq), 
to_sfixed(1885.0/65536.0,1,-nbitq), 
to_sfixed(1053.0/65536.0,1,-nbitq), 
to_sfixed(2583.0/65536.0,1,-nbitq), 
to_sfixed(1389.0/65536.0,1,-nbitq), 
to_sfixed(3431.0/65536.0,1,-nbitq), 
to_sfixed(-973.0/65536.0,1,-nbitq), 
to_sfixed(-177.0/65536.0,1,-nbitq), 
to_sfixed(2628.0/65536.0,1,-nbitq), 
to_sfixed(981.0/65536.0,1,-nbitq), 
to_sfixed(-3636.0/65536.0,1,-nbitq), 
to_sfixed(-2719.0/65536.0,1,-nbitq), 
to_sfixed(2282.0/65536.0,1,-nbitq), 
to_sfixed(-188.0/65536.0,1,-nbitq), 
to_sfixed(1144.0/65536.0,1,-nbitq), 
to_sfixed(-3130.0/65536.0,1,-nbitq), 
to_sfixed(-1238.0/65536.0,1,-nbitq), 
to_sfixed(583.0/65536.0,1,-nbitq), 
to_sfixed(-3479.0/65536.0,1,-nbitq), 
to_sfixed(401.0/65536.0,1,-nbitq), 
to_sfixed(-2516.0/65536.0,1,-nbitq), 
to_sfixed(-522.0/65536.0,1,-nbitq), 
to_sfixed(298.0/65536.0,1,-nbitq), 
to_sfixed(696.0/65536.0,1,-nbitq), 
to_sfixed(-1155.0/65536.0,1,-nbitq), 
to_sfixed(-2090.0/65536.0,1,-nbitq), 
to_sfixed(-1515.0/65536.0,1,-nbitq), 
to_sfixed(-850.0/65536.0,1,-nbitq), 
to_sfixed(-2303.0/65536.0,1,-nbitq), 
to_sfixed(977.0/65536.0,1,-nbitq), 
to_sfixed(-774.0/65536.0,1,-nbitq), 
to_sfixed(-2958.0/65536.0,1,-nbitq), 
to_sfixed(3639.0/65536.0,1,-nbitq), 
to_sfixed(-1242.0/65536.0,1,-nbitq), 
to_sfixed(245.0/65536.0,1,-nbitq), 
to_sfixed(-207.0/65536.0,1,-nbitq), 
to_sfixed(-2513.0/65536.0,1,-nbitq), 
to_sfixed(4848.0/65536.0,1,-nbitq), 
to_sfixed(1083.0/65536.0,1,-nbitq), 
to_sfixed(1990.0/65536.0,1,-nbitq), 
to_sfixed(-1213.0/65536.0,1,-nbitq), 
to_sfixed(-2231.0/65536.0,1,-nbitq), 
to_sfixed(1416.0/65536.0,1,-nbitq), 
to_sfixed(1785.0/65536.0,1,-nbitq), 
to_sfixed(-263.0/65536.0,1,-nbitq), 
to_sfixed(-3054.0/65536.0,1,-nbitq), 
to_sfixed(3074.0/65536.0,1,-nbitq), 
to_sfixed(-3076.0/65536.0,1,-nbitq), 
to_sfixed(-1374.0/65536.0,1,-nbitq), 
to_sfixed(-3633.0/65536.0,1,-nbitq), 
to_sfixed(-1868.0/65536.0,1,-nbitq), 
to_sfixed(418.0/65536.0,1,-nbitq), 
to_sfixed(250.0/65536.0,1,-nbitq), 
to_sfixed(-1104.0/65536.0,1,-nbitq), 
to_sfixed(988.0/65536.0,1,-nbitq), 
to_sfixed(2926.0/65536.0,1,-nbitq), 
to_sfixed(1233.0/65536.0,1,-nbitq), 
to_sfixed(-583.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1636.0/65536.0,1,-nbitq), 
to_sfixed(2574.0/65536.0,1,-nbitq), 
to_sfixed(3175.0/65536.0,1,-nbitq), 
to_sfixed(1763.0/65536.0,1,-nbitq), 
to_sfixed(1224.0/65536.0,1,-nbitq), 
to_sfixed(-1306.0/65536.0,1,-nbitq), 
to_sfixed(-2463.0/65536.0,1,-nbitq), 
to_sfixed(-904.0/65536.0,1,-nbitq), 
to_sfixed(-1813.0/65536.0,1,-nbitq), 
to_sfixed(-2659.0/65536.0,1,-nbitq), 
to_sfixed(1603.0/65536.0,1,-nbitq), 
to_sfixed(-2088.0/65536.0,1,-nbitq), 
to_sfixed(-1307.0/65536.0,1,-nbitq), 
to_sfixed(-2306.0/65536.0,1,-nbitq), 
to_sfixed(1085.0/65536.0,1,-nbitq), 
to_sfixed(1195.0/65536.0,1,-nbitq), 
to_sfixed(-3039.0/65536.0,1,-nbitq), 
to_sfixed(3006.0/65536.0,1,-nbitq), 
to_sfixed(461.0/65536.0,1,-nbitq), 
to_sfixed(2596.0/65536.0,1,-nbitq), 
to_sfixed(-1946.0/65536.0,1,-nbitq), 
to_sfixed(-15.0/65536.0,1,-nbitq), 
to_sfixed(-3679.0/65536.0,1,-nbitq), 
to_sfixed(-871.0/65536.0,1,-nbitq), 
to_sfixed(992.0/65536.0,1,-nbitq), 
to_sfixed(124.0/65536.0,1,-nbitq), 
to_sfixed(1492.0/65536.0,1,-nbitq), 
to_sfixed(-1787.0/65536.0,1,-nbitq), 
to_sfixed(655.0/65536.0,1,-nbitq), 
to_sfixed(-420.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(3523.0/65536.0,1,-nbitq), 
to_sfixed(-1986.0/65536.0,1,-nbitq), 
to_sfixed(-1252.0/65536.0,1,-nbitq), 
to_sfixed(-138.0/65536.0,1,-nbitq), 
to_sfixed(1417.0/65536.0,1,-nbitq), 
to_sfixed(904.0/65536.0,1,-nbitq), 
to_sfixed(-3950.0/65536.0,1,-nbitq), 
to_sfixed(-3926.0/65536.0,1,-nbitq), 
to_sfixed(-995.0/65536.0,1,-nbitq), 
to_sfixed(-3406.0/65536.0,1,-nbitq), 
to_sfixed(-164.0/65536.0,1,-nbitq), 
to_sfixed(-2803.0/65536.0,1,-nbitq), 
to_sfixed(-35.0/65536.0,1,-nbitq), 
to_sfixed(-1384.0/65536.0,1,-nbitq), 
to_sfixed(4995.0/65536.0,1,-nbitq), 
to_sfixed(2212.0/65536.0,1,-nbitq), 
to_sfixed(-358.0/65536.0,1,-nbitq), 
to_sfixed(3042.0/65536.0,1,-nbitq), 
to_sfixed(-1301.0/65536.0,1,-nbitq), 
to_sfixed(1859.0/65536.0,1,-nbitq), 
to_sfixed(1692.0/65536.0,1,-nbitq), 
to_sfixed(640.0/65536.0,1,-nbitq), 
to_sfixed(-5067.0/65536.0,1,-nbitq), 
to_sfixed(2802.0/65536.0,1,-nbitq), 
to_sfixed(-2469.0/65536.0,1,-nbitq), 
to_sfixed(-2153.0/65536.0,1,-nbitq), 
to_sfixed(-1595.0/65536.0,1,-nbitq), 
to_sfixed(2165.0/65536.0,1,-nbitq), 
to_sfixed(2361.0/65536.0,1,-nbitq), 
to_sfixed(-2571.0/65536.0,1,-nbitq), 
to_sfixed(-2812.0/65536.0,1,-nbitq), 
to_sfixed(-180.0/65536.0,1,-nbitq), 
to_sfixed(-3410.0/65536.0,1,-nbitq), 
to_sfixed(3406.0/65536.0,1,-nbitq), 
to_sfixed(-996.0/65536.0,1,-nbitq), 
to_sfixed(-2149.0/65536.0,1,-nbitq), 
to_sfixed(-2497.0/65536.0,1,-nbitq), 
to_sfixed(305.0/65536.0,1,-nbitq), 
to_sfixed(-2826.0/65536.0,1,-nbitq), 
to_sfixed(4002.0/65536.0,1,-nbitq), 
to_sfixed(-2687.0/65536.0,1,-nbitq), 
to_sfixed(-1044.0/65536.0,1,-nbitq), 
to_sfixed(-2907.0/65536.0,1,-nbitq), 
to_sfixed(-1405.0/65536.0,1,-nbitq), 
to_sfixed(-930.0/65536.0,1,-nbitq), 
to_sfixed(-1679.0/65536.0,1,-nbitq), 
to_sfixed(3332.0/65536.0,1,-nbitq), 
to_sfixed(594.0/65536.0,1,-nbitq), 
to_sfixed(-262.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2911.0/65536.0,1,-nbitq), 
to_sfixed(1817.0/65536.0,1,-nbitq), 
to_sfixed(2927.0/65536.0,1,-nbitq), 
to_sfixed(-320.0/65536.0,1,-nbitq), 
to_sfixed(-2907.0/65536.0,1,-nbitq), 
to_sfixed(543.0/65536.0,1,-nbitq), 
to_sfixed(-1269.0/65536.0,1,-nbitq), 
to_sfixed(-1690.0/65536.0,1,-nbitq), 
to_sfixed(1482.0/65536.0,1,-nbitq), 
to_sfixed(-2780.0/65536.0,1,-nbitq), 
to_sfixed(-3713.0/65536.0,1,-nbitq), 
to_sfixed(-22.0/65536.0,1,-nbitq), 
to_sfixed(498.0/65536.0,1,-nbitq), 
to_sfixed(-1488.0/65536.0,1,-nbitq), 
to_sfixed(2980.0/65536.0,1,-nbitq), 
to_sfixed(1549.0/65536.0,1,-nbitq), 
to_sfixed(1623.0/65536.0,1,-nbitq), 
to_sfixed(-641.0/65536.0,1,-nbitq), 
to_sfixed(1631.0/65536.0,1,-nbitq), 
to_sfixed(804.0/65536.0,1,-nbitq), 
to_sfixed(-1705.0/65536.0,1,-nbitq), 
to_sfixed(-2193.0/65536.0,1,-nbitq), 
to_sfixed(874.0/65536.0,1,-nbitq), 
to_sfixed(-53.0/65536.0,1,-nbitq), 
to_sfixed(657.0/65536.0,1,-nbitq), 
to_sfixed(2452.0/65536.0,1,-nbitq), 
to_sfixed(-3308.0/65536.0,1,-nbitq), 
to_sfixed(-2029.0/65536.0,1,-nbitq), 
to_sfixed(-1417.0/65536.0,1,-nbitq), 
to_sfixed(-741.0/65536.0,1,-nbitq), 
to_sfixed(2730.0/65536.0,1,-nbitq), 
to_sfixed(2233.0/65536.0,1,-nbitq), 
to_sfixed(346.0/65536.0,1,-nbitq), 
to_sfixed(-3636.0/65536.0,1,-nbitq), 
to_sfixed(-2514.0/65536.0,1,-nbitq), 
to_sfixed(-2543.0/65536.0,1,-nbitq), 
to_sfixed(926.0/65536.0,1,-nbitq), 
to_sfixed(973.0/65536.0,1,-nbitq), 
to_sfixed(-914.0/65536.0,1,-nbitq), 
to_sfixed(-2264.0/65536.0,1,-nbitq), 
to_sfixed(616.0/65536.0,1,-nbitq), 
to_sfixed(-2668.0/65536.0,1,-nbitq), 
to_sfixed(-4357.0/65536.0,1,-nbitq), 
to_sfixed(2369.0/65536.0,1,-nbitq), 
to_sfixed(-667.0/65536.0,1,-nbitq), 
to_sfixed(3543.0/65536.0,1,-nbitq), 
to_sfixed(2656.0/65536.0,1,-nbitq), 
to_sfixed(338.0/65536.0,1,-nbitq), 
to_sfixed(2021.0/65536.0,1,-nbitq), 
to_sfixed(-323.0/65536.0,1,-nbitq), 
to_sfixed(1797.0/65536.0,1,-nbitq), 
to_sfixed(3232.0/65536.0,1,-nbitq), 
to_sfixed(2351.0/65536.0,1,-nbitq), 
to_sfixed(-5663.0/65536.0,1,-nbitq), 
to_sfixed(1328.0/65536.0,1,-nbitq), 
to_sfixed(-1940.0/65536.0,1,-nbitq), 
to_sfixed(1130.0/65536.0,1,-nbitq), 
to_sfixed(893.0/65536.0,1,-nbitq), 
to_sfixed(1532.0/65536.0,1,-nbitq), 
to_sfixed(4017.0/65536.0,1,-nbitq), 
to_sfixed(-2865.0/65536.0,1,-nbitq), 
to_sfixed(-2626.0/65536.0,1,-nbitq), 
to_sfixed(1817.0/65536.0,1,-nbitq), 
to_sfixed(-2237.0/65536.0,1,-nbitq), 
to_sfixed(461.0/65536.0,1,-nbitq), 
to_sfixed(1198.0/65536.0,1,-nbitq), 
to_sfixed(-1317.0/65536.0,1,-nbitq), 
to_sfixed(-464.0/65536.0,1,-nbitq), 
to_sfixed(644.0/65536.0,1,-nbitq), 
to_sfixed(-2639.0/65536.0,1,-nbitq), 
to_sfixed(2837.0/65536.0,1,-nbitq), 
to_sfixed(-3742.0/65536.0,1,-nbitq), 
to_sfixed(-1112.0/65536.0,1,-nbitq), 
to_sfixed(-1863.0/65536.0,1,-nbitq), 
to_sfixed(-34.0/65536.0,1,-nbitq), 
to_sfixed(-672.0/65536.0,1,-nbitq), 
to_sfixed(-2325.0/65536.0,1,-nbitq), 
to_sfixed(-232.0/65536.0,1,-nbitq), 
to_sfixed(-2522.0/65536.0,1,-nbitq), 
to_sfixed(4215.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1698.0/65536.0,1,-nbitq), 
to_sfixed(847.0/65536.0,1,-nbitq), 
to_sfixed(3569.0/65536.0,1,-nbitq), 
to_sfixed(-1004.0/65536.0,1,-nbitq), 
to_sfixed(21.0/65536.0,1,-nbitq), 
to_sfixed(21.0/65536.0,1,-nbitq), 
to_sfixed(-534.0/65536.0,1,-nbitq), 
to_sfixed(402.0/65536.0,1,-nbitq), 
to_sfixed(-2747.0/65536.0,1,-nbitq), 
to_sfixed(2664.0/65536.0,1,-nbitq), 
to_sfixed(-2842.0/65536.0,1,-nbitq), 
to_sfixed(-2938.0/65536.0,1,-nbitq), 
to_sfixed(1631.0/65536.0,1,-nbitq), 
to_sfixed(-2107.0/65536.0,1,-nbitq), 
to_sfixed(3261.0/65536.0,1,-nbitq), 
to_sfixed(-393.0/65536.0,1,-nbitq), 
to_sfixed(-1517.0/65536.0,1,-nbitq), 
to_sfixed(-2399.0/65536.0,1,-nbitq), 
to_sfixed(1845.0/65536.0,1,-nbitq), 
to_sfixed(47.0/65536.0,1,-nbitq), 
to_sfixed(-1412.0/65536.0,1,-nbitq), 
to_sfixed(1264.0/65536.0,1,-nbitq), 
to_sfixed(-3168.0/65536.0,1,-nbitq), 
to_sfixed(-150.0/65536.0,1,-nbitq), 
to_sfixed(1691.0/65536.0,1,-nbitq), 
to_sfixed(1972.0/65536.0,1,-nbitq), 
to_sfixed(-3257.0/65536.0,1,-nbitq), 
to_sfixed(-2421.0/65536.0,1,-nbitq), 
to_sfixed(-3966.0/65536.0,1,-nbitq), 
to_sfixed(-3626.0/65536.0,1,-nbitq), 
to_sfixed(-13.0/65536.0,1,-nbitq), 
to_sfixed(1225.0/65536.0,1,-nbitq), 
to_sfixed(82.0/65536.0,1,-nbitq), 
to_sfixed(-1006.0/65536.0,1,-nbitq), 
to_sfixed(-2279.0/65536.0,1,-nbitq), 
to_sfixed(653.0/65536.0,1,-nbitq), 
to_sfixed(-3088.0/65536.0,1,-nbitq), 
to_sfixed(-3926.0/65536.0,1,-nbitq), 
to_sfixed(-4139.0/65536.0,1,-nbitq), 
to_sfixed(-2083.0/65536.0,1,-nbitq), 
to_sfixed(-2599.0/65536.0,1,-nbitq), 
to_sfixed(-2146.0/65536.0,1,-nbitq), 
to_sfixed(-3286.0/65536.0,1,-nbitq), 
to_sfixed(-151.0/65536.0,1,-nbitq), 
to_sfixed(-1335.0/65536.0,1,-nbitq), 
to_sfixed(1213.0/65536.0,1,-nbitq), 
to_sfixed(3323.0/65536.0,1,-nbitq), 
to_sfixed(946.0/65536.0,1,-nbitq), 
to_sfixed(928.0/65536.0,1,-nbitq), 
to_sfixed(-367.0/65536.0,1,-nbitq), 
to_sfixed(-1300.0/65536.0,1,-nbitq), 
to_sfixed(-2202.0/65536.0,1,-nbitq), 
to_sfixed(2402.0/65536.0,1,-nbitq), 
to_sfixed(-1667.0/65536.0,1,-nbitq), 
to_sfixed(2416.0/65536.0,1,-nbitq), 
to_sfixed(-2165.0/65536.0,1,-nbitq), 
to_sfixed(-1935.0/65536.0,1,-nbitq), 
to_sfixed(1111.0/65536.0,1,-nbitq), 
to_sfixed(2730.0/65536.0,1,-nbitq), 
to_sfixed(2399.0/65536.0,1,-nbitq), 
to_sfixed(-2605.0/65536.0,1,-nbitq), 
to_sfixed(-819.0/65536.0,1,-nbitq), 
to_sfixed(-2409.0/65536.0,1,-nbitq), 
to_sfixed(675.0/65536.0,1,-nbitq), 
to_sfixed(633.0/65536.0,1,-nbitq), 
to_sfixed(3736.0/65536.0,1,-nbitq), 
to_sfixed(-235.0/65536.0,1,-nbitq), 
to_sfixed(-740.0/65536.0,1,-nbitq), 
to_sfixed(-1099.0/65536.0,1,-nbitq), 
to_sfixed(-1371.0/65536.0,1,-nbitq), 
to_sfixed(-1104.0/65536.0,1,-nbitq), 
to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(2601.0/65536.0,1,-nbitq), 
to_sfixed(-1189.0/65536.0,1,-nbitq), 
to_sfixed(866.0/65536.0,1,-nbitq), 
to_sfixed(412.0/65536.0,1,-nbitq), 
to_sfixed(-1824.0/65536.0,1,-nbitq), 
to_sfixed(4517.0/65536.0,1,-nbitq), 
to_sfixed(403.0/65536.0,1,-nbitq), 
to_sfixed(1613.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1895.0/65536.0,1,-nbitq), 
to_sfixed(-341.0/65536.0,1,-nbitq), 
to_sfixed(564.0/65536.0,1,-nbitq), 
to_sfixed(-1436.0/65536.0,1,-nbitq), 
to_sfixed(-1227.0/65536.0,1,-nbitq), 
to_sfixed(-274.0/65536.0,1,-nbitq), 
to_sfixed(-589.0/65536.0,1,-nbitq), 
to_sfixed(-1025.0/65536.0,1,-nbitq), 
to_sfixed(-2949.0/65536.0,1,-nbitq), 
to_sfixed(-2701.0/65536.0,1,-nbitq), 
to_sfixed(-2342.0/65536.0,1,-nbitq), 
to_sfixed(-3459.0/65536.0,1,-nbitq), 
to_sfixed(777.0/65536.0,1,-nbitq), 
to_sfixed(334.0/65536.0,1,-nbitq), 
to_sfixed(4168.0/65536.0,1,-nbitq), 
to_sfixed(-79.0/65536.0,1,-nbitq), 
to_sfixed(-1730.0/65536.0,1,-nbitq), 
to_sfixed(1801.0/65536.0,1,-nbitq), 
to_sfixed(2489.0/65536.0,1,-nbitq), 
to_sfixed(1933.0/65536.0,1,-nbitq), 
to_sfixed(-122.0/65536.0,1,-nbitq), 
to_sfixed(-1490.0/65536.0,1,-nbitq), 
to_sfixed(741.0/65536.0,1,-nbitq), 
to_sfixed(829.0/65536.0,1,-nbitq), 
to_sfixed(-1660.0/65536.0,1,-nbitq), 
to_sfixed(-1637.0/65536.0,1,-nbitq), 
to_sfixed(899.0/65536.0,1,-nbitq), 
to_sfixed(-2229.0/65536.0,1,-nbitq), 
to_sfixed(-3598.0/65536.0,1,-nbitq), 
to_sfixed(16.0/65536.0,1,-nbitq), 
to_sfixed(2793.0/65536.0,1,-nbitq), 
to_sfixed(266.0/65536.0,1,-nbitq), 
to_sfixed(-315.0/65536.0,1,-nbitq), 
to_sfixed(-2978.0/65536.0,1,-nbitq), 
to_sfixed(2895.0/65536.0,1,-nbitq), 
to_sfixed(147.0/65536.0,1,-nbitq), 
to_sfixed(123.0/65536.0,1,-nbitq), 
to_sfixed(-4609.0/65536.0,1,-nbitq), 
to_sfixed(285.0/65536.0,1,-nbitq), 
to_sfixed(1715.0/65536.0,1,-nbitq), 
to_sfixed(-2853.0/65536.0,1,-nbitq), 
to_sfixed(-146.0/65536.0,1,-nbitq), 
to_sfixed(-3564.0/65536.0,1,-nbitq), 
to_sfixed(812.0/65536.0,1,-nbitq), 
to_sfixed(-250.0/65536.0,1,-nbitq), 
to_sfixed(2378.0/65536.0,1,-nbitq), 
to_sfixed(-1147.0/65536.0,1,-nbitq), 
to_sfixed(-1653.0/65536.0,1,-nbitq), 
to_sfixed(-2254.0/65536.0,1,-nbitq), 
to_sfixed(4195.0/65536.0,1,-nbitq), 
to_sfixed(1316.0/65536.0,1,-nbitq), 
to_sfixed(2829.0/65536.0,1,-nbitq), 
to_sfixed(-2748.0/65536.0,1,-nbitq), 
to_sfixed(-88.0/65536.0,1,-nbitq), 
to_sfixed(3795.0/65536.0,1,-nbitq), 
to_sfixed(-446.0/65536.0,1,-nbitq), 
to_sfixed(-282.0/65536.0,1,-nbitq), 
to_sfixed(-1156.0/65536.0,1,-nbitq), 
to_sfixed(1242.0/65536.0,1,-nbitq), 
to_sfixed(2436.0/65536.0,1,-nbitq), 
to_sfixed(-4346.0/65536.0,1,-nbitq), 
to_sfixed(1354.0/65536.0,1,-nbitq), 
to_sfixed(1204.0/65536.0,1,-nbitq), 
to_sfixed(860.0/65536.0,1,-nbitq), 
to_sfixed(2137.0/65536.0,1,-nbitq), 
to_sfixed(1048.0/65536.0,1,-nbitq), 
to_sfixed(-227.0/65536.0,1,-nbitq), 
to_sfixed(733.0/65536.0,1,-nbitq), 
to_sfixed(-3.0/65536.0,1,-nbitq), 
to_sfixed(1066.0/65536.0,1,-nbitq), 
to_sfixed(2270.0/65536.0,1,-nbitq), 
to_sfixed(2053.0/65536.0,1,-nbitq), 
to_sfixed(497.0/65536.0,1,-nbitq), 
to_sfixed(505.0/65536.0,1,-nbitq), 
to_sfixed(2436.0/65536.0,1,-nbitq), 
to_sfixed(1296.0/65536.0,1,-nbitq), 
to_sfixed(-4717.0/65536.0,1,-nbitq), 
to_sfixed(5390.0/65536.0,1,-nbitq), 
to_sfixed(607.0/65536.0,1,-nbitq), 
to_sfixed(1823.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2243.0/65536.0,1,-nbitq), 
to_sfixed(-1846.0/65536.0,1,-nbitq), 
to_sfixed(2454.0/65536.0,1,-nbitq), 
to_sfixed(34.0/65536.0,1,-nbitq), 
to_sfixed(-2326.0/65536.0,1,-nbitq), 
to_sfixed(-3814.0/65536.0,1,-nbitq), 
to_sfixed(-3012.0/65536.0,1,-nbitq), 
to_sfixed(-1026.0/65536.0,1,-nbitq), 
to_sfixed(-2776.0/65536.0,1,-nbitq), 
to_sfixed(1438.0/65536.0,1,-nbitq), 
to_sfixed(-2177.0/65536.0,1,-nbitq), 
to_sfixed(-721.0/65536.0,1,-nbitq), 
to_sfixed(1253.0/65536.0,1,-nbitq), 
to_sfixed(-2109.0/65536.0,1,-nbitq), 
to_sfixed(-488.0/65536.0,1,-nbitq), 
to_sfixed(2945.0/65536.0,1,-nbitq), 
to_sfixed(-1593.0/65536.0,1,-nbitq), 
to_sfixed(2767.0/65536.0,1,-nbitq), 
to_sfixed(-688.0/65536.0,1,-nbitq), 
to_sfixed(-289.0/65536.0,1,-nbitq), 
to_sfixed(-4117.0/65536.0,1,-nbitq), 
to_sfixed(1961.0/65536.0,1,-nbitq), 
to_sfixed(-1950.0/65536.0,1,-nbitq), 
to_sfixed(-1600.0/65536.0,1,-nbitq), 
to_sfixed(1493.0/65536.0,1,-nbitq), 
to_sfixed(40.0/65536.0,1,-nbitq), 
to_sfixed(-145.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(-727.0/65536.0,1,-nbitq), 
to_sfixed(-3838.0/65536.0,1,-nbitq), 
to_sfixed(3216.0/65536.0,1,-nbitq), 
to_sfixed(2093.0/65536.0,1,-nbitq), 
to_sfixed(-623.0/65536.0,1,-nbitq), 
to_sfixed(693.0/65536.0,1,-nbitq), 
to_sfixed(-532.0/65536.0,1,-nbitq), 
to_sfixed(593.0/65536.0,1,-nbitq), 
to_sfixed(-617.0/65536.0,1,-nbitq), 
to_sfixed(-1683.0/65536.0,1,-nbitq), 
to_sfixed(-3171.0/65536.0,1,-nbitq), 
to_sfixed(-1391.0/65536.0,1,-nbitq), 
to_sfixed(-779.0/65536.0,1,-nbitq), 
to_sfixed(-1957.0/65536.0,1,-nbitq), 
to_sfixed(-657.0/65536.0,1,-nbitq), 
to_sfixed(3543.0/65536.0,1,-nbitq), 
to_sfixed(-2462.0/65536.0,1,-nbitq), 
to_sfixed(3137.0/65536.0,1,-nbitq), 
to_sfixed(-1658.0/65536.0,1,-nbitq), 
to_sfixed(1646.0/65536.0,1,-nbitq), 
to_sfixed(3501.0/65536.0,1,-nbitq), 
to_sfixed(-892.0/65536.0,1,-nbitq), 
to_sfixed(3008.0/65536.0,1,-nbitq), 
to_sfixed(-2893.0/65536.0,1,-nbitq), 
to_sfixed(210.0/65536.0,1,-nbitq), 
to_sfixed(-1098.0/65536.0,1,-nbitq), 
to_sfixed(1922.0/65536.0,1,-nbitq), 
to_sfixed(1751.0/65536.0,1,-nbitq), 
to_sfixed(2446.0/65536.0,1,-nbitq), 
to_sfixed(1143.0/65536.0,1,-nbitq), 
to_sfixed(-2522.0/65536.0,1,-nbitq), 
to_sfixed(2393.0/65536.0,1,-nbitq), 
to_sfixed(-4023.0/65536.0,1,-nbitq), 
to_sfixed(-2894.0/65536.0,1,-nbitq), 
to_sfixed(-2210.0/65536.0,1,-nbitq), 
to_sfixed(257.0/65536.0,1,-nbitq), 
to_sfixed(4093.0/65536.0,1,-nbitq), 
to_sfixed(985.0/65536.0,1,-nbitq), 
to_sfixed(-48.0/65536.0,1,-nbitq), 
to_sfixed(1915.0/65536.0,1,-nbitq), 
to_sfixed(3949.0/65536.0,1,-nbitq), 
to_sfixed(97.0/65536.0,1,-nbitq), 
to_sfixed(3456.0/65536.0,1,-nbitq), 
to_sfixed(2084.0/65536.0,1,-nbitq), 
to_sfixed(-676.0/65536.0,1,-nbitq), 
to_sfixed(664.0/65536.0,1,-nbitq), 
to_sfixed(-1797.0/65536.0,1,-nbitq), 
to_sfixed(260.0/65536.0,1,-nbitq), 
to_sfixed(-921.0/65536.0,1,-nbitq), 
to_sfixed(3640.0/65536.0,1,-nbitq), 
to_sfixed(-714.0/65536.0,1,-nbitq), 
to_sfixed(3395.0/65536.0,1,-nbitq)  ), 
( to_sfixed(899.0/65536.0,1,-nbitq), 
to_sfixed(286.0/65536.0,1,-nbitq), 
to_sfixed(1962.0/65536.0,1,-nbitq), 
to_sfixed(-91.0/65536.0,1,-nbitq), 
to_sfixed(-859.0/65536.0,1,-nbitq), 
to_sfixed(-3680.0/65536.0,1,-nbitq), 
to_sfixed(493.0/65536.0,1,-nbitq), 
to_sfixed(3157.0/65536.0,1,-nbitq), 
to_sfixed(-880.0/65536.0,1,-nbitq), 
to_sfixed(2889.0/65536.0,1,-nbitq), 
to_sfixed(-2548.0/65536.0,1,-nbitq), 
to_sfixed(145.0/65536.0,1,-nbitq), 
to_sfixed(-390.0/65536.0,1,-nbitq), 
to_sfixed(-2341.0/65536.0,1,-nbitq), 
to_sfixed(-62.0/65536.0,1,-nbitq), 
to_sfixed(-2119.0/65536.0,1,-nbitq), 
to_sfixed(-1339.0/65536.0,1,-nbitq), 
to_sfixed(2130.0/65536.0,1,-nbitq), 
to_sfixed(2930.0/65536.0,1,-nbitq), 
to_sfixed(1642.0/65536.0,1,-nbitq), 
to_sfixed(-4117.0/65536.0,1,-nbitq), 
to_sfixed(2719.0/65536.0,1,-nbitq), 
to_sfixed(2692.0/65536.0,1,-nbitq), 
to_sfixed(3451.0/65536.0,1,-nbitq), 
to_sfixed(-2543.0/65536.0,1,-nbitq), 
to_sfixed(603.0/65536.0,1,-nbitq), 
to_sfixed(29.0/65536.0,1,-nbitq), 
to_sfixed(1259.0/65536.0,1,-nbitq), 
to_sfixed(-3079.0/65536.0,1,-nbitq), 
to_sfixed(-2448.0/65536.0,1,-nbitq), 
to_sfixed(2493.0/65536.0,1,-nbitq), 
to_sfixed(501.0/65536.0,1,-nbitq), 
to_sfixed(-1845.0/65536.0,1,-nbitq), 
to_sfixed(-3416.0/65536.0,1,-nbitq), 
to_sfixed(-1841.0/65536.0,1,-nbitq), 
to_sfixed(1719.0/65536.0,1,-nbitq), 
to_sfixed(738.0/65536.0,1,-nbitq), 
to_sfixed(1125.0/65536.0,1,-nbitq), 
to_sfixed(-4730.0/65536.0,1,-nbitq), 
to_sfixed(-1833.0/65536.0,1,-nbitq), 
to_sfixed(-2705.0/65536.0,1,-nbitq), 
to_sfixed(-362.0/65536.0,1,-nbitq), 
to_sfixed(-3809.0/65536.0,1,-nbitq), 
to_sfixed(4210.0/65536.0,1,-nbitq), 
to_sfixed(-2049.0/65536.0,1,-nbitq), 
to_sfixed(-89.0/65536.0,1,-nbitq), 
to_sfixed(1693.0/65536.0,1,-nbitq), 
to_sfixed(997.0/65536.0,1,-nbitq), 
to_sfixed(-553.0/65536.0,1,-nbitq), 
to_sfixed(-463.0/65536.0,1,-nbitq), 
to_sfixed(-549.0/65536.0,1,-nbitq), 
to_sfixed(-1619.0/65536.0,1,-nbitq), 
to_sfixed(181.0/65536.0,1,-nbitq), 
to_sfixed(-1369.0/65536.0,1,-nbitq), 
to_sfixed(2085.0/65536.0,1,-nbitq), 
to_sfixed(-2437.0/65536.0,1,-nbitq), 
to_sfixed(-631.0/65536.0,1,-nbitq), 
to_sfixed(-2425.0/65536.0,1,-nbitq), 
to_sfixed(-212.0/65536.0,1,-nbitq), 
to_sfixed(4162.0/65536.0,1,-nbitq), 
to_sfixed(1242.0/65536.0,1,-nbitq), 
to_sfixed(1613.0/65536.0,1,-nbitq), 
to_sfixed(83.0/65536.0,1,-nbitq), 
to_sfixed(1958.0/65536.0,1,-nbitq), 
to_sfixed(-1019.0/65536.0,1,-nbitq), 
to_sfixed(306.0/65536.0,1,-nbitq), 
to_sfixed(2945.0/65536.0,1,-nbitq), 
to_sfixed(1438.0/65536.0,1,-nbitq), 
to_sfixed(2269.0/65536.0,1,-nbitq), 
to_sfixed(-198.0/65536.0,1,-nbitq), 
to_sfixed(182.0/65536.0,1,-nbitq), 
to_sfixed(2776.0/65536.0,1,-nbitq), 
to_sfixed(-2247.0/65536.0,1,-nbitq), 
to_sfixed(1068.0/65536.0,1,-nbitq), 
to_sfixed(685.0/65536.0,1,-nbitq), 
to_sfixed(3040.0/65536.0,1,-nbitq), 
to_sfixed(-1778.0/65536.0,1,-nbitq), 
to_sfixed(4266.0/65536.0,1,-nbitq), 
to_sfixed(1835.0/65536.0,1,-nbitq), 
to_sfixed(1434.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-35.0/65536.0,1,-nbitq), 
to_sfixed(2657.0/65536.0,1,-nbitq), 
to_sfixed(1606.0/65536.0,1,-nbitq), 
to_sfixed(-1557.0/65536.0,1,-nbitq), 
to_sfixed(213.0/65536.0,1,-nbitq), 
to_sfixed(-1806.0/65536.0,1,-nbitq), 
to_sfixed(349.0/65536.0,1,-nbitq), 
to_sfixed(26.0/65536.0,1,-nbitq), 
to_sfixed(96.0/65536.0,1,-nbitq), 
to_sfixed(1254.0/65536.0,1,-nbitq), 
to_sfixed(1587.0/65536.0,1,-nbitq), 
to_sfixed(-2667.0/65536.0,1,-nbitq), 
to_sfixed(1860.0/65536.0,1,-nbitq), 
to_sfixed(342.0/65536.0,1,-nbitq), 
to_sfixed(4179.0/65536.0,1,-nbitq), 
to_sfixed(-2678.0/65536.0,1,-nbitq), 
to_sfixed(-1058.0/65536.0,1,-nbitq), 
to_sfixed(1932.0/65536.0,1,-nbitq), 
to_sfixed(-57.0/65536.0,1,-nbitq), 
to_sfixed(-1165.0/65536.0,1,-nbitq), 
to_sfixed(144.0/65536.0,1,-nbitq), 
to_sfixed(806.0/65536.0,1,-nbitq), 
to_sfixed(493.0/65536.0,1,-nbitq), 
to_sfixed(2646.0/65536.0,1,-nbitq), 
to_sfixed(-2569.0/65536.0,1,-nbitq), 
to_sfixed(552.0/65536.0,1,-nbitq), 
to_sfixed(-1681.0/65536.0,1,-nbitq), 
to_sfixed(-1448.0/65536.0,1,-nbitq), 
to_sfixed(-180.0/65536.0,1,-nbitq), 
to_sfixed(997.0/65536.0,1,-nbitq), 
to_sfixed(465.0/65536.0,1,-nbitq), 
to_sfixed(2218.0/65536.0,1,-nbitq), 
to_sfixed(-5010.0/65536.0,1,-nbitq), 
to_sfixed(-343.0/65536.0,1,-nbitq), 
to_sfixed(-2107.0/65536.0,1,-nbitq), 
to_sfixed(224.0/65536.0,1,-nbitq), 
to_sfixed(-1608.0/65536.0,1,-nbitq), 
to_sfixed(681.0/65536.0,1,-nbitq), 
to_sfixed(-2317.0/65536.0,1,-nbitq), 
to_sfixed(49.0/65536.0,1,-nbitq), 
to_sfixed(2036.0/65536.0,1,-nbitq), 
to_sfixed(-1192.0/65536.0,1,-nbitq), 
to_sfixed(-2254.0/65536.0,1,-nbitq), 
to_sfixed(5486.0/65536.0,1,-nbitq), 
to_sfixed(-2389.0/65536.0,1,-nbitq), 
to_sfixed(5444.0/65536.0,1,-nbitq), 
to_sfixed(-473.0/65536.0,1,-nbitq), 
to_sfixed(391.0/65536.0,1,-nbitq), 
to_sfixed(1070.0/65536.0,1,-nbitq), 
to_sfixed(2333.0/65536.0,1,-nbitq), 
to_sfixed(-419.0/65536.0,1,-nbitq), 
to_sfixed(1073.0/65536.0,1,-nbitq), 
to_sfixed(2788.0/65536.0,1,-nbitq), 
to_sfixed(-6698.0/65536.0,1,-nbitq), 
to_sfixed(-1430.0/65536.0,1,-nbitq), 
to_sfixed(2947.0/65536.0,1,-nbitq), 
to_sfixed(920.0/65536.0,1,-nbitq), 
to_sfixed(-1324.0/65536.0,1,-nbitq), 
to_sfixed(-780.0/65536.0,1,-nbitq), 
to_sfixed(2338.0/65536.0,1,-nbitq), 
to_sfixed(-2612.0/65536.0,1,-nbitq), 
to_sfixed(-1632.0/65536.0,1,-nbitq), 
to_sfixed(-848.0/65536.0,1,-nbitq), 
to_sfixed(-2520.0/65536.0,1,-nbitq), 
to_sfixed(105.0/65536.0,1,-nbitq), 
to_sfixed(-1643.0/65536.0,1,-nbitq), 
to_sfixed(2670.0/65536.0,1,-nbitq), 
to_sfixed(-3764.0/65536.0,1,-nbitq), 
to_sfixed(3450.0/65536.0,1,-nbitq), 
to_sfixed(-1252.0/65536.0,1,-nbitq), 
to_sfixed(-1371.0/65536.0,1,-nbitq), 
to_sfixed(-1317.0/65536.0,1,-nbitq), 
to_sfixed(1939.0/65536.0,1,-nbitq), 
to_sfixed(1448.0/65536.0,1,-nbitq), 
to_sfixed(97.0/65536.0,1,-nbitq), 
to_sfixed(1608.0/65536.0,1,-nbitq), 
to_sfixed(1663.0/65536.0,1,-nbitq), 
to_sfixed(-335.0/65536.0,1,-nbitq), 
to_sfixed(-1363.0/65536.0,1,-nbitq), 
to_sfixed(-431.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2143.0/65536.0,1,-nbitq), 
to_sfixed(843.0/65536.0,1,-nbitq), 
to_sfixed(2245.0/65536.0,1,-nbitq), 
to_sfixed(1754.0/65536.0,1,-nbitq), 
to_sfixed(699.0/65536.0,1,-nbitq), 
to_sfixed(-3406.0/65536.0,1,-nbitq), 
to_sfixed(1157.0/65536.0,1,-nbitq), 
to_sfixed(2562.0/65536.0,1,-nbitq), 
to_sfixed(-1055.0/65536.0,1,-nbitq), 
to_sfixed(361.0/65536.0,1,-nbitq), 
to_sfixed(1837.0/65536.0,1,-nbitq), 
to_sfixed(347.0/65536.0,1,-nbitq), 
to_sfixed(1865.0/65536.0,1,-nbitq), 
to_sfixed(-1005.0/65536.0,1,-nbitq), 
to_sfixed(1100.0/65536.0,1,-nbitq), 
to_sfixed(525.0/65536.0,1,-nbitq), 
to_sfixed(-1622.0/65536.0,1,-nbitq), 
to_sfixed(2601.0/65536.0,1,-nbitq), 
to_sfixed(1322.0/65536.0,1,-nbitq), 
to_sfixed(1352.0/65536.0,1,-nbitq), 
to_sfixed(-2371.0/65536.0,1,-nbitq), 
to_sfixed(-2386.0/65536.0,1,-nbitq), 
to_sfixed(-354.0/65536.0,1,-nbitq), 
to_sfixed(741.0/65536.0,1,-nbitq), 
to_sfixed(1764.0/65536.0,1,-nbitq), 
to_sfixed(3375.0/65536.0,1,-nbitq), 
to_sfixed(-463.0/65536.0,1,-nbitq), 
to_sfixed(-1672.0/65536.0,1,-nbitq), 
to_sfixed(-4402.0/65536.0,1,-nbitq), 
to_sfixed(-693.0/65536.0,1,-nbitq), 
to_sfixed(732.0/65536.0,1,-nbitq), 
to_sfixed(3557.0/65536.0,1,-nbitq), 
to_sfixed(-41.0/65536.0,1,-nbitq), 
to_sfixed(-3590.0/65536.0,1,-nbitq), 
to_sfixed(1866.0/65536.0,1,-nbitq), 
to_sfixed(2010.0/65536.0,1,-nbitq), 
to_sfixed(-192.0/65536.0,1,-nbitq), 
to_sfixed(1206.0/65536.0,1,-nbitq), 
to_sfixed(94.0/65536.0,1,-nbitq), 
to_sfixed(406.0/65536.0,1,-nbitq), 
to_sfixed(862.0/65536.0,1,-nbitq), 
to_sfixed(172.0/65536.0,1,-nbitq), 
to_sfixed(-4891.0/65536.0,1,-nbitq), 
to_sfixed(2706.0/65536.0,1,-nbitq), 
to_sfixed(1233.0/65536.0,1,-nbitq), 
to_sfixed(2734.0/65536.0,1,-nbitq), 
to_sfixed(658.0/65536.0,1,-nbitq), 
to_sfixed(2396.0/65536.0,1,-nbitq), 
to_sfixed(2522.0/65536.0,1,-nbitq), 
to_sfixed(3344.0/65536.0,1,-nbitq), 
to_sfixed(-351.0/65536.0,1,-nbitq), 
to_sfixed(945.0/65536.0,1,-nbitq), 
to_sfixed(3316.0/65536.0,1,-nbitq), 
to_sfixed(-1307.0/65536.0,1,-nbitq), 
to_sfixed(2118.0/65536.0,1,-nbitq), 
to_sfixed(-1602.0/65536.0,1,-nbitq), 
to_sfixed(936.0/65536.0,1,-nbitq), 
to_sfixed(-2318.0/65536.0,1,-nbitq), 
to_sfixed(-757.0/65536.0,1,-nbitq), 
to_sfixed(5580.0/65536.0,1,-nbitq), 
to_sfixed(1434.0/65536.0,1,-nbitq), 
to_sfixed(1619.0/65536.0,1,-nbitq), 
to_sfixed(78.0/65536.0,1,-nbitq), 
to_sfixed(1161.0/65536.0,1,-nbitq), 
to_sfixed(383.0/65536.0,1,-nbitq), 
to_sfixed(4128.0/65536.0,1,-nbitq), 
to_sfixed(3234.0/65536.0,1,-nbitq), 
to_sfixed(921.0/65536.0,1,-nbitq), 
to_sfixed(-133.0/65536.0,1,-nbitq), 
to_sfixed(-930.0/65536.0,1,-nbitq), 
to_sfixed(-101.0/65536.0,1,-nbitq), 
to_sfixed(1086.0/65536.0,1,-nbitq), 
to_sfixed(2952.0/65536.0,1,-nbitq), 
to_sfixed(2156.0/65536.0,1,-nbitq), 
to_sfixed(187.0/65536.0,1,-nbitq), 
to_sfixed(858.0/65536.0,1,-nbitq), 
to_sfixed(-2492.0/65536.0,1,-nbitq), 
to_sfixed(4578.0/65536.0,1,-nbitq), 
to_sfixed(-480.0/65536.0,1,-nbitq), 
to_sfixed(448.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2180.0/65536.0,1,-nbitq), 
to_sfixed(973.0/65536.0,1,-nbitq), 
to_sfixed(3613.0/65536.0,1,-nbitq), 
to_sfixed(-1860.0/65536.0,1,-nbitq), 
to_sfixed(1527.0/65536.0,1,-nbitq), 
to_sfixed(81.0/65536.0,1,-nbitq), 
to_sfixed(-3394.0/65536.0,1,-nbitq), 
to_sfixed(-183.0/65536.0,1,-nbitq), 
to_sfixed(-1107.0/65536.0,1,-nbitq), 
to_sfixed(1382.0/65536.0,1,-nbitq), 
to_sfixed(-2309.0/65536.0,1,-nbitq), 
to_sfixed(1581.0/65536.0,1,-nbitq), 
to_sfixed(1793.0/65536.0,1,-nbitq), 
to_sfixed(-1211.0/65536.0,1,-nbitq), 
to_sfixed(1322.0/65536.0,1,-nbitq), 
to_sfixed(1463.0/65536.0,1,-nbitq), 
to_sfixed(1893.0/65536.0,1,-nbitq), 
to_sfixed(1818.0/65536.0,1,-nbitq), 
to_sfixed(1743.0/65536.0,1,-nbitq), 
to_sfixed(-589.0/65536.0,1,-nbitq), 
to_sfixed(-1492.0/65536.0,1,-nbitq), 
to_sfixed(1010.0/65536.0,1,-nbitq), 
to_sfixed(2095.0/65536.0,1,-nbitq), 
to_sfixed(2885.0/65536.0,1,-nbitq), 
to_sfixed(-2959.0/65536.0,1,-nbitq), 
to_sfixed(2789.0/65536.0,1,-nbitq), 
to_sfixed(-1632.0/65536.0,1,-nbitq), 
to_sfixed(260.0/65536.0,1,-nbitq), 
to_sfixed(-3804.0/65536.0,1,-nbitq), 
to_sfixed(1043.0/65536.0,1,-nbitq), 
to_sfixed(437.0/65536.0,1,-nbitq), 
to_sfixed(-801.0/65536.0,1,-nbitq), 
to_sfixed(-3814.0/65536.0,1,-nbitq), 
to_sfixed(-3159.0/65536.0,1,-nbitq), 
to_sfixed(326.0/65536.0,1,-nbitq), 
to_sfixed(52.0/65536.0,1,-nbitq), 
to_sfixed(-1377.0/65536.0,1,-nbitq), 
to_sfixed(-1860.0/65536.0,1,-nbitq), 
to_sfixed(-2580.0/65536.0,1,-nbitq), 
to_sfixed(1082.0/65536.0,1,-nbitq), 
to_sfixed(2008.0/65536.0,1,-nbitq), 
to_sfixed(1060.0/65536.0,1,-nbitq), 
to_sfixed(-2665.0/65536.0,1,-nbitq), 
to_sfixed(4980.0/65536.0,1,-nbitq), 
to_sfixed(-1835.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(-1052.0/65536.0,1,-nbitq), 
to_sfixed(-2108.0/65536.0,1,-nbitq), 
to_sfixed(-481.0/65536.0,1,-nbitq), 
to_sfixed(8.0/65536.0,1,-nbitq), 
to_sfixed(-2489.0/65536.0,1,-nbitq), 
to_sfixed(610.0/65536.0,1,-nbitq), 
to_sfixed(-1475.0/65536.0,1,-nbitq), 
to_sfixed(-5665.0/65536.0,1,-nbitq), 
to_sfixed(1865.0/65536.0,1,-nbitq), 
to_sfixed(2331.0/65536.0,1,-nbitq), 
to_sfixed(2842.0/65536.0,1,-nbitq), 
to_sfixed(805.0/65536.0,1,-nbitq), 
to_sfixed(2834.0/65536.0,1,-nbitq), 
to_sfixed(4917.0/65536.0,1,-nbitq), 
to_sfixed(-1055.0/65536.0,1,-nbitq), 
to_sfixed(-1195.0/65536.0,1,-nbitq), 
to_sfixed(-255.0/65536.0,1,-nbitq), 
to_sfixed(-450.0/65536.0,1,-nbitq), 
to_sfixed(-1735.0/65536.0,1,-nbitq), 
to_sfixed(3596.0/65536.0,1,-nbitq), 
to_sfixed(-2142.0/65536.0,1,-nbitq), 
to_sfixed(-1580.0/65536.0,1,-nbitq), 
to_sfixed(2490.0/65536.0,1,-nbitq), 
to_sfixed(-965.0/65536.0,1,-nbitq), 
to_sfixed(2089.0/65536.0,1,-nbitq), 
to_sfixed(1186.0/65536.0,1,-nbitq), 
to_sfixed(2977.0/65536.0,1,-nbitq), 
to_sfixed(2259.0/65536.0,1,-nbitq), 
to_sfixed(-2009.0/65536.0,1,-nbitq), 
to_sfixed(-816.0/65536.0,1,-nbitq), 
to_sfixed(2209.0/65536.0,1,-nbitq), 
to_sfixed(2772.0/65536.0,1,-nbitq), 
to_sfixed(-161.0/65536.0,1,-nbitq), 
to_sfixed(2978.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1698.0/65536.0,1,-nbitq), 
to_sfixed(-478.0/65536.0,1,-nbitq), 
to_sfixed(-63.0/65536.0,1,-nbitq), 
to_sfixed(-927.0/65536.0,1,-nbitq), 
to_sfixed(157.0/65536.0,1,-nbitq), 
to_sfixed(1814.0/65536.0,1,-nbitq), 
to_sfixed(-232.0/65536.0,1,-nbitq), 
to_sfixed(1128.0/65536.0,1,-nbitq), 
to_sfixed(1547.0/65536.0,1,-nbitq), 
to_sfixed(-798.0/65536.0,1,-nbitq), 
to_sfixed(-892.0/65536.0,1,-nbitq), 
to_sfixed(-569.0/65536.0,1,-nbitq), 
to_sfixed(-2148.0/65536.0,1,-nbitq), 
to_sfixed(-229.0/65536.0,1,-nbitq), 
to_sfixed(2594.0/65536.0,1,-nbitq), 
to_sfixed(-47.0/65536.0,1,-nbitq), 
to_sfixed(1936.0/65536.0,1,-nbitq), 
to_sfixed(2535.0/65536.0,1,-nbitq), 
to_sfixed(412.0/65536.0,1,-nbitq), 
to_sfixed(185.0/65536.0,1,-nbitq), 
to_sfixed(-1906.0/65536.0,1,-nbitq), 
to_sfixed(1397.0/65536.0,1,-nbitq), 
to_sfixed(1196.0/65536.0,1,-nbitq), 
to_sfixed(1151.0/65536.0,1,-nbitq), 
to_sfixed(1078.0/65536.0,1,-nbitq), 
to_sfixed(4436.0/65536.0,1,-nbitq), 
to_sfixed(675.0/65536.0,1,-nbitq), 
to_sfixed(1874.0/65536.0,1,-nbitq), 
to_sfixed(-3826.0/65536.0,1,-nbitq), 
to_sfixed(-1171.0/65536.0,1,-nbitq), 
to_sfixed(1573.0/65536.0,1,-nbitq), 
to_sfixed(405.0/65536.0,1,-nbitq), 
to_sfixed(-5541.0/65536.0,1,-nbitq), 
to_sfixed(-4114.0/65536.0,1,-nbitq), 
to_sfixed(2070.0/65536.0,1,-nbitq), 
to_sfixed(-3144.0/65536.0,1,-nbitq), 
to_sfixed(1562.0/65536.0,1,-nbitq), 
to_sfixed(-3930.0/65536.0,1,-nbitq), 
to_sfixed(-1657.0/65536.0,1,-nbitq), 
to_sfixed(106.0/65536.0,1,-nbitq), 
to_sfixed(-2607.0/65536.0,1,-nbitq), 
to_sfixed(144.0/65536.0,1,-nbitq), 
to_sfixed(-4367.0/65536.0,1,-nbitq), 
to_sfixed(3924.0/65536.0,1,-nbitq), 
to_sfixed(951.0/65536.0,1,-nbitq), 
to_sfixed(-1.0/65536.0,1,-nbitq), 
to_sfixed(-1209.0/65536.0,1,-nbitq), 
to_sfixed(-1994.0/65536.0,1,-nbitq), 
to_sfixed(-2292.0/65536.0,1,-nbitq), 
to_sfixed(725.0/65536.0,1,-nbitq), 
to_sfixed(2370.0/65536.0,1,-nbitq), 
to_sfixed(1086.0/65536.0,1,-nbitq), 
to_sfixed(927.0/65536.0,1,-nbitq), 
to_sfixed(-1030.0/65536.0,1,-nbitq), 
to_sfixed(-1383.0/65536.0,1,-nbitq), 
to_sfixed(2717.0/65536.0,1,-nbitq), 
to_sfixed(-2317.0/65536.0,1,-nbitq), 
to_sfixed(471.0/65536.0,1,-nbitq), 
to_sfixed(-2360.0/65536.0,1,-nbitq), 
to_sfixed(4959.0/65536.0,1,-nbitq), 
to_sfixed(-4072.0/65536.0,1,-nbitq), 
to_sfixed(1355.0/65536.0,1,-nbitq), 
to_sfixed(2276.0/65536.0,1,-nbitq), 
to_sfixed(2131.0/65536.0,1,-nbitq), 
to_sfixed(3726.0/65536.0,1,-nbitq), 
to_sfixed(1062.0/65536.0,1,-nbitq), 
to_sfixed(-941.0/65536.0,1,-nbitq), 
to_sfixed(-3582.0/65536.0,1,-nbitq), 
to_sfixed(686.0/65536.0,1,-nbitq), 
to_sfixed(518.0/65536.0,1,-nbitq), 
to_sfixed(2963.0/65536.0,1,-nbitq), 
to_sfixed(-3278.0/65536.0,1,-nbitq), 
to_sfixed(1597.0/65536.0,1,-nbitq), 
to_sfixed(-204.0/65536.0,1,-nbitq), 
to_sfixed(-2127.0/65536.0,1,-nbitq), 
to_sfixed(3811.0/65536.0,1,-nbitq), 
to_sfixed(371.0/65536.0,1,-nbitq), 
to_sfixed(1908.0/65536.0,1,-nbitq), 
to_sfixed(2473.0/65536.0,1,-nbitq), 
to_sfixed(3253.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-709.0/65536.0,1,-nbitq), 
to_sfixed(1840.0/65536.0,1,-nbitq), 
to_sfixed(1652.0/65536.0,1,-nbitq), 
to_sfixed(-310.0/65536.0,1,-nbitq), 
to_sfixed(399.0/65536.0,1,-nbitq), 
to_sfixed(-2338.0/65536.0,1,-nbitq), 
to_sfixed(-2029.0/65536.0,1,-nbitq), 
to_sfixed(518.0/65536.0,1,-nbitq), 
to_sfixed(1647.0/65536.0,1,-nbitq), 
to_sfixed(-443.0/65536.0,1,-nbitq), 
to_sfixed(-3312.0/65536.0,1,-nbitq), 
to_sfixed(-1300.0/65536.0,1,-nbitq), 
to_sfixed(-1316.0/65536.0,1,-nbitq), 
to_sfixed(-1388.0/65536.0,1,-nbitq), 
to_sfixed(2508.0/65536.0,1,-nbitq), 
to_sfixed(-393.0/65536.0,1,-nbitq), 
to_sfixed(-816.0/65536.0,1,-nbitq), 
to_sfixed(378.0/65536.0,1,-nbitq), 
to_sfixed(-894.0/65536.0,1,-nbitq), 
to_sfixed(-975.0/65536.0,1,-nbitq), 
to_sfixed(-3756.0/65536.0,1,-nbitq), 
to_sfixed(-609.0/65536.0,1,-nbitq), 
to_sfixed(-1601.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(-549.0/65536.0,1,-nbitq), 
to_sfixed(-1323.0/65536.0,1,-nbitq), 
to_sfixed(-1156.0/65536.0,1,-nbitq), 
to_sfixed(1417.0/65536.0,1,-nbitq), 
to_sfixed(-2302.0/65536.0,1,-nbitq), 
to_sfixed(845.0/65536.0,1,-nbitq), 
to_sfixed(-2618.0/65536.0,1,-nbitq), 
to_sfixed(-759.0/65536.0,1,-nbitq), 
to_sfixed(-5741.0/65536.0,1,-nbitq), 
to_sfixed(-4251.0/65536.0,1,-nbitq), 
to_sfixed(-3027.0/65536.0,1,-nbitq), 
to_sfixed(-2124.0/65536.0,1,-nbitq), 
to_sfixed(-2752.0/65536.0,1,-nbitq), 
to_sfixed(-2565.0/65536.0,1,-nbitq), 
to_sfixed(-3420.0/65536.0,1,-nbitq), 
to_sfixed(-2134.0/65536.0,1,-nbitq), 
to_sfixed(-279.0/65536.0,1,-nbitq), 
to_sfixed(2156.0/65536.0,1,-nbitq), 
to_sfixed(540.0/65536.0,1,-nbitq), 
to_sfixed(-497.0/65536.0,1,-nbitq), 
to_sfixed(251.0/65536.0,1,-nbitq), 
to_sfixed(2063.0/65536.0,1,-nbitq), 
to_sfixed(267.0/65536.0,1,-nbitq), 
to_sfixed(-1104.0/65536.0,1,-nbitq), 
to_sfixed(-1995.0/65536.0,1,-nbitq), 
to_sfixed(1320.0/65536.0,1,-nbitq), 
to_sfixed(-1528.0/65536.0,1,-nbitq), 
to_sfixed(-2541.0/65536.0,1,-nbitq), 
to_sfixed(3054.0/65536.0,1,-nbitq), 
to_sfixed(-1186.0/65536.0,1,-nbitq), 
to_sfixed(3958.0/65536.0,1,-nbitq), 
to_sfixed(1815.0/65536.0,1,-nbitq), 
to_sfixed(-2781.0/65536.0,1,-nbitq), 
to_sfixed(1509.0/65536.0,1,-nbitq), 
to_sfixed(1093.0/65536.0,1,-nbitq), 
to_sfixed(3665.0/65536.0,1,-nbitq), 
to_sfixed(-829.0/65536.0,1,-nbitq), 
to_sfixed(-1854.0/65536.0,1,-nbitq), 
to_sfixed(1814.0/65536.0,1,-nbitq), 
to_sfixed(-2052.0/65536.0,1,-nbitq), 
to_sfixed(-178.0/65536.0,1,-nbitq), 
to_sfixed(3399.0/65536.0,1,-nbitq), 
to_sfixed(2476.0/65536.0,1,-nbitq), 
to_sfixed(-1794.0/65536.0,1,-nbitq), 
to_sfixed(-442.0/65536.0,1,-nbitq), 
to_sfixed(877.0/65536.0,1,-nbitq), 
to_sfixed(2762.0/65536.0,1,-nbitq), 
to_sfixed(2802.0/65536.0,1,-nbitq), 
to_sfixed(1901.0/65536.0,1,-nbitq), 
to_sfixed(-1300.0/65536.0,1,-nbitq), 
to_sfixed(1933.0/65536.0,1,-nbitq), 
to_sfixed(783.0/65536.0,1,-nbitq), 
to_sfixed(2276.0/65536.0,1,-nbitq), 
to_sfixed(-340.0/65536.0,1,-nbitq), 
to_sfixed(13.0/65536.0,1,-nbitq), 
to_sfixed(3624.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2421.0/65536.0,1,-nbitq), 
to_sfixed(-676.0/65536.0,1,-nbitq), 
to_sfixed(-289.0/65536.0,1,-nbitq), 
to_sfixed(-1689.0/65536.0,1,-nbitq), 
to_sfixed(-2094.0/65536.0,1,-nbitq), 
to_sfixed(-1439.0/65536.0,1,-nbitq), 
to_sfixed(-2483.0/65536.0,1,-nbitq), 
to_sfixed(-81.0/65536.0,1,-nbitq), 
to_sfixed(-3081.0/65536.0,1,-nbitq), 
to_sfixed(-1419.0/65536.0,1,-nbitq), 
to_sfixed(-2537.0/65536.0,1,-nbitq), 
to_sfixed(-3305.0/65536.0,1,-nbitq), 
to_sfixed(2549.0/65536.0,1,-nbitq), 
to_sfixed(986.0/65536.0,1,-nbitq), 
to_sfixed(2402.0/65536.0,1,-nbitq), 
to_sfixed(1589.0/65536.0,1,-nbitq), 
to_sfixed(-2135.0/65536.0,1,-nbitq), 
to_sfixed(-584.0/65536.0,1,-nbitq), 
to_sfixed(-736.0/65536.0,1,-nbitq), 
to_sfixed(-2542.0/65536.0,1,-nbitq), 
to_sfixed(-2110.0/65536.0,1,-nbitq), 
to_sfixed(1767.0/65536.0,1,-nbitq), 
to_sfixed(610.0/65536.0,1,-nbitq), 
to_sfixed(718.0/65536.0,1,-nbitq), 
to_sfixed(-398.0/65536.0,1,-nbitq), 
to_sfixed(-518.0/65536.0,1,-nbitq), 
to_sfixed(-1166.0/65536.0,1,-nbitq), 
to_sfixed(933.0/65536.0,1,-nbitq), 
to_sfixed(799.0/65536.0,1,-nbitq), 
to_sfixed(-362.0/65536.0,1,-nbitq), 
to_sfixed(1444.0/65536.0,1,-nbitq), 
to_sfixed(788.0/65536.0,1,-nbitq), 
to_sfixed(-4990.0/65536.0,1,-nbitq), 
to_sfixed(-2596.0/65536.0,1,-nbitq), 
to_sfixed(-918.0/65536.0,1,-nbitq), 
to_sfixed(-2590.0/65536.0,1,-nbitq), 
to_sfixed(-2684.0/65536.0,1,-nbitq), 
to_sfixed(-3320.0/65536.0,1,-nbitq), 
to_sfixed(-327.0/65536.0,1,-nbitq), 
to_sfixed(-305.0/65536.0,1,-nbitq), 
to_sfixed(427.0/65536.0,1,-nbitq), 
to_sfixed(-1771.0/65536.0,1,-nbitq), 
to_sfixed(-5085.0/65536.0,1,-nbitq), 
to_sfixed(1073.0/65536.0,1,-nbitq), 
to_sfixed(-968.0/65536.0,1,-nbitq), 
to_sfixed(5520.0/65536.0,1,-nbitq), 
to_sfixed(2518.0/65536.0,1,-nbitq), 
to_sfixed(-479.0/65536.0,1,-nbitq), 
to_sfixed(-2237.0/65536.0,1,-nbitq), 
to_sfixed(2710.0/65536.0,1,-nbitq), 
to_sfixed(2401.0/65536.0,1,-nbitq), 
to_sfixed(3438.0/65536.0,1,-nbitq), 
to_sfixed(-2251.0/65536.0,1,-nbitq), 
to_sfixed(-1107.0/65536.0,1,-nbitq), 
to_sfixed(1660.0/65536.0,1,-nbitq), 
to_sfixed(1343.0/65536.0,1,-nbitq), 
to_sfixed(1458.0/65536.0,1,-nbitq), 
to_sfixed(1295.0/65536.0,1,-nbitq), 
to_sfixed(1117.0/65536.0,1,-nbitq), 
to_sfixed(1960.0/65536.0,1,-nbitq), 
to_sfixed(-638.0/65536.0,1,-nbitq), 
to_sfixed(-2456.0/65536.0,1,-nbitq), 
to_sfixed(-2511.0/65536.0,1,-nbitq), 
to_sfixed(2516.0/65536.0,1,-nbitq), 
to_sfixed(74.0/65536.0,1,-nbitq), 
to_sfixed(1400.0/65536.0,1,-nbitq), 
to_sfixed(3193.0/65536.0,1,-nbitq), 
to_sfixed(-3852.0/65536.0,1,-nbitq), 
to_sfixed(-312.0/65536.0,1,-nbitq), 
to_sfixed(-681.0/65536.0,1,-nbitq), 
to_sfixed(2875.0/65536.0,1,-nbitq), 
to_sfixed(-299.0/65536.0,1,-nbitq), 
to_sfixed(-56.0/65536.0,1,-nbitq), 
to_sfixed(-2374.0/65536.0,1,-nbitq), 
to_sfixed(-889.0/65536.0,1,-nbitq), 
to_sfixed(341.0/65536.0,1,-nbitq), 
to_sfixed(-3994.0/65536.0,1,-nbitq), 
to_sfixed(2172.0/65536.0,1,-nbitq), 
to_sfixed(-2640.0/65536.0,1,-nbitq), 
to_sfixed(3268.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3434.0/65536.0,1,-nbitq), 
to_sfixed(1106.0/65536.0,1,-nbitq), 
to_sfixed(3503.0/65536.0,1,-nbitq), 
to_sfixed(-2229.0/65536.0,1,-nbitq), 
to_sfixed(-2848.0/65536.0,1,-nbitq), 
to_sfixed(-1373.0/65536.0,1,-nbitq), 
to_sfixed(-2618.0/65536.0,1,-nbitq), 
to_sfixed(-272.0/65536.0,1,-nbitq), 
to_sfixed(-457.0/65536.0,1,-nbitq), 
to_sfixed(-1540.0/65536.0,1,-nbitq), 
to_sfixed(996.0/65536.0,1,-nbitq), 
to_sfixed(1238.0/65536.0,1,-nbitq), 
to_sfixed(1903.0/65536.0,1,-nbitq), 
to_sfixed(-1801.0/65536.0,1,-nbitq), 
to_sfixed(-925.0/65536.0,1,-nbitq), 
to_sfixed(1701.0/65536.0,1,-nbitq), 
to_sfixed(-1733.0/65536.0,1,-nbitq), 
to_sfixed(3082.0/65536.0,1,-nbitq), 
to_sfixed(1931.0/65536.0,1,-nbitq), 
to_sfixed(1083.0/65536.0,1,-nbitq), 
to_sfixed(-2921.0/65536.0,1,-nbitq), 
to_sfixed(-1897.0/65536.0,1,-nbitq), 
to_sfixed(-1584.0/65536.0,1,-nbitq), 
to_sfixed(3126.0/65536.0,1,-nbitq), 
to_sfixed(2701.0/65536.0,1,-nbitq), 
to_sfixed(1695.0/65536.0,1,-nbitq), 
to_sfixed(172.0/65536.0,1,-nbitq), 
to_sfixed(-2638.0/65536.0,1,-nbitq), 
to_sfixed(-321.0/65536.0,1,-nbitq), 
to_sfixed(844.0/65536.0,1,-nbitq), 
to_sfixed(-622.0/65536.0,1,-nbitq), 
to_sfixed(2896.0/65536.0,1,-nbitq), 
to_sfixed(-5142.0/65536.0,1,-nbitq), 
to_sfixed(-3670.0/65536.0,1,-nbitq), 
to_sfixed(122.0/65536.0,1,-nbitq), 
to_sfixed(-2813.0/65536.0,1,-nbitq), 
to_sfixed(898.0/65536.0,1,-nbitq), 
to_sfixed(-948.0/65536.0,1,-nbitq), 
to_sfixed(-583.0/65536.0,1,-nbitq), 
to_sfixed(2180.0/65536.0,1,-nbitq), 
to_sfixed(1986.0/65536.0,1,-nbitq), 
to_sfixed(1465.0/65536.0,1,-nbitq), 
to_sfixed(-3077.0/65536.0,1,-nbitq), 
to_sfixed(492.0/65536.0,1,-nbitq), 
to_sfixed(1861.0/65536.0,1,-nbitq), 
to_sfixed(503.0/65536.0,1,-nbitq), 
to_sfixed(-2304.0/65536.0,1,-nbitq), 
to_sfixed(-1905.0/65536.0,1,-nbitq), 
to_sfixed(714.0/65536.0,1,-nbitq), 
to_sfixed(4514.0/65536.0,1,-nbitq), 
to_sfixed(1651.0/65536.0,1,-nbitq), 
to_sfixed(-624.0/65536.0,1,-nbitq), 
to_sfixed(-595.0/65536.0,1,-nbitq), 
to_sfixed(1257.0/65536.0,1,-nbitq), 
to_sfixed(3616.0/65536.0,1,-nbitq), 
to_sfixed(1063.0/65536.0,1,-nbitq), 
to_sfixed(-1305.0/65536.0,1,-nbitq), 
to_sfixed(-2216.0/65536.0,1,-nbitq), 
to_sfixed(1843.0/65536.0,1,-nbitq), 
to_sfixed(3233.0/65536.0,1,-nbitq), 
to_sfixed(1696.0/65536.0,1,-nbitq), 
to_sfixed(-2801.0/65536.0,1,-nbitq), 
to_sfixed(678.0/65536.0,1,-nbitq), 
to_sfixed(-1705.0/65536.0,1,-nbitq), 
to_sfixed(3215.0/65536.0,1,-nbitq), 
to_sfixed(-2278.0/65536.0,1,-nbitq), 
to_sfixed(196.0/65536.0,1,-nbitq), 
to_sfixed(-2652.0/65536.0,1,-nbitq), 
to_sfixed(3700.0/65536.0,1,-nbitq), 
to_sfixed(1303.0/65536.0,1,-nbitq), 
to_sfixed(-1510.0/65536.0,1,-nbitq), 
to_sfixed(-720.0/65536.0,1,-nbitq), 
to_sfixed(-914.0/65536.0,1,-nbitq), 
to_sfixed(716.0/65536.0,1,-nbitq), 
to_sfixed(177.0/65536.0,1,-nbitq), 
to_sfixed(-910.0/65536.0,1,-nbitq), 
to_sfixed(-3961.0/65536.0,1,-nbitq), 
to_sfixed(2505.0/65536.0,1,-nbitq), 
to_sfixed(2274.0/65536.0,1,-nbitq), 
to_sfixed(2900.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3286.0/65536.0,1,-nbitq), 
to_sfixed(-2227.0/65536.0,1,-nbitq), 
to_sfixed(3547.0/65536.0,1,-nbitq), 
to_sfixed(-941.0/65536.0,1,-nbitq), 
to_sfixed(-2964.0/65536.0,1,-nbitq), 
to_sfixed(-5.0/65536.0,1,-nbitq), 
to_sfixed(-1057.0/65536.0,1,-nbitq), 
to_sfixed(87.0/65536.0,1,-nbitq), 
to_sfixed(352.0/65536.0,1,-nbitq), 
to_sfixed(2295.0/65536.0,1,-nbitq), 
to_sfixed(-2026.0/65536.0,1,-nbitq), 
to_sfixed(-734.0/65536.0,1,-nbitq), 
to_sfixed(2657.0/65536.0,1,-nbitq), 
to_sfixed(-4085.0/65536.0,1,-nbitq), 
to_sfixed(981.0/65536.0,1,-nbitq), 
to_sfixed(-330.0/65536.0,1,-nbitq), 
to_sfixed(-1289.0/65536.0,1,-nbitq), 
to_sfixed(-702.0/65536.0,1,-nbitq), 
to_sfixed(2803.0/65536.0,1,-nbitq), 
to_sfixed(3471.0/65536.0,1,-nbitq), 
to_sfixed(-2918.0/65536.0,1,-nbitq), 
to_sfixed(1940.0/65536.0,1,-nbitq), 
to_sfixed(-1952.0/65536.0,1,-nbitq), 
to_sfixed(4286.0/65536.0,1,-nbitq), 
to_sfixed(2023.0/65536.0,1,-nbitq), 
to_sfixed(93.0/65536.0,1,-nbitq), 
to_sfixed(212.0/65536.0,1,-nbitq), 
to_sfixed(-786.0/65536.0,1,-nbitq), 
to_sfixed(1069.0/65536.0,1,-nbitq), 
to_sfixed(-1792.0/65536.0,1,-nbitq), 
to_sfixed(-2614.0/65536.0,1,-nbitq), 
to_sfixed(457.0/65536.0,1,-nbitq), 
to_sfixed(-320.0/65536.0,1,-nbitq), 
to_sfixed(-4413.0/65536.0,1,-nbitq), 
to_sfixed(-360.0/65536.0,1,-nbitq), 
to_sfixed(1182.0/65536.0,1,-nbitq), 
to_sfixed(-3337.0/65536.0,1,-nbitq), 
to_sfixed(1503.0/65536.0,1,-nbitq), 
to_sfixed(788.0/65536.0,1,-nbitq), 
to_sfixed(484.0/65536.0,1,-nbitq), 
to_sfixed(-2179.0/65536.0,1,-nbitq), 
to_sfixed(-305.0/65536.0,1,-nbitq), 
to_sfixed(-1859.0/65536.0,1,-nbitq), 
to_sfixed(3902.0/65536.0,1,-nbitq), 
to_sfixed(2476.0/65536.0,1,-nbitq), 
to_sfixed(5589.0/65536.0,1,-nbitq), 
to_sfixed(1132.0/65536.0,1,-nbitq), 
to_sfixed(-1035.0/65536.0,1,-nbitq), 
to_sfixed(3149.0/65536.0,1,-nbitq), 
to_sfixed(1556.0/65536.0,1,-nbitq), 
to_sfixed(-1184.0/65536.0,1,-nbitq), 
to_sfixed(-164.0/65536.0,1,-nbitq), 
to_sfixed(1862.0/65536.0,1,-nbitq), 
to_sfixed(-478.0/65536.0,1,-nbitq), 
to_sfixed(2685.0/65536.0,1,-nbitq), 
to_sfixed(3169.0/65536.0,1,-nbitq), 
to_sfixed(2905.0/65536.0,1,-nbitq), 
to_sfixed(576.0/65536.0,1,-nbitq), 
to_sfixed(2640.0/65536.0,1,-nbitq), 
to_sfixed(497.0/65536.0,1,-nbitq), 
to_sfixed(-3629.0/65536.0,1,-nbitq), 
to_sfixed(-1375.0/65536.0,1,-nbitq), 
to_sfixed(651.0/65536.0,1,-nbitq), 
to_sfixed(-211.0/65536.0,1,-nbitq), 
to_sfixed(3407.0/65536.0,1,-nbitq), 
to_sfixed(-78.0/65536.0,1,-nbitq), 
to_sfixed(95.0/65536.0,1,-nbitq), 
to_sfixed(-1515.0/65536.0,1,-nbitq), 
to_sfixed(2736.0/65536.0,1,-nbitq), 
to_sfixed(-2646.0/65536.0,1,-nbitq), 
to_sfixed(2080.0/65536.0,1,-nbitq), 
to_sfixed(-1766.0/65536.0,1,-nbitq), 
to_sfixed(1207.0/65536.0,1,-nbitq), 
to_sfixed(-1750.0/65536.0,1,-nbitq), 
to_sfixed(-1000.0/65536.0,1,-nbitq), 
to_sfixed(2124.0/65536.0,1,-nbitq), 
to_sfixed(-3326.0/65536.0,1,-nbitq), 
to_sfixed(1267.0/65536.0,1,-nbitq), 
to_sfixed(-1998.0/65536.0,1,-nbitq), 
to_sfixed(578.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1492.0/65536.0,1,-nbitq), 
to_sfixed(2832.0/65536.0,1,-nbitq), 
to_sfixed(1875.0/65536.0,1,-nbitq), 
to_sfixed(-1273.0/65536.0,1,-nbitq), 
to_sfixed(-4530.0/65536.0,1,-nbitq), 
to_sfixed(817.0/65536.0,1,-nbitq), 
to_sfixed(-1029.0/65536.0,1,-nbitq), 
to_sfixed(1678.0/65536.0,1,-nbitq), 
to_sfixed(-214.0/65536.0,1,-nbitq), 
to_sfixed(-629.0/65536.0,1,-nbitq), 
to_sfixed(1262.0/65536.0,1,-nbitq), 
to_sfixed(-267.0/65536.0,1,-nbitq), 
to_sfixed(-344.0/65536.0,1,-nbitq), 
to_sfixed(-184.0/65536.0,1,-nbitq), 
to_sfixed(2884.0/65536.0,1,-nbitq), 
to_sfixed(-236.0/65536.0,1,-nbitq), 
to_sfixed(-1133.0/65536.0,1,-nbitq), 
to_sfixed(698.0/65536.0,1,-nbitq), 
to_sfixed(3485.0/65536.0,1,-nbitq), 
to_sfixed(1681.0/65536.0,1,-nbitq), 
to_sfixed(-1647.0/65536.0,1,-nbitq), 
to_sfixed(1898.0/65536.0,1,-nbitq), 
to_sfixed(2505.0/65536.0,1,-nbitq), 
to_sfixed(1323.0/65536.0,1,-nbitq), 
to_sfixed(474.0/65536.0,1,-nbitq), 
to_sfixed(-869.0/65536.0,1,-nbitq), 
to_sfixed(-3751.0/65536.0,1,-nbitq), 
to_sfixed(-2987.0/65536.0,1,-nbitq), 
to_sfixed(-3708.0/65536.0,1,-nbitq), 
to_sfixed(-1190.0/65536.0,1,-nbitq), 
to_sfixed(-2930.0/65536.0,1,-nbitq), 
to_sfixed(2507.0/65536.0,1,-nbitq), 
to_sfixed(-1970.0/65536.0,1,-nbitq), 
to_sfixed(-5469.0/65536.0,1,-nbitq), 
to_sfixed(-2680.0/65536.0,1,-nbitq), 
to_sfixed(-1970.0/65536.0,1,-nbitq), 
to_sfixed(-778.0/65536.0,1,-nbitq), 
to_sfixed(-3504.0/65536.0,1,-nbitq), 
to_sfixed(-3658.0/65536.0,1,-nbitq), 
to_sfixed(1331.0/65536.0,1,-nbitq), 
to_sfixed(-708.0/65536.0,1,-nbitq), 
to_sfixed(1412.0/65536.0,1,-nbitq), 
to_sfixed(-2226.0/65536.0,1,-nbitq), 
to_sfixed(981.0/65536.0,1,-nbitq), 
to_sfixed(-2360.0/65536.0,1,-nbitq), 
to_sfixed(108.0/65536.0,1,-nbitq), 
to_sfixed(-2325.0/65536.0,1,-nbitq), 
to_sfixed(-181.0/65536.0,1,-nbitq), 
to_sfixed(-982.0/65536.0,1,-nbitq), 
to_sfixed(3462.0/65536.0,1,-nbitq), 
to_sfixed(2522.0/65536.0,1,-nbitq), 
to_sfixed(3358.0/65536.0,1,-nbitq), 
to_sfixed(814.0/65536.0,1,-nbitq), 
to_sfixed(-2870.0/65536.0,1,-nbitq), 
to_sfixed(-492.0/65536.0,1,-nbitq), 
to_sfixed(478.0/65536.0,1,-nbitq), 
to_sfixed(1711.0/65536.0,1,-nbitq), 
to_sfixed(-741.0/65536.0,1,-nbitq), 
to_sfixed(-438.0/65536.0,1,-nbitq), 
to_sfixed(3735.0/65536.0,1,-nbitq), 
to_sfixed(1663.0/65536.0,1,-nbitq), 
to_sfixed(-2215.0/65536.0,1,-nbitq), 
to_sfixed(1470.0/65536.0,1,-nbitq), 
to_sfixed(68.0/65536.0,1,-nbitq), 
to_sfixed(1112.0/65536.0,1,-nbitq), 
to_sfixed(1877.0/65536.0,1,-nbitq), 
to_sfixed(-147.0/65536.0,1,-nbitq), 
to_sfixed(-3999.0/65536.0,1,-nbitq), 
to_sfixed(2349.0/65536.0,1,-nbitq), 
to_sfixed(847.0/65536.0,1,-nbitq), 
to_sfixed(-749.0/65536.0,1,-nbitq), 
to_sfixed(2378.0/65536.0,1,-nbitq), 
to_sfixed(4400.0/65536.0,1,-nbitq), 
to_sfixed(2560.0/65536.0,1,-nbitq), 
to_sfixed(-2465.0/65536.0,1,-nbitq), 
to_sfixed(-763.0/65536.0,1,-nbitq), 
to_sfixed(-4449.0/65536.0,1,-nbitq), 
to_sfixed(3141.0/65536.0,1,-nbitq), 
to_sfixed(-2531.0/65536.0,1,-nbitq), 
to_sfixed(2123.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1911.0/65536.0,1,-nbitq), 
to_sfixed(809.0/65536.0,1,-nbitq), 
to_sfixed(1458.0/65536.0,1,-nbitq), 
to_sfixed(-2531.0/65536.0,1,-nbitq), 
to_sfixed(-3394.0/65536.0,1,-nbitq), 
to_sfixed(493.0/65536.0,1,-nbitq), 
to_sfixed(-3097.0/65536.0,1,-nbitq), 
to_sfixed(-817.0/65536.0,1,-nbitq), 
to_sfixed(1202.0/65536.0,1,-nbitq), 
to_sfixed(-2606.0/65536.0,1,-nbitq), 
to_sfixed(190.0/65536.0,1,-nbitq), 
to_sfixed(421.0/65536.0,1,-nbitq), 
to_sfixed(-1415.0/65536.0,1,-nbitq), 
to_sfixed(-4801.0/65536.0,1,-nbitq), 
to_sfixed(1513.0/65536.0,1,-nbitq), 
to_sfixed(2696.0/65536.0,1,-nbitq), 
to_sfixed(573.0/65536.0,1,-nbitq), 
to_sfixed(1938.0/65536.0,1,-nbitq), 
to_sfixed(-1075.0/65536.0,1,-nbitq), 
to_sfixed(1976.0/65536.0,1,-nbitq), 
to_sfixed(-1695.0/65536.0,1,-nbitq), 
to_sfixed(160.0/65536.0,1,-nbitq), 
to_sfixed(-2389.0/65536.0,1,-nbitq), 
to_sfixed(2498.0/65536.0,1,-nbitq), 
to_sfixed(1016.0/65536.0,1,-nbitq), 
to_sfixed(1451.0/65536.0,1,-nbitq), 
to_sfixed(672.0/65536.0,1,-nbitq), 
to_sfixed(-4045.0/65536.0,1,-nbitq), 
to_sfixed(680.0/65536.0,1,-nbitq), 
to_sfixed(-1007.0/65536.0,1,-nbitq), 
to_sfixed(1677.0/65536.0,1,-nbitq), 
to_sfixed(1529.0/65536.0,1,-nbitq), 
to_sfixed(-976.0/65536.0,1,-nbitq), 
to_sfixed(-4435.0/65536.0,1,-nbitq), 
to_sfixed(78.0/65536.0,1,-nbitq), 
to_sfixed(446.0/65536.0,1,-nbitq), 
to_sfixed(2074.0/65536.0,1,-nbitq), 
to_sfixed(633.0/65536.0,1,-nbitq), 
to_sfixed(1736.0/65536.0,1,-nbitq), 
to_sfixed(46.0/65536.0,1,-nbitq), 
to_sfixed(1151.0/65536.0,1,-nbitq), 
to_sfixed(1862.0/65536.0,1,-nbitq), 
to_sfixed(-4550.0/65536.0,1,-nbitq), 
to_sfixed(4482.0/65536.0,1,-nbitq), 
to_sfixed(-219.0/65536.0,1,-nbitq), 
to_sfixed(-6.0/65536.0,1,-nbitq), 
to_sfixed(1708.0/65536.0,1,-nbitq), 
to_sfixed(-3255.0/65536.0,1,-nbitq), 
to_sfixed(-1573.0/65536.0,1,-nbitq), 
to_sfixed(1745.0/65536.0,1,-nbitq), 
to_sfixed(-1045.0/65536.0,1,-nbitq), 
to_sfixed(-551.0/65536.0,1,-nbitq), 
to_sfixed(752.0/65536.0,1,-nbitq), 
to_sfixed(-2401.0/65536.0,1,-nbitq), 
to_sfixed(527.0/65536.0,1,-nbitq), 
to_sfixed(926.0/65536.0,1,-nbitq), 
to_sfixed(-1836.0/65536.0,1,-nbitq), 
to_sfixed(-1968.0/65536.0,1,-nbitq), 
to_sfixed(-2701.0/65536.0,1,-nbitq), 
to_sfixed(1964.0/65536.0,1,-nbitq), 
to_sfixed(914.0/65536.0,1,-nbitq), 
to_sfixed(-1794.0/65536.0,1,-nbitq), 
to_sfixed(1623.0/65536.0,1,-nbitq), 
to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(3979.0/65536.0,1,-nbitq), 
to_sfixed(1464.0/65536.0,1,-nbitq), 
to_sfixed(-733.0/65536.0,1,-nbitq), 
to_sfixed(-3403.0/65536.0,1,-nbitq), 
to_sfixed(1585.0/65536.0,1,-nbitq), 
to_sfixed(-1223.0/65536.0,1,-nbitq), 
to_sfixed(2334.0/65536.0,1,-nbitq), 
to_sfixed(3053.0/65536.0,1,-nbitq), 
to_sfixed(1583.0/65536.0,1,-nbitq), 
to_sfixed(-1706.0/65536.0,1,-nbitq), 
to_sfixed(821.0/65536.0,1,-nbitq), 
to_sfixed(-1221.0/65536.0,1,-nbitq), 
to_sfixed(-2185.0/65536.0,1,-nbitq), 
to_sfixed(1687.0/65536.0,1,-nbitq), 
to_sfixed(34.0/65536.0,1,-nbitq), 
to_sfixed(5989.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1083.0/65536.0,1,-nbitq), 
to_sfixed(3700.0/65536.0,1,-nbitq), 
to_sfixed(428.0/65536.0,1,-nbitq), 
to_sfixed(-451.0/65536.0,1,-nbitq), 
to_sfixed(-5914.0/65536.0,1,-nbitq), 
to_sfixed(-620.0/65536.0,1,-nbitq), 
to_sfixed(-503.0/65536.0,1,-nbitq), 
to_sfixed(1582.0/65536.0,1,-nbitq), 
to_sfixed(1990.0/65536.0,1,-nbitq), 
to_sfixed(2615.0/65536.0,1,-nbitq), 
to_sfixed(-1445.0/65536.0,1,-nbitq), 
to_sfixed(-5716.0/65536.0,1,-nbitq), 
to_sfixed(113.0/65536.0,1,-nbitq), 
to_sfixed(-4719.0/65536.0,1,-nbitq), 
to_sfixed(-1633.0/65536.0,1,-nbitq), 
to_sfixed(-871.0/65536.0,1,-nbitq), 
to_sfixed(-2589.0/65536.0,1,-nbitq), 
to_sfixed(994.0/65536.0,1,-nbitq), 
to_sfixed(1923.0/65536.0,1,-nbitq), 
to_sfixed(702.0/65536.0,1,-nbitq), 
to_sfixed(-1552.0/65536.0,1,-nbitq), 
to_sfixed(2947.0/65536.0,1,-nbitq), 
to_sfixed(-111.0/65536.0,1,-nbitq), 
to_sfixed(2918.0/65536.0,1,-nbitq), 
to_sfixed(2701.0/65536.0,1,-nbitq), 
to_sfixed(-1102.0/65536.0,1,-nbitq), 
to_sfixed(-989.0/65536.0,1,-nbitq), 
to_sfixed(-2458.0/65536.0,1,-nbitq), 
to_sfixed(-1441.0/65536.0,1,-nbitq), 
to_sfixed(711.0/65536.0,1,-nbitq), 
to_sfixed(1420.0/65536.0,1,-nbitq), 
to_sfixed(-2271.0/65536.0,1,-nbitq), 
to_sfixed(-474.0/65536.0,1,-nbitq), 
to_sfixed(-4651.0/65536.0,1,-nbitq), 
to_sfixed(-220.0/65536.0,1,-nbitq), 
to_sfixed(1129.0/65536.0,1,-nbitq), 
to_sfixed(1043.0/65536.0,1,-nbitq), 
to_sfixed(-2133.0/65536.0,1,-nbitq), 
to_sfixed(1297.0/65536.0,1,-nbitq), 
to_sfixed(1786.0/65536.0,1,-nbitq), 
to_sfixed(-845.0/65536.0,1,-nbitq), 
to_sfixed(-2554.0/65536.0,1,-nbitq), 
to_sfixed(-2999.0/65536.0,1,-nbitq), 
to_sfixed(1289.0/65536.0,1,-nbitq), 
to_sfixed(-942.0/65536.0,1,-nbitq), 
to_sfixed(5353.0/65536.0,1,-nbitq), 
to_sfixed(-2562.0/65536.0,1,-nbitq), 
to_sfixed(-819.0/65536.0,1,-nbitq), 
to_sfixed(-1471.0/65536.0,1,-nbitq), 
to_sfixed(3196.0/65536.0,1,-nbitq), 
to_sfixed(-1559.0/65536.0,1,-nbitq), 
to_sfixed(318.0/65536.0,1,-nbitq), 
to_sfixed(4469.0/65536.0,1,-nbitq), 
to_sfixed(-2443.0/65536.0,1,-nbitq), 
to_sfixed(-1407.0/65536.0,1,-nbitq), 
to_sfixed(-1579.0/65536.0,1,-nbitq), 
to_sfixed(-453.0/65536.0,1,-nbitq), 
to_sfixed(-1123.0/65536.0,1,-nbitq), 
to_sfixed(-1892.0/65536.0,1,-nbitq), 
to_sfixed(5625.0/65536.0,1,-nbitq), 
to_sfixed(447.0/65536.0,1,-nbitq), 
to_sfixed(2474.0/65536.0,1,-nbitq), 
to_sfixed(-178.0/65536.0,1,-nbitq), 
to_sfixed(2262.0/65536.0,1,-nbitq), 
to_sfixed(-635.0/65536.0,1,-nbitq), 
to_sfixed(93.0/65536.0,1,-nbitq), 
to_sfixed(2231.0/65536.0,1,-nbitq), 
to_sfixed(-3758.0/65536.0,1,-nbitq), 
to_sfixed(4049.0/65536.0,1,-nbitq), 
to_sfixed(1113.0/65536.0,1,-nbitq), 
to_sfixed(2293.0/65536.0,1,-nbitq), 
to_sfixed(1124.0/65536.0,1,-nbitq), 
to_sfixed(2768.0/65536.0,1,-nbitq), 
to_sfixed(-1314.0/65536.0,1,-nbitq), 
to_sfixed(-1921.0/65536.0,1,-nbitq), 
to_sfixed(-649.0/65536.0,1,-nbitq), 
to_sfixed(-2028.0/65536.0,1,-nbitq), 
to_sfixed(4155.0/65536.0,1,-nbitq), 
to_sfixed(-1460.0/65536.0,1,-nbitq), 
to_sfixed(2203.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1606.0/65536.0,1,-nbitq), 
to_sfixed(2192.0/65536.0,1,-nbitq), 
to_sfixed(3416.0/65536.0,1,-nbitq), 
to_sfixed(-2074.0/65536.0,1,-nbitq), 
to_sfixed(-1950.0/65536.0,1,-nbitq), 
to_sfixed(-812.0/65536.0,1,-nbitq), 
to_sfixed(-3092.0/65536.0,1,-nbitq), 
to_sfixed(-794.0/65536.0,1,-nbitq), 
to_sfixed(-1140.0/65536.0,1,-nbitq), 
to_sfixed(662.0/65536.0,1,-nbitq), 
to_sfixed(1023.0/65536.0,1,-nbitq), 
to_sfixed(-4516.0/65536.0,1,-nbitq), 
to_sfixed(1793.0/65536.0,1,-nbitq), 
to_sfixed(-792.0/65536.0,1,-nbitq), 
to_sfixed(-1280.0/65536.0,1,-nbitq), 
to_sfixed(-311.0/65536.0,1,-nbitq), 
to_sfixed(376.0/65536.0,1,-nbitq), 
to_sfixed(980.0/65536.0,1,-nbitq), 
to_sfixed(1096.0/65536.0,1,-nbitq), 
to_sfixed(2015.0/65536.0,1,-nbitq), 
to_sfixed(-1332.0/65536.0,1,-nbitq), 
to_sfixed(1160.0/65536.0,1,-nbitq), 
to_sfixed(2422.0/65536.0,1,-nbitq), 
to_sfixed(254.0/65536.0,1,-nbitq), 
to_sfixed(2711.0/65536.0,1,-nbitq), 
to_sfixed(-2115.0/65536.0,1,-nbitq), 
to_sfixed(-553.0/65536.0,1,-nbitq), 
to_sfixed(-1008.0/65536.0,1,-nbitq), 
to_sfixed(-301.0/65536.0,1,-nbitq), 
to_sfixed(-3521.0/65536.0,1,-nbitq), 
to_sfixed(-456.0/65536.0,1,-nbitq), 
to_sfixed(50.0/65536.0,1,-nbitq), 
to_sfixed(-3405.0/65536.0,1,-nbitq), 
to_sfixed(2805.0/65536.0,1,-nbitq), 
to_sfixed(2673.0/65536.0,1,-nbitq), 
to_sfixed(-440.0/65536.0,1,-nbitq), 
to_sfixed(864.0/65536.0,1,-nbitq), 
to_sfixed(-3411.0/65536.0,1,-nbitq), 
to_sfixed(1481.0/65536.0,1,-nbitq), 
to_sfixed(-2310.0/65536.0,1,-nbitq), 
to_sfixed(173.0/65536.0,1,-nbitq), 
to_sfixed(1791.0/65536.0,1,-nbitq), 
to_sfixed(-2778.0/65536.0,1,-nbitq), 
to_sfixed(884.0/65536.0,1,-nbitq), 
to_sfixed(246.0/65536.0,1,-nbitq), 
to_sfixed(1761.0/65536.0,1,-nbitq), 
to_sfixed(1725.0/65536.0,1,-nbitq), 
to_sfixed(942.0/65536.0,1,-nbitq), 
to_sfixed(-1502.0/65536.0,1,-nbitq), 
to_sfixed(-158.0/65536.0,1,-nbitq), 
to_sfixed(1608.0/65536.0,1,-nbitq), 
to_sfixed(-872.0/65536.0,1,-nbitq), 
to_sfixed(4162.0/65536.0,1,-nbitq), 
to_sfixed(1079.0/65536.0,1,-nbitq), 
to_sfixed(3027.0/65536.0,1,-nbitq), 
to_sfixed(1305.0/65536.0,1,-nbitq), 
to_sfixed(-410.0/65536.0,1,-nbitq), 
to_sfixed(663.0/65536.0,1,-nbitq), 
to_sfixed(2744.0/65536.0,1,-nbitq), 
to_sfixed(2910.0/65536.0,1,-nbitq), 
to_sfixed(1811.0/65536.0,1,-nbitq), 
to_sfixed(1039.0/65536.0,1,-nbitq), 
to_sfixed(126.0/65536.0,1,-nbitq), 
to_sfixed(421.0/65536.0,1,-nbitq), 
to_sfixed(4585.0/65536.0,1,-nbitq), 
to_sfixed(-2235.0/65536.0,1,-nbitq), 
to_sfixed(1.0/65536.0,1,-nbitq), 
to_sfixed(993.0/65536.0,1,-nbitq), 
to_sfixed(346.0/65536.0,1,-nbitq), 
to_sfixed(-1079.0/65536.0,1,-nbitq), 
to_sfixed(2597.0/65536.0,1,-nbitq), 
to_sfixed(3348.0/65536.0,1,-nbitq), 
to_sfixed(1751.0/65536.0,1,-nbitq), 
to_sfixed(-2625.0/65536.0,1,-nbitq), 
to_sfixed(-3043.0/65536.0,1,-nbitq), 
to_sfixed(815.0/65536.0,1,-nbitq), 
to_sfixed(-2498.0/65536.0,1,-nbitq), 
to_sfixed(4453.0/65536.0,1,-nbitq), 
to_sfixed(1279.0/65536.0,1,-nbitq), 
to_sfixed(3513.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-460.0/65536.0,1,-nbitq), 
to_sfixed(908.0/65536.0,1,-nbitq), 
to_sfixed(1961.0/65536.0,1,-nbitq), 
to_sfixed(108.0/65536.0,1,-nbitq), 
to_sfixed(-6550.0/65536.0,1,-nbitq), 
to_sfixed(-1511.0/65536.0,1,-nbitq), 
to_sfixed(-1425.0/65536.0,1,-nbitq), 
to_sfixed(-4121.0/65536.0,1,-nbitq), 
to_sfixed(2389.0/65536.0,1,-nbitq), 
to_sfixed(-928.0/65536.0,1,-nbitq), 
to_sfixed(-3569.0/65536.0,1,-nbitq), 
to_sfixed(-3924.0/65536.0,1,-nbitq), 
to_sfixed(-1148.0/65536.0,1,-nbitq), 
to_sfixed(-3788.0/65536.0,1,-nbitq), 
to_sfixed(843.0/65536.0,1,-nbitq), 
to_sfixed(-2591.0/65536.0,1,-nbitq), 
to_sfixed(-1444.0/65536.0,1,-nbitq), 
to_sfixed(-1070.0/65536.0,1,-nbitq), 
to_sfixed(1369.0/65536.0,1,-nbitq), 
to_sfixed(123.0/65536.0,1,-nbitq), 
to_sfixed(962.0/65536.0,1,-nbitq), 
to_sfixed(3931.0/65536.0,1,-nbitq), 
to_sfixed(2723.0/65536.0,1,-nbitq), 
to_sfixed(-3581.0/65536.0,1,-nbitq), 
to_sfixed(3753.0/65536.0,1,-nbitq), 
to_sfixed(897.0/65536.0,1,-nbitq), 
to_sfixed(-4524.0/65536.0,1,-nbitq), 
to_sfixed(-1664.0/65536.0,1,-nbitq), 
to_sfixed(-5333.0/65536.0,1,-nbitq), 
to_sfixed(-383.0/65536.0,1,-nbitq), 
to_sfixed(-1589.0/65536.0,1,-nbitq), 
to_sfixed(513.0/65536.0,1,-nbitq), 
to_sfixed(65.0/65536.0,1,-nbitq), 
to_sfixed(2988.0/65536.0,1,-nbitq), 
to_sfixed(50.0/65536.0,1,-nbitq), 
to_sfixed(-2494.0/65536.0,1,-nbitq), 
to_sfixed(-485.0/65536.0,1,-nbitq), 
to_sfixed(-1885.0/65536.0,1,-nbitq), 
to_sfixed(-689.0/65536.0,1,-nbitq), 
to_sfixed(-1083.0/65536.0,1,-nbitq), 
to_sfixed(3.0/65536.0,1,-nbitq), 
to_sfixed(8.0/65536.0,1,-nbitq), 
to_sfixed(768.0/65536.0,1,-nbitq), 
to_sfixed(2997.0/65536.0,1,-nbitq), 
to_sfixed(2590.0/65536.0,1,-nbitq), 
to_sfixed(-52.0/65536.0,1,-nbitq), 
to_sfixed(-1345.0/65536.0,1,-nbitq), 
to_sfixed(-3149.0/65536.0,1,-nbitq), 
to_sfixed(3274.0/65536.0,1,-nbitq), 
to_sfixed(3280.0/65536.0,1,-nbitq), 
to_sfixed(126.0/65536.0,1,-nbitq), 
to_sfixed(-1068.0/65536.0,1,-nbitq), 
to_sfixed(-1307.0/65536.0,1,-nbitq), 
to_sfixed(-1222.0/65536.0,1,-nbitq), 
to_sfixed(2799.0/65536.0,1,-nbitq), 
to_sfixed(-3476.0/65536.0,1,-nbitq), 
to_sfixed(-305.0/65536.0,1,-nbitq), 
to_sfixed(-2359.0/65536.0,1,-nbitq), 
to_sfixed(1489.0/65536.0,1,-nbitq), 
to_sfixed(1703.0/65536.0,1,-nbitq), 
to_sfixed(2101.0/65536.0,1,-nbitq), 
to_sfixed(-3113.0/65536.0,1,-nbitq), 
to_sfixed(2225.0/65536.0,1,-nbitq), 
to_sfixed(330.0/65536.0,1,-nbitq), 
to_sfixed(2475.0/65536.0,1,-nbitq), 
to_sfixed(786.0/65536.0,1,-nbitq), 
to_sfixed(2200.0/65536.0,1,-nbitq), 
to_sfixed(-4468.0/65536.0,1,-nbitq), 
to_sfixed(3200.0/65536.0,1,-nbitq), 
to_sfixed(-6301.0/65536.0,1,-nbitq), 
to_sfixed(-944.0/65536.0,1,-nbitq), 
to_sfixed(-1428.0/65536.0,1,-nbitq), 
to_sfixed(2899.0/65536.0,1,-nbitq), 
to_sfixed(-2863.0/65536.0,1,-nbitq), 
to_sfixed(214.0/65536.0,1,-nbitq), 
to_sfixed(-394.0/65536.0,1,-nbitq), 
to_sfixed(-1994.0/65536.0,1,-nbitq), 
to_sfixed(3543.0/65536.0,1,-nbitq), 
to_sfixed(-2872.0/65536.0,1,-nbitq), 
to_sfixed(4685.0/65536.0,1,-nbitq)  ), 
( to_sfixed(298.0/65536.0,1,-nbitq), 
to_sfixed(4331.0/65536.0,1,-nbitq), 
to_sfixed(-3850.0/65536.0,1,-nbitq), 
to_sfixed(87.0/65536.0,1,-nbitq), 
to_sfixed(-1599.0/65536.0,1,-nbitq), 
to_sfixed(24.0/65536.0,1,-nbitq), 
to_sfixed(-1851.0/65536.0,1,-nbitq), 
to_sfixed(-4424.0/65536.0,1,-nbitq), 
to_sfixed(-2123.0/65536.0,1,-nbitq), 
to_sfixed(840.0/65536.0,1,-nbitq), 
to_sfixed(-799.0/65536.0,1,-nbitq), 
to_sfixed(200.0/65536.0,1,-nbitq), 
to_sfixed(-856.0/65536.0,1,-nbitq), 
to_sfixed(599.0/65536.0,1,-nbitq), 
to_sfixed(367.0/65536.0,1,-nbitq), 
to_sfixed(2823.0/65536.0,1,-nbitq), 
to_sfixed(-2682.0/65536.0,1,-nbitq), 
to_sfixed(-1751.0/65536.0,1,-nbitq), 
to_sfixed(249.0/65536.0,1,-nbitq), 
to_sfixed(2954.0/65536.0,1,-nbitq), 
to_sfixed(1351.0/65536.0,1,-nbitq), 
to_sfixed(2622.0/65536.0,1,-nbitq), 
to_sfixed(-199.0/65536.0,1,-nbitq), 
to_sfixed(-381.0/65536.0,1,-nbitq), 
to_sfixed(2539.0/65536.0,1,-nbitq), 
to_sfixed(-2855.0/65536.0,1,-nbitq), 
to_sfixed(-4420.0/65536.0,1,-nbitq), 
to_sfixed(-2508.0/65536.0,1,-nbitq), 
to_sfixed(-3055.0/65536.0,1,-nbitq), 
to_sfixed(746.0/65536.0,1,-nbitq), 
to_sfixed(928.0/65536.0,1,-nbitq), 
to_sfixed(854.0/65536.0,1,-nbitq), 
to_sfixed(-1709.0/65536.0,1,-nbitq), 
to_sfixed(4196.0/65536.0,1,-nbitq), 
to_sfixed(2168.0/65536.0,1,-nbitq), 
to_sfixed(-92.0/65536.0,1,-nbitq), 
to_sfixed(-545.0/65536.0,1,-nbitq), 
to_sfixed(-969.0/65536.0,1,-nbitq), 
to_sfixed(1286.0/65536.0,1,-nbitq), 
to_sfixed(416.0/65536.0,1,-nbitq), 
to_sfixed(2611.0/65536.0,1,-nbitq), 
to_sfixed(2179.0/65536.0,1,-nbitq), 
to_sfixed(327.0/65536.0,1,-nbitq), 
to_sfixed(871.0/65536.0,1,-nbitq), 
to_sfixed(1505.0/65536.0,1,-nbitq), 
to_sfixed(42.0/65536.0,1,-nbitq), 
to_sfixed(-1507.0/65536.0,1,-nbitq), 
to_sfixed(-5072.0/65536.0,1,-nbitq), 
to_sfixed(-1514.0/65536.0,1,-nbitq), 
to_sfixed(1722.0/65536.0,1,-nbitq), 
to_sfixed(-2116.0/65536.0,1,-nbitq), 
to_sfixed(2145.0/65536.0,1,-nbitq), 
to_sfixed(3404.0/65536.0,1,-nbitq), 
to_sfixed(-952.0/65536.0,1,-nbitq), 
to_sfixed(3008.0/65536.0,1,-nbitq), 
to_sfixed(-1498.0/65536.0,1,-nbitq), 
to_sfixed(2384.0/65536.0,1,-nbitq), 
to_sfixed(-244.0/65536.0,1,-nbitq), 
to_sfixed(-1255.0/65536.0,1,-nbitq), 
to_sfixed(6319.0/65536.0,1,-nbitq), 
to_sfixed(-2856.0/65536.0,1,-nbitq), 
to_sfixed(-1322.0/65536.0,1,-nbitq), 
to_sfixed(3102.0/65536.0,1,-nbitq), 
to_sfixed(-1244.0/65536.0,1,-nbitq), 
to_sfixed(952.0/65536.0,1,-nbitq), 
to_sfixed(-2556.0/65536.0,1,-nbitq), 
to_sfixed(3206.0/65536.0,1,-nbitq), 
to_sfixed(-4069.0/65536.0,1,-nbitq), 
to_sfixed(228.0/65536.0,1,-nbitq), 
to_sfixed(-496.0/65536.0,1,-nbitq), 
to_sfixed(1018.0/65536.0,1,-nbitq), 
to_sfixed(-765.0/65536.0,1,-nbitq), 
to_sfixed(75.0/65536.0,1,-nbitq), 
to_sfixed(886.0/65536.0,1,-nbitq), 
to_sfixed(-3092.0/65536.0,1,-nbitq), 
to_sfixed(-1687.0/65536.0,1,-nbitq), 
to_sfixed(-5707.0/65536.0,1,-nbitq), 
to_sfixed(2925.0/65536.0,1,-nbitq), 
to_sfixed(-1167.0/65536.0,1,-nbitq), 
to_sfixed(5098.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-604.0/65536.0,1,-nbitq), 
to_sfixed(3991.0/65536.0,1,-nbitq), 
to_sfixed(515.0/65536.0,1,-nbitq), 
to_sfixed(-2762.0/65536.0,1,-nbitq), 
to_sfixed(-5281.0/65536.0,1,-nbitq), 
to_sfixed(-5216.0/65536.0,1,-nbitq), 
to_sfixed(29.0/65536.0,1,-nbitq), 
to_sfixed(-1388.0/65536.0,1,-nbitq), 
to_sfixed(-1496.0/65536.0,1,-nbitq), 
to_sfixed(1833.0/65536.0,1,-nbitq), 
to_sfixed(-1713.0/65536.0,1,-nbitq), 
to_sfixed(-3035.0/65536.0,1,-nbitq), 
to_sfixed(-2448.0/65536.0,1,-nbitq), 
to_sfixed(-4030.0/65536.0,1,-nbitq), 
to_sfixed(2378.0/65536.0,1,-nbitq), 
to_sfixed(-2421.0/65536.0,1,-nbitq), 
to_sfixed(-1674.0/65536.0,1,-nbitq), 
to_sfixed(-2352.0/65536.0,1,-nbitq), 
to_sfixed(-4065.0/65536.0,1,-nbitq), 
to_sfixed(2603.0/65536.0,1,-nbitq), 
to_sfixed(771.0/65536.0,1,-nbitq), 
to_sfixed(4601.0/65536.0,1,-nbitq), 
to_sfixed(2452.0/65536.0,1,-nbitq), 
to_sfixed(-2191.0/65536.0,1,-nbitq), 
to_sfixed(-543.0/65536.0,1,-nbitq), 
to_sfixed(-850.0/65536.0,1,-nbitq), 
to_sfixed(-4020.0/65536.0,1,-nbitq), 
to_sfixed(-3314.0/65536.0,1,-nbitq), 
to_sfixed(-6404.0/65536.0,1,-nbitq), 
to_sfixed(1632.0/65536.0,1,-nbitq), 
to_sfixed(2332.0/65536.0,1,-nbitq), 
to_sfixed(-2283.0/65536.0,1,-nbitq), 
to_sfixed(13.0/65536.0,1,-nbitq), 
to_sfixed(3925.0/65536.0,1,-nbitq), 
to_sfixed(-926.0/65536.0,1,-nbitq), 
to_sfixed(1614.0/65536.0,1,-nbitq), 
to_sfixed(-407.0/65536.0,1,-nbitq), 
to_sfixed(-1171.0/65536.0,1,-nbitq), 
to_sfixed(74.0/65536.0,1,-nbitq), 
to_sfixed(1045.0/65536.0,1,-nbitq), 
to_sfixed(2180.0/65536.0,1,-nbitq), 
to_sfixed(1090.0/65536.0,1,-nbitq), 
to_sfixed(-2019.0/65536.0,1,-nbitq), 
to_sfixed(3816.0/65536.0,1,-nbitq), 
to_sfixed(-1092.0/65536.0,1,-nbitq), 
to_sfixed(2147.0/65536.0,1,-nbitq), 
to_sfixed(3087.0/65536.0,1,-nbitq), 
to_sfixed(-4320.0/65536.0,1,-nbitq), 
to_sfixed(-851.0/65536.0,1,-nbitq), 
to_sfixed(3579.0/65536.0,1,-nbitq), 
to_sfixed(-2150.0/65536.0,1,-nbitq), 
to_sfixed(-1103.0/65536.0,1,-nbitq), 
to_sfixed(1910.0/65536.0,1,-nbitq), 
to_sfixed(-4535.0/65536.0,1,-nbitq), 
to_sfixed(3674.0/65536.0,1,-nbitq), 
to_sfixed(-689.0/65536.0,1,-nbitq), 
to_sfixed(72.0/65536.0,1,-nbitq), 
to_sfixed(552.0/65536.0,1,-nbitq), 
to_sfixed(1967.0/65536.0,1,-nbitq), 
to_sfixed(2659.0/65536.0,1,-nbitq), 
to_sfixed(365.0/65536.0,1,-nbitq), 
to_sfixed(-2570.0/65536.0,1,-nbitq), 
to_sfixed(328.0/65536.0,1,-nbitq), 
to_sfixed(1646.0/65536.0,1,-nbitq), 
to_sfixed(3831.0/65536.0,1,-nbitq), 
to_sfixed(-22.0/65536.0,1,-nbitq), 
to_sfixed(-1020.0/65536.0,1,-nbitq), 
to_sfixed(-296.0/65536.0,1,-nbitq), 
to_sfixed(3785.0/65536.0,1,-nbitq), 
to_sfixed(-2390.0/65536.0,1,-nbitq), 
to_sfixed(4355.0/65536.0,1,-nbitq), 
to_sfixed(-4601.0/65536.0,1,-nbitq), 
to_sfixed(-3115.0/65536.0,1,-nbitq), 
to_sfixed(-1485.0/65536.0,1,-nbitq), 
to_sfixed(-894.0/65536.0,1,-nbitq), 
to_sfixed(-1068.0/65536.0,1,-nbitq), 
to_sfixed(-3911.0/65536.0,1,-nbitq), 
to_sfixed(1979.0/65536.0,1,-nbitq), 
to_sfixed(-2666.0/65536.0,1,-nbitq), 
to_sfixed(2265.0/65536.0,1,-nbitq)  ), 
( to_sfixed(273.0/65536.0,1,-nbitq), 
to_sfixed(2265.0/65536.0,1,-nbitq), 
to_sfixed(-3995.0/65536.0,1,-nbitq), 
to_sfixed(522.0/65536.0,1,-nbitq), 
to_sfixed(-3199.0/65536.0,1,-nbitq), 
to_sfixed(-3490.0/65536.0,1,-nbitq), 
to_sfixed(-4107.0/65536.0,1,-nbitq), 
to_sfixed(-3269.0/65536.0,1,-nbitq), 
to_sfixed(1259.0/65536.0,1,-nbitq), 
to_sfixed(2276.0/65536.0,1,-nbitq), 
to_sfixed(-4434.0/65536.0,1,-nbitq), 
to_sfixed(2672.0/65536.0,1,-nbitq), 
to_sfixed(-2134.0/65536.0,1,-nbitq), 
to_sfixed(601.0/65536.0,1,-nbitq), 
to_sfixed(2742.0/65536.0,1,-nbitq), 
to_sfixed(2646.0/65536.0,1,-nbitq), 
to_sfixed(-2313.0/65536.0,1,-nbitq), 
to_sfixed(-1533.0/65536.0,1,-nbitq), 
to_sfixed(-2384.0/65536.0,1,-nbitq), 
to_sfixed(-1562.0/65536.0,1,-nbitq), 
to_sfixed(-702.0/65536.0,1,-nbitq), 
to_sfixed(2544.0/65536.0,1,-nbitq), 
to_sfixed(-462.0/65536.0,1,-nbitq), 
to_sfixed(-1650.0/65536.0,1,-nbitq), 
to_sfixed(3222.0/65536.0,1,-nbitq), 
to_sfixed(-1927.0/65536.0,1,-nbitq), 
to_sfixed(496.0/65536.0,1,-nbitq), 
to_sfixed(-1471.0/65536.0,1,-nbitq), 
to_sfixed(-4873.0/65536.0,1,-nbitq), 
to_sfixed(-1891.0/65536.0,1,-nbitq), 
to_sfixed(542.0/65536.0,1,-nbitq), 
to_sfixed(-1216.0/65536.0,1,-nbitq), 
to_sfixed(-2303.0/65536.0,1,-nbitq), 
to_sfixed(2590.0/65536.0,1,-nbitq), 
to_sfixed(-505.0/65536.0,1,-nbitq), 
to_sfixed(1385.0/65536.0,1,-nbitq), 
to_sfixed(-1194.0/65536.0,1,-nbitq), 
to_sfixed(1129.0/65536.0,1,-nbitq), 
to_sfixed(2211.0/65536.0,1,-nbitq), 
to_sfixed(-2259.0/65536.0,1,-nbitq), 
to_sfixed(-3005.0/65536.0,1,-nbitq), 
to_sfixed(1660.0/65536.0,1,-nbitq), 
to_sfixed(-1023.0/65536.0,1,-nbitq), 
to_sfixed(-2089.0/65536.0,1,-nbitq), 
to_sfixed(2748.0/65536.0,1,-nbitq), 
to_sfixed(2281.0/65536.0,1,-nbitq), 
to_sfixed(335.0/65536.0,1,-nbitq), 
to_sfixed(-1962.0/65536.0,1,-nbitq), 
to_sfixed(2213.0/65536.0,1,-nbitq), 
to_sfixed(2984.0/65536.0,1,-nbitq), 
to_sfixed(-306.0/65536.0,1,-nbitq), 
to_sfixed(-2596.0/65536.0,1,-nbitq), 
to_sfixed(2376.0/65536.0,1,-nbitq), 
to_sfixed(-2839.0/65536.0,1,-nbitq), 
to_sfixed(4607.0/65536.0,1,-nbitq), 
to_sfixed(-2502.0/65536.0,1,-nbitq), 
to_sfixed(2049.0/65536.0,1,-nbitq), 
to_sfixed(-2266.0/65536.0,1,-nbitq), 
to_sfixed(-2034.0/65536.0,1,-nbitq), 
to_sfixed(7236.0/65536.0,1,-nbitq), 
to_sfixed(-3074.0/65536.0,1,-nbitq), 
to_sfixed(792.0/65536.0,1,-nbitq), 
to_sfixed(1642.0/65536.0,1,-nbitq), 
to_sfixed(-787.0/65536.0,1,-nbitq), 
to_sfixed(235.0/65536.0,1,-nbitq), 
to_sfixed(3696.0/65536.0,1,-nbitq), 
to_sfixed(-1010.0/65536.0,1,-nbitq), 
to_sfixed(-1174.0/65536.0,1,-nbitq), 
to_sfixed(-1136.0/65536.0,1,-nbitq), 
to_sfixed(-3759.0/65536.0,1,-nbitq), 
to_sfixed(717.0/65536.0,1,-nbitq), 
to_sfixed(-589.0/65536.0,1,-nbitq), 
to_sfixed(-2418.0/65536.0,1,-nbitq), 
to_sfixed(-1391.0/65536.0,1,-nbitq), 
to_sfixed(-809.0/65536.0,1,-nbitq), 
to_sfixed(1590.0/65536.0,1,-nbitq), 
to_sfixed(-4153.0/65536.0,1,-nbitq), 
to_sfixed(3025.0/65536.0,1,-nbitq), 
to_sfixed(-2726.0/65536.0,1,-nbitq), 
to_sfixed(2469.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1356.0/65536.0,1,-nbitq), 
to_sfixed(3484.0/65536.0,1,-nbitq), 
to_sfixed(474.0/65536.0,1,-nbitq), 
to_sfixed(-1433.0/65536.0,1,-nbitq), 
to_sfixed(-712.0/65536.0,1,-nbitq), 
to_sfixed(109.0/65536.0,1,-nbitq), 
to_sfixed(922.0/65536.0,1,-nbitq), 
to_sfixed(-1350.0/65536.0,1,-nbitq), 
to_sfixed(2491.0/65536.0,1,-nbitq), 
to_sfixed(-381.0/65536.0,1,-nbitq), 
to_sfixed(-1481.0/65536.0,1,-nbitq), 
to_sfixed(-1073.0/65536.0,1,-nbitq), 
to_sfixed(-1496.0/65536.0,1,-nbitq), 
to_sfixed(1428.0/65536.0,1,-nbitq), 
to_sfixed(845.0/65536.0,1,-nbitq), 
to_sfixed(-1444.0/65536.0,1,-nbitq), 
to_sfixed(-527.0/65536.0,1,-nbitq), 
to_sfixed(-131.0/65536.0,1,-nbitq), 
to_sfixed(-2448.0/65536.0,1,-nbitq), 
to_sfixed(-1518.0/65536.0,1,-nbitq), 
to_sfixed(43.0/65536.0,1,-nbitq), 
to_sfixed(845.0/65536.0,1,-nbitq), 
to_sfixed(825.0/65536.0,1,-nbitq), 
to_sfixed(-1528.0/65536.0,1,-nbitq), 
to_sfixed(-1499.0/65536.0,1,-nbitq), 
to_sfixed(-1663.0/65536.0,1,-nbitq), 
to_sfixed(-194.0/65536.0,1,-nbitq), 
to_sfixed(672.0/65536.0,1,-nbitq), 
to_sfixed(-3519.0/65536.0,1,-nbitq), 
to_sfixed(1534.0/65536.0,1,-nbitq), 
to_sfixed(-945.0/65536.0,1,-nbitq), 
to_sfixed(-2866.0/65536.0,1,-nbitq), 
to_sfixed(2306.0/65536.0,1,-nbitq), 
to_sfixed(16.0/65536.0,1,-nbitq), 
to_sfixed(933.0/65536.0,1,-nbitq), 
to_sfixed(42.0/65536.0,1,-nbitq), 
to_sfixed(-4510.0/65536.0,1,-nbitq), 
to_sfixed(-4069.0/65536.0,1,-nbitq), 
to_sfixed(1046.0/65536.0,1,-nbitq), 
to_sfixed(1352.0/65536.0,1,-nbitq), 
to_sfixed(-1349.0/65536.0,1,-nbitq), 
to_sfixed(-2984.0/65536.0,1,-nbitq), 
to_sfixed(-1908.0/65536.0,1,-nbitq), 
to_sfixed(-1740.0/65536.0,1,-nbitq), 
to_sfixed(1746.0/65536.0,1,-nbitq), 
to_sfixed(3145.0/65536.0,1,-nbitq), 
to_sfixed(-1972.0/65536.0,1,-nbitq), 
to_sfixed(468.0/65536.0,1,-nbitq), 
to_sfixed(2174.0/65536.0,1,-nbitq), 
to_sfixed(3381.0/65536.0,1,-nbitq), 
to_sfixed(-2182.0/65536.0,1,-nbitq), 
to_sfixed(-2579.0/65536.0,1,-nbitq), 
to_sfixed(948.0/65536.0,1,-nbitq), 
to_sfixed(1348.0/65536.0,1,-nbitq), 
to_sfixed(4010.0/65536.0,1,-nbitq), 
to_sfixed(-1021.0/65536.0,1,-nbitq), 
to_sfixed(-271.0/65536.0,1,-nbitq), 
to_sfixed(586.0/65536.0,1,-nbitq), 
to_sfixed(2284.0/65536.0,1,-nbitq), 
to_sfixed(5812.0/65536.0,1,-nbitq), 
to_sfixed(-785.0/65536.0,1,-nbitq), 
to_sfixed(-1435.0/65536.0,1,-nbitq), 
to_sfixed(1456.0/65536.0,1,-nbitq), 
to_sfixed(-1115.0/65536.0,1,-nbitq), 
to_sfixed(1170.0/65536.0,1,-nbitq), 
to_sfixed(4502.0/65536.0,1,-nbitq), 
to_sfixed(1032.0/65536.0,1,-nbitq), 
to_sfixed(1852.0/65536.0,1,-nbitq), 
to_sfixed(2620.0/65536.0,1,-nbitq), 
to_sfixed(-1029.0/65536.0,1,-nbitq), 
to_sfixed(-1658.0/65536.0,1,-nbitq), 
to_sfixed(-3785.0/65536.0,1,-nbitq), 
to_sfixed(-2951.0/65536.0,1,-nbitq), 
to_sfixed(-1679.0/65536.0,1,-nbitq), 
to_sfixed(-3115.0/65536.0,1,-nbitq), 
to_sfixed(938.0/65536.0,1,-nbitq), 
to_sfixed(-2460.0/65536.0,1,-nbitq), 
to_sfixed(1455.0/65536.0,1,-nbitq), 
to_sfixed(2348.0/65536.0,1,-nbitq), 
to_sfixed(1833.0/65536.0,1,-nbitq)  ), 
( to_sfixed(479.0/65536.0,1,-nbitq), 
to_sfixed(2312.0/65536.0,1,-nbitq), 
to_sfixed(-1585.0/65536.0,1,-nbitq), 
to_sfixed(-1771.0/65536.0,1,-nbitq), 
to_sfixed(-1210.0/65536.0,1,-nbitq), 
to_sfixed(2845.0/65536.0,1,-nbitq), 
to_sfixed(-2005.0/65536.0,1,-nbitq), 
to_sfixed(89.0/65536.0,1,-nbitq), 
to_sfixed(174.0/65536.0,1,-nbitq), 
to_sfixed(-199.0/65536.0,1,-nbitq), 
to_sfixed(204.0/65536.0,1,-nbitq), 
to_sfixed(157.0/65536.0,1,-nbitq), 
to_sfixed(-2568.0/65536.0,1,-nbitq), 
to_sfixed(-2085.0/65536.0,1,-nbitq), 
to_sfixed(1017.0/65536.0,1,-nbitq), 
to_sfixed(613.0/65536.0,1,-nbitq), 
to_sfixed(2193.0/65536.0,1,-nbitq), 
to_sfixed(-1489.0/65536.0,1,-nbitq), 
to_sfixed(-1908.0/65536.0,1,-nbitq), 
to_sfixed(1891.0/65536.0,1,-nbitq), 
to_sfixed(-2844.0/65536.0,1,-nbitq), 
to_sfixed(1043.0/65536.0,1,-nbitq), 
to_sfixed(1298.0/65536.0,1,-nbitq), 
to_sfixed(1934.0/65536.0,1,-nbitq), 
to_sfixed(166.0/65536.0,1,-nbitq), 
to_sfixed(-2923.0/65536.0,1,-nbitq), 
to_sfixed(-1944.0/65536.0,1,-nbitq), 
to_sfixed(-3003.0/65536.0,1,-nbitq), 
to_sfixed(1285.0/65536.0,1,-nbitq), 
to_sfixed(-1783.0/65536.0,1,-nbitq), 
to_sfixed(859.0/65536.0,1,-nbitq), 
to_sfixed(942.0/65536.0,1,-nbitq), 
to_sfixed(2042.0/65536.0,1,-nbitq), 
to_sfixed(4381.0/65536.0,1,-nbitq), 
to_sfixed(-1832.0/65536.0,1,-nbitq), 
to_sfixed(-971.0/65536.0,1,-nbitq), 
to_sfixed(-398.0/65536.0,1,-nbitq), 
to_sfixed(-640.0/65536.0,1,-nbitq), 
to_sfixed(721.0/65536.0,1,-nbitq), 
to_sfixed(-312.0/65536.0,1,-nbitq), 
to_sfixed(-3638.0/65536.0,1,-nbitq), 
to_sfixed(460.0/65536.0,1,-nbitq), 
to_sfixed(-4422.0/65536.0,1,-nbitq), 
to_sfixed(503.0/65536.0,1,-nbitq), 
to_sfixed(1723.0/65536.0,1,-nbitq), 
to_sfixed(3439.0/65536.0,1,-nbitq), 
to_sfixed(168.0/65536.0,1,-nbitq), 
to_sfixed(-2007.0/65536.0,1,-nbitq), 
to_sfixed(-933.0/65536.0,1,-nbitq), 
to_sfixed(762.0/65536.0,1,-nbitq), 
to_sfixed(-2543.0/65536.0,1,-nbitq), 
to_sfixed(-443.0/65536.0,1,-nbitq), 
to_sfixed(821.0/65536.0,1,-nbitq), 
to_sfixed(-2037.0/65536.0,1,-nbitq), 
to_sfixed(-309.0/65536.0,1,-nbitq), 
to_sfixed(1705.0/65536.0,1,-nbitq), 
to_sfixed(-1332.0/65536.0,1,-nbitq), 
to_sfixed(-2973.0/65536.0,1,-nbitq), 
to_sfixed(1850.0/65536.0,1,-nbitq), 
to_sfixed(2839.0/65536.0,1,-nbitq), 
to_sfixed(251.0/65536.0,1,-nbitq), 
to_sfixed(-2588.0/65536.0,1,-nbitq), 
to_sfixed(-683.0/65536.0,1,-nbitq), 
to_sfixed(165.0/65536.0,1,-nbitq), 
to_sfixed(1070.0/65536.0,1,-nbitq), 
to_sfixed(4565.0/65536.0,1,-nbitq), 
to_sfixed(-191.0/65536.0,1,-nbitq), 
to_sfixed(-607.0/65536.0,1,-nbitq), 
to_sfixed(-2456.0/65536.0,1,-nbitq), 
to_sfixed(-950.0/65536.0,1,-nbitq), 
to_sfixed(-513.0/65536.0,1,-nbitq), 
to_sfixed(950.0/65536.0,1,-nbitq), 
to_sfixed(2064.0/65536.0,1,-nbitq), 
to_sfixed(-2729.0/65536.0,1,-nbitq), 
to_sfixed(2558.0/65536.0,1,-nbitq), 
to_sfixed(-901.0/65536.0,1,-nbitq), 
to_sfixed(518.0/65536.0,1,-nbitq), 
to_sfixed(3997.0/65536.0,1,-nbitq), 
to_sfixed(-2918.0/65536.0,1,-nbitq), 
to_sfixed(4005.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3952.0/65536.0,1,-nbitq), 
to_sfixed(-310.0/65536.0,1,-nbitq), 
to_sfixed(1195.0/65536.0,1,-nbitq), 
to_sfixed(488.0/65536.0,1,-nbitq), 
to_sfixed(546.0/65536.0,1,-nbitq), 
to_sfixed(1964.0/65536.0,1,-nbitq), 
to_sfixed(-3126.0/65536.0,1,-nbitq), 
to_sfixed(-1797.0/65536.0,1,-nbitq), 
to_sfixed(-243.0/65536.0,1,-nbitq), 
to_sfixed(40.0/65536.0,1,-nbitq), 
to_sfixed(3571.0/65536.0,1,-nbitq), 
to_sfixed(-1683.0/65536.0,1,-nbitq), 
to_sfixed(250.0/65536.0,1,-nbitq), 
to_sfixed(-2145.0/65536.0,1,-nbitq), 
to_sfixed(117.0/65536.0,1,-nbitq), 
to_sfixed(2488.0/65536.0,1,-nbitq), 
to_sfixed(-464.0/65536.0,1,-nbitq), 
to_sfixed(710.0/65536.0,1,-nbitq), 
to_sfixed(-3168.0/65536.0,1,-nbitq), 
to_sfixed(2604.0/65536.0,1,-nbitq), 
to_sfixed(-4414.0/65536.0,1,-nbitq), 
to_sfixed(993.0/65536.0,1,-nbitq), 
to_sfixed(2624.0/65536.0,1,-nbitq), 
to_sfixed(1621.0/65536.0,1,-nbitq), 
to_sfixed(-1761.0/65536.0,1,-nbitq), 
to_sfixed(-3109.0/65536.0,1,-nbitq), 
to_sfixed(1590.0/65536.0,1,-nbitq), 
to_sfixed(1155.0/65536.0,1,-nbitq), 
to_sfixed(-2631.0/65536.0,1,-nbitq), 
to_sfixed(1449.0/65536.0,1,-nbitq), 
to_sfixed(2044.0/65536.0,1,-nbitq), 
to_sfixed(-1352.0/65536.0,1,-nbitq), 
to_sfixed(523.0/65536.0,1,-nbitq), 
to_sfixed(320.0/65536.0,1,-nbitq), 
to_sfixed(-1444.0/65536.0,1,-nbitq), 
to_sfixed(1327.0/65536.0,1,-nbitq), 
to_sfixed(-1878.0/65536.0,1,-nbitq), 
to_sfixed(-2935.0/65536.0,1,-nbitq), 
to_sfixed(-1970.0/65536.0,1,-nbitq), 
to_sfixed(-643.0/65536.0,1,-nbitq), 
to_sfixed(-2996.0/65536.0,1,-nbitq), 
to_sfixed(-3189.0/65536.0,1,-nbitq), 
to_sfixed(-2427.0/65536.0,1,-nbitq), 
to_sfixed(-1543.0/65536.0,1,-nbitq), 
to_sfixed(-587.0/65536.0,1,-nbitq), 
to_sfixed(583.0/65536.0,1,-nbitq), 
to_sfixed(-2254.0/65536.0,1,-nbitq), 
to_sfixed(-1949.0/65536.0,1,-nbitq), 
to_sfixed(1709.0/65536.0,1,-nbitq), 
to_sfixed(-186.0/65536.0,1,-nbitq), 
to_sfixed(1332.0/65536.0,1,-nbitq), 
to_sfixed(-1120.0/65536.0,1,-nbitq), 
to_sfixed(-2139.0/65536.0,1,-nbitq), 
to_sfixed(-1873.0/65536.0,1,-nbitq), 
to_sfixed(255.0/65536.0,1,-nbitq), 
to_sfixed(416.0/65536.0,1,-nbitq), 
to_sfixed(-1220.0/65536.0,1,-nbitq), 
to_sfixed(913.0/65536.0,1,-nbitq), 
to_sfixed(2606.0/65536.0,1,-nbitq), 
to_sfixed(5551.0/65536.0,1,-nbitq), 
to_sfixed(-1583.0/65536.0,1,-nbitq), 
to_sfixed(2473.0/65536.0,1,-nbitq), 
to_sfixed(1869.0/65536.0,1,-nbitq), 
to_sfixed(242.0/65536.0,1,-nbitq), 
to_sfixed(2738.0/65536.0,1,-nbitq), 
to_sfixed(949.0/65536.0,1,-nbitq), 
to_sfixed(-2133.0/65536.0,1,-nbitq), 
to_sfixed(3175.0/65536.0,1,-nbitq), 
to_sfixed(2052.0/65536.0,1,-nbitq), 
to_sfixed(-1428.0/65536.0,1,-nbitq), 
to_sfixed(2144.0/65536.0,1,-nbitq), 
to_sfixed(-1573.0/65536.0,1,-nbitq), 
to_sfixed(-902.0/65536.0,1,-nbitq), 
to_sfixed(-1967.0/65536.0,1,-nbitq), 
to_sfixed(-993.0/65536.0,1,-nbitq), 
to_sfixed(-434.0/65536.0,1,-nbitq), 
to_sfixed(-2508.0/65536.0,1,-nbitq), 
to_sfixed(1717.0/65536.0,1,-nbitq), 
to_sfixed(2674.0/65536.0,1,-nbitq), 
to_sfixed(3628.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2795.0/65536.0,1,-nbitq), 
to_sfixed(37.0/65536.0,1,-nbitq), 
to_sfixed(357.0/65536.0,1,-nbitq), 
to_sfixed(1331.0/65536.0,1,-nbitq), 
to_sfixed(2412.0/65536.0,1,-nbitq), 
to_sfixed(84.0/65536.0,1,-nbitq), 
to_sfixed(1909.0/65536.0,1,-nbitq), 
to_sfixed(1041.0/65536.0,1,-nbitq), 
to_sfixed(-1029.0/65536.0,1,-nbitq), 
to_sfixed(2854.0/65536.0,1,-nbitq), 
to_sfixed(2412.0/65536.0,1,-nbitq), 
to_sfixed(-451.0/65536.0,1,-nbitq), 
to_sfixed(662.0/65536.0,1,-nbitq), 
to_sfixed(-2452.0/65536.0,1,-nbitq), 
to_sfixed(1801.0/65536.0,1,-nbitq), 
to_sfixed(2677.0/65536.0,1,-nbitq), 
to_sfixed(-3131.0/65536.0,1,-nbitq), 
to_sfixed(-3286.0/65536.0,1,-nbitq), 
to_sfixed(-109.0/65536.0,1,-nbitq), 
to_sfixed(707.0/65536.0,1,-nbitq), 
to_sfixed(-3754.0/65536.0,1,-nbitq), 
to_sfixed(-520.0/65536.0,1,-nbitq), 
to_sfixed(2001.0/65536.0,1,-nbitq), 
to_sfixed(-1386.0/65536.0,1,-nbitq), 
to_sfixed(108.0/65536.0,1,-nbitq), 
to_sfixed(-2119.0/65536.0,1,-nbitq), 
to_sfixed(2234.0/65536.0,1,-nbitq), 
to_sfixed(-423.0/65536.0,1,-nbitq), 
to_sfixed(-1562.0/65536.0,1,-nbitq), 
to_sfixed(-2239.0/65536.0,1,-nbitq), 
to_sfixed(880.0/65536.0,1,-nbitq), 
to_sfixed(1864.0/65536.0,1,-nbitq), 
to_sfixed(637.0/65536.0,1,-nbitq), 
to_sfixed(2256.0/65536.0,1,-nbitq), 
to_sfixed(-1540.0/65536.0,1,-nbitq), 
to_sfixed(12.0/65536.0,1,-nbitq), 
to_sfixed(-16.0/65536.0,1,-nbitq), 
to_sfixed(-3789.0/65536.0,1,-nbitq), 
to_sfixed(52.0/65536.0,1,-nbitq), 
to_sfixed(2452.0/65536.0,1,-nbitq), 
to_sfixed(-2021.0/65536.0,1,-nbitq), 
to_sfixed(-2874.0/65536.0,1,-nbitq), 
to_sfixed(-2383.0/65536.0,1,-nbitq), 
to_sfixed(2209.0/65536.0,1,-nbitq), 
to_sfixed(184.0/65536.0,1,-nbitq), 
to_sfixed(1116.0/65536.0,1,-nbitq), 
to_sfixed(47.0/65536.0,1,-nbitq), 
to_sfixed(-3651.0/65536.0,1,-nbitq), 
to_sfixed(-1647.0/65536.0,1,-nbitq), 
to_sfixed(4007.0/65536.0,1,-nbitq), 
to_sfixed(962.0/65536.0,1,-nbitq), 
to_sfixed(-1655.0/65536.0,1,-nbitq), 
to_sfixed(1213.0/65536.0,1,-nbitq), 
to_sfixed(-3578.0/65536.0,1,-nbitq), 
to_sfixed(1736.0/65536.0,1,-nbitq), 
to_sfixed(1297.0/65536.0,1,-nbitq), 
to_sfixed(-815.0/65536.0,1,-nbitq), 
to_sfixed(134.0/65536.0,1,-nbitq), 
to_sfixed(53.0/65536.0,1,-nbitq), 
to_sfixed(6515.0/65536.0,1,-nbitq), 
to_sfixed(-1105.0/65536.0,1,-nbitq), 
to_sfixed(-2761.0/65536.0,1,-nbitq), 
to_sfixed(-1144.0/65536.0,1,-nbitq), 
to_sfixed(-1178.0/65536.0,1,-nbitq), 
to_sfixed(2827.0/65536.0,1,-nbitq), 
to_sfixed(2637.0/65536.0,1,-nbitq), 
to_sfixed(-2046.0/65536.0,1,-nbitq), 
to_sfixed(1037.0/65536.0,1,-nbitq), 
to_sfixed(696.0/65536.0,1,-nbitq), 
to_sfixed(884.0/65536.0,1,-nbitq), 
to_sfixed(3741.0/65536.0,1,-nbitq), 
to_sfixed(1462.0/65536.0,1,-nbitq), 
to_sfixed(1276.0/65536.0,1,-nbitq), 
to_sfixed(1175.0/65536.0,1,-nbitq), 
to_sfixed(2074.0/65536.0,1,-nbitq), 
to_sfixed(-798.0/65536.0,1,-nbitq), 
to_sfixed(-3347.0/65536.0,1,-nbitq), 
to_sfixed(40.0/65536.0,1,-nbitq), 
to_sfixed(1793.0/65536.0,1,-nbitq), 
to_sfixed(3214.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-632.0/65536.0,1,-nbitq), 
to_sfixed(-1185.0/65536.0,1,-nbitq), 
to_sfixed(572.0/65536.0,1,-nbitq), 
to_sfixed(-1940.0/65536.0,1,-nbitq), 
to_sfixed(-2910.0/65536.0,1,-nbitq), 
to_sfixed(-2953.0/65536.0,1,-nbitq), 
to_sfixed(-3561.0/65536.0,1,-nbitq), 
to_sfixed(-90.0/65536.0,1,-nbitq), 
to_sfixed(-3015.0/65536.0,1,-nbitq), 
to_sfixed(-248.0/65536.0,1,-nbitq), 
to_sfixed(2484.0/65536.0,1,-nbitq), 
to_sfixed(-2926.0/65536.0,1,-nbitq), 
to_sfixed(-2428.0/65536.0,1,-nbitq), 
to_sfixed(-1143.0/65536.0,1,-nbitq), 
to_sfixed(3738.0/65536.0,1,-nbitq), 
to_sfixed(-804.0/65536.0,1,-nbitq), 
to_sfixed(-2971.0/65536.0,1,-nbitq), 
to_sfixed(-2652.0/65536.0,1,-nbitq), 
to_sfixed(-1984.0/65536.0,1,-nbitq), 
to_sfixed(1916.0/65536.0,1,-nbitq), 
to_sfixed(-912.0/65536.0,1,-nbitq), 
to_sfixed(-769.0/65536.0,1,-nbitq), 
to_sfixed(377.0/65536.0,1,-nbitq), 
to_sfixed(1667.0/65536.0,1,-nbitq), 
to_sfixed(1129.0/65536.0,1,-nbitq), 
to_sfixed(2012.0/65536.0,1,-nbitq), 
to_sfixed(-746.0/65536.0,1,-nbitq), 
to_sfixed(1418.0/65536.0,1,-nbitq), 
to_sfixed(-1144.0/65536.0,1,-nbitq), 
to_sfixed(-2387.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(1202.0/65536.0,1,-nbitq), 
to_sfixed(-2641.0/65536.0,1,-nbitq), 
to_sfixed(474.0/65536.0,1,-nbitq), 
to_sfixed(1054.0/65536.0,1,-nbitq), 
to_sfixed(-31.0/65536.0,1,-nbitq), 
to_sfixed(159.0/65536.0,1,-nbitq), 
to_sfixed(-770.0/65536.0,1,-nbitq), 
to_sfixed(-1278.0/65536.0,1,-nbitq), 
to_sfixed(31.0/65536.0,1,-nbitq), 
to_sfixed(2718.0/65536.0,1,-nbitq), 
to_sfixed(-974.0/65536.0,1,-nbitq), 
to_sfixed(-4029.0/65536.0,1,-nbitq), 
to_sfixed(-603.0/65536.0,1,-nbitq), 
to_sfixed(1470.0/65536.0,1,-nbitq), 
to_sfixed(3535.0/65536.0,1,-nbitq), 
to_sfixed(2998.0/65536.0,1,-nbitq), 
to_sfixed(-3273.0/65536.0,1,-nbitq), 
to_sfixed(2102.0/65536.0,1,-nbitq), 
to_sfixed(2382.0/65536.0,1,-nbitq), 
to_sfixed(-210.0/65536.0,1,-nbitq), 
to_sfixed(314.0/65536.0,1,-nbitq), 
to_sfixed(580.0/65536.0,1,-nbitq), 
to_sfixed(-1203.0/65536.0,1,-nbitq), 
to_sfixed(3549.0/65536.0,1,-nbitq), 
to_sfixed(-1291.0/65536.0,1,-nbitq), 
to_sfixed(-2293.0/65536.0,1,-nbitq), 
to_sfixed(2758.0/65536.0,1,-nbitq), 
to_sfixed(-760.0/65536.0,1,-nbitq), 
to_sfixed(5328.0/65536.0,1,-nbitq), 
to_sfixed(-3707.0/65536.0,1,-nbitq), 
to_sfixed(-2526.0/65536.0,1,-nbitq), 
to_sfixed(2641.0/65536.0,1,-nbitq), 
to_sfixed(1842.0/65536.0,1,-nbitq), 
to_sfixed(3887.0/65536.0,1,-nbitq), 
to_sfixed(3833.0/65536.0,1,-nbitq), 
to_sfixed(-2870.0/65536.0,1,-nbitq), 
to_sfixed(273.0/65536.0,1,-nbitq), 
to_sfixed(3701.0/65536.0,1,-nbitq), 
to_sfixed(-1254.0/65536.0,1,-nbitq), 
to_sfixed(3077.0/65536.0,1,-nbitq), 
to_sfixed(-2796.0/65536.0,1,-nbitq), 
to_sfixed(3469.0/65536.0,1,-nbitq), 
to_sfixed(2227.0/65536.0,1,-nbitq), 
to_sfixed(132.0/65536.0,1,-nbitq), 
to_sfixed(517.0/65536.0,1,-nbitq), 
to_sfixed(-2722.0/65536.0,1,-nbitq), 
to_sfixed(3666.0/65536.0,1,-nbitq), 
to_sfixed(-3102.0/65536.0,1,-nbitq), 
to_sfixed(1957.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2222.0/65536.0,1,-nbitq), 
to_sfixed(644.0/65536.0,1,-nbitq), 
to_sfixed(488.0/65536.0,1,-nbitq), 
to_sfixed(-518.0/65536.0,1,-nbitq), 
to_sfixed(-1787.0/65536.0,1,-nbitq), 
to_sfixed(1644.0/65536.0,1,-nbitq), 
to_sfixed(1851.0/65536.0,1,-nbitq), 
to_sfixed(1041.0/65536.0,1,-nbitq), 
to_sfixed(2423.0/65536.0,1,-nbitq), 
to_sfixed(-174.0/65536.0,1,-nbitq), 
to_sfixed(-1622.0/65536.0,1,-nbitq), 
to_sfixed(-3728.0/65536.0,1,-nbitq), 
to_sfixed(-1965.0/65536.0,1,-nbitq), 
to_sfixed(558.0/65536.0,1,-nbitq), 
to_sfixed(2617.0/65536.0,1,-nbitq), 
to_sfixed(273.0/65536.0,1,-nbitq), 
to_sfixed(1886.0/65536.0,1,-nbitq), 
to_sfixed(500.0/65536.0,1,-nbitq), 
to_sfixed(1313.0/65536.0,1,-nbitq), 
to_sfixed(-1263.0/65536.0,1,-nbitq), 
to_sfixed(-234.0/65536.0,1,-nbitq), 
to_sfixed(-3607.0/65536.0,1,-nbitq), 
to_sfixed(-3035.0/65536.0,1,-nbitq), 
to_sfixed(2141.0/65536.0,1,-nbitq), 
to_sfixed(1042.0/65536.0,1,-nbitq), 
to_sfixed(-1057.0/65536.0,1,-nbitq), 
to_sfixed(-3074.0/65536.0,1,-nbitq), 
to_sfixed(-33.0/65536.0,1,-nbitq), 
to_sfixed(-1977.0/65536.0,1,-nbitq), 
to_sfixed(-2876.0/65536.0,1,-nbitq), 
to_sfixed(356.0/65536.0,1,-nbitq), 
to_sfixed(-3001.0/65536.0,1,-nbitq), 
to_sfixed(-3012.0/65536.0,1,-nbitq), 
to_sfixed(-1581.0/65536.0,1,-nbitq), 
to_sfixed(-1963.0/65536.0,1,-nbitq), 
to_sfixed(825.0/65536.0,1,-nbitq), 
to_sfixed(-3739.0/65536.0,1,-nbitq), 
to_sfixed(-2972.0/65536.0,1,-nbitq), 
to_sfixed(2036.0/65536.0,1,-nbitq), 
to_sfixed(3053.0/65536.0,1,-nbitq), 
to_sfixed(-2320.0/65536.0,1,-nbitq), 
to_sfixed(-341.0/65536.0,1,-nbitq), 
to_sfixed(426.0/65536.0,1,-nbitq), 
to_sfixed(51.0/65536.0,1,-nbitq), 
to_sfixed(2359.0/65536.0,1,-nbitq), 
to_sfixed(3363.0/65536.0,1,-nbitq), 
to_sfixed(1387.0/65536.0,1,-nbitq), 
to_sfixed(-4809.0/65536.0,1,-nbitq), 
to_sfixed(-178.0/65536.0,1,-nbitq), 
to_sfixed(4176.0/65536.0,1,-nbitq), 
to_sfixed(1449.0/65536.0,1,-nbitq), 
to_sfixed(-283.0/65536.0,1,-nbitq), 
to_sfixed(1962.0/65536.0,1,-nbitq), 
to_sfixed(-4866.0/65536.0,1,-nbitq), 
to_sfixed(1887.0/65536.0,1,-nbitq), 
to_sfixed(2852.0/65536.0,1,-nbitq), 
to_sfixed(2188.0/65536.0,1,-nbitq), 
to_sfixed(-722.0/65536.0,1,-nbitq), 
to_sfixed(916.0/65536.0,1,-nbitq), 
to_sfixed(2902.0/65536.0,1,-nbitq), 
to_sfixed(1673.0/65536.0,1,-nbitq), 
to_sfixed(-2670.0/65536.0,1,-nbitq), 
to_sfixed(-1325.0/65536.0,1,-nbitq), 
to_sfixed(1451.0/65536.0,1,-nbitq), 
to_sfixed(-1076.0/65536.0,1,-nbitq), 
to_sfixed(1139.0/65536.0,1,-nbitq), 
to_sfixed(2103.0/65536.0,1,-nbitq), 
to_sfixed(58.0/65536.0,1,-nbitq), 
to_sfixed(-1270.0/65536.0,1,-nbitq), 
to_sfixed(-1529.0/65536.0,1,-nbitq), 
to_sfixed(-352.0/65536.0,1,-nbitq), 
to_sfixed(643.0/65536.0,1,-nbitq), 
to_sfixed(1390.0/65536.0,1,-nbitq), 
to_sfixed(-2407.0/65536.0,1,-nbitq), 
to_sfixed(2204.0/65536.0,1,-nbitq), 
to_sfixed(695.0/65536.0,1,-nbitq), 
to_sfixed(-3662.0/65536.0,1,-nbitq), 
to_sfixed(2498.0/65536.0,1,-nbitq), 
to_sfixed(2429.0/65536.0,1,-nbitq), 
to_sfixed(4369.0/65536.0,1,-nbitq)  ), 
( to_sfixed(842.0/65536.0,1,-nbitq), 
to_sfixed(-393.0/65536.0,1,-nbitq), 
to_sfixed(-993.0/65536.0,1,-nbitq), 
to_sfixed(-67.0/65536.0,1,-nbitq), 
to_sfixed(-1335.0/65536.0,1,-nbitq), 
to_sfixed(-1890.0/65536.0,1,-nbitq), 
to_sfixed(1104.0/65536.0,1,-nbitq), 
to_sfixed(3554.0/65536.0,1,-nbitq), 
to_sfixed(1727.0/65536.0,1,-nbitq), 
to_sfixed(2604.0/65536.0,1,-nbitq), 
to_sfixed(-3301.0/65536.0,1,-nbitq), 
to_sfixed(-1324.0/65536.0,1,-nbitq), 
to_sfixed(588.0/65536.0,1,-nbitq), 
to_sfixed(1559.0/65536.0,1,-nbitq), 
to_sfixed(2128.0/65536.0,1,-nbitq), 
to_sfixed(-585.0/65536.0,1,-nbitq), 
to_sfixed(1308.0/65536.0,1,-nbitq), 
to_sfixed(2986.0/65536.0,1,-nbitq), 
to_sfixed(1831.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(1536.0/65536.0,1,-nbitq), 
to_sfixed(-3922.0/65536.0,1,-nbitq), 
to_sfixed(63.0/65536.0,1,-nbitq), 
to_sfixed(-1402.0/65536.0,1,-nbitq), 
to_sfixed(-511.0/65536.0,1,-nbitq), 
to_sfixed(3368.0/65536.0,1,-nbitq), 
to_sfixed(-3753.0/65536.0,1,-nbitq), 
to_sfixed(2355.0/65536.0,1,-nbitq), 
to_sfixed(-1109.0/65536.0,1,-nbitq), 
to_sfixed(-1688.0/65536.0,1,-nbitq), 
to_sfixed(1373.0/65536.0,1,-nbitq), 
to_sfixed(-878.0/65536.0,1,-nbitq), 
to_sfixed(-1445.0/65536.0,1,-nbitq), 
to_sfixed(-4932.0/65536.0,1,-nbitq), 
to_sfixed(1172.0/65536.0,1,-nbitq), 
to_sfixed(479.0/65536.0,1,-nbitq), 
to_sfixed(590.0/65536.0,1,-nbitq), 
to_sfixed(2424.0/65536.0,1,-nbitq), 
to_sfixed(-2411.0/65536.0,1,-nbitq), 
to_sfixed(-1377.0/65536.0,1,-nbitq), 
to_sfixed(2311.0/65536.0,1,-nbitq), 
to_sfixed(1562.0/65536.0,1,-nbitq), 
to_sfixed(-2025.0/65536.0,1,-nbitq), 
to_sfixed(340.0/65536.0,1,-nbitq), 
to_sfixed(743.0/65536.0,1,-nbitq), 
to_sfixed(-420.0/65536.0,1,-nbitq), 
to_sfixed(1437.0/65536.0,1,-nbitq), 
to_sfixed(-1928.0/65536.0,1,-nbitq), 
to_sfixed(-578.0/65536.0,1,-nbitq), 
to_sfixed(2751.0/65536.0,1,-nbitq), 
to_sfixed(490.0/65536.0,1,-nbitq), 
to_sfixed(2211.0/65536.0,1,-nbitq), 
to_sfixed(-235.0/65536.0,1,-nbitq), 
to_sfixed(-3081.0/65536.0,1,-nbitq), 
to_sfixed(-1336.0/65536.0,1,-nbitq), 
to_sfixed(1748.0/65536.0,1,-nbitq), 
to_sfixed(1104.0/65536.0,1,-nbitq), 
to_sfixed(3228.0/65536.0,1,-nbitq), 
to_sfixed(-2720.0/65536.0,1,-nbitq), 
to_sfixed(6675.0/65536.0,1,-nbitq), 
to_sfixed(-966.0/65536.0,1,-nbitq), 
to_sfixed(464.0/65536.0,1,-nbitq), 
to_sfixed(-938.0/65536.0,1,-nbitq), 
to_sfixed(-2979.0/65536.0,1,-nbitq), 
to_sfixed(3256.0/65536.0,1,-nbitq), 
to_sfixed(-670.0/65536.0,1,-nbitq), 
to_sfixed(-208.0/65536.0,1,-nbitq), 
to_sfixed(-719.0/65536.0,1,-nbitq), 
to_sfixed(3518.0/65536.0,1,-nbitq), 
to_sfixed(-562.0/65536.0,1,-nbitq), 
to_sfixed(4078.0/65536.0,1,-nbitq), 
to_sfixed(-1352.0/65536.0,1,-nbitq), 
to_sfixed(-79.0/65536.0,1,-nbitq), 
to_sfixed(866.0/65536.0,1,-nbitq), 
to_sfixed(-2789.0/65536.0,1,-nbitq), 
to_sfixed(1227.0/65536.0,1,-nbitq), 
to_sfixed(-1624.0/65536.0,1,-nbitq), 
to_sfixed(3846.0/65536.0,1,-nbitq), 
to_sfixed(-896.0/65536.0,1,-nbitq), 
to_sfixed(1011.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2728.0/65536.0,1,-nbitq), 
to_sfixed(893.0/65536.0,1,-nbitq), 
to_sfixed(489.0/65536.0,1,-nbitq), 
to_sfixed(-2960.0/65536.0,1,-nbitq), 
to_sfixed(1814.0/65536.0,1,-nbitq), 
to_sfixed(-106.0/65536.0,1,-nbitq), 
to_sfixed(-3834.0/65536.0,1,-nbitq), 
to_sfixed(-1548.0/65536.0,1,-nbitq), 
to_sfixed(2885.0/65536.0,1,-nbitq), 
to_sfixed(80.0/65536.0,1,-nbitq), 
to_sfixed(-3910.0/65536.0,1,-nbitq), 
to_sfixed(-4057.0/65536.0,1,-nbitq), 
to_sfixed(-2276.0/65536.0,1,-nbitq), 
to_sfixed(1394.0/65536.0,1,-nbitq), 
to_sfixed(980.0/65536.0,1,-nbitq), 
to_sfixed(585.0/65536.0,1,-nbitq), 
to_sfixed(-191.0/65536.0,1,-nbitq), 
to_sfixed(-1435.0/65536.0,1,-nbitq), 
to_sfixed(3668.0/65536.0,1,-nbitq), 
to_sfixed(-813.0/65536.0,1,-nbitq), 
to_sfixed(-2410.0/65536.0,1,-nbitq), 
to_sfixed(258.0/65536.0,1,-nbitq), 
to_sfixed(-267.0/65536.0,1,-nbitq), 
to_sfixed(121.0/65536.0,1,-nbitq), 
to_sfixed(1023.0/65536.0,1,-nbitq), 
to_sfixed(4186.0/65536.0,1,-nbitq), 
to_sfixed(-1019.0/65536.0,1,-nbitq), 
to_sfixed(-866.0/65536.0,1,-nbitq), 
to_sfixed(-3677.0/65536.0,1,-nbitq), 
to_sfixed(-1253.0/65536.0,1,-nbitq), 
to_sfixed(-868.0/65536.0,1,-nbitq), 
to_sfixed(3107.0/65536.0,1,-nbitq), 
to_sfixed(-2263.0/65536.0,1,-nbitq), 
to_sfixed(-4126.0/65536.0,1,-nbitq), 
to_sfixed(155.0/65536.0,1,-nbitq), 
to_sfixed(-2886.0/65536.0,1,-nbitq), 
to_sfixed(1467.0/65536.0,1,-nbitq), 
to_sfixed(-1146.0/65536.0,1,-nbitq), 
to_sfixed(-1816.0/65536.0,1,-nbitq), 
to_sfixed(516.0/65536.0,1,-nbitq), 
to_sfixed(732.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(-4285.0/65536.0,1,-nbitq), 
to_sfixed(2810.0/65536.0,1,-nbitq), 
to_sfixed(-2353.0/65536.0,1,-nbitq), 
to_sfixed(3684.0/65536.0,1,-nbitq), 
to_sfixed(-1402.0/65536.0,1,-nbitq), 
to_sfixed(2208.0/65536.0,1,-nbitq), 
to_sfixed(1972.0/65536.0,1,-nbitq), 
to_sfixed(3836.0/65536.0,1,-nbitq), 
to_sfixed(483.0/65536.0,1,-nbitq), 
to_sfixed(-1208.0/65536.0,1,-nbitq), 
to_sfixed(18.0/65536.0,1,-nbitq), 
to_sfixed(-2241.0/65536.0,1,-nbitq), 
to_sfixed(3993.0/65536.0,1,-nbitq), 
to_sfixed(-804.0/65536.0,1,-nbitq), 
to_sfixed(1527.0/65536.0,1,-nbitq), 
to_sfixed(-2092.0/65536.0,1,-nbitq), 
to_sfixed(391.0/65536.0,1,-nbitq), 
to_sfixed(4020.0/65536.0,1,-nbitq), 
to_sfixed(485.0/65536.0,1,-nbitq), 
to_sfixed(-1606.0/65536.0,1,-nbitq), 
to_sfixed(-2281.0/65536.0,1,-nbitq), 
to_sfixed(-694.0/65536.0,1,-nbitq), 
to_sfixed(1911.0/65536.0,1,-nbitq), 
to_sfixed(-989.0/65536.0,1,-nbitq), 
to_sfixed(287.0/65536.0,1,-nbitq), 
to_sfixed(-473.0/65536.0,1,-nbitq), 
to_sfixed(2637.0/65536.0,1,-nbitq), 
to_sfixed(-1508.0/65536.0,1,-nbitq), 
to_sfixed(734.0/65536.0,1,-nbitq), 
to_sfixed(1772.0/65536.0,1,-nbitq), 
to_sfixed(1839.0/65536.0,1,-nbitq), 
to_sfixed(-1840.0/65536.0,1,-nbitq), 
to_sfixed(1377.0/65536.0,1,-nbitq), 
to_sfixed(-1092.0/65536.0,1,-nbitq), 
to_sfixed(-2461.0/65536.0,1,-nbitq), 
to_sfixed(-707.0/65536.0,1,-nbitq), 
to_sfixed(-933.0/65536.0,1,-nbitq), 
to_sfixed(1784.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1451.0/65536.0,1,-nbitq), 
to_sfixed(-1887.0/65536.0,1,-nbitq), 
to_sfixed(82.0/65536.0,1,-nbitq), 
to_sfixed(1914.0/65536.0,1,-nbitq), 
to_sfixed(2511.0/65536.0,1,-nbitq), 
to_sfixed(-1406.0/65536.0,1,-nbitq), 
to_sfixed(-1092.0/65536.0,1,-nbitq), 
to_sfixed(529.0/65536.0,1,-nbitq), 
to_sfixed(151.0/65536.0,1,-nbitq), 
to_sfixed(-1255.0/65536.0,1,-nbitq), 
to_sfixed(1901.0/65536.0,1,-nbitq), 
to_sfixed(-3042.0/65536.0,1,-nbitq), 
to_sfixed(1928.0/65536.0,1,-nbitq), 
to_sfixed(-3450.0/65536.0,1,-nbitq), 
to_sfixed(314.0/65536.0,1,-nbitq), 
to_sfixed(1911.0/65536.0,1,-nbitq), 
to_sfixed(765.0/65536.0,1,-nbitq), 
to_sfixed(-803.0/65536.0,1,-nbitq), 
to_sfixed(4008.0/65536.0,1,-nbitq), 
to_sfixed(728.0/65536.0,1,-nbitq), 
to_sfixed(-2691.0/65536.0,1,-nbitq), 
to_sfixed(284.0/65536.0,1,-nbitq), 
to_sfixed(2339.0/65536.0,1,-nbitq), 
to_sfixed(3826.0/65536.0,1,-nbitq), 
to_sfixed(-163.0/65536.0,1,-nbitq), 
to_sfixed(1303.0/65536.0,1,-nbitq), 
to_sfixed(-2414.0/65536.0,1,-nbitq), 
to_sfixed(-2027.0/65536.0,1,-nbitq), 
to_sfixed(-259.0/65536.0,1,-nbitq), 
to_sfixed(-2702.0/65536.0,1,-nbitq), 
to_sfixed(399.0/65536.0,1,-nbitq), 
to_sfixed(37.0/65536.0,1,-nbitq), 
to_sfixed(-558.0/65536.0,1,-nbitq), 
to_sfixed(-5316.0/65536.0,1,-nbitq), 
to_sfixed(2128.0/65536.0,1,-nbitq), 
to_sfixed(-1535.0/65536.0,1,-nbitq), 
to_sfixed(-2206.0/65536.0,1,-nbitq), 
to_sfixed(-1168.0/65536.0,1,-nbitq), 
to_sfixed(-1030.0/65536.0,1,-nbitq), 
to_sfixed(-1748.0/65536.0,1,-nbitq), 
to_sfixed(-2390.0/65536.0,1,-nbitq), 
to_sfixed(2605.0/65536.0,1,-nbitq), 
to_sfixed(-1397.0/65536.0,1,-nbitq), 
to_sfixed(1769.0/65536.0,1,-nbitq), 
to_sfixed(3158.0/65536.0,1,-nbitq), 
to_sfixed(4673.0/65536.0,1,-nbitq), 
to_sfixed(-440.0/65536.0,1,-nbitq), 
to_sfixed(-3247.0/65536.0,1,-nbitq), 
to_sfixed(1753.0/65536.0,1,-nbitq), 
to_sfixed(3334.0/65536.0,1,-nbitq), 
to_sfixed(-1857.0/65536.0,1,-nbitq), 
to_sfixed(-2465.0/65536.0,1,-nbitq), 
to_sfixed(1924.0/65536.0,1,-nbitq), 
to_sfixed(-2675.0/65536.0,1,-nbitq), 
to_sfixed(1197.0/65536.0,1,-nbitq), 
to_sfixed(-2668.0/65536.0,1,-nbitq), 
to_sfixed(1146.0/65536.0,1,-nbitq), 
to_sfixed(3104.0/65536.0,1,-nbitq), 
to_sfixed(2082.0/65536.0,1,-nbitq), 
to_sfixed(2210.0/65536.0,1,-nbitq), 
to_sfixed(-1879.0/65536.0,1,-nbitq), 
to_sfixed(-1721.0/65536.0,1,-nbitq), 
to_sfixed(534.0/65536.0,1,-nbitq), 
to_sfixed(288.0/65536.0,1,-nbitq), 
to_sfixed(-250.0/65536.0,1,-nbitq), 
to_sfixed(2885.0/65536.0,1,-nbitq), 
to_sfixed(2182.0/65536.0,1,-nbitq), 
to_sfixed(460.0/65536.0,1,-nbitq), 
to_sfixed(-232.0/65536.0,1,-nbitq), 
to_sfixed(-2677.0/65536.0,1,-nbitq), 
to_sfixed(2605.0/65536.0,1,-nbitq), 
to_sfixed(2373.0/65536.0,1,-nbitq), 
to_sfixed(-1491.0/65536.0,1,-nbitq), 
to_sfixed(-2604.0/65536.0,1,-nbitq), 
to_sfixed(2303.0/65536.0,1,-nbitq), 
to_sfixed(638.0/65536.0,1,-nbitq), 
to_sfixed(1759.0/65536.0,1,-nbitq), 
to_sfixed(4198.0/65536.0,1,-nbitq), 
to_sfixed(-2069.0/65536.0,1,-nbitq), 
to_sfixed(409.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3175.0/65536.0,1,-nbitq), 
to_sfixed(421.0/65536.0,1,-nbitq), 
to_sfixed(2978.0/65536.0,1,-nbitq), 
to_sfixed(-607.0/65536.0,1,-nbitq), 
to_sfixed(-4373.0/65536.0,1,-nbitq), 
to_sfixed(1991.0/65536.0,1,-nbitq), 
to_sfixed(-534.0/65536.0,1,-nbitq), 
to_sfixed(-517.0/65536.0,1,-nbitq), 
to_sfixed(-2328.0/65536.0,1,-nbitq), 
to_sfixed(843.0/65536.0,1,-nbitq), 
to_sfixed(-562.0/65536.0,1,-nbitq), 
to_sfixed(585.0/65536.0,1,-nbitq), 
to_sfixed(-2375.0/65536.0,1,-nbitq), 
to_sfixed(-1510.0/65536.0,1,-nbitq), 
to_sfixed(-1705.0/65536.0,1,-nbitq), 
to_sfixed(2355.0/65536.0,1,-nbitq), 
to_sfixed(-1125.0/65536.0,1,-nbitq), 
to_sfixed(-133.0/65536.0,1,-nbitq), 
to_sfixed(-1719.0/65536.0,1,-nbitq), 
to_sfixed(2309.0/65536.0,1,-nbitq), 
to_sfixed(-1359.0/65536.0,1,-nbitq), 
to_sfixed(38.0/65536.0,1,-nbitq), 
to_sfixed(2173.0/65536.0,1,-nbitq), 
to_sfixed(2954.0/65536.0,1,-nbitq), 
to_sfixed(942.0/65536.0,1,-nbitq), 
to_sfixed(-901.0/65536.0,1,-nbitq), 
to_sfixed(-1261.0/65536.0,1,-nbitq), 
to_sfixed(2876.0/65536.0,1,-nbitq), 
to_sfixed(-913.0/65536.0,1,-nbitq), 
to_sfixed(942.0/65536.0,1,-nbitq), 
to_sfixed(3666.0/65536.0,1,-nbitq), 
to_sfixed(2463.0/65536.0,1,-nbitq), 
to_sfixed(-4282.0/65536.0,1,-nbitq), 
to_sfixed(-5376.0/65536.0,1,-nbitq), 
to_sfixed(-308.0/65536.0,1,-nbitq), 
to_sfixed(-3117.0/65536.0,1,-nbitq), 
to_sfixed(-790.0/65536.0,1,-nbitq), 
to_sfixed(2063.0/65536.0,1,-nbitq), 
to_sfixed(-3024.0/65536.0,1,-nbitq), 
to_sfixed(-598.0/65536.0,1,-nbitq), 
to_sfixed(-924.0/65536.0,1,-nbitq), 
to_sfixed(1726.0/65536.0,1,-nbitq), 
to_sfixed(-82.0/65536.0,1,-nbitq), 
to_sfixed(1145.0/65536.0,1,-nbitq), 
to_sfixed(-359.0/65536.0,1,-nbitq), 
to_sfixed(4345.0/65536.0,1,-nbitq), 
to_sfixed(1731.0/65536.0,1,-nbitq), 
to_sfixed(1264.0/65536.0,1,-nbitq), 
to_sfixed(3038.0/65536.0,1,-nbitq), 
to_sfixed(1759.0/65536.0,1,-nbitq), 
to_sfixed(2134.0/65536.0,1,-nbitq), 
to_sfixed(65.0/65536.0,1,-nbitq), 
to_sfixed(3725.0/65536.0,1,-nbitq), 
to_sfixed(-2061.0/65536.0,1,-nbitq), 
to_sfixed(2599.0/65536.0,1,-nbitq), 
to_sfixed(2939.0/65536.0,1,-nbitq), 
to_sfixed(281.0/65536.0,1,-nbitq), 
to_sfixed(-170.0/65536.0,1,-nbitq), 
to_sfixed(-1949.0/65536.0,1,-nbitq), 
to_sfixed(1783.0/65536.0,1,-nbitq), 
to_sfixed(-3261.0/65536.0,1,-nbitq), 
to_sfixed(-935.0/65536.0,1,-nbitq), 
to_sfixed(-857.0/65536.0,1,-nbitq), 
to_sfixed(-1348.0/65536.0,1,-nbitq), 
to_sfixed(2787.0/65536.0,1,-nbitq), 
to_sfixed(1279.0/65536.0,1,-nbitq), 
to_sfixed(712.0/65536.0,1,-nbitq), 
to_sfixed(401.0/65536.0,1,-nbitq), 
to_sfixed(-1495.0/65536.0,1,-nbitq), 
to_sfixed(775.0/65536.0,1,-nbitq), 
to_sfixed(-686.0/65536.0,1,-nbitq), 
to_sfixed(-148.0/65536.0,1,-nbitq), 
to_sfixed(1698.0/65536.0,1,-nbitq), 
to_sfixed(1861.0/65536.0,1,-nbitq), 
to_sfixed(-1983.0/65536.0,1,-nbitq), 
to_sfixed(1286.0/65536.0,1,-nbitq), 
to_sfixed(2206.0/65536.0,1,-nbitq), 
to_sfixed(711.0/65536.0,1,-nbitq), 
to_sfixed(-1390.0/65536.0,1,-nbitq), 
to_sfixed(1417.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1604.0/65536.0,1,-nbitq), 
to_sfixed(-222.0/65536.0,1,-nbitq), 
to_sfixed(-2.0/65536.0,1,-nbitq), 
to_sfixed(-378.0/65536.0,1,-nbitq), 
to_sfixed(-2521.0/65536.0,1,-nbitq), 
to_sfixed(-1519.0/65536.0,1,-nbitq), 
to_sfixed(-3359.0/65536.0,1,-nbitq), 
to_sfixed(1617.0/65536.0,1,-nbitq), 
to_sfixed(-428.0/65536.0,1,-nbitq), 
to_sfixed(-598.0/65536.0,1,-nbitq), 
to_sfixed(-3604.0/65536.0,1,-nbitq), 
to_sfixed(-1959.0/65536.0,1,-nbitq), 
to_sfixed(-1894.0/65536.0,1,-nbitq), 
to_sfixed(-2398.0/65536.0,1,-nbitq), 
to_sfixed(2128.0/65536.0,1,-nbitq), 
to_sfixed(-456.0/65536.0,1,-nbitq), 
to_sfixed(-2876.0/65536.0,1,-nbitq), 
to_sfixed(450.0/65536.0,1,-nbitq), 
to_sfixed(2988.0/65536.0,1,-nbitq), 
to_sfixed(-1540.0/65536.0,1,-nbitq), 
to_sfixed(1096.0/65536.0,1,-nbitq), 
to_sfixed(-1133.0/65536.0,1,-nbitq), 
to_sfixed(-883.0/65536.0,1,-nbitq), 
to_sfixed(-130.0/65536.0,1,-nbitq), 
to_sfixed(1531.0/65536.0,1,-nbitq), 
to_sfixed(-1652.0/65536.0,1,-nbitq), 
to_sfixed(951.0/65536.0,1,-nbitq), 
to_sfixed(-1938.0/65536.0,1,-nbitq), 
to_sfixed(-2725.0/65536.0,1,-nbitq), 
to_sfixed(203.0/65536.0,1,-nbitq), 
to_sfixed(-1151.0/65536.0,1,-nbitq), 
to_sfixed(322.0/65536.0,1,-nbitq), 
to_sfixed(-1327.0/65536.0,1,-nbitq), 
to_sfixed(-266.0/65536.0,1,-nbitq), 
to_sfixed(1400.0/65536.0,1,-nbitq), 
to_sfixed(1216.0/65536.0,1,-nbitq), 
to_sfixed(-1115.0/65536.0,1,-nbitq), 
to_sfixed(-2138.0/65536.0,1,-nbitq), 
to_sfixed(-1177.0/65536.0,1,-nbitq), 
to_sfixed(-1618.0/65536.0,1,-nbitq), 
to_sfixed(1659.0/65536.0,1,-nbitq), 
to_sfixed(704.0/65536.0,1,-nbitq), 
to_sfixed(-305.0/65536.0,1,-nbitq), 
to_sfixed(2849.0/65536.0,1,-nbitq), 
to_sfixed(172.0/65536.0,1,-nbitq), 
to_sfixed(673.0/65536.0,1,-nbitq), 
to_sfixed(1238.0/65536.0,1,-nbitq), 
to_sfixed(2874.0/65536.0,1,-nbitq), 
to_sfixed(1989.0/65536.0,1,-nbitq), 
to_sfixed(3740.0/65536.0,1,-nbitq), 
to_sfixed(1627.0/65536.0,1,-nbitq), 
to_sfixed(947.0/65536.0,1,-nbitq), 
to_sfixed(3244.0/65536.0,1,-nbitq), 
to_sfixed(-1357.0/65536.0,1,-nbitq), 
to_sfixed(3207.0/65536.0,1,-nbitq), 
to_sfixed(-2406.0/65536.0,1,-nbitq), 
to_sfixed(2952.0/65536.0,1,-nbitq), 
to_sfixed(-2260.0/65536.0,1,-nbitq), 
to_sfixed(121.0/65536.0,1,-nbitq), 
to_sfixed(1997.0/65536.0,1,-nbitq), 
to_sfixed(-2966.0/65536.0,1,-nbitq), 
to_sfixed(1109.0/65536.0,1,-nbitq), 
to_sfixed(858.0/65536.0,1,-nbitq), 
to_sfixed(1332.0/65536.0,1,-nbitq), 
to_sfixed(1673.0/65536.0,1,-nbitq), 
to_sfixed(2916.0/65536.0,1,-nbitq), 
to_sfixed(1322.0/65536.0,1,-nbitq), 
to_sfixed(1280.0/65536.0,1,-nbitq), 
to_sfixed(3581.0/65536.0,1,-nbitq), 
to_sfixed(-235.0/65536.0,1,-nbitq), 
to_sfixed(1402.0/65536.0,1,-nbitq), 
to_sfixed(836.0/65536.0,1,-nbitq), 
to_sfixed(3367.0/65536.0,1,-nbitq), 
to_sfixed(-1359.0/65536.0,1,-nbitq), 
to_sfixed(2669.0/65536.0,1,-nbitq), 
to_sfixed(-1583.0/65536.0,1,-nbitq), 
to_sfixed(-2876.0/65536.0,1,-nbitq), 
to_sfixed(4207.0/65536.0,1,-nbitq), 
to_sfixed(1817.0/65536.0,1,-nbitq), 
to_sfixed(4103.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2121.0/65536.0,1,-nbitq), 
to_sfixed(1540.0/65536.0,1,-nbitq), 
to_sfixed(1867.0/65536.0,1,-nbitq), 
to_sfixed(-674.0/65536.0,1,-nbitq), 
to_sfixed(-1300.0/65536.0,1,-nbitq), 
to_sfixed(1094.0/65536.0,1,-nbitq), 
to_sfixed(-2999.0/65536.0,1,-nbitq), 
to_sfixed(1093.0/65536.0,1,-nbitq), 
to_sfixed(-2160.0/65536.0,1,-nbitq), 
to_sfixed(-491.0/65536.0,1,-nbitq), 
to_sfixed(-2396.0/65536.0,1,-nbitq), 
to_sfixed(1003.0/65536.0,1,-nbitq), 
to_sfixed(2791.0/65536.0,1,-nbitq), 
to_sfixed(5.0/65536.0,1,-nbitq), 
to_sfixed(1354.0/65536.0,1,-nbitq), 
to_sfixed(2847.0/65536.0,1,-nbitq), 
to_sfixed(1046.0/65536.0,1,-nbitq), 
to_sfixed(1581.0/65536.0,1,-nbitq), 
to_sfixed(574.0/65536.0,1,-nbitq), 
to_sfixed(1290.0/65536.0,1,-nbitq), 
to_sfixed(-2113.0/65536.0,1,-nbitq), 
to_sfixed(-457.0/65536.0,1,-nbitq), 
to_sfixed(-511.0/65536.0,1,-nbitq), 
to_sfixed(1300.0/65536.0,1,-nbitq), 
to_sfixed(-69.0/65536.0,1,-nbitq), 
to_sfixed(3425.0/65536.0,1,-nbitq), 
to_sfixed(-3283.0/65536.0,1,-nbitq), 
to_sfixed(-831.0/65536.0,1,-nbitq), 
to_sfixed(-404.0/65536.0,1,-nbitq), 
to_sfixed(-886.0/65536.0,1,-nbitq), 
to_sfixed(-698.0/65536.0,1,-nbitq), 
to_sfixed(887.0/65536.0,1,-nbitq), 
to_sfixed(-673.0/65536.0,1,-nbitq), 
to_sfixed(-5406.0/65536.0,1,-nbitq), 
to_sfixed(-335.0/65536.0,1,-nbitq), 
to_sfixed(-2683.0/65536.0,1,-nbitq), 
to_sfixed(-20.0/65536.0,1,-nbitq), 
to_sfixed(-834.0/65536.0,1,-nbitq), 
to_sfixed(333.0/65536.0,1,-nbitq), 
to_sfixed(-1507.0/65536.0,1,-nbitq), 
to_sfixed(-185.0/65536.0,1,-nbitq), 
to_sfixed(-536.0/65536.0,1,-nbitq), 
to_sfixed(-185.0/65536.0,1,-nbitq), 
to_sfixed(1882.0/65536.0,1,-nbitq), 
to_sfixed(-521.0/65536.0,1,-nbitq), 
to_sfixed(1892.0/65536.0,1,-nbitq), 
to_sfixed(-1361.0/65536.0,1,-nbitq), 
to_sfixed(3135.0/65536.0,1,-nbitq), 
to_sfixed(-624.0/65536.0,1,-nbitq), 
to_sfixed(-332.0/65536.0,1,-nbitq), 
to_sfixed(-416.0/65536.0,1,-nbitq), 
to_sfixed(1846.0/65536.0,1,-nbitq), 
to_sfixed(1872.0/65536.0,1,-nbitq), 
to_sfixed(-58.0/65536.0,1,-nbitq), 
to_sfixed(-2177.0/65536.0,1,-nbitq), 
to_sfixed(-457.0/65536.0,1,-nbitq), 
to_sfixed(2546.0/65536.0,1,-nbitq), 
to_sfixed(-798.0/65536.0,1,-nbitq), 
to_sfixed(425.0/65536.0,1,-nbitq), 
to_sfixed(1526.0/65536.0,1,-nbitq), 
to_sfixed(-2664.0/65536.0,1,-nbitq), 
to_sfixed(-857.0/65536.0,1,-nbitq), 
to_sfixed(2084.0/65536.0,1,-nbitq), 
to_sfixed(2525.0/65536.0,1,-nbitq), 
to_sfixed(3594.0/65536.0,1,-nbitq), 
to_sfixed(-1679.0/65536.0,1,-nbitq), 
to_sfixed(74.0/65536.0,1,-nbitq), 
to_sfixed(-3040.0/65536.0,1,-nbitq), 
to_sfixed(766.0/65536.0,1,-nbitq), 
to_sfixed(2461.0/65536.0,1,-nbitq), 
to_sfixed(-311.0/65536.0,1,-nbitq), 
to_sfixed(1882.0/65536.0,1,-nbitq), 
to_sfixed(3460.0/65536.0,1,-nbitq), 
to_sfixed(-2285.0/65536.0,1,-nbitq), 
to_sfixed(2232.0/65536.0,1,-nbitq), 
to_sfixed(-2183.0/65536.0,1,-nbitq), 
to_sfixed(1071.0/65536.0,1,-nbitq), 
to_sfixed(4219.0/65536.0,1,-nbitq), 
to_sfixed(1128.0/65536.0,1,-nbitq), 
to_sfixed(42.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-789.0/65536.0,1,-nbitq), 
to_sfixed(368.0/65536.0,1,-nbitq), 
to_sfixed(1788.0/65536.0,1,-nbitq), 
to_sfixed(1525.0/65536.0,1,-nbitq), 
to_sfixed(-446.0/65536.0,1,-nbitq), 
to_sfixed(89.0/65536.0,1,-nbitq), 
to_sfixed(376.0/65536.0,1,-nbitq), 
to_sfixed(2338.0/65536.0,1,-nbitq), 
to_sfixed(-4326.0/65536.0,1,-nbitq), 
to_sfixed(350.0/65536.0,1,-nbitq), 
to_sfixed(-2308.0/65536.0,1,-nbitq), 
to_sfixed(-1236.0/65536.0,1,-nbitq), 
to_sfixed(951.0/65536.0,1,-nbitq), 
to_sfixed(-3301.0/65536.0,1,-nbitq), 
to_sfixed(1103.0/65536.0,1,-nbitq), 
to_sfixed(-865.0/65536.0,1,-nbitq), 
to_sfixed(2217.0/65536.0,1,-nbitq), 
to_sfixed(-1922.0/65536.0,1,-nbitq), 
to_sfixed(-1265.0/65536.0,1,-nbitq), 
to_sfixed(3252.0/65536.0,1,-nbitq), 
to_sfixed(-3093.0/65536.0,1,-nbitq), 
to_sfixed(-1484.0/65536.0,1,-nbitq), 
to_sfixed(-2207.0/65536.0,1,-nbitq), 
to_sfixed(-1991.0/65536.0,1,-nbitq), 
to_sfixed(-305.0/65536.0,1,-nbitq), 
to_sfixed(1798.0/65536.0,1,-nbitq), 
to_sfixed(820.0/65536.0,1,-nbitq), 
to_sfixed(1102.0/65536.0,1,-nbitq), 
to_sfixed(500.0/65536.0,1,-nbitq), 
to_sfixed(-962.0/65536.0,1,-nbitq), 
to_sfixed(1209.0/65536.0,1,-nbitq), 
to_sfixed(2708.0/65536.0,1,-nbitq), 
to_sfixed(-2736.0/65536.0,1,-nbitq), 
to_sfixed(-3761.0/65536.0,1,-nbitq), 
to_sfixed(1759.0/65536.0,1,-nbitq), 
to_sfixed(-1746.0/65536.0,1,-nbitq), 
to_sfixed(-2152.0/65536.0,1,-nbitq), 
to_sfixed(-1719.0/65536.0,1,-nbitq), 
to_sfixed(-646.0/65536.0,1,-nbitq), 
to_sfixed(838.0/65536.0,1,-nbitq), 
to_sfixed(-3063.0/65536.0,1,-nbitq), 
to_sfixed(-2581.0/65536.0,1,-nbitq), 
to_sfixed(-3423.0/65536.0,1,-nbitq), 
to_sfixed(2300.0/65536.0,1,-nbitq), 
to_sfixed(-178.0/65536.0,1,-nbitq), 
to_sfixed(4818.0/65536.0,1,-nbitq), 
to_sfixed(2690.0/65536.0,1,-nbitq), 
to_sfixed(-440.0/65536.0,1,-nbitq), 
to_sfixed(-2074.0/65536.0,1,-nbitq), 
to_sfixed(2113.0/65536.0,1,-nbitq), 
to_sfixed(1871.0/65536.0,1,-nbitq), 
to_sfixed(-555.0/65536.0,1,-nbitq), 
to_sfixed(349.0/65536.0,1,-nbitq), 
to_sfixed(-2472.0/65536.0,1,-nbitq), 
to_sfixed(3811.0/65536.0,1,-nbitq), 
to_sfixed(141.0/65536.0,1,-nbitq), 
to_sfixed(390.0/65536.0,1,-nbitq), 
to_sfixed(-1388.0/65536.0,1,-nbitq), 
to_sfixed(-2723.0/65536.0,1,-nbitq), 
to_sfixed(99.0/65536.0,1,-nbitq), 
to_sfixed(774.0/65536.0,1,-nbitq), 
to_sfixed(1382.0/65536.0,1,-nbitq), 
to_sfixed(-1675.0/65536.0,1,-nbitq), 
to_sfixed(2002.0/65536.0,1,-nbitq), 
to_sfixed(2463.0/65536.0,1,-nbitq), 
to_sfixed(1778.0/65536.0,1,-nbitq), 
to_sfixed(3357.0/65536.0,1,-nbitq), 
to_sfixed(-4758.0/65536.0,1,-nbitq), 
to_sfixed(1068.0/65536.0,1,-nbitq), 
to_sfixed(204.0/65536.0,1,-nbitq), 
to_sfixed(768.0/65536.0,1,-nbitq), 
to_sfixed(-2119.0/65536.0,1,-nbitq), 
to_sfixed(2329.0/65536.0,1,-nbitq), 
to_sfixed(-2967.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(2416.0/65536.0,1,-nbitq), 
to_sfixed(-1819.0/65536.0,1,-nbitq), 
to_sfixed(3269.0/65536.0,1,-nbitq), 
to_sfixed(-1904.0/65536.0,1,-nbitq), 
to_sfixed(3462.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1188.0/65536.0,1,-nbitq), 
to_sfixed(-2088.0/65536.0,1,-nbitq), 
to_sfixed(861.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(-3073.0/65536.0,1,-nbitq), 
to_sfixed(-997.0/65536.0,1,-nbitq), 
to_sfixed(327.0/65536.0,1,-nbitq), 
to_sfixed(-918.0/65536.0,1,-nbitq), 
to_sfixed(-3422.0/65536.0,1,-nbitq), 
to_sfixed(2220.0/65536.0,1,-nbitq), 
to_sfixed(1139.0/65536.0,1,-nbitq), 
to_sfixed(-2483.0/65536.0,1,-nbitq), 
to_sfixed(542.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(3242.0/65536.0,1,-nbitq), 
to_sfixed(2757.0/65536.0,1,-nbitq), 
to_sfixed(-844.0/65536.0,1,-nbitq), 
to_sfixed(-1749.0/65536.0,1,-nbitq), 
to_sfixed(2982.0/65536.0,1,-nbitq), 
to_sfixed(-1861.0/65536.0,1,-nbitq), 
to_sfixed(-3058.0/65536.0,1,-nbitq), 
to_sfixed(-276.0/65536.0,1,-nbitq), 
to_sfixed(1944.0/65536.0,1,-nbitq), 
to_sfixed(956.0/65536.0,1,-nbitq), 
to_sfixed(491.0/65536.0,1,-nbitq), 
to_sfixed(3357.0/65536.0,1,-nbitq), 
to_sfixed(-724.0/65536.0,1,-nbitq), 
to_sfixed(-3494.0/65536.0,1,-nbitq), 
to_sfixed(1082.0/65536.0,1,-nbitq), 
to_sfixed(-172.0/65536.0,1,-nbitq), 
to_sfixed(-166.0/65536.0,1,-nbitq), 
to_sfixed(-1530.0/65536.0,1,-nbitq), 
to_sfixed(-4195.0/65536.0,1,-nbitq), 
to_sfixed(-2732.0/65536.0,1,-nbitq), 
to_sfixed(-1644.0/65536.0,1,-nbitq), 
to_sfixed(-2845.0/65536.0,1,-nbitq), 
to_sfixed(-2552.0/65536.0,1,-nbitq), 
to_sfixed(-2958.0/65536.0,1,-nbitq), 
to_sfixed(-3191.0/65536.0,1,-nbitq), 
to_sfixed(778.0/65536.0,1,-nbitq), 
to_sfixed(1216.0/65536.0,1,-nbitq), 
to_sfixed(1599.0/65536.0,1,-nbitq), 
to_sfixed(-291.0/65536.0,1,-nbitq), 
to_sfixed(2133.0/65536.0,1,-nbitq), 
to_sfixed(2507.0/65536.0,1,-nbitq), 
to_sfixed(4532.0/65536.0,1,-nbitq), 
to_sfixed(-1697.0/65536.0,1,-nbitq), 
to_sfixed(3229.0/65536.0,1,-nbitq), 
to_sfixed(-1828.0/65536.0,1,-nbitq), 
to_sfixed(2586.0/65536.0,1,-nbitq), 
to_sfixed(-1282.0/65536.0,1,-nbitq), 
to_sfixed(-1023.0/65536.0,1,-nbitq), 
to_sfixed(-565.0/65536.0,1,-nbitq), 
to_sfixed(-2614.0/65536.0,1,-nbitq), 
to_sfixed(1205.0/65536.0,1,-nbitq), 
to_sfixed(2896.0/65536.0,1,-nbitq), 
to_sfixed(-476.0/65536.0,1,-nbitq), 
to_sfixed(884.0/65536.0,1,-nbitq), 
to_sfixed(384.0/65536.0,1,-nbitq), 
to_sfixed(3983.0/65536.0,1,-nbitq), 
to_sfixed(-1707.0/65536.0,1,-nbitq), 
to_sfixed(1893.0/65536.0,1,-nbitq), 
to_sfixed(2710.0/65536.0,1,-nbitq), 
to_sfixed(1125.0/65536.0,1,-nbitq), 
to_sfixed(79.0/65536.0,1,-nbitq), 
to_sfixed(2634.0/65536.0,1,-nbitq), 
to_sfixed(-1569.0/65536.0,1,-nbitq), 
to_sfixed(-1953.0/65536.0,1,-nbitq), 
to_sfixed(2180.0/65536.0,1,-nbitq), 
to_sfixed(1479.0/65536.0,1,-nbitq), 
to_sfixed(-439.0/65536.0,1,-nbitq), 
to_sfixed(1701.0/65536.0,1,-nbitq), 
to_sfixed(3729.0/65536.0,1,-nbitq), 
to_sfixed(-2946.0/65536.0,1,-nbitq), 
to_sfixed(-2438.0/65536.0,1,-nbitq), 
to_sfixed(3345.0/65536.0,1,-nbitq), 
to_sfixed(-2222.0/65536.0,1,-nbitq), 
to_sfixed(2030.0/65536.0,1,-nbitq), 
to_sfixed(2581.0/65536.0,1,-nbitq), 
to_sfixed(4115.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2490.0/65536.0,1,-nbitq), 
to_sfixed(-1232.0/65536.0,1,-nbitq), 
to_sfixed(-812.0/65536.0,1,-nbitq), 
to_sfixed(-1317.0/65536.0,1,-nbitq), 
to_sfixed(-1699.0/65536.0,1,-nbitq), 
to_sfixed(-1329.0/65536.0,1,-nbitq), 
to_sfixed(3016.0/65536.0,1,-nbitq), 
to_sfixed(-449.0/65536.0,1,-nbitq), 
to_sfixed(-2335.0/65536.0,1,-nbitq), 
to_sfixed(3024.0/65536.0,1,-nbitq), 
to_sfixed(-2429.0/65536.0,1,-nbitq), 
to_sfixed(-167.0/65536.0,1,-nbitq), 
to_sfixed(2595.0/65536.0,1,-nbitq), 
to_sfixed(-663.0/65536.0,1,-nbitq), 
to_sfixed(-803.0/65536.0,1,-nbitq), 
to_sfixed(386.0/65536.0,1,-nbitq), 
to_sfixed(-3207.0/65536.0,1,-nbitq), 
to_sfixed(2452.0/65536.0,1,-nbitq), 
to_sfixed(558.0/65536.0,1,-nbitq), 
to_sfixed(-729.0/65536.0,1,-nbitq), 
to_sfixed(1733.0/65536.0,1,-nbitq), 
to_sfixed(375.0/65536.0,1,-nbitq), 
to_sfixed(-1420.0/65536.0,1,-nbitq), 
to_sfixed(-2030.0/65536.0,1,-nbitq), 
to_sfixed(504.0/65536.0,1,-nbitq), 
to_sfixed(-1385.0/65536.0,1,-nbitq), 
to_sfixed(-3751.0/65536.0,1,-nbitq), 
to_sfixed(-237.0/65536.0,1,-nbitq), 
to_sfixed(-2079.0/65536.0,1,-nbitq), 
to_sfixed(-1624.0/65536.0,1,-nbitq), 
to_sfixed(1310.0/65536.0,1,-nbitq), 
to_sfixed(2100.0/65536.0,1,-nbitq), 
to_sfixed(-3655.0/65536.0,1,-nbitq), 
to_sfixed(77.0/65536.0,1,-nbitq), 
to_sfixed(2758.0/65536.0,1,-nbitq), 
to_sfixed(-1922.0/65536.0,1,-nbitq), 
to_sfixed(1133.0/65536.0,1,-nbitq), 
to_sfixed(-806.0/65536.0,1,-nbitq), 
to_sfixed(1239.0/65536.0,1,-nbitq), 
to_sfixed(753.0/65536.0,1,-nbitq), 
to_sfixed(563.0/65536.0,1,-nbitq), 
to_sfixed(1191.0/65536.0,1,-nbitq), 
to_sfixed(-2788.0/65536.0,1,-nbitq), 
to_sfixed(-616.0/65536.0,1,-nbitq), 
to_sfixed(-2423.0/65536.0,1,-nbitq), 
to_sfixed(2682.0/65536.0,1,-nbitq), 
to_sfixed(947.0/65536.0,1,-nbitq), 
to_sfixed(-1289.0/65536.0,1,-nbitq), 
to_sfixed(693.0/65536.0,1,-nbitq), 
to_sfixed(152.0/65536.0,1,-nbitq), 
to_sfixed(-794.0/65536.0,1,-nbitq), 
to_sfixed(1483.0/65536.0,1,-nbitq), 
to_sfixed(2770.0/65536.0,1,-nbitq), 
to_sfixed(1333.0/65536.0,1,-nbitq), 
to_sfixed(-590.0/65536.0,1,-nbitq), 
to_sfixed(-347.0/65536.0,1,-nbitq), 
to_sfixed(2461.0/65536.0,1,-nbitq), 
to_sfixed(-1176.0/65536.0,1,-nbitq), 
to_sfixed(2576.0/65536.0,1,-nbitq), 
to_sfixed(3423.0/65536.0,1,-nbitq), 
to_sfixed(-3080.0/65536.0,1,-nbitq), 
to_sfixed(1699.0/65536.0,1,-nbitq), 
to_sfixed(1108.0/65536.0,1,-nbitq), 
to_sfixed(-117.0/65536.0,1,-nbitq), 
to_sfixed(-88.0/65536.0,1,-nbitq), 
to_sfixed(-2166.0/65536.0,1,-nbitq), 
to_sfixed(-1037.0/65536.0,1,-nbitq), 
to_sfixed(-2863.0/65536.0,1,-nbitq), 
to_sfixed(2403.0/65536.0,1,-nbitq), 
to_sfixed(3164.0/65536.0,1,-nbitq), 
to_sfixed(-1501.0/65536.0,1,-nbitq), 
to_sfixed(1853.0/65536.0,1,-nbitq), 
to_sfixed(3722.0/65536.0,1,-nbitq), 
to_sfixed(-469.0/65536.0,1,-nbitq), 
to_sfixed(-2317.0/65536.0,1,-nbitq), 
to_sfixed(3022.0/65536.0,1,-nbitq), 
to_sfixed(-2010.0/65536.0,1,-nbitq), 
to_sfixed(255.0/65536.0,1,-nbitq), 
to_sfixed(2078.0/65536.0,1,-nbitq), 
to_sfixed(3421.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2925.0/65536.0,1,-nbitq), 
to_sfixed(3111.0/65536.0,1,-nbitq), 
to_sfixed(-996.0/65536.0,1,-nbitq), 
to_sfixed(-3395.0/65536.0,1,-nbitq), 
to_sfixed(223.0/65536.0,1,-nbitq), 
to_sfixed(-730.0/65536.0,1,-nbitq), 
to_sfixed(-774.0/65536.0,1,-nbitq), 
to_sfixed(-440.0/65536.0,1,-nbitq), 
to_sfixed(-41.0/65536.0,1,-nbitq), 
to_sfixed(-2557.0/65536.0,1,-nbitq), 
to_sfixed(385.0/65536.0,1,-nbitq), 
to_sfixed(-482.0/65536.0,1,-nbitq), 
to_sfixed(-373.0/65536.0,1,-nbitq), 
to_sfixed(-1755.0/65536.0,1,-nbitq), 
to_sfixed(-570.0/65536.0,1,-nbitq), 
to_sfixed(-1814.0/65536.0,1,-nbitq), 
to_sfixed(-731.0/65536.0,1,-nbitq), 
to_sfixed(2281.0/65536.0,1,-nbitq), 
to_sfixed(-982.0/65536.0,1,-nbitq), 
to_sfixed(-392.0/65536.0,1,-nbitq), 
to_sfixed(-1770.0/65536.0,1,-nbitq), 
to_sfixed(-1963.0/65536.0,1,-nbitq), 
to_sfixed(-246.0/65536.0,1,-nbitq), 
to_sfixed(2340.0/65536.0,1,-nbitq), 
to_sfixed(2690.0/65536.0,1,-nbitq), 
to_sfixed(1759.0/65536.0,1,-nbitq), 
to_sfixed(-1869.0/65536.0,1,-nbitq), 
to_sfixed(-2417.0/65536.0,1,-nbitq), 
to_sfixed(-7.0/65536.0,1,-nbitq), 
to_sfixed(1262.0/65536.0,1,-nbitq), 
to_sfixed(2536.0/65536.0,1,-nbitq), 
to_sfixed(-2582.0/65536.0,1,-nbitq), 
to_sfixed(-2760.0/65536.0,1,-nbitq), 
to_sfixed(-4813.0/65536.0,1,-nbitq), 
to_sfixed(-1401.0/65536.0,1,-nbitq), 
to_sfixed(2050.0/65536.0,1,-nbitq), 
to_sfixed(-2415.0/65536.0,1,-nbitq), 
to_sfixed(-3732.0/65536.0,1,-nbitq), 
to_sfixed(-758.0/65536.0,1,-nbitq), 
to_sfixed(-1181.0/65536.0,1,-nbitq), 
to_sfixed(-910.0/65536.0,1,-nbitq), 
to_sfixed(1476.0/65536.0,1,-nbitq), 
to_sfixed(228.0/65536.0,1,-nbitq), 
to_sfixed(2576.0/65536.0,1,-nbitq), 
to_sfixed(-149.0/65536.0,1,-nbitq), 
to_sfixed(3665.0/65536.0,1,-nbitq), 
to_sfixed(-1565.0/65536.0,1,-nbitq), 
to_sfixed(22.0/65536.0,1,-nbitq), 
to_sfixed(1617.0/65536.0,1,-nbitq), 
to_sfixed(1811.0/65536.0,1,-nbitq), 
to_sfixed(-505.0/65536.0,1,-nbitq), 
to_sfixed(-157.0/65536.0,1,-nbitq), 
to_sfixed(-1141.0/65536.0,1,-nbitq), 
to_sfixed(787.0/65536.0,1,-nbitq), 
to_sfixed(1075.0/65536.0,1,-nbitq), 
to_sfixed(-569.0/65536.0,1,-nbitq), 
to_sfixed(1786.0/65536.0,1,-nbitq), 
to_sfixed(-1483.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(4870.0/65536.0,1,-nbitq), 
to_sfixed(1196.0/65536.0,1,-nbitq), 
to_sfixed(-1001.0/65536.0,1,-nbitq), 
to_sfixed(-544.0/65536.0,1,-nbitq), 
to_sfixed(1787.0/65536.0,1,-nbitq), 
to_sfixed(1420.0/65536.0,1,-nbitq), 
to_sfixed(2.0/65536.0,1,-nbitq), 
to_sfixed(1581.0/65536.0,1,-nbitq), 
to_sfixed(368.0/65536.0,1,-nbitq), 
to_sfixed(2432.0/65536.0,1,-nbitq), 
to_sfixed(1090.0/65536.0,1,-nbitq), 
to_sfixed(755.0/65536.0,1,-nbitq), 
to_sfixed(2514.0/65536.0,1,-nbitq), 
to_sfixed(3551.0/65536.0,1,-nbitq), 
to_sfixed(-2269.0/65536.0,1,-nbitq), 
to_sfixed(-2216.0/65536.0,1,-nbitq), 
to_sfixed(-499.0/65536.0,1,-nbitq), 
to_sfixed(-1131.0/65536.0,1,-nbitq), 
to_sfixed(446.0/65536.0,1,-nbitq), 
to_sfixed(2709.0/65536.0,1,-nbitq), 
to_sfixed(4047.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2452.0/65536.0,1,-nbitq), 
to_sfixed(2864.0/65536.0,1,-nbitq), 
to_sfixed(4315.0/65536.0,1,-nbitq), 
to_sfixed(1923.0/65536.0,1,-nbitq), 
to_sfixed(-2715.0/65536.0,1,-nbitq), 
to_sfixed(-1731.0/65536.0,1,-nbitq), 
to_sfixed(-2442.0/65536.0,1,-nbitq), 
to_sfixed(-474.0/65536.0,1,-nbitq), 
to_sfixed(-1128.0/65536.0,1,-nbitq), 
to_sfixed(-1899.0/65536.0,1,-nbitq), 
to_sfixed(-990.0/65536.0,1,-nbitq), 
to_sfixed(-2277.0/65536.0,1,-nbitq), 
to_sfixed(-1913.0/65536.0,1,-nbitq), 
to_sfixed(-1916.0/65536.0,1,-nbitq), 
to_sfixed(-2613.0/65536.0,1,-nbitq), 
to_sfixed(-910.0/65536.0,1,-nbitq), 
to_sfixed(95.0/65536.0,1,-nbitq), 
to_sfixed(-1571.0/65536.0,1,-nbitq), 
to_sfixed(1347.0/65536.0,1,-nbitq), 
to_sfixed(-397.0/65536.0,1,-nbitq), 
to_sfixed(-2988.0/65536.0,1,-nbitq), 
to_sfixed(3055.0/65536.0,1,-nbitq), 
to_sfixed(518.0/65536.0,1,-nbitq), 
to_sfixed(1115.0/65536.0,1,-nbitq), 
to_sfixed(1341.0/65536.0,1,-nbitq), 
to_sfixed(1581.0/65536.0,1,-nbitq), 
to_sfixed(803.0/65536.0,1,-nbitq), 
to_sfixed(-1555.0/65536.0,1,-nbitq), 
to_sfixed(-4305.0/65536.0,1,-nbitq), 
to_sfixed(-1650.0/65536.0,1,-nbitq), 
to_sfixed(2002.0/65536.0,1,-nbitq), 
to_sfixed(-1998.0/65536.0,1,-nbitq), 
to_sfixed(-3912.0/65536.0,1,-nbitq), 
to_sfixed(432.0/65536.0,1,-nbitq), 
to_sfixed(2252.0/65536.0,1,-nbitq), 
to_sfixed(-1811.0/65536.0,1,-nbitq), 
to_sfixed(2528.0/65536.0,1,-nbitq), 
to_sfixed(-4110.0/65536.0,1,-nbitq), 
to_sfixed(-1230.0/65536.0,1,-nbitq), 
to_sfixed(-1041.0/65536.0,1,-nbitq), 
to_sfixed(-139.0/65536.0,1,-nbitq), 
to_sfixed(-2662.0/65536.0,1,-nbitq), 
to_sfixed(-2343.0/65536.0,1,-nbitq), 
to_sfixed(2854.0/65536.0,1,-nbitq), 
to_sfixed(3265.0/65536.0,1,-nbitq), 
to_sfixed(1082.0/65536.0,1,-nbitq), 
to_sfixed(-666.0/65536.0,1,-nbitq), 
to_sfixed(-2481.0/65536.0,1,-nbitq), 
to_sfixed(-689.0/65536.0,1,-nbitq), 
to_sfixed(-764.0/65536.0,1,-nbitq), 
to_sfixed(-2417.0/65536.0,1,-nbitq), 
to_sfixed(287.0/65536.0,1,-nbitq), 
to_sfixed(-153.0/65536.0,1,-nbitq), 
to_sfixed(351.0/65536.0,1,-nbitq), 
to_sfixed(1359.0/65536.0,1,-nbitq), 
to_sfixed(2718.0/65536.0,1,-nbitq), 
to_sfixed(2970.0/65536.0,1,-nbitq), 
to_sfixed(559.0/65536.0,1,-nbitq), 
to_sfixed(-2600.0/65536.0,1,-nbitq), 
to_sfixed(5500.0/65536.0,1,-nbitq), 
to_sfixed(-253.0/65536.0,1,-nbitq), 
to_sfixed(2005.0/65536.0,1,-nbitq), 
to_sfixed(-291.0/65536.0,1,-nbitq), 
to_sfixed(240.0/65536.0,1,-nbitq), 
to_sfixed(-502.0/65536.0,1,-nbitq), 
to_sfixed(2053.0/65536.0,1,-nbitq), 
to_sfixed(1357.0/65536.0,1,-nbitq), 
to_sfixed(-4841.0/65536.0,1,-nbitq), 
to_sfixed(2886.0/65536.0,1,-nbitq), 
to_sfixed(-824.0/65536.0,1,-nbitq), 
to_sfixed(-2167.0/65536.0,1,-nbitq), 
to_sfixed(-564.0/65536.0,1,-nbitq), 
to_sfixed(-292.0/65536.0,1,-nbitq), 
to_sfixed(-1922.0/65536.0,1,-nbitq), 
to_sfixed(915.0/65536.0,1,-nbitq), 
to_sfixed(1893.0/65536.0,1,-nbitq), 
to_sfixed(-2358.0/65536.0,1,-nbitq), 
to_sfixed(2677.0/65536.0,1,-nbitq), 
to_sfixed(586.0/65536.0,1,-nbitq), 
to_sfixed(5926.0/65536.0,1,-nbitq)  ), 
( to_sfixed(351.0/65536.0,1,-nbitq), 
to_sfixed(1840.0/65536.0,1,-nbitq), 
to_sfixed(4643.0/65536.0,1,-nbitq), 
to_sfixed(-532.0/65536.0,1,-nbitq), 
to_sfixed(-4352.0/65536.0,1,-nbitq), 
to_sfixed(582.0/65536.0,1,-nbitq), 
to_sfixed(-1202.0/65536.0,1,-nbitq), 
to_sfixed(-83.0/65536.0,1,-nbitq), 
to_sfixed(928.0/65536.0,1,-nbitq), 
to_sfixed(1066.0/65536.0,1,-nbitq), 
to_sfixed(-2671.0/65536.0,1,-nbitq), 
to_sfixed(-5788.0/65536.0,1,-nbitq), 
to_sfixed(-1431.0/65536.0,1,-nbitq), 
to_sfixed(-1462.0/65536.0,1,-nbitq), 
to_sfixed(335.0/65536.0,1,-nbitq), 
to_sfixed(-23.0/65536.0,1,-nbitq), 
to_sfixed(-540.0/65536.0,1,-nbitq), 
to_sfixed(354.0/65536.0,1,-nbitq), 
to_sfixed(1544.0/65536.0,1,-nbitq), 
to_sfixed(1384.0/65536.0,1,-nbitq), 
to_sfixed(-2614.0/65536.0,1,-nbitq), 
to_sfixed(698.0/65536.0,1,-nbitq), 
to_sfixed(106.0/65536.0,1,-nbitq), 
to_sfixed(-1578.0/65536.0,1,-nbitq), 
to_sfixed(175.0/65536.0,1,-nbitq), 
to_sfixed(-1436.0/65536.0,1,-nbitq), 
to_sfixed(172.0/65536.0,1,-nbitq), 
to_sfixed(-2853.0/65536.0,1,-nbitq), 
to_sfixed(-1819.0/65536.0,1,-nbitq), 
to_sfixed(-954.0/65536.0,1,-nbitq), 
to_sfixed(1486.0/65536.0,1,-nbitq), 
to_sfixed(2647.0/65536.0,1,-nbitq), 
to_sfixed(-2446.0/65536.0,1,-nbitq), 
to_sfixed(1052.0/65536.0,1,-nbitq), 
to_sfixed(-1025.0/65536.0,1,-nbitq), 
to_sfixed(2003.0/65536.0,1,-nbitq), 
to_sfixed(-2612.0/65536.0,1,-nbitq), 
to_sfixed(-1694.0/65536.0,1,-nbitq), 
to_sfixed(-2929.0/65536.0,1,-nbitq), 
to_sfixed(1185.0/65536.0,1,-nbitq), 
to_sfixed(-1006.0/65536.0,1,-nbitq), 
to_sfixed(-2339.0/65536.0,1,-nbitq), 
to_sfixed(-3613.0/65536.0,1,-nbitq), 
to_sfixed(3605.0/65536.0,1,-nbitq), 
to_sfixed(-1378.0/65536.0,1,-nbitq), 
to_sfixed(1369.0/65536.0,1,-nbitq), 
to_sfixed(1739.0/65536.0,1,-nbitq), 
to_sfixed(-1509.0/65536.0,1,-nbitq), 
to_sfixed(2952.0/65536.0,1,-nbitq), 
to_sfixed(-1458.0/65536.0,1,-nbitq), 
to_sfixed(39.0/65536.0,1,-nbitq), 
to_sfixed(735.0/65536.0,1,-nbitq), 
to_sfixed(2179.0/65536.0,1,-nbitq), 
to_sfixed(-167.0/65536.0,1,-nbitq), 
to_sfixed(-1172.0/65536.0,1,-nbitq), 
to_sfixed(-1048.0/65536.0,1,-nbitq), 
to_sfixed(-2803.0/65536.0,1,-nbitq), 
to_sfixed(2727.0/65536.0,1,-nbitq), 
to_sfixed(1362.0/65536.0,1,-nbitq), 
to_sfixed(3928.0/65536.0,1,-nbitq), 
to_sfixed(-2793.0/65536.0,1,-nbitq), 
to_sfixed(-1120.0/65536.0,1,-nbitq), 
to_sfixed(-1919.0/65536.0,1,-nbitq), 
to_sfixed(-433.0/65536.0,1,-nbitq), 
to_sfixed(4412.0/65536.0,1,-nbitq), 
to_sfixed(160.0/65536.0,1,-nbitq), 
to_sfixed(1920.0/65536.0,1,-nbitq), 
to_sfixed(-1880.0/65536.0,1,-nbitq), 
to_sfixed(2573.0/65536.0,1,-nbitq), 
to_sfixed(968.0/65536.0,1,-nbitq), 
to_sfixed(1010.0/65536.0,1,-nbitq), 
to_sfixed(-609.0/65536.0,1,-nbitq), 
to_sfixed(1441.0/65536.0,1,-nbitq), 
to_sfixed(-2295.0/65536.0,1,-nbitq), 
to_sfixed(2131.0/65536.0,1,-nbitq), 
to_sfixed(-2930.0/65536.0,1,-nbitq), 
to_sfixed(-3867.0/65536.0,1,-nbitq), 
to_sfixed(2668.0/65536.0,1,-nbitq), 
to_sfixed(-359.0/65536.0,1,-nbitq), 
to_sfixed(4899.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-213.0/65536.0,1,-nbitq), 
to_sfixed(687.0/65536.0,1,-nbitq), 
to_sfixed(1448.0/65536.0,1,-nbitq), 
to_sfixed(-2383.0/65536.0,1,-nbitq), 
to_sfixed(-2052.0/65536.0,1,-nbitq), 
to_sfixed(-1079.0/65536.0,1,-nbitq), 
to_sfixed(-2216.0/65536.0,1,-nbitq), 
to_sfixed(-2327.0/65536.0,1,-nbitq), 
to_sfixed(-1330.0/65536.0,1,-nbitq), 
to_sfixed(-2067.0/65536.0,1,-nbitq), 
to_sfixed(-2235.0/65536.0,1,-nbitq), 
to_sfixed(-160.0/65536.0,1,-nbitq), 
to_sfixed(-2865.0/65536.0,1,-nbitq), 
to_sfixed(-760.0/65536.0,1,-nbitq), 
to_sfixed(-3529.0/65536.0,1,-nbitq), 
to_sfixed(3039.0/65536.0,1,-nbitq), 
to_sfixed(-1341.0/65536.0,1,-nbitq), 
to_sfixed(-443.0/65536.0,1,-nbitq), 
to_sfixed(1675.0/65536.0,1,-nbitq), 
to_sfixed(2840.0/65536.0,1,-nbitq), 
to_sfixed(-1713.0/65536.0,1,-nbitq), 
to_sfixed(2749.0/65536.0,1,-nbitq), 
to_sfixed(2690.0/65536.0,1,-nbitq), 
to_sfixed(533.0/65536.0,1,-nbitq), 
to_sfixed(-2191.0/65536.0,1,-nbitq), 
to_sfixed(-3347.0/65536.0,1,-nbitq), 
to_sfixed(27.0/65536.0,1,-nbitq), 
to_sfixed(-4933.0/65536.0,1,-nbitq), 
to_sfixed(-5300.0/65536.0,1,-nbitq), 
to_sfixed(-894.0/65536.0,1,-nbitq), 
to_sfixed(1743.0/65536.0,1,-nbitq), 
to_sfixed(2915.0/65536.0,1,-nbitq), 
to_sfixed(-3085.0/65536.0,1,-nbitq), 
to_sfixed(868.0/65536.0,1,-nbitq), 
to_sfixed(2730.0/65536.0,1,-nbitq), 
to_sfixed(2164.0/65536.0,1,-nbitq), 
to_sfixed(1951.0/65536.0,1,-nbitq), 
to_sfixed(946.0/65536.0,1,-nbitq), 
to_sfixed(2816.0/65536.0,1,-nbitq), 
to_sfixed(-3430.0/65536.0,1,-nbitq), 
to_sfixed(398.0/65536.0,1,-nbitq), 
to_sfixed(-2318.0/65536.0,1,-nbitq), 
to_sfixed(1390.0/65536.0,1,-nbitq), 
to_sfixed(4542.0/65536.0,1,-nbitq), 
to_sfixed(-1628.0/65536.0,1,-nbitq), 
to_sfixed(4269.0/65536.0,1,-nbitq), 
to_sfixed(-826.0/65536.0,1,-nbitq), 
to_sfixed(-2526.0/65536.0,1,-nbitq), 
to_sfixed(-900.0/65536.0,1,-nbitq), 
to_sfixed(3563.0/65536.0,1,-nbitq), 
to_sfixed(1847.0/65536.0,1,-nbitq), 
to_sfixed(-612.0/65536.0,1,-nbitq), 
to_sfixed(2545.0/65536.0,1,-nbitq), 
to_sfixed(1472.0/65536.0,1,-nbitq), 
to_sfixed(-928.0/65536.0,1,-nbitq), 
to_sfixed(-2979.0/65536.0,1,-nbitq), 
to_sfixed(1026.0/65536.0,1,-nbitq), 
to_sfixed(1720.0/65536.0,1,-nbitq), 
to_sfixed(1863.0/65536.0,1,-nbitq), 
to_sfixed(808.0/65536.0,1,-nbitq), 
to_sfixed(-3292.0/65536.0,1,-nbitq), 
to_sfixed(-2675.0/65536.0,1,-nbitq), 
to_sfixed(-600.0/65536.0,1,-nbitq), 
to_sfixed(1593.0/65536.0,1,-nbitq), 
to_sfixed(301.0/65536.0,1,-nbitq), 
to_sfixed(965.0/65536.0,1,-nbitq), 
to_sfixed(2069.0/65536.0,1,-nbitq), 
to_sfixed(-5045.0/65536.0,1,-nbitq), 
to_sfixed(2270.0/65536.0,1,-nbitq), 
to_sfixed(780.0/65536.0,1,-nbitq), 
to_sfixed(-138.0/65536.0,1,-nbitq), 
to_sfixed(1310.0/65536.0,1,-nbitq), 
to_sfixed(-1703.0/65536.0,1,-nbitq), 
to_sfixed(1246.0/65536.0,1,-nbitq), 
to_sfixed(2279.0/65536.0,1,-nbitq), 
to_sfixed(2157.0/65536.0,1,-nbitq), 
to_sfixed(-5779.0/65536.0,1,-nbitq), 
to_sfixed(-302.0/65536.0,1,-nbitq), 
to_sfixed(-95.0/65536.0,1,-nbitq), 
to_sfixed(1949.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-379.0/65536.0,1,-nbitq), 
to_sfixed(7198.0/65536.0,1,-nbitq), 
to_sfixed(-1630.0/65536.0,1,-nbitq), 
to_sfixed(3625.0/65536.0,1,-nbitq), 
to_sfixed(-2984.0/65536.0,1,-nbitq), 
to_sfixed(-4276.0/65536.0,1,-nbitq), 
to_sfixed(2835.0/65536.0,1,-nbitq), 
to_sfixed(1146.0/65536.0,1,-nbitq), 
to_sfixed(650.0/65536.0,1,-nbitq), 
to_sfixed(-2623.0/65536.0,1,-nbitq), 
to_sfixed(-3826.0/65536.0,1,-nbitq), 
to_sfixed(-1167.0/65536.0,1,-nbitq), 
to_sfixed(1163.0/65536.0,1,-nbitq), 
to_sfixed(-5738.0/65536.0,1,-nbitq), 
to_sfixed(210.0/65536.0,1,-nbitq), 
to_sfixed(1327.0/65536.0,1,-nbitq), 
to_sfixed(-2481.0/65536.0,1,-nbitq), 
to_sfixed(-689.0/65536.0,1,-nbitq), 
to_sfixed(308.0/65536.0,1,-nbitq), 
to_sfixed(-1737.0/65536.0,1,-nbitq), 
to_sfixed(3642.0/65536.0,1,-nbitq), 
to_sfixed(7109.0/65536.0,1,-nbitq), 
to_sfixed(-628.0/65536.0,1,-nbitq), 
to_sfixed(-4445.0/65536.0,1,-nbitq), 
to_sfixed(-1956.0/65536.0,1,-nbitq), 
to_sfixed(-2600.0/65536.0,1,-nbitq), 
to_sfixed(-3466.0/65536.0,1,-nbitq), 
to_sfixed(-4841.0/65536.0,1,-nbitq), 
to_sfixed(932.0/65536.0,1,-nbitq), 
to_sfixed(1303.0/65536.0,1,-nbitq), 
to_sfixed(-2375.0/65536.0,1,-nbitq), 
to_sfixed(814.0/65536.0,1,-nbitq), 
to_sfixed(-1026.0/65536.0,1,-nbitq), 
to_sfixed(720.0/65536.0,1,-nbitq), 
to_sfixed(-2551.0/65536.0,1,-nbitq), 
to_sfixed(-217.0/65536.0,1,-nbitq), 
to_sfixed(-1635.0/65536.0,1,-nbitq), 
to_sfixed(1634.0/65536.0,1,-nbitq), 
to_sfixed(3697.0/65536.0,1,-nbitq), 
to_sfixed(1724.0/65536.0,1,-nbitq), 
to_sfixed(1087.0/65536.0,1,-nbitq), 
to_sfixed(192.0/65536.0,1,-nbitq), 
to_sfixed(597.0/65536.0,1,-nbitq), 
to_sfixed(576.0/65536.0,1,-nbitq), 
to_sfixed(-2600.0/65536.0,1,-nbitq), 
to_sfixed(3069.0/65536.0,1,-nbitq), 
to_sfixed(2571.0/65536.0,1,-nbitq), 
to_sfixed(-5645.0/65536.0,1,-nbitq), 
to_sfixed(2332.0/65536.0,1,-nbitq), 
to_sfixed(3419.0/65536.0,1,-nbitq), 
to_sfixed(3359.0/65536.0,1,-nbitq), 
to_sfixed(-1688.0/65536.0,1,-nbitq), 
to_sfixed(2646.0/65536.0,1,-nbitq), 
to_sfixed(1753.0/65536.0,1,-nbitq), 
to_sfixed(-919.0/65536.0,1,-nbitq), 
to_sfixed(-4805.0/65536.0,1,-nbitq), 
to_sfixed(1738.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(-2565.0/65536.0,1,-nbitq), 
to_sfixed(-492.0/65536.0,1,-nbitq), 
to_sfixed(-2681.0/65536.0,1,-nbitq), 
to_sfixed(2214.0/65536.0,1,-nbitq), 
to_sfixed(-827.0/65536.0,1,-nbitq), 
to_sfixed(1761.0/65536.0,1,-nbitq), 
to_sfixed(-1409.0/65536.0,1,-nbitq), 
to_sfixed(1233.0/65536.0,1,-nbitq), 
to_sfixed(-262.0/65536.0,1,-nbitq), 
to_sfixed(-223.0/65536.0,1,-nbitq), 
to_sfixed(-1938.0/65536.0,1,-nbitq), 
to_sfixed(204.0/65536.0,1,-nbitq), 
to_sfixed(-38.0/65536.0,1,-nbitq), 
to_sfixed(-2382.0/65536.0,1,-nbitq), 
to_sfixed(-1765.0/65536.0,1,-nbitq), 
to_sfixed(1426.0/65536.0,1,-nbitq), 
to_sfixed(-2406.0/65536.0,1,-nbitq), 
to_sfixed(73.0/65536.0,1,-nbitq), 
to_sfixed(-7773.0/65536.0,1,-nbitq), 
to_sfixed(-1049.0/65536.0,1,-nbitq), 
to_sfixed(-319.0/65536.0,1,-nbitq), 
to_sfixed(4242.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1184.0/65536.0,1,-nbitq), 
to_sfixed(7204.0/65536.0,1,-nbitq), 
to_sfixed(-2790.0/65536.0,1,-nbitq), 
to_sfixed(-1540.0/65536.0,1,-nbitq), 
to_sfixed(-3138.0/65536.0,1,-nbitq), 
to_sfixed(-2743.0/65536.0,1,-nbitq), 
to_sfixed(-905.0/65536.0,1,-nbitq), 
to_sfixed(135.0/65536.0,1,-nbitq), 
to_sfixed(2341.0/65536.0,1,-nbitq), 
to_sfixed(572.0/65536.0,1,-nbitq), 
to_sfixed(-1841.0/65536.0,1,-nbitq), 
to_sfixed(-1228.0/65536.0,1,-nbitq), 
to_sfixed(73.0/65536.0,1,-nbitq), 
to_sfixed(-6337.0/65536.0,1,-nbitq), 
to_sfixed(-800.0/65536.0,1,-nbitq), 
to_sfixed(316.0/65536.0,1,-nbitq), 
to_sfixed(750.0/65536.0,1,-nbitq), 
to_sfixed(3348.0/65536.0,1,-nbitq), 
to_sfixed(424.0/65536.0,1,-nbitq), 
to_sfixed(-2037.0/65536.0,1,-nbitq), 
to_sfixed(3261.0/65536.0,1,-nbitq), 
to_sfixed(6608.0/65536.0,1,-nbitq), 
to_sfixed(4671.0/65536.0,1,-nbitq), 
to_sfixed(-6173.0/65536.0,1,-nbitq), 
to_sfixed(-394.0/65536.0,1,-nbitq), 
to_sfixed(-2778.0/65536.0,1,-nbitq), 
to_sfixed(1357.0/65536.0,1,-nbitq), 
to_sfixed(-4239.0/65536.0,1,-nbitq), 
to_sfixed(-108.0/65536.0,1,-nbitq), 
to_sfixed(-1402.0/65536.0,1,-nbitq), 
to_sfixed(1380.0/65536.0,1,-nbitq), 
to_sfixed(-2046.0/65536.0,1,-nbitq), 
to_sfixed(1483.0/65536.0,1,-nbitq), 
to_sfixed(-27.0/65536.0,1,-nbitq), 
to_sfixed(334.0/65536.0,1,-nbitq), 
to_sfixed(1569.0/65536.0,1,-nbitq), 
to_sfixed(-796.0/65536.0,1,-nbitq), 
to_sfixed(-1527.0/65536.0,1,-nbitq), 
to_sfixed(5212.0/65536.0,1,-nbitq), 
to_sfixed(-1481.0/65536.0,1,-nbitq), 
to_sfixed(1223.0/65536.0,1,-nbitq), 
to_sfixed(-245.0/65536.0,1,-nbitq), 
to_sfixed(347.0/65536.0,1,-nbitq), 
to_sfixed(947.0/65536.0,1,-nbitq), 
to_sfixed(3161.0/65536.0,1,-nbitq), 
to_sfixed(2101.0/65536.0,1,-nbitq), 
to_sfixed(-1766.0/65536.0,1,-nbitq), 
to_sfixed(-2903.0/65536.0,1,-nbitq), 
to_sfixed(-220.0/65536.0,1,-nbitq), 
to_sfixed(4386.0/65536.0,1,-nbitq), 
to_sfixed(-855.0/65536.0,1,-nbitq), 
to_sfixed(1193.0/65536.0,1,-nbitq), 
to_sfixed(1273.0/65536.0,1,-nbitq), 
to_sfixed(-2160.0/65536.0,1,-nbitq), 
to_sfixed(3405.0/65536.0,1,-nbitq), 
to_sfixed(-7112.0/65536.0,1,-nbitq), 
to_sfixed(-1806.0/65536.0,1,-nbitq), 
to_sfixed(-3108.0/65536.0,1,-nbitq), 
to_sfixed(2519.0/65536.0,1,-nbitq), 
to_sfixed(1994.0/65536.0,1,-nbitq), 
to_sfixed(-2599.0/65536.0,1,-nbitq), 
to_sfixed(-799.0/65536.0,1,-nbitq), 
to_sfixed(-2023.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(1374.0/65536.0,1,-nbitq), 
to_sfixed(-3265.0/65536.0,1,-nbitq), 
to_sfixed(4519.0/65536.0,1,-nbitq), 
to_sfixed(-1082.0/65536.0,1,-nbitq), 
to_sfixed(116.0/65536.0,1,-nbitq), 
to_sfixed(2474.0/65536.0,1,-nbitq), 
to_sfixed(3260.0/65536.0,1,-nbitq), 
to_sfixed(-4139.0/65536.0,1,-nbitq), 
to_sfixed(-3726.0/65536.0,1,-nbitq), 
to_sfixed(-1030.0/65536.0,1,-nbitq), 
to_sfixed(-2299.0/65536.0,1,-nbitq), 
to_sfixed(-2153.0/65536.0,1,-nbitq), 
to_sfixed(-7806.0/65536.0,1,-nbitq), 
to_sfixed(2702.0/65536.0,1,-nbitq), 
to_sfixed(1538.0/65536.0,1,-nbitq), 
to_sfixed(1343.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3833.0/65536.0,1,-nbitq), 
to_sfixed(7625.0/65536.0,1,-nbitq), 
to_sfixed(-4612.0/65536.0,1,-nbitq), 
to_sfixed(451.0/65536.0,1,-nbitq), 
to_sfixed(-2267.0/65536.0,1,-nbitq), 
to_sfixed(-7455.0/65536.0,1,-nbitq), 
to_sfixed(415.0/65536.0,1,-nbitq), 
to_sfixed(-204.0/65536.0,1,-nbitq), 
to_sfixed(366.0/65536.0,1,-nbitq), 
to_sfixed(869.0/65536.0,1,-nbitq), 
to_sfixed(-1857.0/65536.0,1,-nbitq), 
to_sfixed(-832.0/65536.0,1,-nbitq), 
to_sfixed(-1844.0/65536.0,1,-nbitq), 
to_sfixed(-2700.0/65536.0,1,-nbitq), 
to_sfixed(1626.0/65536.0,1,-nbitq), 
to_sfixed(-1846.0/65536.0,1,-nbitq), 
to_sfixed(635.0/65536.0,1,-nbitq), 
to_sfixed(-2557.0/65536.0,1,-nbitq), 
to_sfixed(-2713.0/65536.0,1,-nbitq), 
to_sfixed(2449.0/65536.0,1,-nbitq), 
to_sfixed(2667.0/65536.0,1,-nbitq), 
to_sfixed(2566.0/65536.0,1,-nbitq), 
to_sfixed(1757.0/65536.0,1,-nbitq), 
to_sfixed(-9039.0/65536.0,1,-nbitq), 
to_sfixed(1114.0/65536.0,1,-nbitq), 
to_sfixed(-2071.0/65536.0,1,-nbitq), 
to_sfixed(-1692.0/65536.0,1,-nbitq), 
to_sfixed(-4263.0/65536.0,1,-nbitq), 
to_sfixed(-1987.0/65536.0,1,-nbitq), 
to_sfixed(307.0/65536.0,1,-nbitq), 
to_sfixed(2369.0/65536.0,1,-nbitq), 
to_sfixed(868.0/65536.0,1,-nbitq), 
to_sfixed(4298.0/65536.0,1,-nbitq), 
to_sfixed(4111.0/65536.0,1,-nbitq), 
to_sfixed(-1861.0/65536.0,1,-nbitq), 
to_sfixed(726.0/65536.0,1,-nbitq), 
to_sfixed(-494.0/65536.0,1,-nbitq), 
to_sfixed(-1732.0/65536.0,1,-nbitq), 
to_sfixed(8250.0/65536.0,1,-nbitq), 
to_sfixed(-751.0/65536.0,1,-nbitq), 
to_sfixed(1397.0/65536.0,1,-nbitq), 
to_sfixed(-2973.0/65536.0,1,-nbitq), 
to_sfixed(-918.0/65536.0,1,-nbitq), 
to_sfixed(-1365.0/65536.0,1,-nbitq), 
to_sfixed(-1817.0/65536.0,1,-nbitq), 
to_sfixed(826.0/65536.0,1,-nbitq), 
to_sfixed(-993.0/65536.0,1,-nbitq), 
to_sfixed(-2630.0/65536.0,1,-nbitq), 
to_sfixed(1352.0/65536.0,1,-nbitq), 
to_sfixed(238.0/65536.0,1,-nbitq), 
to_sfixed(-801.0/65536.0,1,-nbitq), 
to_sfixed(-689.0/65536.0,1,-nbitq), 
to_sfixed(4384.0/65536.0,1,-nbitq), 
to_sfixed(-1235.0/65536.0,1,-nbitq), 
to_sfixed(867.0/65536.0,1,-nbitq), 
to_sfixed(-4034.0/65536.0,1,-nbitq), 
to_sfixed(2720.0/65536.0,1,-nbitq), 
to_sfixed(-2242.0/65536.0,1,-nbitq), 
to_sfixed(2454.0/65536.0,1,-nbitq), 
to_sfixed(-2258.0/65536.0,1,-nbitq), 
to_sfixed(-1690.0/65536.0,1,-nbitq), 
to_sfixed(1284.0/65536.0,1,-nbitq), 
to_sfixed(-679.0/65536.0,1,-nbitq), 
to_sfixed(355.0/65536.0,1,-nbitq), 
to_sfixed(-2612.0/65536.0,1,-nbitq), 
to_sfixed(-3207.0/65536.0,1,-nbitq), 
to_sfixed(1602.0/65536.0,1,-nbitq), 
to_sfixed(2496.0/65536.0,1,-nbitq), 
to_sfixed(2715.0/65536.0,1,-nbitq), 
to_sfixed(155.0/65536.0,1,-nbitq), 
to_sfixed(928.0/65536.0,1,-nbitq), 
to_sfixed(-3887.0/65536.0,1,-nbitq), 
to_sfixed(568.0/65536.0,1,-nbitq), 
to_sfixed(-2870.0/65536.0,1,-nbitq), 
to_sfixed(-2706.0/65536.0,1,-nbitq), 
to_sfixed(1040.0/65536.0,1,-nbitq), 
to_sfixed(-3176.0/65536.0,1,-nbitq), 
to_sfixed(3717.0/65536.0,1,-nbitq), 
to_sfixed(-2481.0/65536.0,1,-nbitq), 
to_sfixed(1706.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2964.0/65536.0,1,-nbitq), 
to_sfixed(4129.0/65536.0,1,-nbitq), 
to_sfixed(-1746.0/65536.0,1,-nbitq), 
to_sfixed(-817.0/65536.0,1,-nbitq), 
to_sfixed(-1491.0/65536.0,1,-nbitq), 
to_sfixed(-2425.0/65536.0,1,-nbitq), 
to_sfixed(-1624.0/65536.0,1,-nbitq), 
to_sfixed(963.0/65536.0,1,-nbitq), 
to_sfixed(1857.0/65536.0,1,-nbitq), 
to_sfixed(-458.0/65536.0,1,-nbitq), 
to_sfixed(-3341.0/65536.0,1,-nbitq), 
to_sfixed(-5387.0/65536.0,1,-nbitq), 
to_sfixed(-926.0/65536.0,1,-nbitq), 
to_sfixed(1349.0/65536.0,1,-nbitq), 
to_sfixed(2520.0/65536.0,1,-nbitq), 
to_sfixed(-819.0/65536.0,1,-nbitq), 
to_sfixed(-1413.0/65536.0,1,-nbitq), 
to_sfixed(-952.0/65536.0,1,-nbitq), 
to_sfixed(-656.0/65536.0,1,-nbitq), 
to_sfixed(2889.0/65536.0,1,-nbitq), 
to_sfixed(2044.0/65536.0,1,-nbitq), 
to_sfixed(1381.0/65536.0,1,-nbitq), 
to_sfixed(4725.0/65536.0,1,-nbitq), 
to_sfixed(-8659.0/65536.0,1,-nbitq), 
to_sfixed(-126.0/65536.0,1,-nbitq), 
to_sfixed(-6202.0/65536.0,1,-nbitq), 
to_sfixed(42.0/65536.0,1,-nbitq), 
to_sfixed(-2189.0/65536.0,1,-nbitq), 
to_sfixed(-2935.0/65536.0,1,-nbitq), 
to_sfixed(-3214.0/65536.0,1,-nbitq), 
to_sfixed(4273.0/65536.0,1,-nbitq), 
to_sfixed(491.0/65536.0,1,-nbitq), 
to_sfixed(-1367.0/65536.0,1,-nbitq), 
to_sfixed(-1500.0/65536.0,1,-nbitq), 
to_sfixed(-1316.0/65536.0,1,-nbitq), 
to_sfixed(-2334.0/65536.0,1,-nbitq), 
to_sfixed(-1536.0/65536.0,1,-nbitq), 
to_sfixed(-477.0/65536.0,1,-nbitq), 
to_sfixed(5001.0/65536.0,1,-nbitq), 
to_sfixed(-341.0/65536.0,1,-nbitq), 
to_sfixed(-936.0/65536.0,1,-nbitq), 
to_sfixed(-2538.0/65536.0,1,-nbitq), 
to_sfixed(1961.0/65536.0,1,-nbitq), 
to_sfixed(-22.0/65536.0,1,-nbitq), 
to_sfixed(2383.0/65536.0,1,-nbitq), 
to_sfixed(456.0/65536.0,1,-nbitq), 
to_sfixed(2881.0/65536.0,1,-nbitq), 
to_sfixed(-1151.0/65536.0,1,-nbitq), 
to_sfixed(-1062.0/65536.0,1,-nbitq), 
to_sfixed(1017.0/65536.0,1,-nbitq), 
to_sfixed(1692.0/65536.0,1,-nbitq), 
to_sfixed(840.0/65536.0,1,-nbitq), 
to_sfixed(5402.0/65536.0,1,-nbitq), 
to_sfixed(-2982.0/65536.0,1,-nbitq), 
to_sfixed(-2205.0/65536.0,1,-nbitq), 
to_sfixed(-3580.0/65536.0,1,-nbitq), 
to_sfixed(-1977.0/65536.0,1,-nbitq), 
to_sfixed(-376.0/65536.0,1,-nbitq), 
to_sfixed(124.0/65536.0,1,-nbitq), 
to_sfixed(1595.0/65536.0,1,-nbitq), 
to_sfixed(-2096.0/65536.0,1,-nbitq), 
to_sfixed(-3208.0/65536.0,1,-nbitq), 
to_sfixed(2171.0/65536.0,1,-nbitq), 
to_sfixed(468.0/65536.0,1,-nbitq), 
to_sfixed(-2409.0/65536.0,1,-nbitq), 
to_sfixed(-340.0/65536.0,1,-nbitq), 
to_sfixed(1971.0/65536.0,1,-nbitq), 
to_sfixed(4679.0/65536.0,1,-nbitq), 
to_sfixed(3064.0/65536.0,1,-nbitq), 
to_sfixed(347.0/65536.0,1,-nbitq), 
to_sfixed(4983.0/65536.0,1,-nbitq), 
to_sfixed(-3163.0/65536.0,1,-nbitq), 
to_sfixed(-4845.0/65536.0,1,-nbitq), 
to_sfixed(-1761.0/65536.0,1,-nbitq), 
to_sfixed(1611.0/65536.0,1,-nbitq), 
to_sfixed(12.0/65536.0,1,-nbitq), 
to_sfixed(-2881.0/65536.0,1,-nbitq), 
to_sfixed(3715.0/65536.0,1,-nbitq), 
to_sfixed(2565.0/65536.0,1,-nbitq), 
to_sfixed(4505.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2266.0/65536.0,1,-nbitq), 
to_sfixed(6404.0/65536.0,1,-nbitq), 
to_sfixed(-1760.0/65536.0,1,-nbitq), 
to_sfixed(-1974.0/65536.0,1,-nbitq), 
to_sfixed(58.0/65536.0,1,-nbitq), 
to_sfixed(-4480.0/65536.0,1,-nbitq), 
to_sfixed(-788.0/65536.0,1,-nbitq), 
to_sfixed(-5485.0/65536.0,1,-nbitq), 
to_sfixed(-2541.0/65536.0,1,-nbitq), 
to_sfixed(-1948.0/65536.0,1,-nbitq), 
to_sfixed(4170.0/65536.0,1,-nbitq), 
to_sfixed(-888.0/65536.0,1,-nbitq), 
to_sfixed(1385.0/65536.0,1,-nbitq), 
to_sfixed(3550.0/65536.0,1,-nbitq), 
to_sfixed(4903.0/65536.0,1,-nbitq), 
to_sfixed(3312.0/65536.0,1,-nbitq), 
to_sfixed(-2265.0/65536.0,1,-nbitq), 
to_sfixed(770.0/65536.0,1,-nbitq), 
to_sfixed(-2861.0/65536.0,1,-nbitq), 
to_sfixed(-2276.0/65536.0,1,-nbitq), 
to_sfixed(-1735.0/65536.0,1,-nbitq), 
to_sfixed(2806.0/65536.0,1,-nbitq), 
to_sfixed(6299.0/65536.0,1,-nbitq), 
to_sfixed(-6750.0/65536.0,1,-nbitq), 
to_sfixed(-209.0/65536.0,1,-nbitq), 
to_sfixed(-1702.0/65536.0,1,-nbitq), 
to_sfixed(-131.0/65536.0,1,-nbitq), 
to_sfixed(-4606.0/65536.0,1,-nbitq), 
to_sfixed(-2205.0/65536.0,1,-nbitq), 
to_sfixed(-2307.0/65536.0,1,-nbitq), 
to_sfixed(387.0/65536.0,1,-nbitq), 
to_sfixed(-150.0/65536.0,1,-nbitq), 
to_sfixed(-2944.0/65536.0,1,-nbitq), 
to_sfixed(1104.0/65536.0,1,-nbitq), 
to_sfixed(489.0/65536.0,1,-nbitq), 
to_sfixed(-1454.0/65536.0,1,-nbitq), 
to_sfixed(-3620.0/65536.0,1,-nbitq), 
to_sfixed(-2203.0/65536.0,1,-nbitq), 
to_sfixed(447.0/65536.0,1,-nbitq), 
to_sfixed(-2628.0/65536.0,1,-nbitq), 
to_sfixed(862.0/65536.0,1,-nbitq), 
to_sfixed(-3285.0/65536.0,1,-nbitq), 
to_sfixed(-3275.0/65536.0,1,-nbitq), 
to_sfixed(-2374.0/65536.0,1,-nbitq), 
to_sfixed(-1132.0/65536.0,1,-nbitq), 
to_sfixed(1488.0/65536.0,1,-nbitq), 
to_sfixed(-1248.0/65536.0,1,-nbitq), 
to_sfixed(-5482.0/65536.0,1,-nbitq), 
to_sfixed(707.0/65536.0,1,-nbitq), 
to_sfixed(-1807.0/65536.0,1,-nbitq), 
to_sfixed(2575.0/65536.0,1,-nbitq), 
to_sfixed(2026.0/65536.0,1,-nbitq), 
to_sfixed(5354.0/65536.0,1,-nbitq), 
to_sfixed(2154.0/65536.0,1,-nbitq), 
to_sfixed(1618.0/65536.0,1,-nbitq), 
to_sfixed(2437.0/65536.0,1,-nbitq), 
to_sfixed(1434.0/65536.0,1,-nbitq), 
to_sfixed(628.0/65536.0,1,-nbitq), 
to_sfixed(-843.0/65536.0,1,-nbitq), 
to_sfixed(3448.0/65536.0,1,-nbitq), 
to_sfixed(2202.0/65536.0,1,-nbitq), 
to_sfixed(-2907.0/65536.0,1,-nbitq), 
to_sfixed(265.0/65536.0,1,-nbitq), 
to_sfixed(-780.0/65536.0,1,-nbitq), 
to_sfixed(1653.0/65536.0,1,-nbitq), 
to_sfixed(2637.0/65536.0,1,-nbitq), 
to_sfixed(1743.0/65536.0,1,-nbitq), 
to_sfixed(2926.0/65536.0,1,-nbitq), 
to_sfixed(1678.0/65536.0,1,-nbitq), 
to_sfixed(-797.0/65536.0,1,-nbitq), 
to_sfixed(2821.0/65536.0,1,-nbitq), 
to_sfixed(-5890.0/65536.0,1,-nbitq), 
to_sfixed(-1056.0/65536.0,1,-nbitq), 
to_sfixed(2567.0/65536.0,1,-nbitq), 
to_sfixed(-80.0/65536.0,1,-nbitq), 
to_sfixed(793.0/65536.0,1,-nbitq), 
to_sfixed(1447.0/65536.0,1,-nbitq), 
to_sfixed(-1453.0/65536.0,1,-nbitq), 
to_sfixed(2064.0/65536.0,1,-nbitq), 
to_sfixed(611.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1162.0/65536.0,1,-nbitq), 
to_sfixed(3108.0/65536.0,1,-nbitq), 
to_sfixed(-743.0/65536.0,1,-nbitq), 
to_sfixed(778.0/65536.0,1,-nbitq), 
to_sfixed(-519.0/65536.0,1,-nbitq), 
to_sfixed(-2426.0/65536.0,1,-nbitq), 
to_sfixed(-152.0/65536.0,1,-nbitq), 
to_sfixed(-2456.0/65536.0,1,-nbitq), 
to_sfixed(3128.0/65536.0,1,-nbitq), 
to_sfixed(-2369.0/65536.0,1,-nbitq), 
to_sfixed(1833.0/65536.0,1,-nbitq), 
to_sfixed(-4415.0/65536.0,1,-nbitq), 
to_sfixed(598.0/65536.0,1,-nbitq), 
to_sfixed(3507.0/65536.0,1,-nbitq), 
to_sfixed(-1481.0/65536.0,1,-nbitq), 
to_sfixed(2006.0/65536.0,1,-nbitq), 
to_sfixed(-708.0/65536.0,1,-nbitq), 
to_sfixed(-1008.0/65536.0,1,-nbitq), 
to_sfixed(-3899.0/65536.0,1,-nbitq), 
to_sfixed(-2349.0/65536.0,1,-nbitq), 
to_sfixed(-4458.0/65536.0,1,-nbitq), 
to_sfixed(-1798.0/65536.0,1,-nbitq), 
to_sfixed(7482.0/65536.0,1,-nbitq), 
to_sfixed(-2649.0/65536.0,1,-nbitq), 
to_sfixed(-3192.0/65536.0,1,-nbitq), 
to_sfixed(-5667.0/65536.0,1,-nbitq), 
to_sfixed(-444.0/65536.0,1,-nbitq), 
to_sfixed(-4546.0/65536.0,1,-nbitq), 
to_sfixed(-3011.0/65536.0,1,-nbitq), 
to_sfixed(-123.0/65536.0,1,-nbitq), 
to_sfixed(-2455.0/65536.0,1,-nbitq), 
to_sfixed(-1745.0/65536.0,1,-nbitq), 
to_sfixed(-4462.0/65536.0,1,-nbitq), 
to_sfixed(-245.0/65536.0,1,-nbitq), 
to_sfixed(-1827.0/65536.0,1,-nbitq), 
to_sfixed(670.0/65536.0,1,-nbitq), 
to_sfixed(-2622.0/65536.0,1,-nbitq), 
to_sfixed(-993.0/65536.0,1,-nbitq), 
to_sfixed(3722.0/65536.0,1,-nbitq), 
to_sfixed(1725.0/65536.0,1,-nbitq), 
to_sfixed(-668.0/65536.0,1,-nbitq), 
to_sfixed(-209.0/65536.0,1,-nbitq), 
to_sfixed(-6802.0/65536.0,1,-nbitq), 
to_sfixed(-1955.0/65536.0,1,-nbitq), 
to_sfixed(2403.0/65536.0,1,-nbitq), 
to_sfixed(3191.0/65536.0,1,-nbitq), 
to_sfixed(445.0/65536.0,1,-nbitq), 
to_sfixed(-4474.0/65536.0,1,-nbitq), 
to_sfixed(-1693.0/65536.0,1,-nbitq), 
to_sfixed(703.0/65536.0,1,-nbitq), 
to_sfixed(-728.0/65536.0,1,-nbitq), 
to_sfixed(-804.0/65536.0,1,-nbitq), 
to_sfixed(1170.0/65536.0,1,-nbitq), 
to_sfixed(-746.0/65536.0,1,-nbitq), 
to_sfixed(1289.0/65536.0,1,-nbitq), 
to_sfixed(-1029.0/65536.0,1,-nbitq), 
to_sfixed(-2570.0/65536.0,1,-nbitq), 
to_sfixed(-1772.0/65536.0,1,-nbitq), 
to_sfixed(-2382.0/65536.0,1,-nbitq), 
to_sfixed(7180.0/65536.0,1,-nbitq), 
to_sfixed(2151.0/65536.0,1,-nbitq), 
to_sfixed(-875.0/65536.0,1,-nbitq), 
to_sfixed(-1735.0/65536.0,1,-nbitq), 
to_sfixed(-793.0/65536.0,1,-nbitq), 
to_sfixed(278.0/65536.0,1,-nbitq), 
to_sfixed(3267.0/65536.0,1,-nbitq), 
to_sfixed(-2915.0/65536.0,1,-nbitq), 
to_sfixed(3653.0/65536.0,1,-nbitq), 
to_sfixed(2531.0/65536.0,1,-nbitq), 
to_sfixed(1467.0/65536.0,1,-nbitq), 
to_sfixed(464.0/65536.0,1,-nbitq), 
to_sfixed(-4479.0/65536.0,1,-nbitq), 
to_sfixed(1061.0/65536.0,1,-nbitq), 
to_sfixed(-1901.0/65536.0,1,-nbitq), 
to_sfixed(-2479.0/65536.0,1,-nbitq), 
to_sfixed(502.0/65536.0,1,-nbitq), 
to_sfixed(3358.0/65536.0,1,-nbitq), 
to_sfixed(-448.0/65536.0,1,-nbitq), 
to_sfixed(-1915.0/65536.0,1,-nbitq), 
to_sfixed(2206.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3530.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(-1208.0/65536.0,1,-nbitq), 
to_sfixed(2537.0/65536.0,1,-nbitq), 
to_sfixed(3084.0/65536.0,1,-nbitq), 
to_sfixed(-3113.0/65536.0,1,-nbitq), 
to_sfixed(-2725.0/65536.0,1,-nbitq), 
to_sfixed(-5214.0/65536.0,1,-nbitq), 
to_sfixed(3175.0/65536.0,1,-nbitq), 
to_sfixed(1214.0/65536.0,1,-nbitq), 
to_sfixed(-102.0/65536.0,1,-nbitq), 
to_sfixed(-1307.0/65536.0,1,-nbitq), 
to_sfixed(1224.0/65536.0,1,-nbitq), 
to_sfixed(4443.0/65536.0,1,-nbitq), 
to_sfixed(-138.0/65536.0,1,-nbitq), 
to_sfixed(1056.0/65536.0,1,-nbitq), 
to_sfixed(1038.0/65536.0,1,-nbitq), 
to_sfixed(-2721.0/65536.0,1,-nbitq), 
to_sfixed(-4458.0/65536.0,1,-nbitq), 
to_sfixed(-250.0/65536.0,1,-nbitq), 
to_sfixed(-4520.0/65536.0,1,-nbitq), 
to_sfixed(956.0/65536.0,1,-nbitq), 
to_sfixed(6242.0/65536.0,1,-nbitq), 
to_sfixed(2714.0/65536.0,1,-nbitq), 
to_sfixed(1306.0/65536.0,1,-nbitq), 
to_sfixed(-3218.0/65536.0,1,-nbitq), 
to_sfixed(2121.0/65536.0,1,-nbitq), 
to_sfixed(-2091.0/65536.0,1,-nbitq), 
to_sfixed(-2623.0/65536.0,1,-nbitq), 
to_sfixed(903.0/65536.0,1,-nbitq), 
to_sfixed(69.0/65536.0,1,-nbitq), 
to_sfixed(-2482.0/65536.0,1,-nbitq), 
to_sfixed(-3466.0/65536.0,1,-nbitq), 
to_sfixed(5049.0/65536.0,1,-nbitq), 
to_sfixed(-396.0/65536.0,1,-nbitq), 
to_sfixed(-2672.0/65536.0,1,-nbitq), 
to_sfixed(-4644.0/65536.0,1,-nbitq), 
to_sfixed(3776.0/65536.0,1,-nbitq), 
to_sfixed(773.0/65536.0,1,-nbitq), 
to_sfixed(-590.0/65536.0,1,-nbitq), 
to_sfixed(261.0/65536.0,1,-nbitq), 
to_sfixed(-3178.0/65536.0,1,-nbitq), 
to_sfixed(-6949.0/65536.0,1,-nbitq), 
to_sfixed(3282.0/65536.0,1,-nbitq), 
to_sfixed(-1073.0/65536.0,1,-nbitq), 
to_sfixed(-4258.0/65536.0,1,-nbitq), 
to_sfixed(-2516.0/65536.0,1,-nbitq), 
to_sfixed(-1819.0/65536.0,1,-nbitq), 
to_sfixed(-409.0/65536.0,1,-nbitq), 
to_sfixed(1325.0/65536.0,1,-nbitq), 
to_sfixed(-2605.0/65536.0,1,-nbitq), 
to_sfixed(1070.0/65536.0,1,-nbitq), 
to_sfixed(-1820.0/65536.0,1,-nbitq), 
to_sfixed(-1765.0/65536.0,1,-nbitq), 
to_sfixed(127.0/65536.0,1,-nbitq), 
to_sfixed(1871.0/65536.0,1,-nbitq), 
to_sfixed(2733.0/65536.0,1,-nbitq), 
to_sfixed(2888.0/65536.0,1,-nbitq), 
to_sfixed(2889.0/65536.0,1,-nbitq), 
to_sfixed(7949.0/65536.0,1,-nbitq), 
to_sfixed(1280.0/65536.0,1,-nbitq), 
to_sfixed(1534.0/65536.0,1,-nbitq), 
to_sfixed(600.0/65536.0,1,-nbitq), 
to_sfixed(-864.0/65536.0,1,-nbitq), 
to_sfixed(-465.0/65536.0,1,-nbitq), 
to_sfixed(3644.0/65536.0,1,-nbitq), 
to_sfixed(-1167.0/65536.0,1,-nbitq), 
to_sfixed(-766.0/65536.0,1,-nbitq), 
to_sfixed(2768.0/65536.0,1,-nbitq), 
to_sfixed(-3320.0/65536.0,1,-nbitq), 
to_sfixed(142.0/65536.0,1,-nbitq), 
to_sfixed(-4856.0/65536.0,1,-nbitq), 
to_sfixed(-3129.0/65536.0,1,-nbitq), 
to_sfixed(619.0/65536.0,1,-nbitq), 
to_sfixed(-1368.0/65536.0,1,-nbitq), 
to_sfixed(3071.0/65536.0,1,-nbitq), 
to_sfixed(1418.0/65536.0,1,-nbitq), 
to_sfixed(1210.0/65536.0,1,-nbitq), 
to_sfixed(-3120.0/65536.0,1,-nbitq), 
to_sfixed(5567.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1566.0/65536.0,1,-nbitq), 
to_sfixed(2156.0/65536.0,1,-nbitq), 
to_sfixed(220.0/65536.0,1,-nbitq), 
to_sfixed(3242.0/65536.0,1,-nbitq), 
to_sfixed(4734.0/65536.0,1,-nbitq), 
to_sfixed(-1861.0/65536.0,1,-nbitq), 
to_sfixed(-6025.0/65536.0,1,-nbitq), 
to_sfixed(-431.0/65536.0,1,-nbitq), 
to_sfixed(-1675.0/65536.0,1,-nbitq), 
to_sfixed(-749.0/65536.0,1,-nbitq), 
to_sfixed(772.0/65536.0,1,-nbitq), 
to_sfixed(-834.0/65536.0,1,-nbitq), 
to_sfixed(-2251.0/65536.0,1,-nbitq), 
to_sfixed(2568.0/65536.0,1,-nbitq), 
to_sfixed(1333.0/65536.0,1,-nbitq), 
to_sfixed(476.0/65536.0,1,-nbitq), 
to_sfixed(-1594.0/65536.0,1,-nbitq), 
to_sfixed(-6768.0/65536.0,1,-nbitq), 
to_sfixed(-1256.0/65536.0,1,-nbitq), 
to_sfixed(-2540.0/65536.0,1,-nbitq), 
to_sfixed(-5026.0/65536.0,1,-nbitq), 
to_sfixed(-4835.0/65536.0,1,-nbitq), 
to_sfixed(1247.0/65536.0,1,-nbitq), 
to_sfixed(4268.0/65536.0,1,-nbitq), 
to_sfixed(2635.0/65536.0,1,-nbitq), 
to_sfixed(-2039.0/65536.0,1,-nbitq), 
to_sfixed(-446.0/65536.0,1,-nbitq), 
to_sfixed(-2809.0/65536.0,1,-nbitq), 
to_sfixed(-2385.0/65536.0,1,-nbitq), 
to_sfixed(1851.0/65536.0,1,-nbitq), 
to_sfixed(-3665.0/65536.0,1,-nbitq), 
to_sfixed(-53.0/65536.0,1,-nbitq), 
to_sfixed(-415.0/65536.0,1,-nbitq), 
to_sfixed(6350.0/65536.0,1,-nbitq), 
to_sfixed(1626.0/65536.0,1,-nbitq), 
to_sfixed(-1082.0/65536.0,1,-nbitq), 
to_sfixed(-4450.0/65536.0,1,-nbitq), 
to_sfixed(2929.0/65536.0,1,-nbitq), 
to_sfixed(-805.0/65536.0,1,-nbitq), 
to_sfixed(-1795.0/65536.0,1,-nbitq), 
to_sfixed(-48.0/65536.0,1,-nbitq), 
to_sfixed(797.0/65536.0,1,-nbitq), 
to_sfixed(-4554.0/65536.0,1,-nbitq), 
to_sfixed(5781.0/65536.0,1,-nbitq), 
to_sfixed(315.0/65536.0,1,-nbitq), 
to_sfixed(-4857.0/65536.0,1,-nbitq), 
to_sfixed(-1059.0/65536.0,1,-nbitq), 
to_sfixed(-5904.0/65536.0,1,-nbitq), 
to_sfixed(-35.0/65536.0,1,-nbitq), 
to_sfixed(3416.0/65536.0,1,-nbitq), 
to_sfixed(1937.0/65536.0,1,-nbitq), 
to_sfixed(464.0/65536.0,1,-nbitq), 
to_sfixed(-298.0/65536.0,1,-nbitq), 
to_sfixed(1552.0/65536.0,1,-nbitq), 
to_sfixed(3412.0/65536.0,1,-nbitq), 
to_sfixed(1601.0/65536.0,1,-nbitq), 
to_sfixed(3067.0/65536.0,1,-nbitq), 
to_sfixed(-2060.0/65536.0,1,-nbitq), 
to_sfixed(-787.0/65536.0,1,-nbitq), 
to_sfixed(5148.0/65536.0,1,-nbitq), 
to_sfixed(-4034.0/65536.0,1,-nbitq), 
to_sfixed(-2940.0/65536.0,1,-nbitq), 
to_sfixed(3142.0/65536.0,1,-nbitq), 
to_sfixed(1008.0/65536.0,1,-nbitq), 
to_sfixed(-1467.0/65536.0,1,-nbitq), 
to_sfixed(3407.0/65536.0,1,-nbitq), 
to_sfixed(-1688.0/65536.0,1,-nbitq), 
to_sfixed(694.0/65536.0,1,-nbitq), 
to_sfixed(-2141.0/65536.0,1,-nbitq), 
to_sfixed(-3563.0/65536.0,1,-nbitq), 
to_sfixed(-1001.0/65536.0,1,-nbitq), 
to_sfixed(-185.0/65536.0,1,-nbitq), 
to_sfixed(1157.0/65536.0,1,-nbitq), 
to_sfixed(-3107.0/65536.0,1,-nbitq), 
to_sfixed(631.0/65536.0,1,-nbitq), 
to_sfixed(869.0/65536.0,1,-nbitq), 
to_sfixed(-350.0/65536.0,1,-nbitq), 
to_sfixed(2447.0/65536.0,1,-nbitq), 
to_sfixed(-1437.0/65536.0,1,-nbitq), 
to_sfixed(1103.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1303.0/65536.0,1,-nbitq), 
to_sfixed(2502.0/65536.0,1,-nbitq), 
to_sfixed(777.0/65536.0,1,-nbitq), 
to_sfixed(2143.0/65536.0,1,-nbitq), 
to_sfixed(3742.0/65536.0,1,-nbitq), 
to_sfixed(2802.0/65536.0,1,-nbitq), 
to_sfixed(-5576.0/65536.0,1,-nbitq), 
to_sfixed(-1069.0/65536.0,1,-nbitq), 
to_sfixed(-1380.0/65536.0,1,-nbitq), 
to_sfixed(-259.0/65536.0,1,-nbitq), 
to_sfixed(4369.0/65536.0,1,-nbitq), 
to_sfixed(-3851.0/65536.0,1,-nbitq), 
to_sfixed(227.0/65536.0,1,-nbitq), 
to_sfixed(-1440.0/65536.0,1,-nbitq), 
to_sfixed(-2047.0/65536.0,1,-nbitq), 
to_sfixed(2321.0/65536.0,1,-nbitq), 
to_sfixed(-1941.0/65536.0,1,-nbitq), 
to_sfixed(-1472.0/65536.0,1,-nbitq), 
to_sfixed(-2332.0/65536.0,1,-nbitq), 
to_sfixed(1411.0/65536.0,1,-nbitq), 
to_sfixed(-4383.0/65536.0,1,-nbitq), 
to_sfixed(-3016.0/65536.0,1,-nbitq), 
to_sfixed(-1794.0/65536.0,1,-nbitq), 
to_sfixed(4596.0/65536.0,1,-nbitq), 
to_sfixed(-756.0/65536.0,1,-nbitq), 
to_sfixed(-2615.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(926.0/65536.0,1,-nbitq), 
to_sfixed(-2355.0/65536.0,1,-nbitq), 
to_sfixed(-1800.0/65536.0,1,-nbitq), 
to_sfixed(-1843.0/65536.0,1,-nbitq), 
to_sfixed(-87.0/65536.0,1,-nbitq), 
to_sfixed(-3105.0/65536.0,1,-nbitq), 
to_sfixed(7878.0/65536.0,1,-nbitq), 
to_sfixed(3025.0/65536.0,1,-nbitq), 
to_sfixed(-1218.0/65536.0,1,-nbitq), 
to_sfixed(-1417.0/65536.0,1,-nbitq), 
to_sfixed(-194.0/65536.0,1,-nbitq), 
to_sfixed(-2929.0/65536.0,1,-nbitq), 
to_sfixed(-920.0/65536.0,1,-nbitq), 
to_sfixed(3662.0/65536.0,1,-nbitq), 
to_sfixed(-2682.0/65536.0,1,-nbitq), 
to_sfixed(-1509.0/65536.0,1,-nbitq), 
to_sfixed(4471.0/65536.0,1,-nbitq), 
to_sfixed(-85.0/65536.0,1,-nbitq), 
to_sfixed(-6076.0/65536.0,1,-nbitq), 
to_sfixed(-2421.0/65536.0,1,-nbitq), 
to_sfixed(-3313.0/65536.0,1,-nbitq), 
to_sfixed(753.0/65536.0,1,-nbitq), 
to_sfixed(579.0/65536.0,1,-nbitq), 
to_sfixed(1899.0/65536.0,1,-nbitq), 
to_sfixed(1848.0/65536.0,1,-nbitq), 
to_sfixed(1434.0/65536.0,1,-nbitq), 
to_sfixed(-949.0/65536.0,1,-nbitq), 
to_sfixed(2617.0/65536.0,1,-nbitq), 
to_sfixed(49.0/65536.0,1,-nbitq), 
to_sfixed(-2006.0/65536.0,1,-nbitq), 
to_sfixed(676.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(4970.0/65536.0,1,-nbitq), 
to_sfixed(720.0/65536.0,1,-nbitq), 
to_sfixed(-655.0/65536.0,1,-nbitq), 
to_sfixed(-2546.0/65536.0,1,-nbitq), 
to_sfixed(2237.0/65536.0,1,-nbitq), 
to_sfixed(3269.0/65536.0,1,-nbitq), 
to_sfixed(5077.0/65536.0,1,-nbitq), 
to_sfixed(-3836.0/65536.0,1,-nbitq), 
to_sfixed(2834.0/65536.0,1,-nbitq), 
to_sfixed(-706.0/65536.0,1,-nbitq), 
to_sfixed(-3995.0/65536.0,1,-nbitq), 
to_sfixed(2525.0/65536.0,1,-nbitq), 
to_sfixed(-1834.0/65536.0,1,-nbitq), 
to_sfixed(314.0/65536.0,1,-nbitq), 
to_sfixed(2453.0/65536.0,1,-nbitq), 
to_sfixed(-2678.0/65536.0,1,-nbitq), 
to_sfixed(1353.0/65536.0,1,-nbitq), 
to_sfixed(3400.0/65536.0,1,-nbitq), 
to_sfixed(-2278.0/65536.0,1,-nbitq), 
to_sfixed(-25.0/65536.0,1,-nbitq), 
to_sfixed(4209.0/65536.0,1,-nbitq)  ), 
( to_sfixed(251.0/65536.0,1,-nbitq), 
to_sfixed(1399.0/65536.0,1,-nbitq), 
to_sfixed(2065.0/65536.0,1,-nbitq), 
to_sfixed(262.0/65536.0,1,-nbitq), 
to_sfixed(4428.0/65536.0,1,-nbitq), 
to_sfixed(24.0/65536.0,1,-nbitq), 
to_sfixed(82.0/65536.0,1,-nbitq), 
to_sfixed(485.0/65536.0,1,-nbitq), 
to_sfixed(652.0/65536.0,1,-nbitq), 
to_sfixed(1874.0/65536.0,1,-nbitq), 
to_sfixed(73.0/65536.0,1,-nbitq), 
to_sfixed(-2180.0/65536.0,1,-nbitq), 
to_sfixed(-430.0/65536.0,1,-nbitq), 
to_sfixed(1206.0/65536.0,1,-nbitq), 
to_sfixed(-1124.0/65536.0,1,-nbitq), 
to_sfixed(1763.0/65536.0,1,-nbitq), 
to_sfixed(-2938.0/65536.0,1,-nbitq), 
to_sfixed(-2990.0/65536.0,1,-nbitq), 
to_sfixed(-3295.0/65536.0,1,-nbitq), 
to_sfixed(3268.0/65536.0,1,-nbitq), 
to_sfixed(-372.0/65536.0,1,-nbitq), 
to_sfixed(-3512.0/65536.0,1,-nbitq), 
to_sfixed(-2813.0/65536.0,1,-nbitq), 
to_sfixed(3589.0/65536.0,1,-nbitq), 
to_sfixed(-903.0/65536.0,1,-nbitq), 
to_sfixed(1464.0/65536.0,1,-nbitq), 
to_sfixed(3192.0/65536.0,1,-nbitq), 
to_sfixed(-2094.0/65536.0,1,-nbitq), 
to_sfixed(-1682.0/65536.0,1,-nbitq), 
to_sfixed(1078.0/65536.0,1,-nbitq), 
to_sfixed(203.0/65536.0,1,-nbitq), 
to_sfixed(-1673.0/65536.0,1,-nbitq), 
to_sfixed(-5452.0/65536.0,1,-nbitq), 
to_sfixed(6618.0/65536.0,1,-nbitq), 
to_sfixed(-1233.0/65536.0,1,-nbitq), 
to_sfixed(-1047.0/65536.0,1,-nbitq), 
to_sfixed(1124.0/65536.0,1,-nbitq), 
to_sfixed(-2007.0/65536.0,1,-nbitq), 
to_sfixed(1354.0/65536.0,1,-nbitq), 
to_sfixed(1768.0/65536.0,1,-nbitq), 
to_sfixed(3739.0/65536.0,1,-nbitq), 
to_sfixed(-958.0/65536.0,1,-nbitq), 
to_sfixed(-10.0/65536.0,1,-nbitq), 
to_sfixed(1566.0/65536.0,1,-nbitq), 
to_sfixed(1087.0/65536.0,1,-nbitq), 
to_sfixed(-2419.0/65536.0,1,-nbitq), 
to_sfixed(-2789.0/65536.0,1,-nbitq), 
to_sfixed(-3253.0/65536.0,1,-nbitq), 
to_sfixed(2823.0/65536.0,1,-nbitq), 
to_sfixed(406.0/65536.0,1,-nbitq), 
to_sfixed(-1279.0/65536.0,1,-nbitq), 
to_sfixed(2335.0/65536.0,1,-nbitq), 
to_sfixed(2229.0/65536.0,1,-nbitq), 
to_sfixed(-2599.0/65536.0,1,-nbitq), 
to_sfixed(713.0/65536.0,1,-nbitq), 
to_sfixed(664.0/65536.0,1,-nbitq), 
to_sfixed(558.0/65536.0,1,-nbitq), 
to_sfixed(-384.0/65536.0,1,-nbitq), 
to_sfixed(1118.0/65536.0,1,-nbitq), 
to_sfixed(4831.0/65536.0,1,-nbitq), 
to_sfixed(-2296.0/65536.0,1,-nbitq), 
to_sfixed(-797.0/65536.0,1,-nbitq), 
to_sfixed(-576.0/65536.0,1,-nbitq), 
to_sfixed(1296.0/65536.0,1,-nbitq), 
to_sfixed(-1602.0/65536.0,1,-nbitq), 
to_sfixed(9057.0/65536.0,1,-nbitq), 
to_sfixed(-3181.0/65536.0,1,-nbitq), 
to_sfixed(457.0/65536.0,1,-nbitq), 
to_sfixed(92.0/65536.0,1,-nbitq), 
to_sfixed(-3717.0/65536.0,1,-nbitq), 
to_sfixed(-683.0/65536.0,1,-nbitq), 
to_sfixed(3866.0/65536.0,1,-nbitq), 
to_sfixed(-3843.0/65536.0,1,-nbitq), 
to_sfixed(2435.0/65536.0,1,-nbitq), 
to_sfixed(2056.0/65536.0,1,-nbitq), 
to_sfixed(-1087.0/65536.0,1,-nbitq), 
to_sfixed(2337.0/65536.0,1,-nbitq), 
to_sfixed(3016.0/65536.0,1,-nbitq), 
to_sfixed(-2405.0/65536.0,1,-nbitq), 
to_sfixed(4193.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1985.0/65536.0,1,-nbitq), 
to_sfixed(2292.0/65536.0,1,-nbitq), 
to_sfixed(-839.0/65536.0,1,-nbitq), 
to_sfixed(-950.0/65536.0,1,-nbitq), 
to_sfixed(-1555.0/65536.0,1,-nbitq), 
to_sfixed(-407.0/65536.0,1,-nbitq), 
to_sfixed(-3907.0/65536.0,1,-nbitq), 
to_sfixed(1515.0/65536.0,1,-nbitq), 
to_sfixed(-611.0/65536.0,1,-nbitq), 
to_sfixed(1706.0/65536.0,1,-nbitq), 
to_sfixed(204.0/65536.0,1,-nbitq), 
to_sfixed(-1266.0/65536.0,1,-nbitq), 
to_sfixed(1822.0/65536.0,1,-nbitq), 
to_sfixed(2475.0/65536.0,1,-nbitq), 
to_sfixed(1285.0/65536.0,1,-nbitq), 
to_sfixed(2750.0/65536.0,1,-nbitq), 
to_sfixed(-2811.0/65536.0,1,-nbitq), 
to_sfixed(-415.0/65536.0,1,-nbitq), 
to_sfixed(-795.0/65536.0,1,-nbitq), 
to_sfixed(-1211.0/65536.0,1,-nbitq), 
to_sfixed(1336.0/65536.0,1,-nbitq), 
to_sfixed(-7007.0/65536.0,1,-nbitq), 
to_sfixed(-3281.0/65536.0,1,-nbitq), 
to_sfixed(-2373.0/65536.0,1,-nbitq), 
to_sfixed(3331.0/65536.0,1,-nbitq), 
to_sfixed(593.0/65536.0,1,-nbitq), 
to_sfixed(579.0/65536.0,1,-nbitq), 
to_sfixed(946.0/65536.0,1,-nbitq), 
to_sfixed(-3349.0/65536.0,1,-nbitq), 
to_sfixed(2857.0/65536.0,1,-nbitq), 
to_sfixed(342.0/65536.0,1,-nbitq), 
to_sfixed(2966.0/65536.0,1,-nbitq), 
to_sfixed(-237.0/65536.0,1,-nbitq), 
to_sfixed(1495.0/65536.0,1,-nbitq), 
to_sfixed(-2395.0/65536.0,1,-nbitq), 
to_sfixed(2069.0/65536.0,1,-nbitq), 
to_sfixed(-1838.0/65536.0,1,-nbitq), 
to_sfixed(1740.0/65536.0,1,-nbitq), 
to_sfixed(591.0/65536.0,1,-nbitq), 
to_sfixed(859.0/65536.0,1,-nbitq), 
to_sfixed(-409.0/65536.0,1,-nbitq), 
to_sfixed(-118.0/65536.0,1,-nbitq), 
to_sfixed(-728.0/65536.0,1,-nbitq), 
to_sfixed(474.0/65536.0,1,-nbitq), 
to_sfixed(162.0/65536.0,1,-nbitq), 
to_sfixed(688.0/65536.0,1,-nbitq), 
to_sfixed(-2480.0/65536.0,1,-nbitq), 
to_sfixed(-4299.0/65536.0,1,-nbitq), 
to_sfixed(1399.0/65536.0,1,-nbitq), 
to_sfixed(731.0/65536.0,1,-nbitq), 
to_sfixed(2986.0/65536.0,1,-nbitq), 
to_sfixed(1693.0/65536.0,1,-nbitq), 
to_sfixed(1783.0/65536.0,1,-nbitq), 
to_sfixed(-2702.0/65536.0,1,-nbitq), 
to_sfixed(4853.0/65536.0,1,-nbitq), 
to_sfixed(821.0/65536.0,1,-nbitq), 
to_sfixed(1688.0/65536.0,1,-nbitq), 
to_sfixed(3277.0/65536.0,1,-nbitq), 
to_sfixed(2271.0/65536.0,1,-nbitq), 
to_sfixed(506.0/65536.0,1,-nbitq), 
to_sfixed(-2333.0/65536.0,1,-nbitq), 
to_sfixed(-2330.0/65536.0,1,-nbitq), 
to_sfixed(-2623.0/65536.0,1,-nbitq), 
to_sfixed(-3426.0/65536.0,1,-nbitq), 
to_sfixed(1778.0/65536.0,1,-nbitq), 
to_sfixed(5441.0/65536.0,1,-nbitq), 
to_sfixed(1747.0/65536.0,1,-nbitq), 
to_sfixed(-350.0/65536.0,1,-nbitq), 
to_sfixed(-721.0/65536.0,1,-nbitq), 
to_sfixed(-4652.0/65536.0,1,-nbitq), 
to_sfixed(-630.0/65536.0,1,-nbitq), 
to_sfixed(3659.0/65536.0,1,-nbitq), 
to_sfixed(-2614.0/65536.0,1,-nbitq), 
to_sfixed(1211.0/65536.0,1,-nbitq), 
to_sfixed(1571.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(-1376.0/65536.0,1,-nbitq), 
to_sfixed(1098.0/65536.0,1,-nbitq), 
to_sfixed(-333.0/65536.0,1,-nbitq), 
to_sfixed(-129.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1290.0/65536.0,1,-nbitq), 
to_sfixed(1387.0/65536.0,1,-nbitq), 
to_sfixed(-370.0/65536.0,1,-nbitq), 
to_sfixed(2465.0/65536.0,1,-nbitq), 
to_sfixed(-1823.0/65536.0,1,-nbitq), 
to_sfixed(-1246.0/65536.0,1,-nbitq), 
to_sfixed(-1506.0/65536.0,1,-nbitq), 
to_sfixed(557.0/65536.0,1,-nbitq), 
to_sfixed(-3029.0/65536.0,1,-nbitq), 
to_sfixed(1269.0/65536.0,1,-nbitq), 
to_sfixed(-3033.0/65536.0,1,-nbitq), 
to_sfixed(-1825.0/65536.0,1,-nbitq), 
to_sfixed(-1784.0/65536.0,1,-nbitq), 
to_sfixed(-39.0/65536.0,1,-nbitq), 
to_sfixed(3256.0/65536.0,1,-nbitq), 
to_sfixed(-1390.0/65536.0,1,-nbitq), 
to_sfixed(-3166.0/65536.0,1,-nbitq), 
to_sfixed(2708.0/65536.0,1,-nbitq), 
to_sfixed(2111.0/65536.0,1,-nbitq), 
to_sfixed(555.0/65536.0,1,-nbitq), 
to_sfixed(-641.0/65536.0,1,-nbitq), 
to_sfixed(-6477.0/65536.0,1,-nbitq), 
to_sfixed(2847.0/65536.0,1,-nbitq), 
to_sfixed(-1405.0/65536.0,1,-nbitq), 
to_sfixed(1019.0/65536.0,1,-nbitq), 
to_sfixed(118.0/65536.0,1,-nbitq), 
to_sfixed(-6452.0/65536.0,1,-nbitq), 
to_sfixed(-607.0/65536.0,1,-nbitq), 
to_sfixed(-4397.0/65536.0,1,-nbitq), 
to_sfixed(-1380.0/65536.0,1,-nbitq), 
to_sfixed(1676.0/65536.0,1,-nbitq), 
to_sfixed(2597.0/65536.0,1,-nbitq), 
to_sfixed(-5975.0/65536.0,1,-nbitq), 
to_sfixed(-2045.0/65536.0,1,-nbitq), 
to_sfixed(1888.0/65536.0,1,-nbitq), 
to_sfixed(3085.0/65536.0,1,-nbitq), 
to_sfixed(267.0/65536.0,1,-nbitq), 
to_sfixed(2319.0/65536.0,1,-nbitq), 
to_sfixed(1602.0/65536.0,1,-nbitq), 
to_sfixed(1136.0/65536.0,1,-nbitq), 
to_sfixed(2307.0/65536.0,1,-nbitq), 
to_sfixed(2360.0/65536.0,1,-nbitq), 
to_sfixed(-1788.0/65536.0,1,-nbitq), 
to_sfixed(2235.0/65536.0,1,-nbitq), 
to_sfixed(1381.0/65536.0,1,-nbitq), 
to_sfixed(-1257.0/65536.0,1,-nbitq), 
to_sfixed(-1363.0/65536.0,1,-nbitq), 
to_sfixed(-2809.0/65536.0,1,-nbitq), 
to_sfixed(679.0/65536.0,1,-nbitq), 
to_sfixed(884.0/65536.0,1,-nbitq), 
to_sfixed(-252.0/65536.0,1,-nbitq), 
to_sfixed(2177.0/65536.0,1,-nbitq), 
to_sfixed(3043.0/65536.0,1,-nbitq), 
to_sfixed(-4797.0/65536.0,1,-nbitq), 
to_sfixed(-1710.0/65536.0,1,-nbitq), 
to_sfixed(-818.0/65536.0,1,-nbitq), 
to_sfixed(-217.0/65536.0,1,-nbitq), 
to_sfixed(1715.0/65536.0,1,-nbitq), 
to_sfixed(1137.0/65536.0,1,-nbitq), 
to_sfixed(5871.0/65536.0,1,-nbitq), 
to_sfixed(2407.0/65536.0,1,-nbitq), 
to_sfixed(-2617.0/65536.0,1,-nbitq), 
to_sfixed(2926.0/65536.0,1,-nbitq), 
to_sfixed(-2467.0/65536.0,1,-nbitq), 
to_sfixed(4686.0/65536.0,1,-nbitq), 
to_sfixed(3728.0/65536.0,1,-nbitq), 
to_sfixed(-736.0/65536.0,1,-nbitq), 
to_sfixed(-5739.0/65536.0,1,-nbitq), 
to_sfixed(619.0/65536.0,1,-nbitq), 
to_sfixed(289.0/65536.0,1,-nbitq), 
to_sfixed(-2796.0/65536.0,1,-nbitq), 
to_sfixed(937.0/65536.0,1,-nbitq), 
to_sfixed(-1573.0/65536.0,1,-nbitq), 
to_sfixed(-2322.0/65536.0,1,-nbitq), 
to_sfixed(-2847.0/65536.0,1,-nbitq), 
to_sfixed(-450.0/65536.0,1,-nbitq), 
to_sfixed(-4063.0/65536.0,1,-nbitq), 
to_sfixed(1853.0/65536.0,1,-nbitq), 
to_sfixed(-2114.0/65536.0,1,-nbitq), 
to_sfixed(2836.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-798.0/65536.0,1,-nbitq), 
to_sfixed(-1525.0/65536.0,1,-nbitq), 
to_sfixed(2719.0/65536.0,1,-nbitq), 
to_sfixed(1730.0/65536.0,1,-nbitq), 
to_sfixed(1584.0/65536.0,1,-nbitq), 
to_sfixed(-3318.0/65536.0,1,-nbitq), 
to_sfixed(-337.0/65536.0,1,-nbitq), 
to_sfixed(-1186.0/65536.0,1,-nbitq), 
to_sfixed(-3066.0/65536.0,1,-nbitq), 
to_sfixed(-2223.0/65536.0,1,-nbitq), 
to_sfixed(-1939.0/65536.0,1,-nbitq), 
to_sfixed(-3638.0/65536.0,1,-nbitq), 
to_sfixed(-1334.0/65536.0,1,-nbitq), 
to_sfixed(-1836.0/65536.0,1,-nbitq), 
to_sfixed(-161.0/65536.0,1,-nbitq), 
to_sfixed(-117.0/65536.0,1,-nbitq), 
to_sfixed(782.0/65536.0,1,-nbitq), 
to_sfixed(2887.0/65536.0,1,-nbitq), 
to_sfixed(-273.0/65536.0,1,-nbitq), 
to_sfixed(2558.0/65536.0,1,-nbitq), 
to_sfixed(561.0/65536.0,1,-nbitq), 
to_sfixed(186.0/65536.0,1,-nbitq), 
to_sfixed(-2137.0/65536.0,1,-nbitq), 
to_sfixed(-2617.0/65536.0,1,-nbitq), 
to_sfixed(898.0/65536.0,1,-nbitq), 
to_sfixed(2613.0/65536.0,1,-nbitq), 
to_sfixed(-6003.0/65536.0,1,-nbitq), 
to_sfixed(-2628.0/65536.0,1,-nbitq), 
to_sfixed(-2779.0/65536.0,1,-nbitq), 
to_sfixed(1253.0/65536.0,1,-nbitq), 
to_sfixed(5857.0/65536.0,1,-nbitq), 
to_sfixed(-1626.0/65536.0,1,-nbitq), 
to_sfixed(-1741.0/65536.0,1,-nbitq), 
to_sfixed(-146.0/65536.0,1,-nbitq), 
to_sfixed(-218.0/65536.0,1,-nbitq), 
to_sfixed(-2571.0/65536.0,1,-nbitq), 
to_sfixed(-2958.0/65536.0,1,-nbitq), 
to_sfixed(1848.0/65536.0,1,-nbitq), 
to_sfixed(-3609.0/65536.0,1,-nbitq), 
to_sfixed(-326.0/65536.0,1,-nbitq), 
to_sfixed(1130.0/65536.0,1,-nbitq), 
to_sfixed(2453.0/65536.0,1,-nbitq), 
to_sfixed(-3616.0/65536.0,1,-nbitq), 
to_sfixed(1068.0/65536.0,1,-nbitq), 
to_sfixed(1238.0/65536.0,1,-nbitq), 
to_sfixed(-1960.0/65536.0,1,-nbitq), 
to_sfixed(4047.0/65536.0,1,-nbitq), 
to_sfixed(-3016.0/65536.0,1,-nbitq), 
to_sfixed(1012.0/65536.0,1,-nbitq), 
to_sfixed(3121.0/65536.0,1,-nbitq), 
to_sfixed(2337.0/65536.0,1,-nbitq), 
to_sfixed(492.0/65536.0,1,-nbitq), 
to_sfixed(4370.0/65536.0,1,-nbitq), 
to_sfixed(-1940.0/65536.0,1,-nbitq), 
to_sfixed(2751.0/65536.0,1,-nbitq), 
to_sfixed(-1548.0/65536.0,1,-nbitq), 
to_sfixed(307.0/65536.0,1,-nbitq), 
to_sfixed(2412.0/65536.0,1,-nbitq), 
to_sfixed(-2083.0/65536.0,1,-nbitq), 
to_sfixed(5248.0/65536.0,1,-nbitq), 
to_sfixed(-143.0/65536.0,1,-nbitq), 
to_sfixed(270.0/65536.0,1,-nbitq), 
to_sfixed(-1274.0/65536.0,1,-nbitq), 
to_sfixed(-2916.0/65536.0,1,-nbitq), 
to_sfixed(615.0/65536.0,1,-nbitq), 
to_sfixed(3386.0/65536.0,1,-nbitq), 
to_sfixed(1216.0/65536.0,1,-nbitq), 
to_sfixed(-3575.0/65536.0,1,-nbitq), 
to_sfixed(3767.0/65536.0,1,-nbitq), 
to_sfixed(1571.0/65536.0,1,-nbitq), 
to_sfixed(-2907.0/65536.0,1,-nbitq), 
to_sfixed(2603.0/65536.0,1,-nbitq), 
to_sfixed(3008.0/65536.0,1,-nbitq), 
to_sfixed(-1346.0/65536.0,1,-nbitq), 
to_sfixed(803.0/65536.0,1,-nbitq), 
to_sfixed(-2954.0/65536.0,1,-nbitq), 
to_sfixed(450.0/65536.0,1,-nbitq), 
to_sfixed(769.0/65536.0,1,-nbitq), 
to_sfixed(-2154.0/65536.0,1,-nbitq), 
to_sfixed(3242.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1158.0/65536.0,1,-nbitq), 
to_sfixed(311.0/65536.0,1,-nbitq), 
to_sfixed(3968.0/65536.0,1,-nbitq), 
to_sfixed(-1567.0/65536.0,1,-nbitq), 
to_sfixed(-4694.0/65536.0,1,-nbitq), 
to_sfixed(1267.0/65536.0,1,-nbitq), 
to_sfixed(-1931.0/65536.0,1,-nbitq), 
to_sfixed(1153.0/65536.0,1,-nbitq), 
to_sfixed(-1765.0/65536.0,1,-nbitq), 
to_sfixed(-2396.0/65536.0,1,-nbitq), 
to_sfixed(-3219.0/65536.0,1,-nbitq), 
to_sfixed(587.0/65536.0,1,-nbitq), 
to_sfixed(-1509.0/65536.0,1,-nbitq), 
to_sfixed(-1325.0/65536.0,1,-nbitq), 
to_sfixed(1722.0/65536.0,1,-nbitq), 
to_sfixed(2317.0/65536.0,1,-nbitq), 
to_sfixed(1555.0/65536.0,1,-nbitq), 
to_sfixed(445.0/65536.0,1,-nbitq), 
to_sfixed(-730.0/65536.0,1,-nbitq), 
to_sfixed(1367.0/65536.0,1,-nbitq), 
to_sfixed(-4435.0/65536.0,1,-nbitq), 
to_sfixed(-1546.0/65536.0,1,-nbitq), 
to_sfixed(908.0/65536.0,1,-nbitq), 
to_sfixed(1949.0/65536.0,1,-nbitq), 
to_sfixed(-1050.0/65536.0,1,-nbitq), 
to_sfixed(4535.0/65536.0,1,-nbitq), 
to_sfixed(-4964.0/65536.0,1,-nbitq), 
to_sfixed(1712.0/65536.0,1,-nbitq), 
to_sfixed(-4944.0/65536.0,1,-nbitq), 
to_sfixed(-1123.0/65536.0,1,-nbitq), 
to_sfixed(4732.0/65536.0,1,-nbitq), 
to_sfixed(332.0/65536.0,1,-nbitq), 
to_sfixed(-5396.0/65536.0,1,-nbitq), 
to_sfixed(-2282.0/65536.0,1,-nbitq), 
to_sfixed(-1288.0/65536.0,1,-nbitq), 
to_sfixed(-2338.0/65536.0,1,-nbitq), 
to_sfixed(170.0/65536.0,1,-nbitq), 
to_sfixed(-72.0/65536.0,1,-nbitq), 
to_sfixed(-3287.0/65536.0,1,-nbitq), 
to_sfixed(-2359.0/65536.0,1,-nbitq), 
to_sfixed(-1566.0/65536.0,1,-nbitq), 
to_sfixed(-2525.0/65536.0,1,-nbitq), 
to_sfixed(-3263.0/65536.0,1,-nbitq), 
to_sfixed(5753.0/65536.0,1,-nbitq), 
to_sfixed(553.0/65536.0,1,-nbitq), 
to_sfixed(4.0/65536.0,1,-nbitq), 
to_sfixed(849.0/65536.0,1,-nbitq), 
to_sfixed(333.0/65536.0,1,-nbitq), 
to_sfixed(668.0/65536.0,1,-nbitq), 
to_sfixed(1859.0/65536.0,1,-nbitq), 
to_sfixed(2554.0/65536.0,1,-nbitq), 
to_sfixed(-402.0/65536.0,1,-nbitq), 
to_sfixed(4176.0/65536.0,1,-nbitq), 
to_sfixed(-6003.0/65536.0,1,-nbitq), 
to_sfixed(-1553.0/65536.0,1,-nbitq), 
to_sfixed(-1023.0/65536.0,1,-nbitq), 
to_sfixed(1914.0/65536.0,1,-nbitq), 
to_sfixed(-552.0/65536.0,1,-nbitq), 
to_sfixed(2669.0/65536.0,1,-nbitq), 
to_sfixed(4754.0/65536.0,1,-nbitq), 
to_sfixed(-1327.0/65536.0,1,-nbitq), 
to_sfixed(2291.0/65536.0,1,-nbitq), 
to_sfixed(2583.0/65536.0,1,-nbitq), 
to_sfixed(1746.0/65536.0,1,-nbitq), 
to_sfixed(323.0/65536.0,1,-nbitq), 
to_sfixed(-533.0/65536.0,1,-nbitq), 
to_sfixed(2850.0/65536.0,1,-nbitq), 
to_sfixed(-284.0/65536.0,1,-nbitq), 
to_sfixed(1732.0/65536.0,1,-nbitq), 
to_sfixed(2274.0/65536.0,1,-nbitq), 
to_sfixed(202.0/65536.0,1,-nbitq), 
to_sfixed(3246.0/65536.0,1,-nbitq), 
to_sfixed(681.0/65536.0,1,-nbitq), 
to_sfixed(-281.0/65536.0,1,-nbitq), 
to_sfixed(1423.0/65536.0,1,-nbitq), 
to_sfixed(-1827.0/65536.0,1,-nbitq), 
to_sfixed(-1152.0/65536.0,1,-nbitq), 
to_sfixed(392.0/65536.0,1,-nbitq), 
to_sfixed(1381.0/65536.0,1,-nbitq), 
to_sfixed(1989.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-233.0/65536.0,1,-nbitq), 
to_sfixed(1417.0/65536.0,1,-nbitq), 
to_sfixed(-162.0/65536.0,1,-nbitq), 
to_sfixed(1675.0/65536.0,1,-nbitq), 
to_sfixed(-1025.0/65536.0,1,-nbitq), 
to_sfixed(-2122.0/65536.0,1,-nbitq), 
to_sfixed(714.0/65536.0,1,-nbitq), 
to_sfixed(-609.0/65536.0,1,-nbitq), 
to_sfixed(-1606.0/65536.0,1,-nbitq), 
to_sfixed(-1845.0/65536.0,1,-nbitq), 
to_sfixed(-56.0/65536.0,1,-nbitq), 
to_sfixed(-1064.0/65536.0,1,-nbitq), 
to_sfixed(1627.0/65536.0,1,-nbitq), 
to_sfixed(-2071.0/65536.0,1,-nbitq), 
to_sfixed(-1676.0/65536.0,1,-nbitq), 
to_sfixed(-160.0/65536.0,1,-nbitq), 
to_sfixed(-247.0/65536.0,1,-nbitq), 
to_sfixed(2873.0/65536.0,1,-nbitq), 
to_sfixed(-949.0/65536.0,1,-nbitq), 
to_sfixed(-2230.0/65536.0,1,-nbitq), 
to_sfixed(-780.0/65536.0,1,-nbitq), 
to_sfixed(-2690.0/65536.0,1,-nbitq), 
to_sfixed(-1836.0/65536.0,1,-nbitq), 
to_sfixed(2682.0/65536.0,1,-nbitq), 
to_sfixed(36.0/65536.0,1,-nbitq), 
to_sfixed(1375.0/65536.0,1,-nbitq), 
to_sfixed(-287.0/65536.0,1,-nbitq), 
to_sfixed(1866.0/65536.0,1,-nbitq), 
to_sfixed(-1941.0/65536.0,1,-nbitq), 
to_sfixed(-2144.0/65536.0,1,-nbitq), 
to_sfixed(-526.0/65536.0,1,-nbitq), 
to_sfixed(3097.0/65536.0,1,-nbitq), 
to_sfixed(68.0/65536.0,1,-nbitq), 
to_sfixed(-246.0/65536.0,1,-nbitq), 
to_sfixed(889.0/65536.0,1,-nbitq), 
to_sfixed(-2577.0/65536.0,1,-nbitq), 
to_sfixed(-3321.0/65536.0,1,-nbitq), 
to_sfixed(-2368.0/65536.0,1,-nbitq), 
to_sfixed(-4366.0/65536.0,1,-nbitq), 
to_sfixed(1534.0/65536.0,1,-nbitq), 
to_sfixed(-2358.0/65536.0,1,-nbitq), 
to_sfixed(534.0/65536.0,1,-nbitq), 
to_sfixed(-578.0/65536.0,1,-nbitq), 
to_sfixed(1866.0/65536.0,1,-nbitq), 
to_sfixed(-376.0/65536.0,1,-nbitq), 
to_sfixed(3726.0/65536.0,1,-nbitq), 
to_sfixed(-699.0/65536.0,1,-nbitq), 
to_sfixed(-1416.0/65536.0,1,-nbitq), 
to_sfixed(2084.0/65536.0,1,-nbitq), 
to_sfixed(1642.0/65536.0,1,-nbitq), 
to_sfixed(-1009.0/65536.0,1,-nbitq), 
to_sfixed(1744.0/65536.0,1,-nbitq), 
to_sfixed(81.0/65536.0,1,-nbitq), 
to_sfixed(182.0/65536.0,1,-nbitq), 
to_sfixed(-857.0/65536.0,1,-nbitq), 
to_sfixed(-2314.0/65536.0,1,-nbitq), 
to_sfixed(-2415.0/65536.0,1,-nbitq), 
to_sfixed(1826.0/65536.0,1,-nbitq), 
to_sfixed(1754.0/65536.0,1,-nbitq), 
to_sfixed(4398.0/65536.0,1,-nbitq), 
to_sfixed(1189.0/65536.0,1,-nbitq), 
to_sfixed(2495.0/65536.0,1,-nbitq), 
to_sfixed(-34.0/65536.0,1,-nbitq), 
to_sfixed(1355.0/65536.0,1,-nbitq), 
to_sfixed(1291.0/65536.0,1,-nbitq), 
to_sfixed(3582.0/65536.0,1,-nbitq), 
to_sfixed(-1726.0/65536.0,1,-nbitq), 
to_sfixed(1331.0/65536.0,1,-nbitq), 
to_sfixed(2276.0/65536.0,1,-nbitq), 
to_sfixed(-1606.0/65536.0,1,-nbitq), 
to_sfixed(-121.0/65536.0,1,-nbitq), 
to_sfixed(-340.0/65536.0,1,-nbitq), 
to_sfixed(-907.0/65536.0,1,-nbitq), 
to_sfixed(681.0/65536.0,1,-nbitq), 
to_sfixed(923.0/65536.0,1,-nbitq), 
to_sfixed(1110.0/65536.0,1,-nbitq), 
to_sfixed(-1497.0/65536.0,1,-nbitq), 
to_sfixed(1342.0/65536.0,1,-nbitq), 
to_sfixed(-1108.0/65536.0,1,-nbitq), 
to_sfixed(477.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1453.0/65536.0,1,-nbitq), 
to_sfixed(1271.0/65536.0,1,-nbitq), 
to_sfixed(281.0/65536.0,1,-nbitq), 
to_sfixed(162.0/65536.0,1,-nbitq), 
to_sfixed(-2041.0/65536.0,1,-nbitq), 
to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(1894.0/65536.0,1,-nbitq), 
to_sfixed(671.0/65536.0,1,-nbitq), 
to_sfixed(-3092.0/65536.0,1,-nbitq), 
to_sfixed(-1560.0/65536.0,1,-nbitq), 
to_sfixed(1173.0/65536.0,1,-nbitq), 
to_sfixed(-1779.0/65536.0,1,-nbitq), 
to_sfixed(715.0/65536.0,1,-nbitq), 
to_sfixed(908.0/65536.0,1,-nbitq), 
to_sfixed(-1508.0/65536.0,1,-nbitq), 
to_sfixed(536.0/65536.0,1,-nbitq), 
to_sfixed(-1779.0/65536.0,1,-nbitq), 
to_sfixed(-1727.0/65536.0,1,-nbitq), 
to_sfixed(2937.0/65536.0,1,-nbitq), 
to_sfixed(-2411.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(-1337.0/65536.0,1,-nbitq), 
to_sfixed(-1441.0/65536.0,1,-nbitq), 
to_sfixed(2489.0/65536.0,1,-nbitq), 
to_sfixed(2422.0/65536.0,1,-nbitq), 
to_sfixed(-2052.0/65536.0,1,-nbitq), 
to_sfixed(-393.0/65536.0,1,-nbitq), 
to_sfixed(1824.0/65536.0,1,-nbitq), 
to_sfixed(1159.0/65536.0,1,-nbitq), 
to_sfixed(1894.0/65536.0,1,-nbitq), 
to_sfixed(-1134.0/65536.0,1,-nbitq), 
to_sfixed(606.0/65536.0,1,-nbitq), 
to_sfixed(-887.0/65536.0,1,-nbitq), 
to_sfixed(-2074.0/65536.0,1,-nbitq), 
to_sfixed(2770.0/65536.0,1,-nbitq), 
to_sfixed(2407.0/65536.0,1,-nbitq), 
to_sfixed(2395.0/65536.0,1,-nbitq), 
to_sfixed(-3336.0/65536.0,1,-nbitq), 
to_sfixed(-1628.0/65536.0,1,-nbitq), 
to_sfixed(-968.0/65536.0,1,-nbitq), 
to_sfixed(-2629.0/65536.0,1,-nbitq), 
to_sfixed(-2512.0/65536.0,1,-nbitq), 
to_sfixed(-532.0/65536.0,1,-nbitq), 
to_sfixed(1061.0/65536.0,1,-nbitq), 
to_sfixed(3018.0/65536.0,1,-nbitq), 
to_sfixed(5205.0/65536.0,1,-nbitq), 
to_sfixed(-437.0/65536.0,1,-nbitq), 
to_sfixed(-729.0/65536.0,1,-nbitq), 
to_sfixed(-1155.0/65536.0,1,-nbitq), 
to_sfixed(1433.0/65536.0,1,-nbitq), 
to_sfixed(-978.0/65536.0,1,-nbitq), 
to_sfixed(105.0/65536.0,1,-nbitq), 
to_sfixed(994.0/65536.0,1,-nbitq), 
to_sfixed(-2950.0/65536.0,1,-nbitq), 
to_sfixed(-1388.0/65536.0,1,-nbitq), 
to_sfixed(-277.0/65536.0,1,-nbitq), 
to_sfixed(201.0/65536.0,1,-nbitq), 
to_sfixed(-844.0/65536.0,1,-nbitq), 
to_sfixed(957.0/65536.0,1,-nbitq), 
to_sfixed(2218.0/65536.0,1,-nbitq), 
to_sfixed(-710.0/65536.0,1,-nbitq), 
to_sfixed(1512.0/65536.0,1,-nbitq), 
to_sfixed(2075.0/65536.0,1,-nbitq), 
to_sfixed(1139.0/65536.0,1,-nbitq), 
to_sfixed(3359.0/65536.0,1,-nbitq), 
to_sfixed(797.0/65536.0,1,-nbitq), 
to_sfixed(1448.0/65536.0,1,-nbitq), 
to_sfixed(-768.0/65536.0,1,-nbitq), 
to_sfixed(-459.0/65536.0,1,-nbitq), 
to_sfixed(-2099.0/65536.0,1,-nbitq), 
to_sfixed(-22.0/65536.0,1,-nbitq), 
to_sfixed(-336.0/65536.0,1,-nbitq), 
to_sfixed(3051.0/65536.0,1,-nbitq), 
to_sfixed(-1687.0/65536.0,1,-nbitq), 
to_sfixed(-2935.0/65536.0,1,-nbitq), 
to_sfixed(-1521.0/65536.0,1,-nbitq), 
to_sfixed(-116.0/65536.0,1,-nbitq), 
to_sfixed(5698.0/65536.0,1,-nbitq), 
to_sfixed(961.0/65536.0,1,-nbitq), 
to_sfixed(3245.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-748.0/65536.0,1,-nbitq), 
to_sfixed(-102.0/65536.0,1,-nbitq), 
to_sfixed(3924.0/65536.0,1,-nbitq), 
to_sfixed(-1088.0/65536.0,1,-nbitq), 
to_sfixed(-3506.0/65536.0,1,-nbitq), 
to_sfixed(-3338.0/65536.0,1,-nbitq), 
to_sfixed(1036.0/65536.0,1,-nbitq), 
to_sfixed(118.0/65536.0,1,-nbitq), 
to_sfixed(-1429.0/65536.0,1,-nbitq), 
to_sfixed(1290.0/65536.0,1,-nbitq), 
to_sfixed(-3343.0/65536.0,1,-nbitq), 
to_sfixed(-4285.0/65536.0,1,-nbitq), 
to_sfixed(449.0/65536.0,1,-nbitq), 
to_sfixed(58.0/65536.0,1,-nbitq), 
to_sfixed(589.0/65536.0,1,-nbitq), 
to_sfixed(2710.0/65536.0,1,-nbitq), 
to_sfixed(728.0/65536.0,1,-nbitq), 
to_sfixed(1327.0/65536.0,1,-nbitq), 
to_sfixed(-167.0/65536.0,1,-nbitq), 
to_sfixed(-2239.0/65536.0,1,-nbitq), 
to_sfixed(100.0/65536.0,1,-nbitq), 
to_sfixed(-1876.0/65536.0,1,-nbitq), 
to_sfixed(-1038.0/65536.0,1,-nbitq), 
to_sfixed(51.0/65536.0,1,-nbitq), 
to_sfixed(195.0/65536.0,1,-nbitq), 
to_sfixed(1186.0/65536.0,1,-nbitq), 
to_sfixed(207.0/65536.0,1,-nbitq), 
to_sfixed(2296.0/65536.0,1,-nbitq), 
to_sfixed(852.0/65536.0,1,-nbitq), 
to_sfixed(1913.0/65536.0,1,-nbitq), 
to_sfixed(-1173.0/65536.0,1,-nbitq), 
to_sfixed(3056.0/65536.0,1,-nbitq), 
to_sfixed(-5588.0/65536.0,1,-nbitq), 
to_sfixed(-4362.0/65536.0,1,-nbitq), 
to_sfixed(-2945.0/65536.0,1,-nbitq), 
to_sfixed(754.0/65536.0,1,-nbitq), 
to_sfixed(2081.0/65536.0,1,-nbitq), 
to_sfixed(-635.0/65536.0,1,-nbitq), 
to_sfixed(-3363.0/65536.0,1,-nbitq), 
to_sfixed(168.0/65536.0,1,-nbitq), 
to_sfixed(-261.0/65536.0,1,-nbitq), 
to_sfixed(-2184.0/65536.0,1,-nbitq), 
to_sfixed(-3445.0/65536.0,1,-nbitq), 
to_sfixed(2208.0/65536.0,1,-nbitq), 
to_sfixed(672.0/65536.0,1,-nbitq), 
to_sfixed(687.0/65536.0,1,-nbitq), 
to_sfixed(-602.0/65536.0,1,-nbitq), 
to_sfixed(-297.0/65536.0,1,-nbitq), 
to_sfixed(1033.0/65536.0,1,-nbitq), 
to_sfixed(-1156.0/65536.0,1,-nbitq), 
to_sfixed(865.0/65536.0,1,-nbitq), 
to_sfixed(3015.0/65536.0,1,-nbitq), 
to_sfixed(-1690.0/65536.0,1,-nbitq), 
to_sfixed(111.0/65536.0,1,-nbitq), 
to_sfixed(3633.0/65536.0,1,-nbitq), 
to_sfixed(922.0/65536.0,1,-nbitq), 
to_sfixed(1464.0/65536.0,1,-nbitq), 
to_sfixed(-897.0/65536.0,1,-nbitq), 
to_sfixed(-415.0/65536.0,1,-nbitq), 
to_sfixed(12.0/65536.0,1,-nbitq), 
to_sfixed(-1071.0/65536.0,1,-nbitq), 
to_sfixed(-1014.0/65536.0,1,-nbitq), 
to_sfixed(-1123.0/65536.0,1,-nbitq), 
to_sfixed(1525.0/65536.0,1,-nbitq), 
to_sfixed(1136.0/65536.0,1,-nbitq), 
to_sfixed(2694.0/65536.0,1,-nbitq), 
to_sfixed(2717.0/65536.0,1,-nbitq), 
to_sfixed(-2795.0/65536.0,1,-nbitq), 
to_sfixed(-673.0/65536.0,1,-nbitq), 
to_sfixed(-3113.0/65536.0,1,-nbitq), 
to_sfixed(224.0/65536.0,1,-nbitq), 
to_sfixed(-24.0/65536.0,1,-nbitq), 
to_sfixed(3877.0/65536.0,1,-nbitq), 
to_sfixed(-795.0/65536.0,1,-nbitq), 
to_sfixed(-2249.0/65536.0,1,-nbitq), 
to_sfixed(485.0/65536.0,1,-nbitq), 
to_sfixed(2218.0/65536.0,1,-nbitq), 
to_sfixed(3826.0/65536.0,1,-nbitq), 
to_sfixed(-815.0/65536.0,1,-nbitq), 
to_sfixed(838.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1674.0/65536.0,1,-nbitq), 
to_sfixed(3010.0/65536.0,1,-nbitq), 
to_sfixed(921.0/65536.0,1,-nbitq), 
to_sfixed(-3189.0/65536.0,1,-nbitq), 
to_sfixed(-3460.0/65536.0,1,-nbitq), 
to_sfixed(-1279.0/65536.0,1,-nbitq), 
to_sfixed(-1667.0/65536.0,1,-nbitq), 
to_sfixed(-1666.0/65536.0,1,-nbitq), 
to_sfixed(-2019.0/65536.0,1,-nbitq), 
to_sfixed(-798.0/65536.0,1,-nbitq), 
to_sfixed(-2091.0/65536.0,1,-nbitq), 
to_sfixed(-1524.0/65536.0,1,-nbitq), 
to_sfixed(-1690.0/65536.0,1,-nbitq), 
to_sfixed(-4496.0/65536.0,1,-nbitq), 
to_sfixed(1419.0/65536.0,1,-nbitq), 
to_sfixed(-1887.0/65536.0,1,-nbitq), 
to_sfixed(1735.0/65536.0,1,-nbitq), 
to_sfixed(-356.0/65536.0,1,-nbitq), 
to_sfixed(53.0/65536.0,1,-nbitq), 
to_sfixed(1962.0/65536.0,1,-nbitq), 
to_sfixed(520.0/65536.0,1,-nbitq), 
to_sfixed(-1331.0/65536.0,1,-nbitq), 
to_sfixed(-2446.0/65536.0,1,-nbitq), 
to_sfixed(-1512.0/65536.0,1,-nbitq), 
to_sfixed(755.0/65536.0,1,-nbitq), 
to_sfixed(2850.0/65536.0,1,-nbitq), 
to_sfixed(-1116.0/65536.0,1,-nbitq), 
to_sfixed(-2599.0/65536.0,1,-nbitq), 
to_sfixed(509.0/65536.0,1,-nbitq), 
to_sfixed(1555.0/65536.0,1,-nbitq), 
to_sfixed(-1731.0/65536.0,1,-nbitq), 
to_sfixed(2177.0/65536.0,1,-nbitq), 
to_sfixed(-4472.0/65536.0,1,-nbitq), 
to_sfixed(-653.0/65536.0,1,-nbitq), 
to_sfixed(2179.0/65536.0,1,-nbitq), 
to_sfixed(-67.0/65536.0,1,-nbitq), 
to_sfixed(-647.0/65536.0,1,-nbitq), 
to_sfixed(822.0/65536.0,1,-nbitq), 
to_sfixed(-3981.0/65536.0,1,-nbitq), 
to_sfixed(182.0/65536.0,1,-nbitq), 
to_sfixed(23.0/65536.0,1,-nbitq), 
to_sfixed(1130.0/65536.0,1,-nbitq), 
to_sfixed(-3735.0/65536.0,1,-nbitq), 
to_sfixed(-1982.0/65536.0,1,-nbitq), 
to_sfixed(-1814.0/65536.0,1,-nbitq), 
to_sfixed(4464.0/65536.0,1,-nbitq), 
to_sfixed(2898.0/65536.0,1,-nbitq), 
to_sfixed(-519.0/65536.0,1,-nbitq), 
to_sfixed(3523.0/65536.0,1,-nbitq), 
to_sfixed(655.0/65536.0,1,-nbitq), 
to_sfixed(-1744.0/65536.0,1,-nbitq), 
to_sfixed(-149.0/65536.0,1,-nbitq), 
to_sfixed(826.0/65536.0,1,-nbitq), 
to_sfixed(-155.0/65536.0,1,-nbitq), 
to_sfixed(1412.0/65536.0,1,-nbitq), 
to_sfixed(-841.0/65536.0,1,-nbitq), 
to_sfixed(-1877.0/65536.0,1,-nbitq), 
to_sfixed(-1838.0/65536.0,1,-nbitq), 
to_sfixed(-2476.0/65536.0,1,-nbitq), 
to_sfixed(3914.0/65536.0,1,-nbitq), 
to_sfixed(-1319.0/65536.0,1,-nbitq), 
to_sfixed(-2473.0/65536.0,1,-nbitq), 
to_sfixed(1382.0/65536.0,1,-nbitq), 
to_sfixed(-2343.0/65536.0,1,-nbitq), 
to_sfixed(3266.0/65536.0,1,-nbitq), 
to_sfixed(858.0/65536.0,1,-nbitq), 
to_sfixed(801.0/65536.0,1,-nbitq), 
to_sfixed(-3751.0/65536.0,1,-nbitq), 
to_sfixed(3221.0/65536.0,1,-nbitq), 
to_sfixed(420.0/65536.0,1,-nbitq), 
to_sfixed(692.0/65536.0,1,-nbitq), 
to_sfixed(2.0/65536.0,1,-nbitq), 
to_sfixed(2705.0/65536.0,1,-nbitq), 
to_sfixed(-2843.0/65536.0,1,-nbitq), 
to_sfixed(294.0/65536.0,1,-nbitq), 
to_sfixed(3321.0/65536.0,1,-nbitq), 
to_sfixed(-2088.0/65536.0,1,-nbitq), 
to_sfixed(3493.0/65536.0,1,-nbitq), 
to_sfixed(-1364.0/65536.0,1,-nbitq), 
to_sfixed(3297.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1814.0/65536.0,1,-nbitq), 
to_sfixed(1936.0/65536.0,1,-nbitq), 
to_sfixed(3754.0/65536.0,1,-nbitq), 
to_sfixed(2205.0/65536.0,1,-nbitq), 
to_sfixed(-1925.0/65536.0,1,-nbitq), 
to_sfixed(-1974.0/65536.0,1,-nbitq), 
to_sfixed(532.0/65536.0,1,-nbitq), 
to_sfixed(1543.0/65536.0,1,-nbitq), 
to_sfixed(-4718.0/65536.0,1,-nbitq), 
to_sfixed(-1743.0/65536.0,1,-nbitq), 
to_sfixed(1667.0/65536.0,1,-nbitq), 
to_sfixed(785.0/65536.0,1,-nbitq), 
to_sfixed(-406.0/65536.0,1,-nbitq), 
to_sfixed(-545.0/65536.0,1,-nbitq), 
to_sfixed(3109.0/65536.0,1,-nbitq), 
to_sfixed(1251.0/65536.0,1,-nbitq), 
to_sfixed(-921.0/65536.0,1,-nbitq), 
to_sfixed(-750.0/65536.0,1,-nbitq), 
to_sfixed(90.0/65536.0,1,-nbitq), 
to_sfixed(1529.0/65536.0,1,-nbitq), 
to_sfixed(-845.0/65536.0,1,-nbitq), 
to_sfixed(3126.0/65536.0,1,-nbitq), 
to_sfixed(-1250.0/65536.0,1,-nbitq), 
to_sfixed(-722.0/65536.0,1,-nbitq), 
to_sfixed(2479.0/65536.0,1,-nbitq), 
to_sfixed(1053.0/65536.0,1,-nbitq), 
to_sfixed(357.0/65536.0,1,-nbitq), 
to_sfixed(-2844.0/65536.0,1,-nbitq), 
to_sfixed(-1354.0/65536.0,1,-nbitq), 
to_sfixed(-3296.0/65536.0,1,-nbitq), 
to_sfixed(989.0/65536.0,1,-nbitq), 
to_sfixed(1242.0/65536.0,1,-nbitq), 
to_sfixed(-285.0/65536.0,1,-nbitq), 
to_sfixed(-1701.0/65536.0,1,-nbitq), 
to_sfixed(1185.0/65536.0,1,-nbitq), 
to_sfixed(1864.0/65536.0,1,-nbitq), 
to_sfixed(-701.0/65536.0,1,-nbitq), 
to_sfixed(-1842.0/65536.0,1,-nbitq), 
to_sfixed(351.0/65536.0,1,-nbitq), 
to_sfixed(2033.0/65536.0,1,-nbitq), 
to_sfixed(-2401.0/65536.0,1,-nbitq), 
to_sfixed(-3179.0/65536.0,1,-nbitq), 
to_sfixed(-4568.0/65536.0,1,-nbitq), 
to_sfixed(-469.0/65536.0,1,-nbitq), 
to_sfixed(-1640.0/65536.0,1,-nbitq), 
to_sfixed(3574.0/65536.0,1,-nbitq), 
to_sfixed(-2646.0/65536.0,1,-nbitq), 
to_sfixed(-162.0/65536.0,1,-nbitq), 
to_sfixed(1644.0/65536.0,1,-nbitq), 
to_sfixed(-977.0/65536.0,1,-nbitq), 
to_sfixed(-1155.0/65536.0,1,-nbitq), 
to_sfixed(-646.0/65536.0,1,-nbitq), 
to_sfixed(-1049.0/65536.0,1,-nbitq), 
to_sfixed(-2899.0/65536.0,1,-nbitq), 
to_sfixed(2958.0/65536.0,1,-nbitq), 
to_sfixed(-888.0/65536.0,1,-nbitq), 
to_sfixed(1790.0/65536.0,1,-nbitq), 
to_sfixed(401.0/65536.0,1,-nbitq), 
to_sfixed(36.0/65536.0,1,-nbitq), 
to_sfixed(4082.0/65536.0,1,-nbitq), 
to_sfixed(662.0/65536.0,1,-nbitq), 
to_sfixed(2132.0/65536.0,1,-nbitq), 
to_sfixed(-2026.0/65536.0,1,-nbitq), 
to_sfixed(1382.0/65536.0,1,-nbitq), 
to_sfixed(38.0/65536.0,1,-nbitq), 
to_sfixed(-2362.0/65536.0,1,-nbitq), 
to_sfixed(-1689.0/65536.0,1,-nbitq), 
to_sfixed(-4327.0/65536.0,1,-nbitq), 
to_sfixed(-654.0/65536.0,1,-nbitq), 
to_sfixed(2858.0/65536.0,1,-nbitq), 
to_sfixed(-1044.0/65536.0,1,-nbitq), 
to_sfixed(3451.0/65536.0,1,-nbitq), 
to_sfixed(2167.0/65536.0,1,-nbitq), 
to_sfixed(1912.0/65536.0,1,-nbitq), 
to_sfixed(-1072.0/65536.0,1,-nbitq), 
to_sfixed(-627.0/65536.0,1,-nbitq), 
to_sfixed(-3921.0/65536.0,1,-nbitq), 
to_sfixed(2583.0/65536.0,1,-nbitq), 
to_sfixed(-1663.0/65536.0,1,-nbitq), 
to_sfixed(1805.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3430.0/65536.0,1,-nbitq), 
to_sfixed(754.0/65536.0,1,-nbitq), 
to_sfixed(4832.0/65536.0,1,-nbitq), 
to_sfixed(1350.0/65536.0,1,-nbitq), 
to_sfixed(-4022.0/65536.0,1,-nbitq), 
to_sfixed(-1414.0/65536.0,1,-nbitq), 
to_sfixed(-1025.0/65536.0,1,-nbitq), 
to_sfixed(-3065.0/65536.0,1,-nbitq), 
to_sfixed(-455.0/65536.0,1,-nbitq), 
to_sfixed(-407.0/65536.0,1,-nbitq), 
to_sfixed(-836.0/65536.0,1,-nbitq), 
to_sfixed(-38.0/65536.0,1,-nbitq), 
to_sfixed(-2163.0/65536.0,1,-nbitq), 
to_sfixed(-3197.0/65536.0,1,-nbitq), 
to_sfixed(-2409.0/65536.0,1,-nbitq), 
to_sfixed(-529.0/65536.0,1,-nbitq), 
to_sfixed(1243.0/65536.0,1,-nbitq), 
to_sfixed(-3434.0/65536.0,1,-nbitq), 
to_sfixed(1109.0/65536.0,1,-nbitq), 
to_sfixed(-812.0/65536.0,1,-nbitq), 
to_sfixed(-80.0/65536.0,1,-nbitq), 
to_sfixed(-1655.0/65536.0,1,-nbitq), 
to_sfixed(-749.0/65536.0,1,-nbitq), 
to_sfixed(-3214.0/65536.0,1,-nbitq), 
to_sfixed(-1552.0/65536.0,1,-nbitq), 
to_sfixed(-1390.0/65536.0,1,-nbitq), 
to_sfixed(-1776.0/65536.0,1,-nbitq), 
to_sfixed(-2496.0/65536.0,1,-nbitq), 
to_sfixed(-3144.0/65536.0,1,-nbitq), 
to_sfixed(782.0/65536.0,1,-nbitq), 
to_sfixed(-423.0/65536.0,1,-nbitq), 
to_sfixed(-2881.0/65536.0,1,-nbitq), 
to_sfixed(-3348.0/65536.0,1,-nbitq), 
to_sfixed(-1787.0/65536.0,1,-nbitq), 
to_sfixed(2047.0/65536.0,1,-nbitq), 
to_sfixed(-1334.0/65536.0,1,-nbitq), 
to_sfixed(2119.0/65536.0,1,-nbitq), 
to_sfixed(-1163.0/65536.0,1,-nbitq), 
to_sfixed(-3836.0/65536.0,1,-nbitq), 
to_sfixed(-1368.0/65536.0,1,-nbitq), 
to_sfixed(422.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(-4149.0/65536.0,1,-nbitq), 
to_sfixed(693.0/65536.0,1,-nbitq), 
to_sfixed(1998.0/65536.0,1,-nbitq), 
to_sfixed(3326.0/65536.0,1,-nbitq), 
to_sfixed(-1892.0/65536.0,1,-nbitq), 
to_sfixed(1074.0/65536.0,1,-nbitq), 
to_sfixed(-2.0/65536.0,1,-nbitq), 
to_sfixed(741.0/65536.0,1,-nbitq), 
to_sfixed(1638.0/65536.0,1,-nbitq), 
to_sfixed(203.0/65536.0,1,-nbitq), 
to_sfixed(-1614.0/65536.0,1,-nbitq), 
to_sfixed(-4433.0/65536.0,1,-nbitq), 
to_sfixed(1602.0/65536.0,1,-nbitq), 
to_sfixed(-59.0/65536.0,1,-nbitq), 
to_sfixed(2694.0/65536.0,1,-nbitq), 
to_sfixed(-2404.0/65536.0,1,-nbitq), 
to_sfixed(-1026.0/65536.0,1,-nbitq), 
to_sfixed(2918.0/65536.0,1,-nbitq), 
to_sfixed(-3057.0/65536.0,1,-nbitq), 
to_sfixed(2139.0/65536.0,1,-nbitq), 
to_sfixed(967.0/65536.0,1,-nbitq), 
to_sfixed(2052.0/65536.0,1,-nbitq), 
to_sfixed(2968.0/65536.0,1,-nbitq), 
to_sfixed(-3392.0/65536.0,1,-nbitq), 
to_sfixed(-580.0/65536.0,1,-nbitq), 
to_sfixed(-5429.0/65536.0,1,-nbitq), 
to_sfixed(2636.0/65536.0,1,-nbitq), 
to_sfixed(-2275.0/65536.0,1,-nbitq), 
to_sfixed(1407.0/65536.0,1,-nbitq), 
to_sfixed(-33.0/65536.0,1,-nbitq), 
to_sfixed(93.0/65536.0,1,-nbitq), 
to_sfixed(-208.0/65536.0,1,-nbitq), 
to_sfixed(958.0/65536.0,1,-nbitq), 
to_sfixed(2545.0/65536.0,1,-nbitq), 
to_sfixed(-3548.0/65536.0,1,-nbitq), 
to_sfixed(797.0/65536.0,1,-nbitq), 
to_sfixed(-1137.0/65536.0,1,-nbitq), 
to_sfixed(4372.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1721.0/65536.0,1,-nbitq), 
to_sfixed(2198.0/65536.0,1,-nbitq), 
to_sfixed(4077.0/65536.0,1,-nbitq), 
to_sfixed(694.0/65536.0,1,-nbitq), 
to_sfixed(-1683.0/65536.0,1,-nbitq), 
to_sfixed(-294.0/65536.0,1,-nbitq), 
to_sfixed(2223.0/65536.0,1,-nbitq), 
to_sfixed(805.0/65536.0,1,-nbitq), 
to_sfixed(3844.0/65536.0,1,-nbitq), 
to_sfixed(-2597.0/65536.0,1,-nbitq), 
to_sfixed(-99.0/65536.0,1,-nbitq), 
to_sfixed(-4178.0/65536.0,1,-nbitq), 
to_sfixed(849.0/65536.0,1,-nbitq), 
to_sfixed(-645.0/65536.0,1,-nbitq), 
to_sfixed(-588.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(-2206.0/65536.0,1,-nbitq), 
to_sfixed(-1707.0/65536.0,1,-nbitq), 
to_sfixed(1210.0/65536.0,1,-nbitq), 
to_sfixed(1677.0/65536.0,1,-nbitq), 
to_sfixed(-1982.0/65536.0,1,-nbitq), 
to_sfixed(-1298.0/65536.0,1,-nbitq), 
to_sfixed(2949.0/65536.0,1,-nbitq), 
to_sfixed(-683.0/65536.0,1,-nbitq), 
to_sfixed(-2505.0/65536.0,1,-nbitq), 
to_sfixed(444.0/65536.0,1,-nbitq), 
to_sfixed(-4604.0/65536.0,1,-nbitq), 
to_sfixed(517.0/65536.0,1,-nbitq), 
to_sfixed(-1889.0/65536.0,1,-nbitq), 
to_sfixed(-1286.0/65536.0,1,-nbitq), 
to_sfixed(-1932.0/65536.0,1,-nbitq), 
to_sfixed(1444.0/65536.0,1,-nbitq), 
to_sfixed(-3843.0/65536.0,1,-nbitq), 
to_sfixed(-1434.0/65536.0,1,-nbitq), 
to_sfixed(-1257.0/65536.0,1,-nbitq), 
to_sfixed(-2691.0/65536.0,1,-nbitq), 
to_sfixed(1837.0/65536.0,1,-nbitq), 
to_sfixed(-1963.0/65536.0,1,-nbitq), 
to_sfixed(1123.0/65536.0,1,-nbitq), 
to_sfixed(34.0/65536.0,1,-nbitq), 
to_sfixed(-753.0/65536.0,1,-nbitq), 
to_sfixed(-2965.0/65536.0,1,-nbitq), 
to_sfixed(-4581.0/65536.0,1,-nbitq), 
to_sfixed(3586.0/65536.0,1,-nbitq), 
to_sfixed(-208.0/65536.0,1,-nbitq), 
to_sfixed(4598.0/65536.0,1,-nbitq), 
to_sfixed(-2397.0/65536.0,1,-nbitq), 
to_sfixed(-746.0/65536.0,1,-nbitq), 
to_sfixed(753.0/65536.0,1,-nbitq), 
to_sfixed(-1210.0/65536.0,1,-nbitq), 
to_sfixed(657.0/65536.0,1,-nbitq), 
to_sfixed(2917.0/65536.0,1,-nbitq), 
to_sfixed(176.0/65536.0,1,-nbitq), 
to_sfixed(-4867.0/65536.0,1,-nbitq), 
to_sfixed(-2008.0/65536.0,1,-nbitq), 
to_sfixed(1037.0/65536.0,1,-nbitq), 
to_sfixed(-2697.0/65536.0,1,-nbitq), 
to_sfixed(-984.0/65536.0,1,-nbitq), 
to_sfixed(2684.0/65536.0,1,-nbitq), 
to_sfixed(3532.0/65536.0,1,-nbitq), 
to_sfixed(-2533.0/65536.0,1,-nbitq), 
to_sfixed(826.0/65536.0,1,-nbitq), 
to_sfixed(-2017.0/65536.0,1,-nbitq), 
to_sfixed(379.0/65536.0,1,-nbitq), 
to_sfixed(4393.0/65536.0,1,-nbitq), 
to_sfixed(2073.0/65536.0,1,-nbitq), 
to_sfixed(141.0/65536.0,1,-nbitq), 
to_sfixed(-3660.0/65536.0,1,-nbitq), 
to_sfixed(2007.0/65536.0,1,-nbitq), 
to_sfixed(495.0/65536.0,1,-nbitq), 
to_sfixed(-34.0/65536.0,1,-nbitq), 
to_sfixed(-352.0/65536.0,1,-nbitq), 
to_sfixed(-219.0/65536.0,1,-nbitq), 
to_sfixed(-2824.0/65536.0,1,-nbitq), 
to_sfixed(-604.0/65536.0,1,-nbitq), 
to_sfixed(-3036.0/65536.0,1,-nbitq), 
to_sfixed(-2849.0/65536.0,1,-nbitq), 
to_sfixed(4277.0/65536.0,1,-nbitq), 
to_sfixed(-155.0/65536.0,1,-nbitq), 
to_sfixed(5857.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2786.0/65536.0,1,-nbitq), 
to_sfixed(4648.0/65536.0,1,-nbitq), 
to_sfixed(-1195.0/65536.0,1,-nbitq), 
to_sfixed(-1419.0/65536.0,1,-nbitq), 
to_sfixed(1633.0/65536.0,1,-nbitq), 
to_sfixed(-1453.0/65536.0,1,-nbitq), 
to_sfixed(462.0/65536.0,1,-nbitq), 
to_sfixed(-1546.0/65536.0,1,-nbitq), 
to_sfixed(348.0/65536.0,1,-nbitq), 
to_sfixed(-1378.0/65536.0,1,-nbitq), 
to_sfixed(-2829.0/65536.0,1,-nbitq), 
to_sfixed(-6090.0/65536.0,1,-nbitq), 
to_sfixed(-1979.0/65536.0,1,-nbitq), 
to_sfixed(-1803.0/65536.0,1,-nbitq), 
to_sfixed(2746.0/65536.0,1,-nbitq), 
to_sfixed(-1535.0/65536.0,1,-nbitq), 
to_sfixed(1117.0/65536.0,1,-nbitq), 
to_sfixed(-4088.0/65536.0,1,-nbitq), 
to_sfixed(-505.0/65536.0,1,-nbitq), 
to_sfixed(1398.0/65536.0,1,-nbitq), 
to_sfixed(-1876.0/65536.0,1,-nbitq), 
to_sfixed(-1469.0/65536.0,1,-nbitq), 
to_sfixed(-614.0/65536.0,1,-nbitq), 
to_sfixed(-1809.0/65536.0,1,-nbitq), 
to_sfixed(-1566.0/65536.0,1,-nbitq), 
to_sfixed(-753.0/65536.0,1,-nbitq), 
to_sfixed(-1750.0/65536.0,1,-nbitq), 
to_sfixed(-1116.0/65536.0,1,-nbitq), 
to_sfixed(-3350.0/65536.0,1,-nbitq), 
to_sfixed(-1051.0/65536.0,1,-nbitq), 
to_sfixed(129.0/65536.0,1,-nbitq), 
to_sfixed(3066.0/65536.0,1,-nbitq), 
to_sfixed(-3181.0/65536.0,1,-nbitq), 
to_sfixed(929.0/65536.0,1,-nbitq), 
to_sfixed(2159.0/65536.0,1,-nbitq), 
to_sfixed(199.0/65536.0,1,-nbitq), 
to_sfixed(1037.0/65536.0,1,-nbitq), 
to_sfixed(1001.0/65536.0,1,-nbitq), 
to_sfixed(-824.0/65536.0,1,-nbitq), 
to_sfixed(-1720.0/65536.0,1,-nbitq), 
to_sfixed(3231.0/65536.0,1,-nbitq), 
to_sfixed(664.0/65536.0,1,-nbitq), 
to_sfixed(751.0/65536.0,1,-nbitq), 
to_sfixed(2373.0/65536.0,1,-nbitq), 
to_sfixed(-1812.0/65536.0,1,-nbitq), 
to_sfixed(3732.0/65536.0,1,-nbitq), 
to_sfixed(2326.0/65536.0,1,-nbitq), 
to_sfixed(-1334.0/65536.0,1,-nbitq), 
to_sfixed(2402.0/65536.0,1,-nbitq), 
to_sfixed(367.0/65536.0,1,-nbitq), 
to_sfixed(-371.0/65536.0,1,-nbitq), 
to_sfixed(1900.0/65536.0,1,-nbitq), 
to_sfixed(-527.0/65536.0,1,-nbitq), 
to_sfixed(234.0/65536.0,1,-nbitq), 
to_sfixed(-2775.0/65536.0,1,-nbitq), 
to_sfixed(-2728.0/65536.0,1,-nbitq), 
to_sfixed(-2501.0/65536.0,1,-nbitq), 
to_sfixed(-242.0/65536.0,1,-nbitq), 
to_sfixed(1482.0/65536.0,1,-nbitq), 
to_sfixed(1206.0/65536.0,1,-nbitq), 
to_sfixed(-1401.0/65536.0,1,-nbitq), 
to_sfixed(1559.0/65536.0,1,-nbitq), 
to_sfixed(601.0/65536.0,1,-nbitq), 
to_sfixed(1128.0/65536.0,1,-nbitq), 
to_sfixed(-1070.0/65536.0,1,-nbitq), 
to_sfixed(-1093.0/65536.0,1,-nbitq), 
to_sfixed(353.0/65536.0,1,-nbitq), 
to_sfixed(-4220.0/65536.0,1,-nbitq), 
to_sfixed(3361.0/65536.0,1,-nbitq), 
to_sfixed(-2654.0/65536.0,1,-nbitq), 
to_sfixed(9.0/65536.0,1,-nbitq), 
to_sfixed(-2530.0/65536.0,1,-nbitq), 
to_sfixed(1244.0/65536.0,1,-nbitq), 
to_sfixed(2647.0/65536.0,1,-nbitq), 
to_sfixed(-2454.0/65536.0,1,-nbitq), 
to_sfixed(2427.0/65536.0,1,-nbitq), 
to_sfixed(-6223.0/65536.0,1,-nbitq), 
to_sfixed(-750.0/65536.0,1,-nbitq), 
to_sfixed(628.0/65536.0,1,-nbitq), 
to_sfixed(536.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2663.0/65536.0,1,-nbitq), 
to_sfixed(3739.0/65536.0,1,-nbitq), 
to_sfixed(-4436.0/65536.0,1,-nbitq), 
to_sfixed(4169.0/65536.0,1,-nbitq), 
to_sfixed(-2047.0/65536.0,1,-nbitq), 
to_sfixed(-5192.0/65536.0,1,-nbitq), 
to_sfixed(4484.0/65536.0,1,-nbitq), 
to_sfixed(3872.0/65536.0,1,-nbitq), 
to_sfixed(848.0/65536.0,1,-nbitq), 
to_sfixed(975.0/65536.0,1,-nbitq), 
to_sfixed(158.0/65536.0,1,-nbitq), 
to_sfixed(-5956.0/65536.0,1,-nbitq), 
to_sfixed(1173.0/65536.0,1,-nbitq), 
to_sfixed(-5570.0/65536.0,1,-nbitq), 
to_sfixed(2206.0/65536.0,1,-nbitq), 
to_sfixed(-1583.0/65536.0,1,-nbitq), 
to_sfixed(1707.0/65536.0,1,-nbitq), 
to_sfixed(4460.0/65536.0,1,-nbitq), 
to_sfixed(-4251.0/65536.0,1,-nbitq), 
to_sfixed(1675.0/65536.0,1,-nbitq), 
to_sfixed(3503.0/65536.0,1,-nbitq), 
to_sfixed(3151.0/65536.0,1,-nbitq), 
to_sfixed(3260.0/65536.0,1,-nbitq), 
to_sfixed(-4415.0/65536.0,1,-nbitq), 
to_sfixed(2221.0/65536.0,1,-nbitq), 
to_sfixed(-1275.0/65536.0,1,-nbitq), 
to_sfixed(-1751.0/65536.0,1,-nbitq), 
to_sfixed(-4513.0/65536.0,1,-nbitq), 
to_sfixed(-1205.0/65536.0,1,-nbitq), 
to_sfixed(-697.0/65536.0,1,-nbitq), 
to_sfixed(-1659.0/65536.0,1,-nbitq), 
to_sfixed(2283.0/65536.0,1,-nbitq), 
to_sfixed(3955.0/65536.0,1,-nbitq), 
to_sfixed(2565.0/65536.0,1,-nbitq), 
to_sfixed(-1050.0/65536.0,1,-nbitq), 
to_sfixed(-2869.0/65536.0,1,-nbitq), 
to_sfixed(792.0/65536.0,1,-nbitq), 
to_sfixed(-2983.0/65536.0,1,-nbitq), 
to_sfixed(4297.0/65536.0,1,-nbitq), 
to_sfixed(653.0/65536.0,1,-nbitq), 
to_sfixed(-1453.0/65536.0,1,-nbitq), 
to_sfixed(-2371.0/65536.0,1,-nbitq), 
to_sfixed(2124.0/65536.0,1,-nbitq), 
to_sfixed(60.0/65536.0,1,-nbitq), 
to_sfixed(-1677.0/65536.0,1,-nbitq), 
to_sfixed(151.0/65536.0,1,-nbitq), 
to_sfixed(1919.0/65536.0,1,-nbitq), 
to_sfixed(640.0/65536.0,1,-nbitq), 
to_sfixed(-1201.0/65536.0,1,-nbitq), 
to_sfixed(680.0/65536.0,1,-nbitq), 
to_sfixed(-1474.0/65536.0,1,-nbitq), 
to_sfixed(20.0/65536.0,1,-nbitq), 
to_sfixed(-409.0/65536.0,1,-nbitq), 
to_sfixed(818.0/65536.0,1,-nbitq), 
to_sfixed(3307.0/65536.0,1,-nbitq), 
to_sfixed(-4560.0/65536.0,1,-nbitq), 
to_sfixed(-525.0/65536.0,1,-nbitq), 
to_sfixed(592.0/65536.0,1,-nbitq), 
to_sfixed(-2964.0/65536.0,1,-nbitq), 
to_sfixed(-8052.0/65536.0,1,-nbitq), 
to_sfixed(13.0/65536.0,1,-nbitq), 
to_sfixed(240.0/65536.0,1,-nbitq), 
to_sfixed(-1555.0/65536.0,1,-nbitq), 
to_sfixed(1699.0/65536.0,1,-nbitq), 
to_sfixed(-563.0/65536.0,1,-nbitq), 
to_sfixed(-1412.0/65536.0,1,-nbitq), 
to_sfixed(2606.0/65536.0,1,-nbitq), 
to_sfixed(-4625.0/65536.0,1,-nbitq), 
to_sfixed(-1830.0/65536.0,1,-nbitq), 
to_sfixed(2401.0/65536.0,1,-nbitq), 
to_sfixed(-3638.0/65536.0,1,-nbitq), 
to_sfixed(-2526.0/65536.0,1,-nbitq), 
to_sfixed(717.0/65536.0,1,-nbitq), 
to_sfixed(491.0/65536.0,1,-nbitq), 
to_sfixed(-3038.0/65536.0,1,-nbitq), 
to_sfixed(1743.0/65536.0,1,-nbitq), 
to_sfixed(-7604.0/65536.0,1,-nbitq), 
to_sfixed(1968.0/65536.0,1,-nbitq), 
to_sfixed(381.0/65536.0,1,-nbitq), 
to_sfixed(4314.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1621.0/65536.0,1,-nbitq), 
to_sfixed(6499.0/65536.0,1,-nbitq), 
to_sfixed(-4213.0/65536.0,1,-nbitq), 
to_sfixed(14.0/65536.0,1,-nbitq), 
to_sfixed(-4099.0/65536.0,1,-nbitq), 
to_sfixed(-6261.0/65536.0,1,-nbitq), 
to_sfixed(1087.0/65536.0,1,-nbitq), 
to_sfixed(513.0/65536.0,1,-nbitq), 
to_sfixed(2741.0/65536.0,1,-nbitq), 
to_sfixed(566.0/65536.0,1,-nbitq), 
to_sfixed(543.0/65536.0,1,-nbitq), 
to_sfixed(-4272.0/65536.0,1,-nbitq), 
to_sfixed(3343.0/65536.0,1,-nbitq), 
to_sfixed(-9473.0/65536.0,1,-nbitq), 
to_sfixed(-1513.0/65536.0,1,-nbitq), 
to_sfixed(2536.0/65536.0,1,-nbitq), 
to_sfixed(-1416.0/65536.0,1,-nbitq), 
to_sfixed(2961.0/65536.0,1,-nbitq), 
to_sfixed(-1573.0/65536.0,1,-nbitq), 
to_sfixed(-2125.0/65536.0,1,-nbitq), 
to_sfixed(1318.0/65536.0,1,-nbitq), 
to_sfixed(4196.0/65536.0,1,-nbitq), 
to_sfixed(7610.0/65536.0,1,-nbitq), 
to_sfixed(-7034.0/65536.0,1,-nbitq), 
to_sfixed(-2607.0/65536.0,1,-nbitq), 
to_sfixed(-1695.0/65536.0,1,-nbitq), 
to_sfixed(-1176.0/65536.0,1,-nbitq), 
to_sfixed(-207.0/65536.0,1,-nbitq), 
to_sfixed(-6199.0/65536.0,1,-nbitq), 
to_sfixed(-2839.0/65536.0,1,-nbitq), 
to_sfixed(-2017.0/65536.0,1,-nbitq), 
to_sfixed(1151.0/65536.0,1,-nbitq), 
to_sfixed(6669.0/65536.0,1,-nbitq), 
to_sfixed(5745.0/65536.0,1,-nbitq), 
to_sfixed(-1673.0/65536.0,1,-nbitq), 
to_sfixed(-2389.0/65536.0,1,-nbitq), 
to_sfixed(5885.0/65536.0,1,-nbitq), 
to_sfixed(589.0/65536.0,1,-nbitq), 
to_sfixed(4526.0/65536.0,1,-nbitq), 
to_sfixed(-1119.0/65536.0,1,-nbitq), 
to_sfixed(-529.0/65536.0,1,-nbitq), 
to_sfixed(-986.0/65536.0,1,-nbitq), 
to_sfixed(2405.0/65536.0,1,-nbitq), 
to_sfixed(-2330.0/65536.0,1,-nbitq), 
to_sfixed(-1435.0/65536.0,1,-nbitq), 
to_sfixed(-1925.0/65536.0,1,-nbitq), 
to_sfixed(798.0/65536.0,1,-nbitq), 
to_sfixed(-3458.0/65536.0,1,-nbitq), 
to_sfixed(926.0/65536.0,1,-nbitq), 
to_sfixed(3168.0/65536.0,1,-nbitq), 
to_sfixed(-1951.0/65536.0,1,-nbitq), 
to_sfixed(1338.0/65536.0,1,-nbitq), 
to_sfixed(2122.0/65536.0,1,-nbitq), 
to_sfixed(1445.0/65536.0,1,-nbitq), 
to_sfixed(4178.0/65536.0,1,-nbitq), 
to_sfixed(-5500.0/65536.0,1,-nbitq), 
to_sfixed(715.0/65536.0,1,-nbitq), 
to_sfixed(-1607.0/65536.0,1,-nbitq), 
to_sfixed(-2891.0/65536.0,1,-nbitq), 
to_sfixed(-6434.0/65536.0,1,-nbitq), 
to_sfixed(3153.0/65536.0,1,-nbitq), 
to_sfixed(111.0/65536.0,1,-nbitq), 
to_sfixed(2333.0/65536.0,1,-nbitq), 
to_sfixed(-2155.0/65536.0,1,-nbitq), 
to_sfixed(-1392.0/65536.0,1,-nbitq), 
to_sfixed(-2154.0/65536.0,1,-nbitq), 
to_sfixed(1679.0/65536.0,1,-nbitq), 
to_sfixed(-4415.0/65536.0,1,-nbitq), 
to_sfixed(2009.0/65536.0,1,-nbitq), 
to_sfixed(5485.0/65536.0,1,-nbitq), 
to_sfixed(1349.0/65536.0,1,-nbitq), 
to_sfixed(-1436.0/65536.0,1,-nbitq), 
to_sfixed(-331.0/65536.0,1,-nbitq), 
to_sfixed(-1566.0/65536.0,1,-nbitq), 
to_sfixed(-1797.0/65536.0,1,-nbitq), 
to_sfixed(-2205.0/65536.0,1,-nbitq), 
to_sfixed(-781.0/65536.0,1,-nbitq), 
to_sfixed(-664.0/65536.0,1,-nbitq), 
to_sfixed(-53.0/65536.0,1,-nbitq), 
to_sfixed(-630.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1548.0/65536.0,1,-nbitq), 
to_sfixed(1619.0/65536.0,1,-nbitq), 
to_sfixed(-5979.0/65536.0,1,-nbitq), 
to_sfixed(1060.0/65536.0,1,-nbitq), 
to_sfixed(1322.0/65536.0,1,-nbitq), 
to_sfixed(-5105.0/65536.0,1,-nbitq), 
to_sfixed(1610.0/65536.0,1,-nbitq), 
to_sfixed(3541.0/65536.0,1,-nbitq), 
to_sfixed(5715.0/65536.0,1,-nbitq), 
to_sfixed(-2907.0/65536.0,1,-nbitq), 
to_sfixed(-1962.0/65536.0,1,-nbitq), 
to_sfixed(-9243.0/65536.0,1,-nbitq), 
to_sfixed(-837.0/65536.0,1,-nbitq), 
to_sfixed(-10048.0/65536.0,1,-nbitq), 
to_sfixed(-80.0/65536.0,1,-nbitq), 
to_sfixed(-1216.0/65536.0,1,-nbitq), 
to_sfixed(2695.0/65536.0,1,-nbitq), 
to_sfixed(608.0/65536.0,1,-nbitq), 
to_sfixed(-6140.0/65536.0,1,-nbitq), 
to_sfixed(-301.0/65536.0,1,-nbitq), 
to_sfixed(1283.0/65536.0,1,-nbitq), 
to_sfixed(3783.0/65536.0,1,-nbitq), 
to_sfixed(4851.0/65536.0,1,-nbitq), 
to_sfixed(-13741.0/65536.0,1,-nbitq), 
to_sfixed(-800.0/65536.0,1,-nbitq), 
to_sfixed(-7255.0/65536.0,1,-nbitq), 
to_sfixed(-1677.0/65536.0,1,-nbitq), 
to_sfixed(-5010.0/65536.0,1,-nbitq), 
to_sfixed(-4215.0/65536.0,1,-nbitq), 
to_sfixed(-1053.0/65536.0,1,-nbitq), 
to_sfixed(-652.0/65536.0,1,-nbitq), 
to_sfixed(2604.0/65536.0,1,-nbitq), 
to_sfixed(1578.0/65536.0,1,-nbitq), 
to_sfixed(3983.0/65536.0,1,-nbitq), 
to_sfixed(1899.0/65536.0,1,-nbitq), 
to_sfixed(-1929.0/65536.0,1,-nbitq), 
to_sfixed(5742.0/65536.0,1,-nbitq), 
to_sfixed(1933.0/65536.0,1,-nbitq), 
to_sfixed(5931.0/65536.0,1,-nbitq), 
to_sfixed(2372.0/65536.0,1,-nbitq), 
to_sfixed(-4241.0/65536.0,1,-nbitq), 
to_sfixed(-3205.0/65536.0,1,-nbitq), 
to_sfixed(3782.0/65536.0,1,-nbitq), 
to_sfixed(2105.0/65536.0,1,-nbitq), 
to_sfixed(1775.0/65536.0,1,-nbitq), 
to_sfixed(-989.0/65536.0,1,-nbitq), 
to_sfixed(-2752.0/65536.0,1,-nbitq), 
to_sfixed(-751.0/65536.0,1,-nbitq), 
to_sfixed(23.0/65536.0,1,-nbitq), 
to_sfixed(1574.0/65536.0,1,-nbitq), 
to_sfixed(1857.0/65536.0,1,-nbitq), 
to_sfixed(2955.0/65536.0,1,-nbitq), 
to_sfixed(1216.0/65536.0,1,-nbitq), 
to_sfixed(-1790.0/65536.0,1,-nbitq), 
to_sfixed(1197.0/65536.0,1,-nbitq), 
to_sfixed(-3600.0/65536.0,1,-nbitq), 
to_sfixed(-1435.0/65536.0,1,-nbitq), 
to_sfixed(-2264.0/65536.0,1,-nbitq), 
to_sfixed(477.0/65536.0,1,-nbitq), 
to_sfixed(-5509.0/65536.0,1,-nbitq), 
to_sfixed(-335.0/65536.0,1,-nbitq), 
to_sfixed(2646.0/65536.0,1,-nbitq), 
to_sfixed(-1232.0/65536.0,1,-nbitq), 
to_sfixed(-1511.0/65536.0,1,-nbitq), 
to_sfixed(-3994.0/65536.0,1,-nbitq), 
to_sfixed(-2722.0/65536.0,1,-nbitq), 
to_sfixed(2853.0/65536.0,1,-nbitq), 
to_sfixed(-482.0/65536.0,1,-nbitq), 
to_sfixed(241.0/65536.0,1,-nbitq), 
to_sfixed(6137.0/65536.0,1,-nbitq), 
to_sfixed(3751.0/65536.0,1,-nbitq), 
to_sfixed(-7961.0/65536.0,1,-nbitq), 
to_sfixed(-1312.0/65536.0,1,-nbitq), 
to_sfixed(-1032.0/65536.0,1,-nbitq), 
to_sfixed(1027.0/65536.0,1,-nbitq), 
to_sfixed(-1820.0/65536.0,1,-nbitq), 
to_sfixed(-3333.0/65536.0,1,-nbitq), 
to_sfixed(1990.0/65536.0,1,-nbitq), 
to_sfixed(1882.0/65536.0,1,-nbitq), 
to_sfixed(2340.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-744.0/65536.0,1,-nbitq), 
to_sfixed(-79.0/65536.0,1,-nbitq), 
to_sfixed(-3597.0/65536.0,1,-nbitq), 
to_sfixed(989.0/65536.0,1,-nbitq), 
to_sfixed(-288.0/65536.0,1,-nbitq), 
to_sfixed(-3364.0/65536.0,1,-nbitq), 
to_sfixed(-1714.0/65536.0,1,-nbitq), 
to_sfixed(-250.0/65536.0,1,-nbitq), 
to_sfixed(4213.0/65536.0,1,-nbitq), 
to_sfixed(-699.0/65536.0,1,-nbitq), 
to_sfixed(1274.0/65536.0,1,-nbitq), 
to_sfixed(-9279.0/65536.0,1,-nbitq), 
to_sfixed(625.0/65536.0,1,-nbitq), 
to_sfixed(-7108.0/65536.0,1,-nbitq), 
to_sfixed(1551.0/65536.0,1,-nbitq), 
to_sfixed(2940.0/65536.0,1,-nbitq), 
to_sfixed(2394.0/65536.0,1,-nbitq), 
to_sfixed(1897.0/65536.0,1,-nbitq), 
to_sfixed(-4687.0/65536.0,1,-nbitq), 
to_sfixed(796.0/65536.0,1,-nbitq), 
to_sfixed(3458.0/65536.0,1,-nbitq), 
to_sfixed(1750.0/65536.0,1,-nbitq), 
to_sfixed(2385.0/65536.0,1,-nbitq), 
to_sfixed(-11320.0/65536.0,1,-nbitq), 
to_sfixed(-2220.0/65536.0,1,-nbitq), 
to_sfixed(-4444.0/65536.0,1,-nbitq), 
to_sfixed(1806.0/65536.0,1,-nbitq), 
to_sfixed(-4459.0/65536.0,1,-nbitq), 
to_sfixed(-6309.0/65536.0,1,-nbitq), 
to_sfixed(-2115.0/65536.0,1,-nbitq), 
to_sfixed(3712.0/65536.0,1,-nbitq), 
to_sfixed(599.0/65536.0,1,-nbitq), 
to_sfixed(823.0/65536.0,1,-nbitq), 
to_sfixed(-993.0/65536.0,1,-nbitq), 
to_sfixed(2017.0/65536.0,1,-nbitq), 
to_sfixed(2482.0/65536.0,1,-nbitq), 
to_sfixed(1600.0/65536.0,1,-nbitq), 
to_sfixed(1507.0/65536.0,1,-nbitq), 
to_sfixed(1502.0/65536.0,1,-nbitq), 
to_sfixed(2276.0/65536.0,1,-nbitq), 
to_sfixed(-697.0/65536.0,1,-nbitq), 
to_sfixed(1891.0/65536.0,1,-nbitq), 
to_sfixed(4898.0/65536.0,1,-nbitq), 
to_sfixed(2064.0/65536.0,1,-nbitq), 
to_sfixed(2835.0/65536.0,1,-nbitq), 
to_sfixed(-1155.0/65536.0,1,-nbitq), 
to_sfixed(-546.0/65536.0,1,-nbitq), 
to_sfixed(-2251.0/65536.0,1,-nbitq), 
to_sfixed(-783.0/65536.0,1,-nbitq), 
to_sfixed(766.0/65536.0,1,-nbitq), 
to_sfixed(-2371.0/65536.0,1,-nbitq), 
to_sfixed(4205.0/65536.0,1,-nbitq), 
to_sfixed(4828.0/65536.0,1,-nbitq), 
to_sfixed(-5914.0/65536.0,1,-nbitq), 
to_sfixed(-1623.0/65536.0,1,-nbitq), 
to_sfixed(2922.0/65536.0,1,-nbitq), 
to_sfixed(-2790.0/65536.0,1,-nbitq), 
to_sfixed(-3524.0/65536.0,1,-nbitq), 
to_sfixed(2372.0/65536.0,1,-nbitq), 
to_sfixed(-7344.0/65536.0,1,-nbitq), 
to_sfixed(-378.0/65536.0,1,-nbitq), 
to_sfixed(-46.0/65536.0,1,-nbitq), 
to_sfixed(-1272.0/65536.0,1,-nbitq), 
to_sfixed(-158.0/65536.0,1,-nbitq), 
to_sfixed(398.0/65536.0,1,-nbitq), 
to_sfixed(1937.0/65536.0,1,-nbitq), 
to_sfixed(4767.0/65536.0,1,-nbitq), 
to_sfixed(2625.0/65536.0,1,-nbitq), 
to_sfixed(-642.0/65536.0,1,-nbitq), 
to_sfixed(1014.0/65536.0,1,-nbitq), 
to_sfixed(3014.0/65536.0,1,-nbitq), 
to_sfixed(-7389.0/65536.0,1,-nbitq), 
to_sfixed(-5321.0/65536.0,1,-nbitq), 
to_sfixed(-1208.0/65536.0,1,-nbitq), 
to_sfixed(-2672.0/65536.0,1,-nbitq), 
to_sfixed(-4007.0/65536.0,1,-nbitq), 
to_sfixed(-2041.0/65536.0,1,-nbitq), 
to_sfixed(690.0/65536.0,1,-nbitq), 
to_sfixed(1027.0/65536.0,1,-nbitq), 
to_sfixed(1812.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1699.0/65536.0,1,-nbitq), 
to_sfixed(-1269.0/65536.0,1,-nbitq), 
to_sfixed(-1288.0/65536.0,1,-nbitq), 
to_sfixed(484.0/65536.0,1,-nbitq), 
to_sfixed(-3477.0/65536.0,1,-nbitq), 
to_sfixed(-509.0/65536.0,1,-nbitq), 
to_sfixed(234.0/65536.0,1,-nbitq), 
to_sfixed(-1338.0/65536.0,1,-nbitq), 
to_sfixed(2550.0/65536.0,1,-nbitq), 
to_sfixed(-509.0/65536.0,1,-nbitq), 
to_sfixed(-375.0/65536.0,1,-nbitq), 
to_sfixed(-10407.0/65536.0,1,-nbitq), 
to_sfixed(3329.0/65536.0,1,-nbitq), 
to_sfixed(750.0/65536.0,1,-nbitq), 
to_sfixed(4470.0/65536.0,1,-nbitq), 
to_sfixed(-2327.0/65536.0,1,-nbitq), 
to_sfixed(-1244.0/65536.0,1,-nbitq), 
to_sfixed(413.0/65536.0,1,-nbitq), 
to_sfixed(-5698.0/65536.0,1,-nbitq), 
to_sfixed(619.0/65536.0,1,-nbitq), 
to_sfixed(16.0/65536.0,1,-nbitq), 
to_sfixed(630.0/65536.0,1,-nbitq), 
to_sfixed(4847.0/65536.0,1,-nbitq), 
to_sfixed(-10895.0/65536.0,1,-nbitq), 
to_sfixed(-5514.0/65536.0,1,-nbitq), 
to_sfixed(-4667.0/65536.0,1,-nbitq), 
to_sfixed(6171.0/65536.0,1,-nbitq), 
to_sfixed(-2705.0/65536.0,1,-nbitq), 
to_sfixed(-404.0/65536.0,1,-nbitq), 
to_sfixed(3972.0/65536.0,1,-nbitq), 
to_sfixed(6494.0/65536.0,1,-nbitq), 
to_sfixed(1790.0/65536.0,1,-nbitq), 
to_sfixed(-328.0/65536.0,1,-nbitq), 
to_sfixed(-3972.0/65536.0,1,-nbitq), 
to_sfixed(-403.0/65536.0,1,-nbitq), 
to_sfixed(1277.0/65536.0,1,-nbitq), 
to_sfixed(-1413.0/65536.0,1,-nbitq), 
to_sfixed(-1057.0/65536.0,1,-nbitq), 
to_sfixed(6153.0/65536.0,1,-nbitq), 
to_sfixed(-1133.0/65536.0,1,-nbitq), 
to_sfixed(-1309.0/65536.0,1,-nbitq), 
to_sfixed(2577.0/65536.0,1,-nbitq), 
to_sfixed(2705.0/65536.0,1,-nbitq), 
to_sfixed(-1491.0/65536.0,1,-nbitq), 
to_sfixed(157.0/65536.0,1,-nbitq), 
to_sfixed(2345.0/65536.0,1,-nbitq), 
to_sfixed(2690.0/65536.0,1,-nbitq), 
to_sfixed(-2278.0/65536.0,1,-nbitq), 
to_sfixed(-825.0/65536.0,1,-nbitq), 
to_sfixed(-212.0/65536.0,1,-nbitq), 
to_sfixed(-1051.0/65536.0,1,-nbitq), 
to_sfixed(423.0/65536.0,1,-nbitq), 
to_sfixed(6291.0/65536.0,1,-nbitq), 
to_sfixed(-1833.0/65536.0,1,-nbitq), 
to_sfixed(-1357.0/65536.0,1,-nbitq), 
to_sfixed(3798.0/65536.0,1,-nbitq), 
to_sfixed(-1104.0/65536.0,1,-nbitq), 
to_sfixed(-2546.0/65536.0,1,-nbitq), 
to_sfixed(-137.0/65536.0,1,-nbitq), 
to_sfixed(-7787.0/65536.0,1,-nbitq), 
to_sfixed(-2839.0/65536.0,1,-nbitq), 
to_sfixed(-2401.0/65536.0,1,-nbitq), 
to_sfixed(-2172.0/65536.0,1,-nbitq), 
to_sfixed(1962.0/65536.0,1,-nbitq), 
to_sfixed(-3224.0/65536.0,1,-nbitq), 
to_sfixed(4251.0/65536.0,1,-nbitq), 
to_sfixed(571.0/65536.0,1,-nbitq), 
to_sfixed(2892.0/65536.0,1,-nbitq), 
to_sfixed(-1549.0/65536.0,1,-nbitq), 
to_sfixed(3262.0/65536.0,1,-nbitq), 
to_sfixed(-761.0/65536.0,1,-nbitq), 
to_sfixed(-4.0/65536.0,1,-nbitq), 
to_sfixed(-1191.0/65536.0,1,-nbitq), 
to_sfixed(-361.0/65536.0,1,-nbitq), 
to_sfixed(1915.0/65536.0,1,-nbitq), 
to_sfixed(-1144.0/65536.0,1,-nbitq), 
to_sfixed(1861.0/65536.0,1,-nbitq), 
to_sfixed(1325.0/65536.0,1,-nbitq), 
to_sfixed(2451.0/65536.0,1,-nbitq), 
to_sfixed(108.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3579.0/65536.0,1,-nbitq), 
to_sfixed(660.0/65536.0,1,-nbitq), 
to_sfixed(-4757.0/65536.0,1,-nbitq), 
to_sfixed(5684.0/65536.0,1,-nbitq), 
to_sfixed(4017.0/65536.0,1,-nbitq), 
to_sfixed(-3433.0/65536.0,1,-nbitq), 
to_sfixed(-3553.0/65536.0,1,-nbitq), 
to_sfixed(-258.0/65536.0,1,-nbitq), 
to_sfixed(2325.0/65536.0,1,-nbitq), 
to_sfixed(-748.0/65536.0,1,-nbitq), 
to_sfixed(698.0/65536.0,1,-nbitq), 
to_sfixed(-7829.0/65536.0,1,-nbitq), 
to_sfixed(2589.0/65536.0,1,-nbitq), 
to_sfixed(2578.0/65536.0,1,-nbitq), 
to_sfixed(2863.0/65536.0,1,-nbitq), 
to_sfixed(-1943.0/65536.0,1,-nbitq), 
to_sfixed(-1147.0/65536.0,1,-nbitq), 
to_sfixed(-3090.0/65536.0,1,-nbitq), 
to_sfixed(-3770.0/65536.0,1,-nbitq), 
to_sfixed(-504.0/65536.0,1,-nbitq), 
to_sfixed(-2735.0/65536.0,1,-nbitq), 
to_sfixed(1031.0/65536.0,1,-nbitq), 
to_sfixed(4005.0/65536.0,1,-nbitq), 
to_sfixed(-715.0/65536.0,1,-nbitq), 
to_sfixed(-4912.0/65536.0,1,-nbitq), 
to_sfixed(-1418.0/65536.0,1,-nbitq), 
to_sfixed(8322.0/65536.0,1,-nbitq), 
to_sfixed(-3490.0/65536.0,1,-nbitq), 
to_sfixed(3248.0/65536.0,1,-nbitq), 
to_sfixed(2019.0/65536.0,1,-nbitq), 
to_sfixed(187.0/65536.0,1,-nbitq), 
to_sfixed(4096.0/65536.0,1,-nbitq), 
to_sfixed(-2658.0/65536.0,1,-nbitq), 
to_sfixed(-4148.0/65536.0,1,-nbitq), 
to_sfixed(41.0/65536.0,1,-nbitq), 
to_sfixed(1763.0/65536.0,1,-nbitq), 
to_sfixed(-1952.0/65536.0,1,-nbitq), 
to_sfixed(-2069.0/65536.0,1,-nbitq), 
to_sfixed(7176.0/65536.0,1,-nbitq), 
to_sfixed(751.0/65536.0,1,-nbitq), 
to_sfixed(-1945.0/65536.0,1,-nbitq), 
to_sfixed(-1309.0/65536.0,1,-nbitq), 
to_sfixed(-3782.0/65536.0,1,-nbitq), 
to_sfixed(-123.0/65536.0,1,-nbitq), 
to_sfixed(-2429.0/65536.0,1,-nbitq), 
to_sfixed(97.0/65536.0,1,-nbitq), 
to_sfixed(2090.0/65536.0,1,-nbitq), 
to_sfixed(-1682.0/65536.0,1,-nbitq), 
to_sfixed(1466.0/65536.0,1,-nbitq), 
to_sfixed(-857.0/65536.0,1,-nbitq), 
to_sfixed(1003.0/65536.0,1,-nbitq), 
to_sfixed(-1692.0/65536.0,1,-nbitq), 
to_sfixed(4860.0/65536.0,1,-nbitq), 
to_sfixed(-1021.0/65536.0,1,-nbitq), 
to_sfixed(-627.0/65536.0,1,-nbitq), 
to_sfixed(-1941.0/65536.0,1,-nbitq), 
to_sfixed(2243.0/65536.0,1,-nbitq), 
to_sfixed(-728.0/65536.0,1,-nbitq), 
to_sfixed(1774.0/65536.0,1,-nbitq), 
to_sfixed(-6060.0/65536.0,1,-nbitq), 
to_sfixed(-5873.0/65536.0,1,-nbitq), 
to_sfixed(2326.0/65536.0,1,-nbitq), 
to_sfixed(-286.0/65536.0,1,-nbitq), 
to_sfixed(991.0/65536.0,1,-nbitq), 
to_sfixed(-2088.0/65536.0,1,-nbitq), 
to_sfixed(4627.0/65536.0,1,-nbitq), 
to_sfixed(670.0/65536.0,1,-nbitq), 
to_sfixed(7266.0/65536.0,1,-nbitq), 
to_sfixed(260.0/65536.0,1,-nbitq), 
to_sfixed(957.0/65536.0,1,-nbitq), 
to_sfixed(1108.0/65536.0,1,-nbitq), 
to_sfixed(-2197.0/65536.0,1,-nbitq), 
to_sfixed(-2005.0/65536.0,1,-nbitq), 
to_sfixed(-1068.0/65536.0,1,-nbitq), 
to_sfixed(990.0/65536.0,1,-nbitq), 
to_sfixed(-1178.0/65536.0,1,-nbitq), 
to_sfixed(-1255.0/65536.0,1,-nbitq), 
to_sfixed(716.0/65536.0,1,-nbitq), 
to_sfixed(111.0/65536.0,1,-nbitq), 
to_sfixed(2821.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3080.0/65536.0,1,-nbitq), 
to_sfixed(3553.0/65536.0,1,-nbitq), 
to_sfixed(-5874.0/65536.0,1,-nbitq), 
to_sfixed(5354.0/65536.0,1,-nbitq), 
to_sfixed(7751.0/65536.0,1,-nbitq), 
to_sfixed(993.0/65536.0,1,-nbitq), 
to_sfixed(-4722.0/65536.0,1,-nbitq), 
to_sfixed(1655.0/65536.0,1,-nbitq), 
to_sfixed(-1051.0/65536.0,1,-nbitq), 
to_sfixed(-16.0/65536.0,1,-nbitq), 
to_sfixed(1212.0/65536.0,1,-nbitq), 
to_sfixed(-7690.0/65536.0,1,-nbitq), 
to_sfixed(3.0/65536.0,1,-nbitq), 
to_sfixed(875.0/65536.0,1,-nbitq), 
to_sfixed(-1565.0/65536.0,1,-nbitq), 
to_sfixed(2135.0/65536.0,1,-nbitq), 
to_sfixed(140.0/65536.0,1,-nbitq), 
to_sfixed(-1498.0/65536.0,1,-nbitq), 
to_sfixed(-852.0/65536.0,1,-nbitq), 
to_sfixed(2625.0/65536.0,1,-nbitq), 
to_sfixed(-5074.0/65536.0,1,-nbitq), 
to_sfixed(819.0/65536.0,1,-nbitq), 
to_sfixed(-2640.0/65536.0,1,-nbitq), 
to_sfixed(2915.0/65536.0,1,-nbitq), 
to_sfixed(-100.0/65536.0,1,-nbitq), 
to_sfixed(-8077.0/65536.0,1,-nbitq), 
to_sfixed(4174.0/65536.0,1,-nbitq), 
to_sfixed(-3654.0/65536.0,1,-nbitq), 
to_sfixed(1730.0/65536.0,1,-nbitq), 
to_sfixed(527.0/65536.0,1,-nbitq), 
to_sfixed(1269.0/65536.0,1,-nbitq), 
to_sfixed(-356.0/65536.0,1,-nbitq), 
to_sfixed(-2762.0/65536.0,1,-nbitq), 
to_sfixed(1486.0/65536.0,1,-nbitq), 
to_sfixed(-1811.0/65536.0,1,-nbitq), 
to_sfixed(1676.0/65536.0,1,-nbitq), 
to_sfixed(405.0/65536.0,1,-nbitq), 
to_sfixed(64.0/65536.0,1,-nbitq), 
to_sfixed(5570.0/65536.0,1,-nbitq), 
to_sfixed(-467.0/65536.0,1,-nbitq), 
to_sfixed(2129.0/65536.0,1,-nbitq), 
to_sfixed(-2265.0/65536.0,1,-nbitq), 
to_sfixed(-3765.0/65536.0,1,-nbitq), 
to_sfixed(2.0/65536.0,1,-nbitq), 
to_sfixed(-2425.0/65536.0,1,-nbitq), 
to_sfixed(-3390.0/65536.0,1,-nbitq), 
to_sfixed(2034.0/65536.0,1,-nbitq), 
to_sfixed(214.0/65536.0,1,-nbitq), 
to_sfixed(2019.0/65536.0,1,-nbitq), 
to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(812.0/65536.0,1,-nbitq), 
to_sfixed(501.0/65536.0,1,-nbitq), 
to_sfixed(-1273.0/65536.0,1,-nbitq), 
to_sfixed(-5639.0/65536.0,1,-nbitq), 
to_sfixed(-2108.0/65536.0,1,-nbitq), 
to_sfixed(-2376.0/65536.0,1,-nbitq), 
to_sfixed(918.0/65536.0,1,-nbitq), 
to_sfixed(1528.0/65536.0,1,-nbitq), 
to_sfixed(673.0/65536.0,1,-nbitq), 
to_sfixed(-1640.0/65536.0,1,-nbitq), 
to_sfixed(-720.0/65536.0,1,-nbitq), 
to_sfixed(1625.0/65536.0,1,-nbitq), 
to_sfixed(1220.0/65536.0,1,-nbitq), 
to_sfixed(-299.0/65536.0,1,-nbitq), 
to_sfixed(223.0/65536.0,1,-nbitq), 
to_sfixed(4475.0/65536.0,1,-nbitq), 
to_sfixed(-4533.0/65536.0,1,-nbitq), 
to_sfixed(5955.0/65536.0,1,-nbitq), 
to_sfixed(901.0/65536.0,1,-nbitq), 
to_sfixed(130.0/65536.0,1,-nbitq), 
to_sfixed(808.0/65536.0,1,-nbitq), 
to_sfixed(-4028.0/65536.0,1,-nbitq), 
to_sfixed(-1752.0/65536.0,1,-nbitq), 
to_sfixed(-1046.0/65536.0,1,-nbitq), 
to_sfixed(2361.0/65536.0,1,-nbitq), 
to_sfixed(2764.0/65536.0,1,-nbitq), 
to_sfixed(1846.0/65536.0,1,-nbitq), 
to_sfixed(-4009.0/65536.0,1,-nbitq), 
to_sfixed(-954.0/65536.0,1,-nbitq), 
to_sfixed(2458.0/65536.0,1,-nbitq)  ), 
( to_sfixed(197.0/65536.0,1,-nbitq), 
to_sfixed(-999.0/65536.0,1,-nbitq), 
to_sfixed(-10642.0/65536.0,1,-nbitq), 
to_sfixed(5566.0/65536.0,1,-nbitq), 
to_sfixed(7408.0/65536.0,1,-nbitq), 
to_sfixed(-2581.0/65536.0,1,-nbitq), 
to_sfixed(-4287.0/65536.0,1,-nbitq), 
to_sfixed(2274.0/65536.0,1,-nbitq), 
to_sfixed(5726.0/65536.0,1,-nbitq), 
to_sfixed(2394.0/65536.0,1,-nbitq), 
to_sfixed(-35.0/65536.0,1,-nbitq), 
to_sfixed(-46.0/65536.0,1,-nbitq), 
to_sfixed(-588.0/65536.0,1,-nbitq), 
to_sfixed(4223.0/65536.0,1,-nbitq), 
to_sfixed(-3034.0/65536.0,1,-nbitq), 
to_sfixed(1675.0/65536.0,1,-nbitq), 
to_sfixed(1697.0/65536.0,1,-nbitq), 
to_sfixed(-6373.0/65536.0,1,-nbitq), 
to_sfixed(-2802.0/65536.0,1,-nbitq), 
to_sfixed(-1520.0/65536.0,1,-nbitq), 
to_sfixed(-4369.0/65536.0,1,-nbitq), 
to_sfixed(4722.0/65536.0,1,-nbitq), 
to_sfixed(-135.0/65536.0,1,-nbitq), 
to_sfixed(2202.0/65536.0,1,-nbitq), 
to_sfixed(-4708.0/65536.0,1,-nbitq), 
to_sfixed(-5064.0/65536.0,1,-nbitq), 
to_sfixed(6544.0/65536.0,1,-nbitq), 
to_sfixed(-3150.0/65536.0,1,-nbitq), 
to_sfixed(-4031.0/65536.0,1,-nbitq), 
to_sfixed(1742.0/65536.0,1,-nbitq), 
to_sfixed(-5530.0/65536.0,1,-nbitq), 
to_sfixed(2308.0/65536.0,1,-nbitq), 
to_sfixed(-1465.0/65536.0,1,-nbitq), 
to_sfixed(1850.0/65536.0,1,-nbitq), 
to_sfixed(184.0/65536.0,1,-nbitq), 
to_sfixed(3397.0/65536.0,1,-nbitq), 
to_sfixed(572.0/65536.0,1,-nbitq), 
to_sfixed(399.0/65536.0,1,-nbitq), 
to_sfixed(6682.0/65536.0,1,-nbitq), 
to_sfixed(1087.0/65536.0,1,-nbitq), 
to_sfixed(4232.0/65536.0,1,-nbitq), 
to_sfixed(2481.0/65536.0,1,-nbitq), 
to_sfixed(-12846.0/65536.0,1,-nbitq), 
to_sfixed(4313.0/65536.0,1,-nbitq), 
to_sfixed(701.0/65536.0,1,-nbitq), 
to_sfixed(-4182.0/65536.0,1,-nbitq), 
to_sfixed(-1653.0/65536.0,1,-nbitq), 
to_sfixed(1797.0/65536.0,1,-nbitq), 
to_sfixed(1913.0/65536.0,1,-nbitq), 
to_sfixed(1231.0/65536.0,1,-nbitq), 
to_sfixed(3110.0/65536.0,1,-nbitq), 
to_sfixed(4361.0/65536.0,1,-nbitq), 
to_sfixed(-4283.0/65536.0,1,-nbitq), 
to_sfixed(-4877.0/65536.0,1,-nbitq), 
to_sfixed(-1713.0/65536.0,1,-nbitq), 
to_sfixed(-4435.0/65536.0,1,-nbitq), 
to_sfixed(1187.0/65536.0,1,-nbitq), 
to_sfixed(-601.0/65536.0,1,-nbitq), 
to_sfixed(-845.0/65536.0,1,-nbitq), 
to_sfixed(1617.0/65536.0,1,-nbitq), 
to_sfixed(-685.0/65536.0,1,-nbitq), 
to_sfixed(1626.0/65536.0,1,-nbitq), 
to_sfixed(-363.0/65536.0,1,-nbitq), 
to_sfixed(1128.0/65536.0,1,-nbitq), 
to_sfixed(697.0/65536.0,1,-nbitq), 
to_sfixed(3504.0/65536.0,1,-nbitq), 
to_sfixed(-907.0/65536.0,1,-nbitq), 
to_sfixed(3270.0/65536.0,1,-nbitq), 
to_sfixed(-1452.0/65536.0,1,-nbitq), 
to_sfixed(-4034.0/65536.0,1,-nbitq), 
to_sfixed(-3117.0/65536.0,1,-nbitq), 
to_sfixed(-6361.0/65536.0,1,-nbitq), 
to_sfixed(-6257.0/65536.0,1,-nbitq), 
to_sfixed(617.0/65536.0,1,-nbitq), 
to_sfixed(-756.0/65536.0,1,-nbitq), 
to_sfixed(470.0/65536.0,1,-nbitq), 
to_sfixed(3762.0/65536.0,1,-nbitq), 
to_sfixed(-1487.0/65536.0,1,-nbitq), 
to_sfixed(2696.0/65536.0,1,-nbitq), 
to_sfixed(7926.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3428.0/65536.0,1,-nbitq), 
to_sfixed(821.0/65536.0,1,-nbitq), 
to_sfixed(-1329.0/65536.0,1,-nbitq), 
to_sfixed(4640.0/65536.0,1,-nbitq), 
to_sfixed(3949.0/65536.0,1,-nbitq), 
to_sfixed(-2049.0/65536.0,1,-nbitq), 
to_sfixed(-2560.0/65536.0,1,-nbitq), 
to_sfixed(-3605.0/65536.0,1,-nbitq), 
to_sfixed(2706.0/65536.0,1,-nbitq), 
to_sfixed(1150.0/65536.0,1,-nbitq), 
to_sfixed(-723.0/65536.0,1,-nbitq), 
to_sfixed(3224.0/65536.0,1,-nbitq), 
to_sfixed(-1624.0/65536.0,1,-nbitq), 
to_sfixed(3780.0/65536.0,1,-nbitq), 
to_sfixed(-698.0/65536.0,1,-nbitq), 
to_sfixed(-998.0/65536.0,1,-nbitq), 
to_sfixed(841.0/65536.0,1,-nbitq), 
to_sfixed(-4194.0/65536.0,1,-nbitq), 
to_sfixed(-2291.0/65536.0,1,-nbitq), 
to_sfixed(580.0/65536.0,1,-nbitq), 
to_sfixed(-3532.0/65536.0,1,-nbitq), 
to_sfixed(2398.0/65536.0,1,-nbitq), 
to_sfixed(3513.0/65536.0,1,-nbitq), 
to_sfixed(3804.0/65536.0,1,-nbitq), 
to_sfixed(-4054.0/65536.0,1,-nbitq), 
to_sfixed(-4833.0/65536.0,1,-nbitq), 
to_sfixed(4039.0/65536.0,1,-nbitq), 
to_sfixed(-4009.0/65536.0,1,-nbitq), 
to_sfixed(-8135.0/65536.0,1,-nbitq), 
to_sfixed(-460.0/65536.0,1,-nbitq), 
to_sfixed(-9021.0/65536.0,1,-nbitq), 
to_sfixed(4473.0/65536.0,1,-nbitq), 
to_sfixed(-1915.0/65536.0,1,-nbitq), 
to_sfixed(7571.0/65536.0,1,-nbitq), 
to_sfixed(305.0/65536.0,1,-nbitq), 
to_sfixed(364.0/65536.0,1,-nbitq), 
to_sfixed(-436.0/65536.0,1,-nbitq), 
to_sfixed(2749.0/65536.0,1,-nbitq), 
to_sfixed(5660.0/65536.0,1,-nbitq), 
to_sfixed(-403.0/65536.0,1,-nbitq), 
to_sfixed(640.0/65536.0,1,-nbitq), 
to_sfixed(228.0/65536.0,1,-nbitq), 
to_sfixed(-6815.0/65536.0,1,-nbitq), 
to_sfixed(2671.0/65536.0,1,-nbitq), 
to_sfixed(478.0/65536.0,1,-nbitq), 
to_sfixed(1788.0/65536.0,1,-nbitq), 
to_sfixed(2627.0/65536.0,1,-nbitq), 
to_sfixed(-2843.0/65536.0,1,-nbitq), 
to_sfixed(3509.0/65536.0,1,-nbitq), 
to_sfixed(-260.0/65536.0,1,-nbitq), 
to_sfixed(-2527.0/65536.0,1,-nbitq), 
to_sfixed(-423.0/65536.0,1,-nbitq), 
to_sfixed(-1207.0/65536.0,1,-nbitq), 
to_sfixed(-4133.0/65536.0,1,-nbitq), 
to_sfixed(-1155.0/65536.0,1,-nbitq), 
to_sfixed(-2052.0/65536.0,1,-nbitq), 
to_sfixed(-121.0/65536.0,1,-nbitq), 
to_sfixed(155.0/65536.0,1,-nbitq), 
to_sfixed(1403.0/65536.0,1,-nbitq), 
to_sfixed(5842.0/65536.0,1,-nbitq), 
to_sfixed(1683.0/65536.0,1,-nbitq), 
to_sfixed(2339.0/65536.0,1,-nbitq), 
to_sfixed(3211.0/65536.0,1,-nbitq), 
to_sfixed(2213.0/65536.0,1,-nbitq), 
to_sfixed(2887.0/65536.0,1,-nbitq), 
to_sfixed(6724.0/65536.0,1,-nbitq), 
to_sfixed(-2722.0/65536.0,1,-nbitq), 
to_sfixed(2780.0/65536.0,1,-nbitq), 
to_sfixed(-597.0/65536.0,1,-nbitq), 
to_sfixed(-3669.0/65536.0,1,-nbitq), 
to_sfixed(-1805.0/65536.0,1,-nbitq), 
to_sfixed(74.0/65536.0,1,-nbitq), 
to_sfixed(-2419.0/65536.0,1,-nbitq), 
to_sfixed(823.0/65536.0,1,-nbitq), 
to_sfixed(-1348.0/65536.0,1,-nbitq), 
to_sfixed(-4194.0/65536.0,1,-nbitq), 
to_sfixed(102.0/65536.0,1,-nbitq), 
to_sfixed(-5740.0/65536.0,1,-nbitq), 
to_sfixed(-1459.0/65536.0,1,-nbitq), 
to_sfixed(6880.0/65536.0,1,-nbitq)  ), 
( to_sfixed(319.0/65536.0,1,-nbitq), 
to_sfixed(1376.0/65536.0,1,-nbitq), 
to_sfixed(1717.0/65536.0,1,-nbitq), 
to_sfixed(2683.0/65536.0,1,-nbitq), 
to_sfixed(5174.0/65536.0,1,-nbitq), 
to_sfixed(1856.0/65536.0,1,-nbitq), 
to_sfixed(-7131.0/65536.0,1,-nbitq), 
to_sfixed(1453.0/65536.0,1,-nbitq), 
to_sfixed(1831.0/65536.0,1,-nbitq), 
to_sfixed(1750.0/65536.0,1,-nbitq), 
to_sfixed(2042.0/65536.0,1,-nbitq), 
to_sfixed(-2351.0/65536.0,1,-nbitq), 
to_sfixed(778.0/65536.0,1,-nbitq), 
to_sfixed(1832.0/65536.0,1,-nbitq), 
to_sfixed(-4648.0/65536.0,1,-nbitq), 
to_sfixed(-2281.0/65536.0,1,-nbitq), 
to_sfixed(-695.0/65536.0,1,-nbitq), 
to_sfixed(-6984.0/65536.0,1,-nbitq), 
to_sfixed(-2282.0/65536.0,1,-nbitq), 
to_sfixed(1998.0/65536.0,1,-nbitq), 
to_sfixed(-6787.0/65536.0,1,-nbitq), 
to_sfixed(-134.0/65536.0,1,-nbitq), 
to_sfixed(-444.0/65536.0,1,-nbitq), 
to_sfixed(6234.0/65536.0,1,-nbitq), 
to_sfixed(941.0/65536.0,1,-nbitq), 
to_sfixed(1502.0/65536.0,1,-nbitq), 
to_sfixed(4314.0/65536.0,1,-nbitq), 
to_sfixed(-4015.0/65536.0,1,-nbitq), 
to_sfixed(-8242.0/65536.0,1,-nbitq), 
to_sfixed(-529.0/65536.0,1,-nbitq), 
to_sfixed(-6273.0/65536.0,1,-nbitq), 
to_sfixed(-324.0/65536.0,1,-nbitq), 
to_sfixed(-3946.0/65536.0,1,-nbitq), 
to_sfixed(9586.0/65536.0,1,-nbitq), 
to_sfixed(-859.0/65536.0,1,-nbitq), 
to_sfixed(1674.0/65536.0,1,-nbitq), 
to_sfixed(-2717.0/65536.0,1,-nbitq), 
to_sfixed(-1713.0/65536.0,1,-nbitq), 
to_sfixed(5356.0/65536.0,1,-nbitq), 
to_sfixed(-1098.0/65536.0,1,-nbitq), 
to_sfixed(887.0/65536.0,1,-nbitq), 
to_sfixed(-1587.0/65536.0,1,-nbitq), 
to_sfixed(-6357.0/65536.0,1,-nbitq), 
to_sfixed(3752.0/65536.0,1,-nbitq), 
to_sfixed(-2275.0/65536.0,1,-nbitq), 
to_sfixed(-399.0/65536.0,1,-nbitq), 
to_sfixed(-1267.0/65536.0,1,-nbitq), 
to_sfixed(-1189.0/65536.0,1,-nbitq), 
to_sfixed(1625.0/65536.0,1,-nbitq), 
to_sfixed(2956.0/65536.0,1,-nbitq), 
to_sfixed(110.0/65536.0,1,-nbitq), 
to_sfixed(-2133.0/65536.0,1,-nbitq), 
to_sfixed(471.0/65536.0,1,-nbitq), 
to_sfixed(-4471.0/65536.0,1,-nbitq), 
to_sfixed(2117.0/65536.0,1,-nbitq), 
to_sfixed(2502.0/65536.0,1,-nbitq), 
to_sfixed(-1784.0/65536.0,1,-nbitq), 
to_sfixed(-2863.0/65536.0,1,-nbitq), 
to_sfixed(1204.0/65536.0,1,-nbitq), 
to_sfixed(2412.0/65536.0,1,-nbitq), 
to_sfixed(196.0/65536.0,1,-nbitq), 
to_sfixed(-2162.0/65536.0,1,-nbitq), 
to_sfixed(-421.0/65536.0,1,-nbitq), 
to_sfixed(2014.0/65536.0,1,-nbitq), 
to_sfixed(5836.0/65536.0,1,-nbitq), 
to_sfixed(6579.0/65536.0,1,-nbitq), 
to_sfixed(-1111.0/65536.0,1,-nbitq), 
to_sfixed(1508.0/65536.0,1,-nbitq), 
to_sfixed(1229.0/65536.0,1,-nbitq), 
to_sfixed(-9473.0/65536.0,1,-nbitq), 
to_sfixed(-915.0/65536.0,1,-nbitq), 
to_sfixed(160.0/65536.0,1,-nbitq), 
to_sfixed(-3028.0/65536.0,1,-nbitq), 
to_sfixed(-1421.0/65536.0,1,-nbitq), 
to_sfixed(-2724.0/65536.0,1,-nbitq), 
to_sfixed(-5097.0/65536.0,1,-nbitq), 
to_sfixed(1801.0/65536.0,1,-nbitq), 
to_sfixed(-261.0/65536.0,1,-nbitq), 
to_sfixed(1541.0/65536.0,1,-nbitq), 
to_sfixed(8239.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2207.0/65536.0,1,-nbitq), 
to_sfixed(31.0/65536.0,1,-nbitq), 
to_sfixed(3773.0/65536.0,1,-nbitq), 
to_sfixed(-2351.0/65536.0,1,-nbitq), 
to_sfixed(2812.0/65536.0,1,-nbitq), 
to_sfixed(1184.0/65536.0,1,-nbitq), 
to_sfixed(-1742.0/65536.0,1,-nbitq), 
to_sfixed(-356.0/65536.0,1,-nbitq), 
to_sfixed(3087.0/65536.0,1,-nbitq), 
to_sfixed(-2402.0/65536.0,1,-nbitq), 
to_sfixed(3909.0/65536.0,1,-nbitq), 
to_sfixed(-419.0/65536.0,1,-nbitq), 
to_sfixed(-1076.0/65536.0,1,-nbitq), 
to_sfixed(1702.0/65536.0,1,-nbitq), 
to_sfixed(-1563.0/65536.0,1,-nbitq), 
to_sfixed(-2058.0/65536.0,1,-nbitq), 
to_sfixed(202.0/65536.0,1,-nbitq), 
to_sfixed(-2484.0/65536.0,1,-nbitq), 
to_sfixed(1765.0/65536.0,1,-nbitq), 
to_sfixed(3035.0/65536.0,1,-nbitq), 
to_sfixed(-2828.0/65536.0,1,-nbitq), 
to_sfixed(-5204.0/65536.0,1,-nbitq), 
to_sfixed(-4416.0/65536.0,1,-nbitq), 
to_sfixed(2093.0/65536.0,1,-nbitq), 
to_sfixed(-375.0/65536.0,1,-nbitq), 
to_sfixed(-962.0/65536.0,1,-nbitq), 
to_sfixed(2116.0/65536.0,1,-nbitq), 
to_sfixed(-4601.0/65536.0,1,-nbitq), 
to_sfixed(-4541.0/65536.0,1,-nbitq), 
to_sfixed(3697.0/65536.0,1,-nbitq), 
to_sfixed(-4953.0/65536.0,1,-nbitq), 
to_sfixed(2227.0/65536.0,1,-nbitq), 
to_sfixed(-3878.0/65536.0,1,-nbitq), 
to_sfixed(11021.0/65536.0,1,-nbitq), 
to_sfixed(2445.0/65536.0,1,-nbitq), 
to_sfixed(1115.0/65536.0,1,-nbitq), 
to_sfixed(-2815.0/65536.0,1,-nbitq), 
to_sfixed(512.0/65536.0,1,-nbitq), 
to_sfixed(4188.0/65536.0,1,-nbitq), 
to_sfixed(1564.0/65536.0,1,-nbitq), 
to_sfixed(2869.0/65536.0,1,-nbitq), 
to_sfixed(-121.0/65536.0,1,-nbitq), 
to_sfixed(-445.0/65536.0,1,-nbitq), 
to_sfixed(5051.0/65536.0,1,-nbitq), 
to_sfixed(1928.0/65536.0,1,-nbitq), 
to_sfixed(-2609.0/65536.0,1,-nbitq), 
to_sfixed(-809.0/65536.0,1,-nbitq), 
to_sfixed(-4225.0/65536.0,1,-nbitq), 
to_sfixed(1598.0/65536.0,1,-nbitq), 
to_sfixed(-487.0/65536.0,1,-nbitq), 
to_sfixed(-1464.0/65536.0,1,-nbitq), 
to_sfixed(2660.0/65536.0,1,-nbitq), 
to_sfixed(2054.0/65536.0,1,-nbitq), 
to_sfixed(1262.0/65536.0,1,-nbitq), 
to_sfixed(3163.0/65536.0,1,-nbitq), 
to_sfixed(6.0/65536.0,1,-nbitq), 
to_sfixed(1651.0/65536.0,1,-nbitq), 
to_sfixed(-1789.0/65536.0,1,-nbitq), 
to_sfixed(-2487.0/65536.0,1,-nbitq), 
to_sfixed(4833.0/65536.0,1,-nbitq), 
to_sfixed(-612.0/65536.0,1,-nbitq), 
to_sfixed(761.0/65536.0,1,-nbitq), 
to_sfixed(2653.0/65536.0,1,-nbitq), 
to_sfixed(-1752.0/65536.0,1,-nbitq), 
to_sfixed(3624.0/65536.0,1,-nbitq), 
to_sfixed(10893.0/65536.0,1,-nbitq), 
to_sfixed(-733.0/65536.0,1,-nbitq), 
to_sfixed(3359.0/65536.0,1,-nbitq), 
to_sfixed(-1354.0/65536.0,1,-nbitq), 
to_sfixed(-6163.0/65536.0,1,-nbitq), 
to_sfixed(3691.0/65536.0,1,-nbitq), 
to_sfixed(2668.0/65536.0,1,-nbitq), 
to_sfixed(-1379.0/65536.0,1,-nbitq), 
to_sfixed(2811.0/65536.0,1,-nbitq), 
to_sfixed(1518.0/65536.0,1,-nbitq), 
to_sfixed(2236.0/65536.0,1,-nbitq), 
to_sfixed(2631.0/65536.0,1,-nbitq), 
to_sfixed(546.0/65536.0,1,-nbitq), 
to_sfixed(-1113.0/65536.0,1,-nbitq), 
to_sfixed(1971.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1646.0/65536.0,1,-nbitq), 
to_sfixed(-4007.0/65536.0,1,-nbitq), 
to_sfixed(3556.0/65536.0,1,-nbitq), 
to_sfixed(-1665.0/65536.0,1,-nbitq), 
to_sfixed(3720.0/65536.0,1,-nbitq), 
to_sfixed(2351.0/65536.0,1,-nbitq), 
to_sfixed(199.0/65536.0,1,-nbitq), 
to_sfixed(2933.0/65536.0,1,-nbitq), 
to_sfixed(-1157.0/65536.0,1,-nbitq), 
to_sfixed(-292.0/65536.0,1,-nbitq), 
to_sfixed(2788.0/65536.0,1,-nbitq), 
to_sfixed(-4618.0/65536.0,1,-nbitq), 
to_sfixed(-1962.0/65536.0,1,-nbitq), 
to_sfixed(-1404.0/65536.0,1,-nbitq), 
to_sfixed(2609.0/65536.0,1,-nbitq), 
to_sfixed(-539.0/65536.0,1,-nbitq), 
to_sfixed(682.0/65536.0,1,-nbitq), 
to_sfixed(-4909.0/65536.0,1,-nbitq), 
to_sfixed(-1673.0/65536.0,1,-nbitq), 
to_sfixed(-769.0/65536.0,1,-nbitq), 
to_sfixed(-1359.0/65536.0,1,-nbitq), 
to_sfixed(-1259.0/65536.0,1,-nbitq), 
to_sfixed(1697.0/65536.0,1,-nbitq), 
to_sfixed(-3699.0/65536.0,1,-nbitq), 
to_sfixed(64.0/65536.0,1,-nbitq), 
to_sfixed(-6183.0/65536.0,1,-nbitq), 
to_sfixed(1344.0/65536.0,1,-nbitq), 
to_sfixed(-1581.0/65536.0,1,-nbitq), 
to_sfixed(-1252.0/65536.0,1,-nbitq), 
to_sfixed(2125.0/65536.0,1,-nbitq), 
to_sfixed(-2734.0/65536.0,1,-nbitq), 
to_sfixed(4083.0/65536.0,1,-nbitq), 
to_sfixed(159.0/65536.0,1,-nbitq), 
to_sfixed(5252.0/65536.0,1,-nbitq), 
to_sfixed(2590.0/65536.0,1,-nbitq), 
to_sfixed(154.0/65536.0,1,-nbitq), 
to_sfixed(-2612.0/65536.0,1,-nbitq), 
to_sfixed(1304.0/65536.0,1,-nbitq), 
to_sfixed(-433.0/65536.0,1,-nbitq), 
to_sfixed(-841.0/65536.0,1,-nbitq), 
to_sfixed(-45.0/65536.0,1,-nbitq), 
to_sfixed(1594.0/65536.0,1,-nbitq), 
to_sfixed(-654.0/65536.0,1,-nbitq), 
to_sfixed(2946.0/65536.0,1,-nbitq), 
to_sfixed(2789.0/65536.0,1,-nbitq), 
to_sfixed(-1960.0/65536.0,1,-nbitq), 
to_sfixed(36.0/65536.0,1,-nbitq), 
to_sfixed(-5286.0/65536.0,1,-nbitq), 
to_sfixed(-1808.0/65536.0,1,-nbitq), 
to_sfixed(1663.0/65536.0,1,-nbitq), 
to_sfixed(2991.0/65536.0,1,-nbitq), 
to_sfixed(2709.0/65536.0,1,-nbitq), 
to_sfixed(5631.0/65536.0,1,-nbitq), 
to_sfixed(5638.0/65536.0,1,-nbitq), 
to_sfixed(2356.0/65536.0,1,-nbitq), 
to_sfixed(-2217.0/65536.0,1,-nbitq), 
to_sfixed(1892.0/65536.0,1,-nbitq), 
to_sfixed(-1866.0/65536.0,1,-nbitq), 
to_sfixed(3216.0/65536.0,1,-nbitq), 
to_sfixed(3479.0/65536.0,1,-nbitq), 
to_sfixed(-115.0/65536.0,1,-nbitq), 
to_sfixed(-1167.0/65536.0,1,-nbitq), 
to_sfixed(1395.0/65536.0,1,-nbitq), 
to_sfixed(926.0/65536.0,1,-nbitq), 
to_sfixed(1403.0/65536.0,1,-nbitq), 
to_sfixed(8857.0/65536.0,1,-nbitq), 
to_sfixed(-4394.0/65536.0,1,-nbitq), 
to_sfixed(-578.0/65536.0,1,-nbitq), 
to_sfixed(-3564.0/65536.0,1,-nbitq), 
to_sfixed(-1456.0/65536.0,1,-nbitq), 
to_sfixed(1841.0/65536.0,1,-nbitq), 
to_sfixed(5200.0/65536.0,1,-nbitq), 
to_sfixed(-5611.0/65536.0,1,-nbitq), 
to_sfixed(1101.0/65536.0,1,-nbitq), 
to_sfixed(1088.0/65536.0,1,-nbitq), 
to_sfixed(-31.0/65536.0,1,-nbitq), 
to_sfixed(-2375.0/65536.0,1,-nbitq), 
to_sfixed(977.0/65536.0,1,-nbitq), 
to_sfixed(1503.0/65536.0,1,-nbitq), 
to_sfixed(2766.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1527.0/65536.0,1,-nbitq), 
to_sfixed(1558.0/65536.0,1,-nbitq), 
to_sfixed(2910.0/65536.0,1,-nbitq), 
to_sfixed(1686.0/65536.0,1,-nbitq), 
to_sfixed(-758.0/65536.0,1,-nbitq), 
to_sfixed(-2305.0/65536.0,1,-nbitq), 
to_sfixed(-2015.0/65536.0,1,-nbitq), 
to_sfixed(4060.0/65536.0,1,-nbitq), 
to_sfixed(-1702.0/65536.0,1,-nbitq), 
to_sfixed(-2101.0/65536.0,1,-nbitq), 
to_sfixed(2268.0/65536.0,1,-nbitq), 
to_sfixed(-2099.0/65536.0,1,-nbitq), 
to_sfixed(2553.0/65536.0,1,-nbitq), 
to_sfixed(-3781.0/65536.0,1,-nbitq), 
to_sfixed(2255.0/65536.0,1,-nbitq), 
to_sfixed(532.0/65536.0,1,-nbitq), 
to_sfixed(609.0/65536.0,1,-nbitq), 
to_sfixed(-4857.0/65536.0,1,-nbitq), 
to_sfixed(1703.0/65536.0,1,-nbitq), 
to_sfixed(1264.0/65536.0,1,-nbitq), 
to_sfixed(-239.0/65536.0,1,-nbitq), 
to_sfixed(-5537.0/65536.0,1,-nbitq), 
to_sfixed(1264.0/65536.0,1,-nbitq), 
to_sfixed(-4571.0/65536.0,1,-nbitq), 
to_sfixed(1354.0/65536.0,1,-nbitq), 
to_sfixed(-3053.0/65536.0,1,-nbitq), 
to_sfixed(-76.0/65536.0,1,-nbitq), 
to_sfixed(-999.0/65536.0,1,-nbitq), 
to_sfixed(-4263.0/65536.0,1,-nbitq), 
to_sfixed(3088.0/65536.0,1,-nbitq), 
to_sfixed(-365.0/65536.0,1,-nbitq), 
to_sfixed(1861.0/65536.0,1,-nbitq), 
to_sfixed(-308.0/65536.0,1,-nbitq), 
to_sfixed(1701.0/65536.0,1,-nbitq), 
to_sfixed(1671.0/65536.0,1,-nbitq), 
to_sfixed(-333.0/65536.0,1,-nbitq), 
to_sfixed(3014.0/65536.0,1,-nbitq), 
to_sfixed(3839.0/65536.0,1,-nbitq), 
to_sfixed(1484.0/65536.0,1,-nbitq), 
to_sfixed(-76.0/65536.0,1,-nbitq), 
to_sfixed(-1854.0/65536.0,1,-nbitq), 
to_sfixed(-1981.0/65536.0,1,-nbitq), 
to_sfixed(-939.0/65536.0,1,-nbitq), 
to_sfixed(4468.0/65536.0,1,-nbitq), 
to_sfixed(-585.0/65536.0,1,-nbitq), 
to_sfixed(-3876.0/65536.0,1,-nbitq), 
to_sfixed(2330.0/65536.0,1,-nbitq), 
to_sfixed(-2106.0/65536.0,1,-nbitq), 
to_sfixed(2998.0/65536.0,1,-nbitq), 
to_sfixed(645.0/65536.0,1,-nbitq), 
to_sfixed(1448.0/65536.0,1,-nbitq), 
to_sfixed(-2436.0/65536.0,1,-nbitq), 
to_sfixed(3906.0/65536.0,1,-nbitq), 
to_sfixed(-2265.0/65536.0,1,-nbitq), 
to_sfixed(695.0/65536.0,1,-nbitq), 
to_sfixed(3068.0/65536.0,1,-nbitq), 
to_sfixed(1665.0/65536.0,1,-nbitq), 
to_sfixed(-1094.0/65536.0,1,-nbitq), 
to_sfixed(1154.0/65536.0,1,-nbitq), 
to_sfixed(431.0/65536.0,1,-nbitq), 
to_sfixed(1900.0/65536.0,1,-nbitq), 
to_sfixed(2457.0/65536.0,1,-nbitq), 
to_sfixed(889.0/65536.0,1,-nbitq), 
to_sfixed(-2551.0/65536.0,1,-nbitq), 
to_sfixed(4320.0/65536.0,1,-nbitq), 
to_sfixed(7463.0/65536.0,1,-nbitq), 
to_sfixed(-2925.0/65536.0,1,-nbitq), 
to_sfixed(-6456.0/65536.0,1,-nbitq), 
to_sfixed(1970.0/65536.0,1,-nbitq), 
to_sfixed(-3711.0/65536.0,1,-nbitq), 
to_sfixed(-293.0/65536.0,1,-nbitq), 
to_sfixed(683.0/65536.0,1,-nbitq), 
to_sfixed(-2015.0/65536.0,1,-nbitq), 
to_sfixed(1516.0/65536.0,1,-nbitq), 
to_sfixed(-1617.0/65536.0,1,-nbitq), 
to_sfixed(1622.0/65536.0,1,-nbitq), 
to_sfixed(-4104.0/65536.0,1,-nbitq), 
to_sfixed(791.0/65536.0,1,-nbitq), 
to_sfixed(-1064.0/65536.0,1,-nbitq), 
to_sfixed(3717.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3426.0/65536.0,1,-nbitq), 
to_sfixed(496.0/65536.0,1,-nbitq), 
to_sfixed(1227.0/65536.0,1,-nbitq), 
to_sfixed(-1024.0/65536.0,1,-nbitq), 
to_sfixed(-3026.0/65536.0,1,-nbitq), 
to_sfixed(-6.0/65536.0,1,-nbitq), 
to_sfixed(1271.0/65536.0,1,-nbitq), 
to_sfixed(4673.0/65536.0,1,-nbitq), 
to_sfixed(-1370.0/65536.0,1,-nbitq), 
to_sfixed(-1757.0/65536.0,1,-nbitq), 
to_sfixed(-1075.0/65536.0,1,-nbitq), 
to_sfixed(-5207.0/65536.0,1,-nbitq), 
to_sfixed(-933.0/65536.0,1,-nbitq), 
to_sfixed(1658.0/65536.0,1,-nbitq), 
to_sfixed(-1362.0/65536.0,1,-nbitq), 
to_sfixed(3075.0/65536.0,1,-nbitq), 
to_sfixed(-799.0/65536.0,1,-nbitq), 
to_sfixed(1392.0/65536.0,1,-nbitq), 
to_sfixed(2220.0/65536.0,1,-nbitq), 
to_sfixed(-1923.0/65536.0,1,-nbitq), 
to_sfixed(-1341.0/65536.0,1,-nbitq), 
to_sfixed(209.0/65536.0,1,-nbitq), 
to_sfixed(-2140.0/65536.0,1,-nbitq), 
to_sfixed(-1746.0/65536.0,1,-nbitq), 
to_sfixed(-1955.0/65536.0,1,-nbitq), 
to_sfixed(-3045.0/65536.0,1,-nbitq), 
to_sfixed(-4992.0/65536.0,1,-nbitq), 
to_sfixed(1205.0/65536.0,1,-nbitq), 
to_sfixed(-4991.0/65536.0,1,-nbitq), 
to_sfixed(1470.0/65536.0,1,-nbitq), 
to_sfixed(2261.0/65536.0,1,-nbitq), 
to_sfixed(761.0/65536.0,1,-nbitq), 
to_sfixed(-1052.0/65536.0,1,-nbitq), 
to_sfixed(-2754.0/65536.0,1,-nbitq), 
to_sfixed(-2569.0/65536.0,1,-nbitq), 
to_sfixed(2547.0/65536.0,1,-nbitq), 
to_sfixed(4350.0/65536.0,1,-nbitq), 
to_sfixed(-1120.0/65536.0,1,-nbitq), 
to_sfixed(3271.0/65536.0,1,-nbitq), 
to_sfixed(-1942.0/65536.0,1,-nbitq), 
to_sfixed(1647.0/65536.0,1,-nbitq), 
to_sfixed(455.0/65536.0,1,-nbitq), 
to_sfixed(-5484.0/65536.0,1,-nbitq), 
to_sfixed(5410.0/65536.0,1,-nbitq), 
to_sfixed(3279.0/65536.0,1,-nbitq), 
to_sfixed(-1435.0/65536.0,1,-nbitq), 
to_sfixed(-426.0/65536.0,1,-nbitq), 
to_sfixed(-4650.0/65536.0,1,-nbitq), 
to_sfixed(-1162.0/65536.0,1,-nbitq), 
to_sfixed(2089.0/65536.0,1,-nbitq), 
to_sfixed(932.0/65536.0,1,-nbitq), 
to_sfixed(-1044.0/65536.0,1,-nbitq), 
to_sfixed(3930.0/65536.0,1,-nbitq), 
to_sfixed(-5670.0/65536.0,1,-nbitq), 
to_sfixed(2928.0/65536.0,1,-nbitq), 
to_sfixed(-1313.0/65536.0,1,-nbitq), 
to_sfixed(-872.0/65536.0,1,-nbitq), 
to_sfixed(1675.0/65536.0,1,-nbitq), 
to_sfixed(106.0/65536.0,1,-nbitq), 
to_sfixed(1173.0/65536.0,1,-nbitq), 
to_sfixed(30.0/65536.0,1,-nbitq), 
to_sfixed(1359.0/65536.0,1,-nbitq), 
to_sfixed(-1134.0/65536.0,1,-nbitq), 
to_sfixed(528.0/65536.0,1,-nbitq), 
to_sfixed(5023.0/65536.0,1,-nbitq), 
to_sfixed(991.0/65536.0,1,-nbitq), 
to_sfixed(3379.0/65536.0,1,-nbitq), 
to_sfixed(-3025.0/65536.0,1,-nbitq), 
to_sfixed(2500.0/65536.0,1,-nbitq), 
to_sfixed(-3108.0/65536.0,1,-nbitq), 
to_sfixed(-2996.0/65536.0,1,-nbitq), 
to_sfixed(4237.0/65536.0,1,-nbitq), 
to_sfixed(-67.0/65536.0,1,-nbitq), 
to_sfixed(794.0/65536.0,1,-nbitq), 
to_sfixed(-3161.0/65536.0,1,-nbitq), 
to_sfixed(-4610.0/65536.0,1,-nbitq), 
to_sfixed(-638.0/65536.0,1,-nbitq), 
to_sfixed(3000.0/65536.0,1,-nbitq), 
to_sfixed(1339.0/65536.0,1,-nbitq), 
to_sfixed(5053.0/65536.0,1,-nbitq)  ), 
( to_sfixed(956.0/65536.0,1,-nbitq), 
to_sfixed(-2304.0/65536.0,1,-nbitq), 
to_sfixed(1022.0/65536.0,1,-nbitq), 
to_sfixed(1767.0/65536.0,1,-nbitq), 
to_sfixed(-2839.0/65536.0,1,-nbitq), 
to_sfixed(156.0/65536.0,1,-nbitq), 
to_sfixed(-362.0/65536.0,1,-nbitq), 
to_sfixed(2609.0/65536.0,1,-nbitq), 
to_sfixed(-3950.0/65536.0,1,-nbitq), 
to_sfixed(51.0/65536.0,1,-nbitq), 
to_sfixed(-2398.0/65536.0,1,-nbitq), 
to_sfixed(-3862.0/65536.0,1,-nbitq), 
to_sfixed(-187.0/65536.0,1,-nbitq), 
to_sfixed(1180.0/65536.0,1,-nbitq), 
to_sfixed(-1058.0/65536.0,1,-nbitq), 
to_sfixed(415.0/65536.0,1,-nbitq), 
to_sfixed(-2360.0/65536.0,1,-nbitq), 
to_sfixed(-556.0/65536.0,1,-nbitq), 
to_sfixed(256.0/65536.0,1,-nbitq), 
to_sfixed(199.0/65536.0,1,-nbitq), 
to_sfixed(-2774.0/65536.0,1,-nbitq), 
to_sfixed(-2489.0/65536.0,1,-nbitq), 
to_sfixed(2175.0/65536.0,1,-nbitq), 
to_sfixed(1204.0/65536.0,1,-nbitq), 
to_sfixed(2628.0/65536.0,1,-nbitq), 
to_sfixed(1258.0/65536.0,1,-nbitq), 
to_sfixed(-5606.0/65536.0,1,-nbitq), 
to_sfixed(-2962.0/65536.0,1,-nbitq), 
to_sfixed(-2465.0/65536.0,1,-nbitq), 
to_sfixed(-1441.0/65536.0,1,-nbitq), 
to_sfixed(5360.0/65536.0,1,-nbitq), 
to_sfixed(2667.0/65536.0,1,-nbitq), 
to_sfixed(-3598.0/65536.0,1,-nbitq), 
to_sfixed(-2120.0/65536.0,1,-nbitq), 
to_sfixed(-1700.0/65536.0,1,-nbitq), 
to_sfixed(3003.0/65536.0,1,-nbitq), 
to_sfixed(-886.0/65536.0,1,-nbitq), 
to_sfixed(-536.0/65536.0,1,-nbitq), 
to_sfixed(-1827.0/65536.0,1,-nbitq), 
to_sfixed(2970.0/65536.0,1,-nbitq), 
to_sfixed(2130.0/65536.0,1,-nbitq), 
to_sfixed(960.0/65536.0,1,-nbitq), 
to_sfixed(-1644.0/65536.0,1,-nbitq), 
to_sfixed(4701.0/65536.0,1,-nbitq), 
to_sfixed(847.0/65536.0,1,-nbitq), 
to_sfixed(468.0/65536.0,1,-nbitq), 
to_sfixed(2887.0/65536.0,1,-nbitq), 
to_sfixed(-1994.0/65536.0,1,-nbitq), 
to_sfixed(-1107.0/65536.0,1,-nbitq), 
to_sfixed(194.0/65536.0,1,-nbitq), 
to_sfixed(2772.0/65536.0,1,-nbitq), 
to_sfixed(1657.0/65536.0,1,-nbitq), 
to_sfixed(5148.0/65536.0,1,-nbitq), 
to_sfixed(-4189.0/65536.0,1,-nbitq), 
to_sfixed(1045.0/65536.0,1,-nbitq), 
to_sfixed(-2069.0/65536.0,1,-nbitq), 
to_sfixed(2600.0/65536.0,1,-nbitq), 
to_sfixed(362.0/65536.0,1,-nbitq), 
to_sfixed(-33.0/65536.0,1,-nbitq), 
to_sfixed(3890.0/65536.0,1,-nbitq), 
to_sfixed(-994.0/65536.0,1,-nbitq), 
to_sfixed(532.0/65536.0,1,-nbitq), 
to_sfixed(-873.0/65536.0,1,-nbitq), 
to_sfixed(-1514.0/65536.0,1,-nbitq), 
to_sfixed(3283.0/65536.0,1,-nbitq), 
to_sfixed(-147.0/65536.0,1,-nbitq), 
to_sfixed(512.0/65536.0,1,-nbitq), 
to_sfixed(-4206.0/65536.0,1,-nbitq), 
to_sfixed(6634.0/65536.0,1,-nbitq), 
to_sfixed(474.0/65536.0,1,-nbitq), 
to_sfixed(-935.0/65536.0,1,-nbitq), 
to_sfixed(965.0/65536.0,1,-nbitq), 
to_sfixed(-1911.0/65536.0,1,-nbitq), 
to_sfixed(124.0/65536.0,1,-nbitq), 
to_sfixed(-2973.0/65536.0,1,-nbitq), 
to_sfixed(-3849.0/65536.0,1,-nbitq), 
to_sfixed(-3713.0/65536.0,1,-nbitq), 
to_sfixed(2361.0/65536.0,1,-nbitq), 
to_sfixed(1459.0/65536.0,1,-nbitq), 
to_sfixed(2679.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3011.0/65536.0,1,-nbitq), 
to_sfixed(-1634.0/65536.0,1,-nbitq), 
to_sfixed(-1382.0/65536.0,1,-nbitq), 
to_sfixed(-2152.0/65536.0,1,-nbitq), 
to_sfixed(-3082.0/65536.0,1,-nbitq), 
to_sfixed(-3124.0/65536.0,1,-nbitq), 
to_sfixed(1967.0/65536.0,1,-nbitq), 
to_sfixed(116.0/65536.0,1,-nbitq), 
to_sfixed(-3428.0/65536.0,1,-nbitq), 
to_sfixed(522.0/65536.0,1,-nbitq), 
to_sfixed(877.0/65536.0,1,-nbitq), 
to_sfixed(-2920.0/65536.0,1,-nbitq), 
to_sfixed(1253.0/65536.0,1,-nbitq), 
to_sfixed(441.0/65536.0,1,-nbitq), 
to_sfixed(469.0/65536.0,1,-nbitq), 
to_sfixed(-503.0/65536.0,1,-nbitq), 
to_sfixed(-740.0/65536.0,1,-nbitq), 
to_sfixed(828.0/65536.0,1,-nbitq), 
to_sfixed(887.0/65536.0,1,-nbitq), 
to_sfixed(-1205.0/65536.0,1,-nbitq), 
to_sfixed(-1541.0/65536.0,1,-nbitq), 
to_sfixed(-2459.0/65536.0,1,-nbitq), 
to_sfixed(1042.0/65536.0,1,-nbitq), 
to_sfixed(-1233.0/65536.0,1,-nbitq), 
to_sfixed(2186.0/65536.0,1,-nbitq), 
to_sfixed(3274.0/65536.0,1,-nbitq), 
to_sfixed(-4036.0/65536.0,1,-nbitq), 
to_sfixed(2480.0/65536.0,1,-nbitq), 
to_sfixed(756.0/65536.0,1,-nbitq), 
to_sfixed(1403.0/65536.0,1,-nbitq), 
to_sfixed(1168.0/65536.0,1,-nbitq), 
to_sfixed(-2023.0/65536.0,1,-nbitq), 
to_sfixed(-4188.0/65536.0,1,-nbitq), 
to_sfixed(-4034.0/65536.0,1,-nbitq), 
to_sfixed(-1525.0/65536.0,1,-nbitq), 
to_sfixed(1558.0/65536.0,1,-nbitq), 
to_sfixed(-3104.0/65536.0,1,-nbitq), 
to_sfixed(-128.0/65536.0,1,-nbitq), 
to_sfixed(-2718.0/65536.0,1,-nbitq), 
to_sfixed(-836.0/65536.0,1,-nbitq), 
to_sfixed(3125.0/65536.0,1,-nbitq), 
to_sfixed(-3264.0/65536.0,1,-nbitq), 
to_sfixed(-4628.0/65536.0,1,-nbitq), 
to_sfixed(1046.0/65536.0,1,-nbitq), 
to_sfixed(2402.0/65536.0,1,-nbitq), 
to_sfixed(-15.0/65536.0,1,-nbitq), 
to_sfixed(2897.0/65536.0,1,-nbitq), 
to_sfixed(2153.0/65536.0,1,-nbitq), 
to_sfixed(-328.0/65536.0,1,-nbitq), 
to_sfixed(4612.0/65536.0,1,-nbitq), 
to_sfixed(-1830.0/65536.0,1,-nbitq), 
to_sfixed(1968.0/65536.0,1,-nbitq), 
to_sfixed(3331.0/65536.0,1,-nbitq), 
to_sfixed(-1846.0/65536.0,1,-nbitq), 
to_sfixed(517.0/65536.0,1,-nbitq), 
to_sfixed(-1654.0/65536.0,1,-nbitq), 
to_sfixed(-1984.0/65536.0,1,-nbitq), 
to_sfixed(924.0/65536.0,1,-nbitq), 
to_sfixed(1642.0/65536.0,1,-nbitq), 
to_sfixed(3505.0/65536.0,1,-nbitq), 
to_sfixed(-538.0/65536.0,1,-nbitq), 
to_sfixed(2399.0/65536.0,1,-nbitq), 
to_sfixed(725.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(3667.0/65536.0,1,-nbitq), 
to_sfixed(-833.0/65536.0,1,-nbitq), 
to_sfixed(3814.0/65536.0,1,-nbitq), 
to_sfixed(1140.0/65536.0,1,-nbitq), 
to_sfixed(1301.0/65536.0,1,-nbitq), 
to_sfixed(1432.0/65536.0,1,-nbitq), 
to_sfixed(-251.0/65536.0,1,-nbitq), 
to_sfixed(-1034.0/65536.0,1,-nbitq), 
to_sfixed(-132.0/65536.0,1,-nbitq), 
to_sfixed(2286.0/65536.0,1,-nbitq), 
to_sfixed(-305.0/65536.0,1,-nbitq), 
to_sfixed(468.0/65536.0,1,-nbitq), 
to_sfixed(602.0/65536.0,1,-nbitq), 
to_sfixed(471.0/65536.0,1,-nbitq), 
to_sfixed(1462.0/65536.0,1,-nbitq), 
to_sfixed(2806.0/65536.0,1,-nbitq)  ), 
( to_sfixed(572.0/65536.0,1,-nbitq), 
to_sfixed(195.0/65536.0,1,-nbitq), 
to_sfixed(2046.0/65536.0,1,-nbitq), 
to_sfixed(-2774.0/65536.0,1,-nbitq), 
to_sfixed(-6054.0/65536.0,1,-nbitq), 
to_sfixed(-3714.0/65536.0,1,-nbitq), 
to_sfixed(-827.0/65536.0,1,-nbitq), 
to_sfixed(-821.0/65536.0,1,-nbitq), 
to_sfixed(-2079.0/65536.0,1,-nbitq), 
to_sfixed(79.0/65536.0,1,-nbitq), 
to_sfixed(-2962.0/65536.0,1,-nbitq), 
to_sfixed(1266.0/65536.0,1,-nbitq), 
to_sfixed(2389.0/65536.0,1,-nbitq), 
to_sfixed(-185.0/65536.0,1,-nbitq), 
to_sfixed(-3261.0/65536.0,1,-nbitq), 
to_sfixed(2652.0/65536.0,1,-nbitq), 
to_sfixed(1026.0/65536.0,1,-nbitq), 
to_sfixed(-1350.0/65536.0,1,-nbitq), 
to_sfixed(4332.0/65536.0,1,-nbitq), 
to_sfixed(-635.0/65536.0,1,-nbitq), 
to_sfixed(394.0/65536.0,1,-nbitq), 
to_sfixed(39.0/65536.0,1,-nbitq), 
to_sfixed(1166.0/65536.0,1,-nbitq), 
to_sfixed(1351.0/65536.0,1,-nbitq), 
to_sfixed(249.0/65536.0,1,-nbitq), 
to_sfixed(-1045.0/65536.0,1,-nbitq), 
to_sfixed(-1967.0/65536.0,1,-nbitq), 
to_sfixed(-2235.0/65536.0,1,-nbitq), 
to_sfixed(-2346.0/65536.0,1,-nbitq), 
to_sfixed(-1162.0/65536.0,1,-nbitq), 
to_sfixed(2477.0/65536.0,1,-nbitq), 
to_sfixed(2917.0/65536.0,1,-nbitq), 
to_sfixed(75.0/65536.0,1,-nbitq), 
to_sfixed(-287.0/65536.0,1,-nbitq), 
to_sfixed(1565.0/65536.0,1,-nbitq), 
to_sfixed(-1834.0/65536.0,1,-nbitq), 
to_sfixed(-3808.0/65536.0,1,-nbitq), 
to_sfixed(-1796.0/65536.0,1,-nbitq), 
to_sfixed(-701.0/65536.0,1,-nbitq), 
to_sfixed(906.0/65536.0,1,-nbitq), 
to_sfixed(-685.0/65536.0,1,-nbitq), 
to_sfixed(537.0/65536.0,1,-nbitq), 
to_sfixed(-165.0/65536.0,1,-nbitq), 
to_sfixed(327.0/65536.0,1,-nbitq), 
to_sfixed(-922.0/65536.0,1,-nbitq), 
to_sfixed(-400.0/65536.0,1,-nbitq), 
to_sfixed(229.0/65536.0,1,-nbitq), 
to_sfixed(1452.0/65536.0,1,-nbitq), 
to_sfixed(-725.0/65536.0,1,-nbitq), 
to_sfixed(3530.0/65536.0,1,-nbitq), 
to_sfixed(38.0/65536.0,1,-nbitq), 
to_sfixed(660.0/65536.0,1,-nbitq), 
to_sfixed(5590.0/65536.0,1,-nbitq), 
to_sfixed(-913.0/65536.0,1,-nbitq), 
to_sfixed(3692.0/65536.0,1,-nbitq), 
to_sfixed(-2433.0/65536.0,1,-nbitq), 
to_sfixed(2535.0/65536.0,1,-nbitq), 
to_sfixed(-2629.0/65536.0,1,-nbitq), 
to_sfixed(-2465.0/65536.0,1,-nbitq), 
to_sfixed(3182.0/65536.0,1,-nbitq), 
to_sfixed(-1192.0/65536.0,1,-nbitq), 
to_sfixed(-1262.0/65536.0,1,-nbitq), 
to_sfixed(1958.0/65536.0,1,-nbitq), 
to_sfixed(-1595.0/65536.0,1,-nbitq), 
to_sfixed(2976.0/65536.0,1,-nbitq), 
to_sfixed(213.0/65536.0,1,-nbitq), 
to_sfixed(740.0/65536.0,1,-nbitq), 
to_sfixed(282.0/65536.0,1,-nbitq), 
to_sfixed(2896.0/65536.0,1,-nbitq), 
to_sfixed(-3593.0/65536.0,1,-nbitq), 
to_sfixed(-2604.0/65536.0,1,-nbitq), 
to_sfixed(-912.0/65536.0,1,-nbitq), 
to_sfixed(1867.0/65536.0,1,-nbitq), 
to_sfixed(-2073.0/65536.0,1,-nbitq), 
to_sfixed(-228.0/65536.0,1,-nbitq), 
to_sfixed(285.0/65536.0,1,-nbitq), 
to_sfixed(2144.0/65536.0,1,-nbitq), 
to_sfixed(4930.0/65536.0,1,-nbitq), 
to_sfixed(-2698.0/65536.0,1,-nbitq), 
to_sfixed(4602.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1652.0/65536.0,1,-nbitq), 
to_sfixed(347.0/65536.0,1,-nbitq), 
to_sfixed(4244.0/65536.0,1,-nbitq), 
to_sfixed(-1447.0/65536.0,1,-nbitq), 
to_sfixed(-1012.0/65536.0,1,-nbitq), 
to_sfixed(-4374.0/65536.0,1,-nbitq), 
to_sfixed(-593.0/65536.0,1,-nbitq), 
to_sfixed(-2164.0/65536.0,1,-nbitq), 
to_sfixed(-1839.0/65536.0,1,-nbitq), 
to_sfixed(-1834.0/65536.0,1,-nbitq), 
to_sfixed(-481.0/65536.0,1,-nbitq), 
to_sfixed(-243.0/65536.0,1,-nbitq), 
to_sfixed(-999.0/65536.0,1,-nbitq), 
to_sfixed(-3490.0/65536.0,1,-nbitq), 
to_sfixed(-2739.0/65536.0,1,-nbitq), 
to_sfixed(-2510.0/65536.0,1,-nbitq), 
to_sfixed(-2755.0/65536.0,1,-nbitq), 
to_sfixed(-1685.0/65536.0,1,-nbitq), 
to_sfixed(4196.0/65536.0,1,-nbitq), 
to_sfixed(1899.0/65536.0,1,-nbitq), 
to_sfixed(203.0/65536.0,1,-nbitq), 
to_sfixed(-2650.0/65536.0,1,-nbitq), 
to_sfixed(-1961.0/65536.0,1,-nbitq), 
to_sfixed(89.0/65536.0,1,-nbitq), 
to_sfixed(2294.0/65536.0,1,-nbitq), 
to_sfixed(3785.0/65536.0,1,-nbitq), 
to_sfixed(1312.0/65536.0,1,-nbitq), 
to_sfixed(-880.0/65536.0,1,-nbitq), 
to_sfixed(-2500.0/65536.0,1,-nbitq), 
to_sfixed(-2893.0/65536.0,1,-nbitq), 
to_sfixed(2874.0/65536.0,1,-nbitq), 
to_sfixed(1819.0/65536.0,1,-nbitq), 
to_sfixed(-4749.0/65536.0,1,-nbitq), 
to_sfixed(-3255.0/65536.0,1,-nbitq), 
to_sfixed(-2699.0/65536.0,1,-nbitq), 
to_sfixed(673.0/65536.0,1,-nbitq), 
to_sfixed(1022.0/65536.0,1,-nbitq), 
to_sfixed(1528.0/65536.0,1,-nbitq), 
to_sfixed(457.0/65536.0,1,-nbitq), 
to_sfixed(-284.0/65536.0,1,-nbitq), 
to_sfixed(-1430.0/65536.0,1,-nbitq), 
to_sfixed(-2995.0/65536.0,1,-nbitq), 
to_sfixed(-489.0/65536.0,1,-nbitq), 
to_sfixed(-920.0/65536.0,1,-nbitq), 
to_sfixed(-2604.0/65536.0,1,-nbitq), 
to_sfixed(1261.0/65536.0,1,-nbitq), 
to_sfixed(2755.0/65536.0,1,-nbitq), 
to_sfixed(1114.0/65536.0,1,-nbitq), 
to_sfixed(-107.0/65536.0,1,-nbitq), 
to_sfixed(3864.0/65536.0,1,-nbitq), 
to_sfixed(1443.0/65536.0,1,-nbitq), 
to_sfixed(1028.0/65536.0,1,-nbitq), 
to_sfixed(903.0/65536.0,1,-nbitq), 
to_sfixed(1353.0/65536.0,1,-nbitq), 
to_sfixed(2834.0/65536.0,1,-nbitq), 
to_sfixed(-2732.0/65536.0,1,-nbitq), 
to_sfixed(-1976.0/65536.0,1,-nbitq), 
to_sfixed(181.0/65536.0,1,-nbitq), 
to_sfixed(324.0/65536.0,1,-nbitq), 
to_sfixed(1414.0/65536.0,1,-nbitq), 
to_sfixed(-873.0/65536.0,1,-nbitq), 
to_sfixed(-800.0/65536.0,1,-nbitq), 
to_sfixed(-2031.0/65536.0,1,-nbitq), 
to_sfixed(2353.0/65536.0,1,-nbitq), 
to_sfixed(743.0/65536.0,1,-nbitq), 
to_sfixed(2794.0/65536.0,1,-nbitq), 
to_sfixed(-1338.0/65536.0,1,-nbitq), 
to_sfixed(-1991.0/65536.0,1,-nbitq), 
to_sfixed(-517.0/65536.0,1,-nbitq), 
to_sfixed(-1681.0/65536.0,1,-nbitq), 
to_sfixed(2041.0/65536.0,1,-nbitq), 
to_sfixed(2594.0/65536.0,1,-nbitq), 
to_sfixed(-610.0/65536.0,1,-nbitq), 
to_sfixed(-89.0/65536.0,1,-nbitq), 
to_sfixed(-1407.0/65536.0,1,-nbitq), 
to_sfixed(2459.0/65536.0,1,-nbitq), 
to_sfixed(-3012.0/65536.0,1,-nbitq), 
to_sfixed(4778.0/65536.0,1,-nbitq), 
to_sfixed(-2138.0/65536.0,1,-nbitq), 
to_sfixed(3699.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2056.0/65536.0,1,-nbitq), 
to_sfixed(-1994.0/65536.0,1,-nbitq), 
to_sfixed(-266.0/65536.0,1,-nbitq), 
to_sfixed(2216.0/65536.0,1,-nbitq), 
to_sfixed(-1396.0/65536.0,1,-nbitq), 
to_sfixed(-745.0/65536.0,1,-nbitq), 
to_sfixed(-3171.0/65536.0,1,-nbitq), 
to_sfixed(-1563.0/65536.0,1,-nbitq), 
to_sfixed(1695.0/65536.0,1,-nbitq), 
to_sfixed(-129.0/65536.0,1,-nbitq), 
to_sfixed(-3964.0/65536.0,1,-nbitq), 
to_sfixed(-1167.0/65536.0,1,-nbitq), 
to_sfixed(1766.0/65536.0,1,-nbitq), 
to_sfixed(1385.0/65536.0,1,-nbitq), 
to_sfixed(-775.0/65536.0,1,-nbitq), 
to_sfixed(-1416.0/65536.0,1,-nbitq), 
to_sfixed(1908.0/65536.0,1,-nbitq), 
to_sfixed(834.0/65536.0,1,-nbitq), 
to_sfixed(1350.0/65536.0,1,-nbitq), 
to_sfixed(-1427.0/65536.0,1,-nbitq), 
to_sfixed(-3367.0/65536.0,1,-nbitq), 
to_sfixed(2228.0/65536.0,1,-nbitq), 
to_sfixed(2809.0/65536.0,1,-nbitq), 
to_sfixed(927.0/65536.0,1,-nbitq), 
to_sfixed(1880.0/65536.0,1,-nbitq), 
to_sfixed(3745.0/65536.0,1,-nbitq), 
to_sfixed(1246.0/65536.0,1,-nbitq), 
to_sfixed(2210.0/65536.0,1,-nbitq), 
to_sfixed(344.0/65536.0,1,-nbitq), 
to_sfixed(-2713.0/65536.0,1,-nbitq), 
to_sfixed(-1635.0/65536.0,1,-nbitq), 
to_sfixed(-511.0/65536.0,1,-nbitq), 
to_sfixed(-5613.0/65536.0,1,-nbitq), 
to_sfixed(-3970.0/65536.0,1,-nbitq), 
to_sfixed(2894.0/65536.0,1,-nbitq), 
to_sfixed(-1402.0/65536.0,1,-nbitq), 
to_sfixed(-113.0/65536.0,1,-nbitq), 
to_sfixed(-500.0/65536.0,1,-nbitq), 
to_sfixed(968.0/65536.0,1,-nbitq), 
to_sfixed(-533.0/65536.0,1,-nbitq), 
to_sfixed(294.0/65536.0,1,-nbitq), 
to_sfixed(-2083.0/65536.0,1,-nbitq), 
to_sfixed(-4762.0/65536.0,1,-nbitq), 
to_sfixed(1923.0/65536.0,1,-nbitq), 
to_sfixed(1481.0/65536.0,1,-nbitq), 
to_sfixed(1589.0/65536.0,1,-nbitq), 
to_sfixed(554.0/65536.0,1,-nbitq), 
to_sfixed(-787.0/65536.0,1,-nbitq), 
to_sfixed(2413.0/65536.0,1,-nbitq), 
to_sfixed(898.0/65536.0,1,-nbitq), 
to_sfixed(1581.0/65536.0,1,-nbitq), 
to_sfixed(1182.0/65536.0,1,-nbitq), 
to_sfixed(3113.0/65536.0,1,-nbitq), 
to_sfixed(-2558.0/65536.0,1,-nbitq), 
to_sfixed(1768.0/65536.0,1,-nbitq), 
to_sfixed(-2176.0/65536.0,1,-nbitq), 
to_sfixed(416.0/65536.0,1,-nbitq), 
to_sfixed(2548.0/65536.0,1,-nbitq), 
to_sfixed(-2955.0/65536.0,1,-nbitq), 
to_sfixed(1792.0/65536.0,1,-nbitq), 
to_sfixed(103.0/65536.0,1,-nbitq), 
to_sfixed(1907.0/65536.0,1,-nbitq), 
to_sfixed(172.0/65536.0,1,-nbitq), 
to_sfixed(2607.0/65536.0,1,-nbitq), 
to_sfixed(168.0/65536.0,1,-nbitq), 
to_sfixed(-414.0/65536.0,1,-nbitq), 
to_sfixed(248.0/65536.0,1,-nbitq), 
to_sfixed(-3234.0/65536.0,1,-nbitq), 
to_sfixed(-1392.0/65536.0,1,-nbitq), 
to_sfixed(-1153.0/65536.0,1,-nbitq), 
to_sfixed(1839.0/65536.0,1,-nbitq), 
to_sfixed(1027.0/65536.0,1,-nbitq), 
to_sfixed(4214.0/65536.0,1,-nbitq), 
to_sfixed(1322.0/65536.0,1,-nbitq), 
to_sfixed(257.0/65536.0,1,-nbitq), 
to_sfixed(831.0/65536.0,1,-nbitq), 
to_sfixed(-1486.0/65536.0,1,-nbitq), 
to_sfixed(3982.0/65536.0,1,-nbitq), 
to_sfixed(-2623.0/65536.0,1,-nbitq), 
to_sfixed(-187.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1005.0/65536.0,1,-nbitq), 
to_sfixed(-1288.0/65536.0,1,-nbitq), 
to_sfixed(1909.0/65536.0,1,-nbitq), 
to_sfixed(-1992.0/65536.0,1,-nbitq), 
to_sfixed(1066.0/65536.0,1,-nbitq), 
to_sfixed(-2626.0/65536.0,1,-nbitq), 
to_sfixed(501.0/65536.0,1,-nbitq), 
to_sfixed(3009.0/65536.0,1,-nbitq), 
to_sfixed(-2469.0/65536.0,1,-nbitq), 
to_sfixed(-81.0/65536.0,1,-nbitq), 
to_sfixed(-3424.0/65536.0,1,-nbitq), 
to_sfixed(422.0/65536.0,1,-nbitq), 
to_sfixed(2284.0/65536.0,1,-nbitq), 
to_sfixed(-3246.0/65536.0,1,-nbitq), 
to_sfixed(496.0/65536.0,1,-nbitq), 
to_sfixed(518.0/65536.0,1,-nbitq), 
to_sfixed(1004.0/65536.0,1,-nbitq), 
to_sfixed(-68.0/65536.0,1,-nbitq), 
to_sfixed(1905.0/65536.0,1,-nbitq), 
to_sfixed(-1348.0/65536.0,1,-nbitq), 
to_sfixed(-343.0/65536.0,1,-nbitq), 
to_sfixed(998.0/65536.0,1,-nbitq), 
to_sfixed(-349.0/65536.0,1,-nbitq), 
to_sfixed(-402.0/65536.0,1,-nbitq), 
to_sfixed(-739.0/65536.0,1,-nbitq), 
to_sfixed(1034.0/65536.0,1,-nbitq), 
to_sfixed(-2341.0/65536.0,1,-nbitq), 
to_sfixed(2173.0/65536.0,1,-nbitq), 
to_sfixed(-3451.0/65536.0,1,-nbitq), 
to_sfixed(-2425.0/65536.0,1,-nbitq), 
to_sfixed(2575.0/65536.0,1,-nbitq), 
to_sfixed(1024.0/65536.0,1,-nbitq), 
to_sfixed(-1339.0/65536.0,1,-nbitq), 
to_sfixed(382.0/65536.0,1,-nbitq), 
to_sfixed(-2740.0/65536.0,1,-nbitq), 
to_sfixed(-834.0/65536.0,1,-nbitq), 
to_sfixed(1130.0/65536.0,1,-nbitq), 
to_sfixed(-3272.0/65536.0,1,-nbitq), 
to_sfixed(-1062.0/65536.0,1,-nbitq), 
to_sfixed(-1085.0/65536.0,1,-nbitq), 
to_sfixed(1037.0/65536.0,1,-nbitq), 
to_sfixed(1764.0/65536.0,1,-nbitq), 
to_sfixed(-2676.0/65536.0,1,-nbitq), 
to_sfixed(677.0/65536.0,1,-nbitq), 
to_sfixed(3121.0/65536.0,1,-nbitq), 
to_sfixed(-241.0/65536.0,1,-nbitq), 
to_sfixed(-485.0/65536.0,1,-nbitq), 
to_sfixed(756.0/65536.0,1,-nbitq), 
to_sfixed(1274.0/65536.0,1,-nbitq), 
to_sfixed(-864.0/65536.0,1,-nbitq), 
to_sfixed(-1712.0/65536.0,1,-nbitq), 
to_sfixed(1301.0/65536.0,1,-nbitq), 
to_sfixed(-1339.0/65536.0,1,-nbitq), 
to_sfixed(-3171.0/65536.0,1,-nbitq), 
to_sfixed(-1574.0/65536.0,1,-nbitq), 
to_sfixed(-1695.0/65536.0,1,-nbitq), 
to_sfixed(219.0/65536.0,1,-nbitq), 
to_sfixed(2764.0/65536.0,1,-nbitq), 
to_sfixed(1426.0/65536.0,1,-nbitq), 
to_sfixed(665.0/65536.0,1,-nbitq), 
to_sfixed(-4078.0/65536.0,1,-nbitq), 
to_sfixed(807.0/65536.0,1,-nbitq), 
to_sfixed(58.0/65536.0,1,-nbitq), 
to_sfixed(-427.0/65536.0,1,-nbitq), 
to_sfixed(-977.0/65536.0,1,-nbitq), 
to_sfixed(-50.0/65536.0,1,-nbitq), 
to_sfixed(2780.0/65536.0,1,-nbitq), 
to_sfixed(-1157.0/65536.0,1,-nbitq), 
to_sfixed(2399.0/65536.0,1,-nbitq), 
to_sfixed(-1668.0/65536.0,1,-nbitq), 
to_sfixed(-2168.0/65536.0,1,-nbitq), 
to_sfixed(-1378.0/65536.0,1,-nbitq), 
to_sfixed(1736.0/65536.0,1,-nbitq), 
to_sfixed(658.0/65536.0,1,-nbitq), 
to_sfixed(2449.0/65536.0,1,-nbitq), 
to_sfixed(-1156.0/65536.0,1,-nbitq), 
to_sfixed(-1868.0/65536.0,1,-nbitq), 
to_sfixed(2147.0/65536.0,1,-nbitq), 
to_sfixed(-1232.0/65536.0,1,-nbitq), 
to_sfixed(-269.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1391.0/65536.0,1,-nbitq), 
to_sfixed(-1379.0/65536.0,1,-nbitq), 
to_sfixed(2743.0/65536.0,1,-nbitq), 
to_sfixed(-677.0/65536.0,1,-nbitq), 
to_sfixed(-2478.0/65536.0,1,-nbitq), 
to_sfixed(-1612.0/65536.0,1,-nbitq), 
to_sfixed(-2500.0/65536.0,1,-nbitq), 
to_sfixed(-1692.0/65536.0,1,-nbitq), 
to_sfixed(558.0/65536.0,1,-nbitq), 
to_sfixed(828.0/65536.0,1,-nbitq), 
to_sfixed(813.0/65536.0,1,-nbitq), 
to_sfixed(-1518.0/65536.0,1,-nbitq), 
to_sfixed(-2929.0/65536.0,1,-nbitq), 
to_sfixed(-140.0/65536.0,1,-nbitq), 
to_sfixed(-1221.0/65536.0,1,-nbitq), 
to_sfixed(2171.0/65536.0,1,-nbitq), 
to_sfixed(1025.0/65536.0,1,-nbitq), 
to_sfixed(671.0/65536.0,1,-nbitq), 
to_sfixed(-41.0/65536.0,1,-nbitq), 
to_sfixed(-2174.0/65536.0,1,-nbitq), 
to_sfixed(2092.0/65536.0,1,-nbitq), 
to_sfixed(1120.0/65536.0,1,-nbitq), 
to_sfixed(-1791.0/65536.0,1,-nbitq), 
to_sfixed(-1355.0/65536.0,1,-nbitq), 
to_sfixed(-2176.0/65536.0,1,-nbitq), 
to_sfixed(1424.0/65536.0,1,-nbitq), 
to_sfixed(-3344.0/65536.0,1,-nbitq), 
to_sfixed(-227.0/65536.0,1,-nbitq), 
to_sfixed(-15.0/65536.0,1,-nbitq), 
to_sfixed(-3215.0/65536.0,1,-nbitq), 
to_sfixed(-330.0/65536.0,1,-nbitq), 
to_sfixed(1329.0/65536.0,1,-nbitq), 
to_sfixed(-2286.0/65536.0,1,-nbitq), 
to_sfixed(2547.0/65536.0,1,-nbitq), 
to_sfixed(-1382.0/65536.0,1,-nbitq), 
to_sfixed(-806.0/65536.0,1,-nbitq), 
to_sfixed(2386.0/65536.0,1,-nbitq), 
to_sfixed(1434.0/65536.0,1,-nbitq), 
to_sfixed(-3116.0/65536.0,1,-nbitq), 
to_sfixed(182.0/65536.0,1,-nbitq), 
to_sfixed(-1520.0/65536.0,1,-nbitq), 
to_sfixed(-1464.0/65536.0,1,-nbitq), 
to_sfixed(-4295.0/65536.0,1,-nbitq), 
to_sfixed(-146.0/65536.0,1,-nbitq), 
to_sfixed(-1666.0/65536.0,1,-nbitq), 
to_sfixed(2406.0/65536.0,1,-nbitq), 
to_sfixed(-2310.0/65536.0,1,-nbitq), 
to_sfixed(4527.0/65536.0,1,-nbitq), 
to_sfixed(-1515.0/65536.0,1,-nbitq), 
to_sfixed(-589.0/65536.0,1,-nbitq), 
to_sfixed(1697.0/65536.0,1,-nbitq), 
to_sfixed(1591.0/65536.0,1,-nbitq), 
to_sfixed(-110.0/65536.0,1,-nbitq), 
to_sfixed(-4337.0/65536.0,1,-nbitq), 
to_sfixed(-1796.0/65536.0,1,-nbitq), 
to_sfixed(-454.0/65536.0,1,-nbitq), 
to_sfixed(1869.0/65536.0,1,-nbitq), 
to_sfixed(151.0/65536.0,1,-nbitq), 
to_sfixed(-2787.0/65536.0,1,-nbitq), 
to_sfixed(4646.0/65536.0,1,-nbitq), 
to_sfixed(-1338.0/65536.0,1,-nbitq), 
to_sfixed(-489.0/65536.0,1,-nbitq), 
to_sfixed(364.0/65536.0,1,-nbitq), 
to_sfixed(-242.0/65536.0,1,-nbitq), 
to_sfixed(640.0/65536.0,1,-nbitq), 
to_sfixed(1560.0/65536.0,1,-nbitq), 
to_sfixed(-1346.0/65536.0,1,-nbitq), 
to_sfixed(1218.0/65536.0,1,-nbitq), 
to_sfixed(252.0/65536.0,1,-nbitq), 
to_sfixed(-356.0/65536.0,1,-nbitq), 
to_sfixed(-1106.0/65536.0,1,-nbitq), 
to_sfixed(-799.0/65536.0,1,-nbitq), 
to_sfixed(-1574.0/65536.0,1,-nbitq), 
to_sfixed(2244.0/65536.0,1,-nbitq), 
to_sfixed(-107.0/65536.0,1,-nbitq), 
to_sfixed(2687.0/65536.0,1,-nbitq), 
to_sfixed(277.0/65536.0,1,-nbitq), 
to_sfixed(1556.0/65536.0,1,-nbitq), 
to_sfixed(-1198.0/65536.0,1,-nbitq), 
to_sfixed(5922.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-664.0/65536.0,1,-nbitq), 
to_sfixed(756.0/65536.0,1,-nbitq), 
to_sfixed(3473.0/65536.0,1,-nbitq), 
to_sfixed(713.0/65536.0,1,-nbitq), 
to_sfixed(-12.0/65536.0,1,-nbitq), 
to_sfixed(-4161.0/65536.0,1,-nbitq), 
to_sfixed(45.0/65536.0,1,-nbitq), 
to_sfixed(-2514.0/65536.0,1,-nbitq), 
to_sfixed(3150.0/65536.0,1,-nbitq), 
to_sfixed(-1885.0/65536.0,1,-nbitq), 
to_sfixed(1758.0/65536.0,1,-nbitq), 
to_sfixed(-2034.0/65536.0,1,-nbitq), 
to_sfixed(-2226.0/65536.0,1,-nbitq), 
to_sfixed(-1009.0/65536.0,1,-nbitq), 
to_sfixed(2815.0/65536.0,1,-nbitq), 
to_sfixed(593.0/65536.0,1,-nbitq), 
to_sfixed(-769.0/65536.0,1,-nbitq), 
to_sfixed(-1628.0/65536.0,1,-nbitq), 
to_sfixed(847.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(-3440.0/65536.0,1,-nbitq), 
to_sfixed(2930.0/65536.0,1,-nbitq), 
to_sfixed(2984.0/65536.0,1,-nbitq), 
to_sfixed(2103.0/65536.0,1,-nbitq), 
to_sfixed(2561.0/65536.0,1,-nbitq), 
to_sfixed(-1137.0/65536.0,1,-nbitq), 
to_sfixed(-4539.0/65536.0,1,-nbitq), 
to_sfixed(-338.0/65536.0,1,-nbitq), 
to_sfixed(-2270.0/65536.0,1,-nbitq), 
to_sfixed(-76.0/65536.0,1,-nbitq), 
to_sfixed(2341.0/65536.0,1,-nbitq), 
to_sfixed(1808.0/65536.0,1,-nbitq), 
to_sfixed(-2107.0/65536.0,1,-nbitq), 
to_sfixed(302.0/65536.0,1,-nbitq), 
to_sfixed(-938.0/65536.0,1,-nbitq), 
to_sfixed(1641.0/65536.0,1,-nbitq), 
to_sfixed(561.0/65536.0,1,-nbitq), 
to_sfixed(-3756.0/65536.0,1,-nbitq), 
to_sfixed(-307.0/65536.0,1,-nbitq), 
to_sfixed(667.0/65536.0,1,-nbitq), 
to_sfixed(-2598.0/65536.0,1,-nbitq), 
to_sfixed(-3306.0/65536.0,1,-nbitq), 
to_sfixed(-2244.0/65536.0,1,-nbitq), 
to_sfixed(2315.0/65536.0,1,-nbitq), 
to_sfixed(-468.0/65536.0,1,-nbitq), 
to_sfixed(1878.0/65536.0,1,-nbitq), 
to_sfixed(375.0/65536.0,1,-nbitq), 
to_sfixed(155.0/65536.0,1,-nbitq), 
to_sfixed(451.0/65536.0,1,-nbitq), 
to_sfixed(-1928.0/65536.0,1,-nbitq), 
to_sfixed(-1532.0/65536.0,1,-nbitq), 
to_sfixed(-416.0/65536.0,1,-nbitq), 
to_sfixed(3194.0/65536.0,1,-nbitq), 
to_sfixed(-2998.0/65536.0,1,-nbitq), 
to_sfixed(2284.0/65536.0,1,-nbitq), 
to_sfixed(2010.0/65536.0,1,-nbitq), 
to_sfixed(2254.0/65536.0,1,-nbitq), 
to_sfixed(-2161.0/65536.0,1,-nbitq), 
to_sfixed(665.0/65536.0,1,-nbitq), 
to_sfixed(3908.0/65536.0,1,-nbitq), 
to_sfixed(-371.0/65536.0,1,-nbitq), 
to_sfixed(398.0/65536.0,1,-nbitq), 
to_sfixed(-2635.0/65536.0,1,-nbitq), 
to_sfixed(-2263.0/65536.0,1,-nbitq), 
to_sfixed(378.0/65536.0,1,-nbitq), 
to_sfixed(694.0/65536.0,1,-nbitq), 
to_sfixed(-1201.0/65536.0,1,-nbitq), 
to_sfixed(-4506.0/65536.0,1,-nbitq), 
to_sfixed(4992.0/65536.0,1,-nbitq), 
to_sfixed(-1295.0/65536.0,1,-nbitq), 
to_sfixed(3391.0/65536.0,1,-nbitq), 
to_sfixed(1575.0/65536.0,1,-nbitq), 
to_sfixed(-173.0/65536.0,1,-nbitq), 
to_sfixed(-199.0/65536.0,1,-nbitq), 
to_sfixed(1049.0/65536.0,1,-nbitq), 
to_sfixed(317.0/65536.0,1,-nbitq), 
to_sfixed(-2505.0/65536.0,1,-nbitq), 
to_sfixed(2219.0/65536.0,1,-nbitq), 
to_sfixed(-1888.0/65536.0,1,-nbitq), 
to_sfixed(2630.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2368.0/65536.0,1,-nbitq), 
to_sfixed(-1465.0/65536.0,1,-nbitq), 
to_sfixed(5582.0/65536.0,1,-nbitq), 
to_sfixed(-2347.0/65536.0,1,-nbitq), 
to_sfixed(1078.0/65536.0,1,-nbitq), 
to_sfixed(-4994.0/65536.0,1,-nbitq), 
to_sfixed(-2719.0/65536.0,1,-nbitq), 
to_sfixed(1610.0/65536.0,1,-nbitq), 
to_sfixed(3762.0/65536.0,1,-nbitq), 
to_sfixed(240.0/65536.0,1,-nbitq), 
to_sfixed(-2384.0/65536.0,1,-nbitq), 
to_sfixed(-827.0/65536.0,1,-nbitq), 
to_sfixed(-2237.0/65536.0,1,-nbitq), 
to_sfixed(-1447.0/65536.0,1,-nbitq), 
to_sfixed(-318.0/65536.0,1,-nbitq), 
to_sfixed(2763.0/65536.0,1,-nbitq), 
to_sfixed(-4.0/65536.0,1,-nbitq), 
to_sfixed(-1126.0/65536.0,1,-nbitq), 
to_sfixed(-1552.0/65536.0,1,-nbitq), 
to_sfixed(-268.0/65536.0,1,-nbitq), 
to_sfixed(228.0/65536.0,1,-nbitq), 
to_sfixed(2885.0/65536.0,1,-nbitq), 
to_sfixed(-1055.0/65536.0,1,-nbitq), 
to_sfixed(-3874.0/65536.0,1,-nbitq), 
to_sfixed(-1361.0/65536.0,1,-nbitq), 
to_sfixed(-1487.0/65536.0,1,-nbitq), 
to_sfixed(-882.0/65536.0,1,-nbitq), 
to_sfixed(-1361.0/65536.0,1,-nbitq), 
to_sfixed(-4753.0/65536.0,1,-nbitq), 
to_sfixed(920.0/65536.0,1,-nbitq), 
to_sfixed(-790.0/65536.0,1,-nbitq), 
to_sfixed(-2545.0/65536.0,1,-nbitq), 
to_sfixed(-2895.0/65536.0,1,-nbitq), 
to_sfixed(1345.0/65536.0,1,-nbitq), 
to_sfixed(1135.0/65536.0,1,-nbitq), 
to_sfixed(-2620.0/65536.0,1,-nbitq), 
to_sfixed(1794.0/65536.0,1,-nbitq), 
to_sfixed(-773.0/65536.0,1,-nbitq), 
to_sfixed(-1142.0/65536.0,1,-nbitq), 
to_sfixed(1251.0/65536.0,1,-nbitq), 
to_sfixed(79.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(-2836.0/65536.0,1,-nbitq), 
to_sfixed(2986.0/65536.0,1,-nbitq), 
to_sfixed(684.0/65536.0,1,-nbitq), 
to_sfixed(179.0/65536.0,1,-nbitq), 
to_sfixed(1652.0/65536.0,1,-nbitq), 
to_sfixed(642.0/65536.0,1,-nbitq), 
to_sfixed(-1917.0/65536.0,1,-nbitq), 
to_sfixed(-430.0/65536.0,1,-nbitq), 
to_sfixed(-759.0/65536.0,1,-nbitq), 
to_sfixed(-1786.0/65536.0,1,-nbitq), 
to_sfixed(225.0/65536.0,1,-nbitq), 
to_sfixed(-1712.0/65536.0,1,-nbitq), 
to_sfixed(1433.0/65536.0,1,-nbitq), 
to_sfixed(1930.0/65536.0,1,-nbitq), 
to_sfixed(-1186.0/65536.0,1,-nbitq), 
to_sfixed(3226.0/65536.0,1,-nbitq), 
to_sfixed(-1926.0/65536.0,1,-nbitq), 
to_sfixed(4012.0/65536.0,1,-nbitq), 
to_sfixed(-1900.0/65536.0,1,-nbitq), 
to_sfixed(-1805.0/65536.0,1,-nbitq), 
to_sfixed(2090.0/65536.0,1,-nbitq), 
to_sfixed(-1258.0/65536.0,1,-nbitq), 
to_sfixed(1826.0/65536.0,1,-nbitq), 
to_sfixed(-74.0/65536.0,1,-nbitq), 
to_sfixed(2719.0/65536.0,1,-nbitq), 
to_sfixed(-4202.0/65536.0,1,-nbitq), 
to_sfixed(64.0/65536.0,1,-nbitq), 
to_sfixed(62.0/65536.0,1,-nbitq), 
to_sfixed(2064.0/65536.0,1,-nbitq), 
to_sfixed(1567.0/65536.0,1,-nbitq), 
to_sfixed(1708.0/65536.0,1,-nbitq), 
to_sfixed(2289.0/65536.0,1,-nbitq), 
to_sfixed(370.0/65536.0,1,-nbitq), 
to_sfixed(4222.0/65536.0,1,-nbitq), 
to_sfixed(1129.0/65536.0,1,-nbitq), 
to_sfixed(-532.0/65536.0,1,-nbitq), 
to_sfixed(-120.0/65536.0,1,-nbitq), 
to_sfixed(5084.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1652.0/65536.0,1,-nbitq), 
to_sfixed(636.0/65536.0,1,-nbitq), 
to_sfixed(6295.0/65536.0,1,-nbitq), 
to_sfixed(-3348.0/65536.0,1,-nbitq), 
to_sfixed(1017.0/65536.0,1,-nbitq), 
to_sfixed(-2175.0/65536.0,1,-nbitq), 
to_sfixed(-2377.0/65536.0,1,-nbitq), 
to_sfixed(-2508.0/65536.0,1,-nbitq), 
to_sfixed(717.0/65536.0,1,-nbitq), 
to_sfixed(763.0/65536.0,1,-nbitq), 
to_sfixed(-2017.0/65536.0,1,-nbitq), 
to_sfixed(-4604.0/65536.0,1,-nbitq), 
to_sfixed(665.0/65536.0,1,-nbitq), 
to_sfixed(-4802.0/65536.0,1,-nbitq), 
to_sfixed(1376.0/65536.0,1,-nbitq), 
to_sfixed(-2559.0/65536.0,1,-nbitq), 
to_sfixed(277.0/65536.0,1,-nbitq), 
to_sfixed(726.0/65536.0,1,-nbitq), 
to_sfixed(-2891.0/65536.0,1,-nbitq), 
to_sfixed(681.0/65536.0,1,-nbitq), 
to_sfixed(3829.0/65536.0,1,-nbitq), 
to_sfixed(-949.0/65536.0,1,-nbitq), 
to_sfixed(3888.0/65536.0,1,-nbitq), 
to_sfixed(-4319.0/65536.0,1,-nbitq), 
to_sfixed(2002.0/65536.0,1,-nbitq), 
to_sfixed(-2403.0/65536.0,1,-nbitq), 
to_sfixed(689.0/65536.0,1,-nbitq), 
to_sfixed(1310.0/65536.0,1,-nbitq), 
to_sfixed(-4216.0/65536.0,1,-nbitq), 
to_sfixed(1217.0/65536.0,1,-nbitq), 
to_sfixed(-1108.0/65536.0,1,-nbitq), 
to_sfixed(2285.0/65536.0,1,-nbitq), 
to_sfixed(463.0/65536.0,1,-nbitq), 
to_sfixed(4089.0/65536.0,1,-nbitq), 
to_sfixed(2639.0/65536.0,1,-nbitq), 
to_sfixed(-2750.0/65536.0,1,-nbitq), 
to_sfixed(1641.0/65536.0,1,-nbitq), 
to_sfixed(1186.0/65536.0,1,-nbitq), 
to_sfixed(-3453.0/65536.0,1,-nbitq), 
to_sfixed(2471.0/65536.0,1,-nbitq), 
to_sfixed(3518.0/65536.0,1,-nbitq), 
to_sfixed(-2622.0/65536.0,1,-nbitq), 
to_sfixed(-1714.0/65536.0,1,-nbitq), 
to_sfixed(2143.0/65536.0,1,-nbitq), 
to_sfixed(1897.0/65536.0,1,-nbitq), 
to_sfixed(-17.0/65536.0,1,-nbitq), 
to_sfixed(2235.0/65536.0,1,-nbitq), 
to_sfixed(-1227.0/65536.0,1,-nbitq), 
to_sfixed(2466.0/65536.0,1,-nbitq), 
to_sfixed(3680.0/65536.0,1,-nbitq), 
to_sfixed(-1403.0/65536.0,1,-nbitq), 
to_sfixed(-2171.0/65536.0,1,-nbitq), 
to_sfixed(2444.0/65536.0,1,-nbitq), 
to_sfixed(-8174.0/65536.0,1,-nbitq), 
to_sfixed(2114.0/65536.0,1,-nbitq), 
to_sfixed(1260.0/65536.0,1,-nbitq), 
to_sfixed(1389.0/65536.0,1,-nbitq), 
to_sfixed(-1304.0/65536.0,1,-nbitq), 
to_sfixed(181.0/65536.0,1,-nbitq), 
to_sfixed(1705.0/65536.0,1,-nbitq), 
to_sfixed(-321.0/65536.0,1,-nbitq), 
to_sfixed(370.0/65536.0,1,-nbitq), 
to_sfixed(1957.0/65536.0,1,-nbitq), 
to_sfixed(1647.0/65536.0,1,-nbitq), 
to_sfixed(1947.0/65536.0,1,-nbitq), 
to_sfixed(-3958.0/65536.0,1,-nbitq), 
to_sfixed(306.0/65536.0,1,-nbitq), 
to_sfixed(-2233.0/65536.0,1,-nbitq), 
to_sfixed(892.0/65536.0,1,-nbitq), 
to_sfixed(1952.0/65536.0,1,-nbitq), 
to_sfixed(-2621.0/65536.0,1,-nbitq), 
to_sfixed(567.0/65536.0,1,-nbitq), 
to_sfixed(-907.0/65536.0,1,-nbitq), 
to_sfixed(-1832.0/65536.0,1,-nbitq), 
to_sfixed(1170.0/65536.0,1,-nbitq), 
to_sfixed(338.0/65536.0,1,-nbitq), 
to_sfixed(-3035.0/65536.0,1,-nbitq), 
to_sfixed(71.0/65536.0,1,-nbitq), 
to_sfixed(-1939.0/65536.0,1,-nbitq), 
to_sfixed(5642.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1015.0/65536.0,1,-nbitq), 
to_sfixed(2293.0/65536.0,1,-nbitq), 
to_sfixed(4990.0/65536.0,1,-nbitq), 
to_sfixed(-586.0/65536.0,1,-nbitq), 
to_sfixed(4402.0/65536.0,1,-nbitq), 
to_sfixed(-1545.0/65536.0,1,-nbitq), 
to_sfixed(1370.0/65536.0,1,-nbitq), 
to_sfixed(313.0/65536.0,1,-nbitq), 
to_sfixed(-184.0/65536.0,1,-nbitq), 
to_sfixed(1950.0/65536.0,1,-nbitq), 
to_sfixed(-1675.0/65536.0,1,-nbitq), 
to_sfixed(-11383.0/65536.0,1,-nbitq), 
to_sfixed(3255.0/65536.0,1,-nbitq), 
to_sfixed(-2084.0/65536.0,1,-nbitq), 
to_sfixed(-1733.0/65536.0,1,-nbitq), 
to_sfixed(-2719.0/65536.0,1,-nbitq), 
to_sfixed(-2195.0/65536.0,1,-nbitq), 
to_sfixed(-58.0/65536.0,1,-nbitq), 
to_sfixed(-1045.0/65536.0,1,-nbitq), 
to_sfixed(2067.0/65536.0,1,-nbitq), 
to_sfixed(5053.0/65536.0,1,-nbitq), 
to_sfixed(3764.0/65536.0,1,-nbitq), 
to_sfixed(2320.0/65536.0,1,-nbitq), 
to_sfixed(-5144.0/65536.0,1,-nbitq), 
to_sfixed(-649.0/65536.0,1,-nbitq), 
to_sfixed(-2880.0/65536.0,1,-nbitq), 
to_sfixed(-855.0/65536.0,1,-nbitq), 
to_sfixed(923.0/65536.0,1,-nbitq), 
to_sfixed(-2762.0/65536.0,1,-nbitq), 
to_sfixed(783.0/65536.0,1,-nbitq), 
to_sfixed(-697.0/65536.0,1,-nbitq), 
to_sfixed(-2465.0/65536.0,1,-nbitq), 
to_sfixed(-258.0/65536.0,1,-nbitq), 
to_sfixed(3683.0/65536.0,1,-nbitq), 
to_sfixed(2646.0/65536.0,1,-nbitq), 
to_sfixed(-1820.0/65536.0,1,-nbitq), 
to_sfixed(6113.0/65536.0,1,-nbitq), 
to_sfixed(-2942.0/65536.0,1,-nbitq), 
to_sfixed(4899.0/65536.0,1,-nbitq), 
to_sfixed(-2524.0/65536.0,1,-nbitq), 
to_sfixed(-1296.0/65536.0,1,-nbitq), 
to_sfixed(1868.0/65536.0,1,-nbitq), 
to_sfixed(2621.0/65536.0,1,-nbitq), 
to_sfixed(3555.0/65536.0,1,-nbitq), 
to_sfixed(3169.0/65536.0,1,-nbitq), 
to_sfixed(-1169.0/65536.0,1,-nbitq), 
to_sfixed(2583.0/65536.0,1,-nbitq), 
to_sfixed(1443.0/65536.0,1,-nbitq), 
to_sfixed(2158.0/65536.0,1,-nbitq), 
to_sfixed(-1478.0/65536.0,1,-nbitq), 
to_sfixed(-1775.0/65536.0,1,-nbitq), 
to_sfixed(2633.0/65536.0,1,-nbitq), 
to_sfixed(690.0/65536.0,1,-nbitq), 
to_sfixed(-1257.0/65536.0,1,-nbitq), 
to_sfixed(201.0/65536.0,1,-nbitq), 
to_sfixed(-5688.0/65536.0,1,-nbitq), 
to_sfixed(-505.0/65536.0,1,-nbitq), 
to_sfixed(-1856.0/65536.0,1,-nbitq), 
to_sfixed(549.0/65536.0,1,-nbitq), 
to_sfixed(-7275.0/65536.0,1,-nbitq), 
to_sfixed(-6594.0/65536.0,1,-nbitq), 
to_sfixed(-738.0/65536.0,1,-nbitq), 
to_sfixed(-175.0/65536.0,1,-nbitq), 
to_sfixed(611.0/65536.0,1,-nbitq), 
to_sfixed(-1972.0/65536.0,1,-nbitq), 
to_sfixed(-5052.0/65536.0,1,-nbitq), 
to_sfixed(3324.0/65536.0,1,-nbitq), 
to_sfixed(230.0/65536.0,1,-nbitq), 
to_sfixed(2685.0/65536.0,1,-nbitq), 
to_sfixed(4575.0/65536.0,1,-nbitq), 
to_sfixed(-1799.0/65536.0,1,-nbitq), 
to_sfixed(-1326.0/65536.0,1,-nbitq), 
to_sfixed(-1063.0/65536.0,1,-nbitq), 
to_sfixed(1486.0/65536.0,1,-nbitq), 
to_sfixed(1055.0/65536.0,1,-nbitq), 
to_sfixed(4898.0/65536.0,1,-nbitq), 
to_sfixed(-1283.0/65536.0,1,-nbitq), 
to_sfixed(3954.0/65536.0,1,-nbitq), 
to_sfixed(-621.0/65536.0,1,-nbitq), 
to_sfixed(3350.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3523.0/65536.0,1,-nbitq), 
to_sfixed(5240.0/65536.0,1,-nbitq), 
to_sfixed(1470.0/65536.0,1,-nbitq), 
to_sfixed(-1682.0/65536.0,1,-nbitq), 
to_sfixed(-933.0/65536.0,1,-nbitq), 
to_sfixed(-6340.0/65536.0,1,-nbitq), 
to_sfixed(673.0/65536.0,1,-nbitq), 
to_sfixed(897.0/65536.0,1,-nbitq), 
to_sfixed(2515.0/65536.0,1,-nbitq), 
to_sfixed(-297.0/65536.0,1,-nbitq), 
to_sfixed(-842.0/65536.0,1,-nbitq), 
to_sfixed(-7760.0/65536.0,1,-nbitq), 
to_sfixed(2370.0/65536.0,1,-nbitq), 
to_sfixed(-8327.0/65536.0,1,-nbitq), 
to_sfixed(-1779.0/65536.0,1,-nbitq), 
to_sfixed(1796.0/65536.0,1,-nbitq), 
to_sfixed(2292.0/65536.0,1,-nbitq), 
to_sfixed(445.0/65536.0,1,-nbitq), 
to_sfixed(-3552.0/65536.0,1,-nbitq), 
to_sfixed(-2701.0/65536.0,1,-nbitq), 
to_sfixed(5357.0/65536.0,1,-nbitq), 
to_sfixed(-1386.0/65536.0,1,-nbitq), 
to_sfixed(637.0/65536.0,1,-nbitq), 
to_sfixed(-9488.0/65536.0,1,-nbitq), 
to_sfixed(447.0/65536.0,1,-nbitq), 
to_sfixed(-8668.0/65536.0,1,-nbitq), 
to_sfixed(52.0/65536.0,1,-nbitq), 
to_sfixed(-4318.0/65536.0,1,-nbitq), 
to_sfixed(-5636.0/65536.0,1,-nbitq), 
to_sfixed(-897.0/65536.0,1,-nbitq), 
to_sfixed(-2302.0/65536.0,1,-nbitq), 
to_sfixed(-617.0/65536.0,1,-nbitq), 
to_sfixed(7760.0/65536.0,1,-nbitq), 
to_sfixed(4112.0/65536.0,1,-nbitq), 
to_sfixed(275.0/65536.0,1,-nbitq), 
to_sfixed(785.0/65536.0,1,-nbitq), 
to_sfixed(6711.0/65536.0,1,-nbitq), 
to_sfixed(-2437.0/65536.0,1,-nbitq), 
to_sfixed(5182.0/65536.0,1,-nbitq), 
to_sfixed(-2551.0/65536.0,1,-nbitq), 
to_sfixed(-2031.0/65536.0,1,-nbitq), 
to_sfixed(991.0/65536.0,1,-nbitq), 
to_sfixed(6964.0/65536.0,1,-nbitq), 
to_sfixed(-2151.0/65536.0,1,-nbitq), 
to_sfixed(-2275.0/65536.0,1,-nbitq), 
to_sfixed(-702.0/65536.0,1,-nbitq), 
to_sfixed(988.0/65536.0,1,-nbitq), 
to_sfixed(3337.0/65536.0,1,-nbitq), 
to_sfixed(-99.0/65536.0,1,-nbitq), 
to_sfixed(931.0/65536.0,1,-nbitq), 
to_sfixed(-624.0/65536.0,1,-nbitq), 
to_sfixed(196.0/65536.0,1,-nbitq), 
to_sfixed(3390.0/65536.0,1,-nbitq), 
to_sfixed(3982.0/65536.0,1,-nbitq), 
to_sfixed(-628.0/65536.0,1,-nbitq), 
to_sfixed(-1688.0/65536.0,1,-nbitq), 
to_sfixed(-2006.0/65536.0,1,-nbitq), 
to_sfixed(-1711.0/65536.0,1,-nbitq), 
to_sfixed(-762.0/65536.0,1,-nbitq), 
to_sfixed(-9074.0/65536.0,1,-nbitq), 
to_sfixed(-393.0/65536.0,1,-nbitq), 
to_sfixed(-2254.0/65536.0,1,-nbitq), 
to_sfixed(1354.0/65536.0,1,-nbitq), 
to_sfixed(-1228.0/65536.0,1,-nbitq), 
to_sfixed(-3870.0/65536.0,1,-nbitq), 
to_sfixed(-2510.0/65536.0,1,-nbitq), 
to_sfixed(5106.0/65536.0,1,-nbitq), 
to_sfixed(-1330.0/65536.0,1,-nbitq), 
to_sfixed(2595.0/65536.0,1,-nbitq), 
to_sfixed(7955.0/65536.0,1,-nbitq), 
to_sfixed(-1535.0/65536.0,1,-nbitq), 
to_sfixed(550.0/65536.0,1,-nbitq), 
to_sfixed(1472.0/65536.0,1,-nbitq), 
to_sfixed(231.0/65536.0,1,-nbitq), 
to_sfixed(-3080.0/65536.0,1,-nbitq), 
to_sfixed(4189.0/65536.0,1,-nbitq), 
to_sfixed(-5033.0/65536.0,1,-nbitq), 
to_sfixed(3892.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(1161.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3879.0/65536.0,1,-nbitq), 
to_sfixed(815.0/65536.0,1,-nbitq), 
to_sfixed(1036.0/65536.0,1,-nbitq), 
to_sfixed(2091.0/65536.0,1,-nbitq), 
to_sfixed(669.0/65536.0,1,-nbitq), 
to_sfixed(-10927.0/65536.0,1,-nbitq), 
to_sfixed(2697.0/65536.0,1,-nbitq), 
to_sfixed(-1556.0/65536.0,1,-nbitq), 
to_sfixed(1240.0/65536.0,1,-nbitq), 
to_sfixed(-1022.0/65536.0,1,-nbitq), 
to_sfixed(1558.0/65536.0,1,-nbitq), 
to_sfixed(-10752.0/65536.0,1,-nbitq), 
to_sfixed(3597.0/65536.0,1,-nbitq), 
to_sfixed(-8828.0/65536.0,1,-nbitq), 
to_sfixed(-1613.0/65536.0,1,-nbitq), 
to_sfixed(-2775.0/65536.0,1,-nbitq), 
to_sfixed(716.0/65536.0,1,-nbitq), 
to_sfixed(6230.0/65536.0,1,-nbitq), 
to_sfixed(-8095.0/65536.0,1,-nbitq), 
to_sfixed(1737.0/65536.0,1,-nbitq), 
to_sfixed(5059.0/65536.0,1,-nbitq), 
to_sfixed(-3084.0/65536.0,1,-nbitq), 
to_sfixed(658.0/65536.0,1,-nbitq), 
to_sfixed(-15436.0/65536.0,1,-nbitq), 
to_sfixed(2104.0/65536.0,1,-nbitq), 
to_sfixed(-10994.0/65536.0,1,-nbitq), 
to_sfixed(867.0/65536.0,1,-nbitq), 
to_sfixed(-2358.0/65536.0,1,-nbitq), 
to_sfixed(-5020.0/65536.0,1,-nbitq), 
to_sfixed(-1797.0/65536.0,1,-nbitq), 
to_sfixed(-91.0/65536.0,1,-nbitq), 
to_sfixed(-3461.0/65536.0,1,-nbitq), 
to_sfixed(4858.0/65536.0,1,-nbitq), 
to_sfixed(-1115.0/65536.0,1,-nbitq), 
to_sfixed(2429.0/65536.0,1,-nbitq), 
to_sfixed(-324.0/65536.0,1,-nbitq), 
to_sfixed(8837.0/65536.0,1,-nbitq), 
to_sfixed(2723.0/65536.0,1,-nbitq), 
to_sfixed(2423.0/65536.0,1,-nbitq), 
to_sfixed(-5183.0/65536.0,1,-nbitq), 
to_sfixed(-887.0/65536.0,1,-nbitq), 
to_sfixed(505.0/65536.0,1,-nbitq), 
to_sfixed(7916.0/65536.0,1,-nbitq), 
to_sfixed(1305.0/65536.0,1,-nbitq), 
to_sfixed(-880.0/65536.0,1,-nbitq), 
to_sfixed(-1606.0/65536.0,1,-nbitq), 
to_sfixed(-696.0/65536.0,1,-nbitq), 
to_sfixed(3638.0/65536.0,1,-nbitq), 
to_sfixed(-1113.0/65536.0,1,-nbitq), 
to_sfixed(2547.0/65536.0,1,-nbitq), 
to_sfixed(2202.0/65536.0,1,-nbitq), 
to_sfixed(-1322.0/65536.0,1,-nbitq), 
to_sfixed(5064.0/65536.0,1,-nbitq), 
to_sfixed(-1735.0/65536.0,1,-nbitq), 
to_sfixed(292.0/65536.0,1,-nbitq), 
to_sfixed(-3243.0/65536.0,1,-nbitq), 
to_sfixed(869.0/65536.0,1,-nbitq), 
to_sfixed(3422.0/65536.0,1,-nbitq), 
to_sfixed(1336.0/65536.0,1,-nbitq), 
to_sfixed(-7622.0/65536.0,1,-nbitq), 
to_sfixed(6781.0/65536.0,1,-nbitq), 
to_sfixed(1237.0/65536.0,1,-nbitq), 
to_sfixed(-24.0/65536.0,1,-nbitq), 
to_sfixed(1786.0/65536.0,1,-nbitq), 
to_sfixed(-3979.0/65536.0,1,-nbitq), 
to_sfixed(681.0/65536.0,1,-nbitq), 
to_sfixed(5997.0/65536.0,1,-nbitq), 
to_sfixed(-2564.0/65536.0,1,-nbitq), 
to_sfixed(-1247.0/65536.0,1,-nbitq), 
to_sfixed(3410.0/65536.0,1,-nbitq), 
to_sfixed(1557.0/65536.0,1,-nbitq), 
to_sfixed(-5319.0/65536.0,1,-nbitq), 
to_sfixed(-1203.0/65536.0,1,-nbitq), 
to_sfixed(2691.0/65536.0,1,-nbitq), 
to_sfixed(859.0/65536.0,1,-nbitq), 
to_sfixed(1695.0/65536.0,1,-nbitq), 
to_sfixed(333.0/65536.0,1,-nbitq), 
to_sfixed(612.0/65536.0,1,-nbitq), 
to_sfixed(-1807.0/65536.0,1,-nbitq), 
to_sfixed(3658.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3174.0/65536.0,1,-nbitq), 
to_sfixed(3977.0/65536.0,1,-nbitq), 
to_sfixed(5740.0/65536.0,1,-nbitq), 
to_sfixed(-4222.0/65536.0,1,-nbitq), 
to_sfixed(-1208.0/65536.0,1,-nbitq), 
to_sfixed(-5844.0/65536.0,1,-nbitq), 
to_sfixed(-4616.0/65536.0,1,-nbitq), 
to_sfixed(-1207.0/65536.0,1,-nbitq), 
to_sfixed(-1202.0/65536.0,1,-nbitq), 
to_sfixed(845.0/65536.0,1,-nbitq), 
to_sfixed(4965.0/65536.0,1,-nbitq), 
to_sfixed(-10065.0/65536.0,1,-nbitq), 
to_sfixed(-1499.0/65536.0,1,-nbitq), 
to_sfixed(-5280.0/65536.0,1,-nbitq), 
to_sfixed(2519.0/65536.0,1,-nbitq), 
to_sfixed(1580.0/65536.0,1,-nbitq), 
to_sfixed(1018.0/65536.0,1,-nbitq), 
to_sfixed(2321.0/65536.0,1,-nbitq), 
to_sfixed(-3649.0/65536.0,1,-nbitq), 
to_sfixed(1001.0/65536.0,1,-nbitq), 
to_sfixed(5942.0/65536.0,1,-nbitq), 
to_sfixed(-3170.0/65536.0,1,-nbitq), 
to_sfixed(-764.0/65536.0,1,-nbitq), 
to_sfixed(-14682.0/65536.0,1,-nbitq), 
to_sfixed(-1205.0/65536.0,1,-nbitq), 
to_sfixed(-9540.0/65536.0,1,-nbitq), 
to_sfixed(5910.0/65536.0,1,-nbitq), 
to_sfixed(-509.0/65536.0,1,-nbitq), 
to_sfixed(-2213.0/65536.0,1,-nbitq), 
to_sfixed(-805.0/65536.0,1,-nbitq), 
to_sfixed(3320.0/65536.0,1,-nbitq), 
to_sfixed(-3441.0/65536.0,1,-nbitq), 
to_sfixed(1105.0/65536.0,1,-nbitq), 
to_sfixed(-1608.0/65536.0,1,-nbitq), 
to_sfixed(466.0/65536.0,1,-nbitq), 
to_sfixed(-480.0/65536.0,1,-nbitq), 
to_sfixed(5252.0/65536.0,1,-nbitq), 
to_sfixed(-363.0/65536.0,1,-nbitq), 
to_sfixed(719.0/65536.0,1,-nbitq), 
to_sfixed(-3539.0/65536.0,1,-nbitq), 
to_sfixed(-4659.0/65536.0,1,-nbitq), 
to_sfixed(2422.0/65536.0,1,-nbitq), 
to_sfixed(8327.0/65536.0,1,-nbitq), 
to_sfixed(3835.0/65536.0,1,-nbitq), 
to_sfixed(-880.0/65536.0,1,-nbitq), 
to_sfixed(-7973.0/65536.0,1,-nbitq), 
to_sfixed(996.0/65536.0,1,-nbitq), 
to_sfixed(-963.0/65536.0,1,-nbitq), 
to_sfixed(1081.0/65536.0,1,-nbitq), 
to_sfixed(2478.0/65536.0,1,-nbitq), 
to_sfixed(-2017.0/65536.0,1,-nbitq), 
to_sfixed(1419.0/65536.0,1,-nbitq), 
to_sfixed(8305.0/65536.0,1,-nbitq), 
to_sfixed(-4949.0/65536.0,1,-nbitq), 
to_sfixed(-65.0/65536.0,1,-nbitq), 
to_sfixed(3742.0/65536.0,1,-nbitq), 
to_sfixed(-1909.0/65536.0,1,-nbitq), 
to_sfixed(864.0/65536.0,1,-nbitq), 
to_sfixed(423.0/65536.0,1,-nbitq), 
to_sfixed(-11213.0/65536.0,1,-nbitq), 
to_sfixed(3939.0/65536.0,1,-nbitq), 
to_sfixed(1785.0/65536.0,1,-nbitq), 
to_sfixed(-352.0/65536.0,1,-nbitq), 
to_sfixed(-804.0/65536.0,1,-nbitq), 
to_sfixed(-4449.0/65536.0,1,-nbitq), 
to_sfixed(2145.0/65536.0,1,-nbitq), 
to_sfixed(6093.0/65536.0,1,-nbitq), 
to_sfixed(-24.0/65536.0,1,-nbitq), 
to_sfixed(-4229.0/65536.0,1,-nbitq), 
to_sfixed(-250.0/65536.0,1,-nbitq), 
to_sfixed(4166.0/65536.0,1,-nbitq), 
to_sfixed(-2150.0/65536.0,1,-nbitq), 
to_sfixed(-1175.0/65536.0,1,-nbitq), 
to_sfixed(-277.0/65536.0,1,-nbitq), 
to_sfixed(-1380.0/65536.0,1,-nbitq), 
to_sfixed(270.0/65536.0,1,-nbitq), 
to_sfixed(3480.0/65536.0,1,-nbitq), 
to_sfixed(5625.0/65536.0,1,-nbitq), 
to_sfixed(-2096.0/65536.0,1,-nbitq), 
to_sfixed(1588.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1556.0/65536.0,1,-nbitq), 
to_sfixed(3332.0/65536.0,1,-nbitq), 
to_sfixed(11230.0/65536.0,1,-nbitq), 
to_sfixed(-5277.0/65536.0,1,-nbitq), 
to_sfixed(619.0/65536.0,1,-nbitq), 
to_sfixed(-3362.0/65536.0,1,-nbitq), 
to_sfixed(-5661.0/65536.0,1,-nbitq), 
to_sfixed(-3866.0/65536.0,1,-nbitq), 
to_sfixed(4230.0/65536.0,1,-nbitq), 
to_sfixed(-1603.0/65536.0,1,-nbitq), 
to_sfixed(1944.0/65536.0,1,-nbitq), 
to_sfixed(-10453.0/65536.0,1,-nbitq), 
to_sfixed(-1428.0/65536.0,1,-nbitq), 
to_sfixed(-3851.0/65536.0,1,-nbitq), 
to_sfixed(297.0/65536.0,1,-nbitq), 
to_sfixed(2704.0/65536.0,1,-nbitq), 
to_sfixed(-2314.0/65536.0,1,-nbitq), 
to_sfixed(4008.0/65536.0,1,-nbitq), 
to_sfixed(-813.0/65536.0,1,-nbitq), 
to_sfixed(-2736.0/65536.0,1,-nbitq), 
to_sfixed(-232.0/65536.0,1,-nbitq), 
to_sfixed(961.0/65536.0,1,-nbitq), 
to_sfixed(7350.0/65536.0,1,-nbitq), 
to_sfixed(-13332.0/65536.0,1,-nbitq), 
to_sfixed(-1147.0/65536.0,1,-nbitq), 
to_sfixed(-11205.0/65536.0,1,-nbitq), 
to_sfixed(9067.0/65536.0,1,-nbitq), 
to_sfixed(-3854.0/65536.0,1,-nbitq), 
to_sfixed(-5466.0/65536.0,1,-nbitq), 
to_sfixed(2132.0/65536.0,1,-nbitq), 
to_sfixed(5086.0/65536.0,1,-nbitq), 
to_sfixed(177.0/65536.0,1,-nbitq), 
to_sfixed(858.0/65536.0,1,-nbitq), 
to_sfixed(-1776.0/65536.0,1,-nbitq), 
to_sfixed(-1247.0/65536.0,1,-nbitq), 
to_sfixed(2868.0/65536.0,1,-nbitq), 
to_sfixed(5620.0/65536.0,1,-nbitq), 
to_sfixed(-3119.0/65536.0,1,-nbitq), 
to_sfixed(5002.0/65536.0,1,-nbitq), 
to_sfixed(60.0/65536.0,1,-nbitq), 
to_sfixed(-6379.0/65536.0,1,-nbitq), 
to_sfixed(-2641.0/65536.0,1,-nbitq), 
to_sfixed(478.0/65536.0,1,-nbitq), 
to_sfixed(1275.0/65536.0,1,-nbitq), 
to_sfixed(-1351.0/65536.0,1,-nbitq), 
to_sfixed(-5801.0/65536.0,1,-nbitq), 
to_sfixed(654.0/65536.0,1,-nbitq), 
to_sfixed(3730.0/65536.0,1,-nbitq), 
to_sfixed(1519.0/65536.0,1,-nbitq), 
to_sfixed(2099.0/65536.0,1,-nbitq), 
to_sfixed(-1242.0/65536.0,1,-nbitq), 
to_sfixed(-2443.0/65536.0,1,-nbitq), 
to_sfixed(2219.0/65536.0,1,-nbitq), 
to_sfixed(-86.0/65536.0,1,-nbitq), 
to_sfixed(-407.0/65536.0,1,-nbitq), 
to_sfixed(2154.0/65536.0,1,-nbitq), 
to_sfixed(2142.0/65536.0,1,-nbitq), 
to_sfixed(2109.0/65536.0,1,-nbitq), 
to_sfixed(1454.0/65536.0,1,-nbitq), 
to_sfixed(-9658.0/65536.0,1,-nbitq), 
to_sfixed(1613.0/65536.0,1,-nbitq), 
to_sfixed(1369.0/65536.0,1,-nbitq), 
to_sfixed(802.0/65536.0,1,-nbitq), 
to_sfixed(1534.0/65536.0,1,-nbitq), 
to_sfixed(2344.0/65536.0,1,-nbitq), 
to_sfixed(6145.0/65536.0,1,-nbitq), 
to_sfixed(274.0/65536.0,1,-nbitq), 
to_sfixed(308.0/65536.0,1,-nbitq), 
to_sfixed(-8189.0/65536.0,1,-nbitq), 
to_sfixed(2075.0/65536.0,1,-nbitq), 
to_sfixed(2305.0/65536.0,1,-nbitq), 
to_sfixed(1025.0/65536.0,1,-nbitq), 
to_sfixed(-3180.0/65536.0,1,-nbitq), 
to_sfixed(-122.0/65536.0,1,-nbitq), 
to_sfixed(-678.0/65536.0,1,-nbitq), 
to_sfixed(211.0/65536.0,1,-nbitq), 
to_sfixed(5812.0/65536.0,1,-nbitq), 
to_sfixed(3672.0/65536.0,1,-nbitq), 
to_sfixed(-1096.0/65536.0,1,-nbitq), 
to_sfixed(-1278.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-609.0/65536.0,1,-nbitq), 
to_sfixed(986.0/65536.0,1,-nbitq), 
to_sfixed(3464.0/65536.0,1,-nbitq), 
to_sfixed(648.0/65536.0,1,-nbitq), 
to_sfixed(1011.0/65536.0,1,-nbitq), 
to_sfixed(-4509.0/65536.0,1,-nbitq), 
to_sfixed(-3582.0/65536.0,1,-nbitq), 
to_sfixed(1807.0/65536.0,1,-nbitq), 
to_sfixed(2231.0/65536.0,1,-nbitq), 
to_sfixed(-1085.0/65536.0,1,-nbitq), 
to_sfixed(88.0/65536.0,1,-nbitq), 
to_sfixed(-9656.0/65536.0,1,-nbitq), 
to_sfixed(547.0/65536.0,1,-nbitq), 
to_sfixed(4723.0/65536.0,1,-nbitq), 
to_sfixed(-835.0/65536.0,1,-nbitq), 
to_sfixed(1901.0/65536.0,1,-nbitq), 
to_sfixed(2539.0/65536.0,1,-nbitq), 
to_sfixed(4089.0/65536.0,1,-nbitq), 
to_sfixed(226.0/65536.0,1,-nbitq), 
to_sfixed(1680.0/65536.0,1,-nbitq), 
to_sfixed(-2018.0/65536.0,1,-nbitq), 
to_sfixed(6076.0/65536.0,1,-nbitq), 
to_sfixed(5580.0/65536.0,1,-nbitq), 
to_sfixed(-1370.0/65536.0,1,-nbitq), 
to_sfixed(-2837.0/65536.0,1,-nbitq), 
to_sfixed(-7310.0/65536.0,1,-nbitq), 
to_sfixed(7781.0/65536.0,1,-nbitq), 
to_sfixed(-3262.0/65536.0,1,-nbitq), 
to_sfixed(-9641.0/65536.0,1,-nbitq), 
to_sfixed(6356.0/65536.0,1,-nbitq), 
to_sfixed(3312.0/65536.0,1,-nbitq), 
to_sfixed(-1371.0/65536.0,1,-nbitq), 
to_sfixed(-6590.0/65536.0,1,-nbitq), 
to_sfixed(-5540.0/65536.0,1,-nbitq), 
to_sfixed(1167.0/65536.0,1,-nbitq), 
to_sfixed(1072.0/65536.0,1,-nbitq), 
to_sfixed(1466.0/65536.0,1,-nbitq), 
to_sfixed(427.0/65536.0,1,-nbitq), 
to_sfixed(5731.0/65536.0,1,-nbitq), 
to_sfixed(1870.0/65536.0,1,-nbitq), 
to_sfixed(-5665.0/65536.0,1,-nbitq), 
to_sfixed(1009.0/65536.0,1,-nbitq), 
to_sfixed(-2995.0/65536.0,1,-nbitq), 
to_sfixed(3243.0/65536.0,1,-nbitq), 
to_sfixed(1137.0/65536.0,1,-nbitq), 
to_sfixed(-1411.0/65536.0,1,-nbitq), 
to_sfixed(-2968.0/65536.0,1,-nbitq), 
to_sfixed(1424.0/65536.0,1,-nbitq), 
to_sfixed(-986.0/65536.0,1,-nbitq), 
to_sfixed(4263.0/65536.0,1,-nbitq), 
to_sfixed(414.0/65536.0,1,-nbitq), 
to_sfixed(1758.0/65536.0,1,-nbitq), 
to_sfixed(971.0/65536.0,1,-nbitq), 
to_sfixed(-5481.0/65536.0,1,-nbitq), 
to_sfixed(-2526.0/65536.0,1,-nbitq), 
to_sfixed(-378.0/65536.0,1,-nbitq), 
to_sfixed(2506.0/65536.0,1,-nbitq), 
to_sfixed(-3626.0/65536.0,1,-nbitq), 
to_sfixed(-1833.0/65536.0,1,-nbitq), 
to_sfixed(-6470.0/65536.0,1,-nbitq), 
to_sfixed(-1337.0/65536.0,1,-nbitq), 
to_sfixed(1094.0/65536.0,1,-nbitq), 
to_sfixed(2308.0/65536.0,1,-nbitq), 
to_sfixed(928.0/65536.0,1,-nbitq), 
to_sfixed(-1665.0/65536.0,1,-nbitq), 
to_sfixed(7075.0/65536.0,1,-nbitq), 
to_sfixed(4102.0/65536.0,1,-nbitq), 
to_sfixed(2495.0/65536.0,1,-nbitq), 
to_sfixed(-6970.0/65536.0,1,-nbitq), 
to_sfixed(-544.0/65536.0,1,-nbitq), 
to_sfixed(-2247.0/65536.0,1,-nbitq), 
to_sfixed(1400.0/65536.0,1,-nbitq), 
to_sfixed(-4429.0/65536.0,1,-nbitq), 
to_sfixed(1350.0/65536.0,1,-nbitq), 
to_sfixed(-1288.0/65536.0,1,-nbitq), 
to_sfixed(-2495.0/65536.0,1,-nbitq), 
to_sfixed(8456.0/65536.0,1,-nbitq), 
to_sfixed(1370.0/65536.0,1,-nbitq), 
to_sfixed(2086.0/65536.0,1,-nbitq), 
to_sfixed(2376.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4259.0/65536.0,1,-nbitq), 
to_sfixed(-49.0/65536.0,1,-nbitq), 
to_sfixed(-6944.0/65536.0,1,-nbitq), 
to_sfixed(3615.0/65536.0,1,-nbitq), 
to_sfixed(3020.0/65536.0,1,-nbitq), 
to_sfixed(2120.0/65536.0,1,-nbitq), 
to_sfixed(-6115.0/65536.0,1,-nbitq), 
to_sfixed(5600.0/65536.0,1,-nbitq), 
to_sfixed(4925.0/65536.0,1,-nbitq), 
to_sfixed(-1323.0/65536.0,1,-nbitq), 
to_sfixed(-2714.0/65536.0,1,-nbitq), 
to_sfixed(-6038.0/65536.0,1,-nbitq), 
to_sfixed(-1468.0/65536.0,1,-nbitq), 
to_sfixed(10073.0/65536.0,1,-nbitq), 
to_sfixed(-2974.0/65536.0,1,-nbitq), 
to_sfixed(550.0/65536.0,1,-nbitq), 
to_sfixed(315.0/65536.0,1,-nbitq), 
to_sfixed(-3026.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(2276.0/65536.0,1,-nbitq), 
to_sfixed(-1301.0/65536.0,1,-nbitq), 
to_sfixed(9687.0/65536.0,1,-nbitq), 
to_sfixed(692.0/65536.0,1,-nbitq), 
to_sfixed(-1939.0/65536.0,1,-nbitq), 
to_sfixed(-4185.0/65536.0,1,-nbitq), 
to_sfixed(-6633.0/65536.0,1,-nbitq), 
to_sfixed(14586.0/65536.0,1,-nbitq), 
to_sfixed(-6140.0/65536.0,1,-nbitq), 
to_sfixed(370.0/65536.0,1,-nbitq), 
to_sfixed(131.0/65536.0,1,-nbitq), 
to_sfixed(2281.0/65536.0,1,-nbitq), 
to_sfixed(607.0/65536.0,1,-nbitq), 
to_sfixed(-4327.0/65536.0,1,-nbitq), 
to_sfixed(-2381.0/65536.0,1,-nbitq), 
to_sfixed(-1586.0/65536.0,1,-nbitq), 
to_sfixed(-1831.0/65536.0,1,-nbitq), 
to_sfixed(-6786.0/65536.0,1,-nbitq), 
to_sfixed(-1877.0/65536.0,1,-nbitq), 
to_sfixed(4450.0/65536.0,1,-nbitq), 
to_sfixed(1690.0/65536.0,1,-nbitq), 
to_sfixed(11.0/65536.0,1,-nbitq), 
to_sfixed(2717.0/65536.0,1,-nbitq), 
to_sfixed(15.0/65536.0,1,-nbitq), 
to_sfixed(3892.0/65536.0,1,-nbitq), 
to_sfixed(2970.0/65536.0,1,-nbitq), 
to_sfixed(-3443.0/65536.0,1,-nbitq), 
to_sfixed(-2127.0/65536.0,1,-nbitq), 
to_sfixed(5088.0/65536.0,1,-nbitq), 
to_sfixed(-2093.0/65536.0,1,-nbitq), 
to_sfixed(-625.0/65536.0,1,-nbitq), 
to_sfixed(-1518.0/65536.0,1,-nbitq), 
to_sfixed(-883.0/65536.0,1,-nbitq), 
to_sfixed(-720.0/65536.0,1,-nbitq), 
to_sfixed(-3566.0/65536.0,1,-nbitq), 
to_sfixed(2330.0/65536.0,1,-nbitq), 
to_sfixed(-6038.0/65536.0,1,-nbitq), 
to_sfixed(2037.0/65536.0,1,-nbitq), 
to_sfixed(-1392.0/65536.0,1,-nbitq), 
to_sfixed(-61.0/65536.0,1,-nbitq), 
to_sfixed(-7480.0/65536.0,1,-nbitq), 
to_sfixed(-3253.0/65536.0,1,-nbitq), 
to_sfixed(-283.0/65536.0,1,-nbitq), 
to_sfixed(-464.0/65536.0,1,-nbitq), 
to_sfixed(-2870.0/65536.0,1,-nbitq), 
to_sfixed(-4897.0/65536.0,1,-nbitq), 
to_sfixed(10487.0/65536.0,1,-nbitq), 
to_sfixed(-268.0/65536.0,1,-nbitq), 
to_sfixed(8753.0/65536.0,1,-nbitq), 
to_sfixed(-9859.0/65536.0,1,-nbitq), 
to_sfixed(-2031.0/65536.0,1,-nbitq), 
to_sfixed(13.0/65536.0,1,-nbitq), 
to_sfixed(-1749.0/65536.0,1,-nbitq), 
to_sfixed(-2543.0/65536.0,1,-nbitq), 
to_sfixed(-1558.0/65536.0,1,-nbitq), 
to_sfixed(1473.0/65536.0,1,-nbitq), 
to_sfixed(2092.0/65536.0,1,-nbitq), 
to_sfixed(625.0/65536.0,1,-nbitq), 
to_sfixed(-1524.0/65536.0,1,-nbitq), 
to_sfixed(-2850.0/65536.0,1,-nbitq), 
to_sfixed(1504.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5353.0/65536.0,1,-nbitq), 
to_sfixed(-960.0/65536.0,1,-nbitq), 
to_sfixed(-5897.0/65536.0,1,-nbitq), 
to_sfixed(5046.0/65536.0,1,-nbitq), 
to_sfixed(5929.0/65536.0,1,-nbitq), 
to_sfixed(4476.0/65536.0,1,-nbitq), 
to_sfixed(-3333.0/65536.0,1,-nbitq), 
to_sfixed(7914.0/65536.0,1,-nbitq), 
to_sfixed(-865.0/65536.0,1,-nbitq), 
to_sfixed(-425.0/65536.0,1,-nbitq), 
to_sfixed(-4977.0/65536.0,1,-nbitq), 
to_sfixed(-2709.0/65536.0,1,-nbitq), 
to_sfixed(552.0/65536.0,1,-nbitq), 
to_sfixed(2566.0/65536.0,1,-nbitq), 
to_sfixed(-1741.0/65536.0,1,-nbitq), 
to_sfixed(-2125.0/65536.0,1,-nbitq), 
to_sfixed(-1257.0/65536.0,1,-nbitq), 
to_sfixed(-4859.0/65536.0,1,-nbitq), 
to_sfixed(-1579.0/65536.0,1,-nbitq), 
to_sfixed(2422.0/65536.0,1,-nbitq), 
to_sfixed(-549.0/65536.0,1,-nbitq), 
to_sfixed(5866.0/65536.0,1,-nbitq), 
to_sfixed(-5753.0/65536.0,1,-nbitq), 
to_sfixed(2208.0/65536.0,1,-nbitq), 
to_sfixed(-4743.0/65536.0,1,-nbitq), 
to_sfixed(-3193.0/65536.0,1,-nbitq), 
to_sfixed(12854.0/65536.0,1,-nbitq), 
to_sfixed(-2290.0/65536.0,1,-nbitq), 
to_sfixed(4675.0/65536.0,1,-nbitq), 
to_sfixed(3456.0/65536.0,1,-nbitq), 
to_sfixed(-790.0/65536.0,1,-nbitq), 
to_sfixed(-1674.0/65536.0,1,-nbitq), 
to_sfixed(-3404.0/65536.0,1,-nbitq), 
to_sfixed(-1601.0/65536.0,1,-nbitq), 
to_sfixed(-2976.0/65536.0,1,-nbitq), 
to_sfixed(619.0/65536.0,1,-nbitq), 
to_sfixed(-4871.0/65536.0,1,-nbitq), 
to_sfixed(531.0/65536.0,1,-nbitq), 
to_sfixed(3690.0/65536.0,1,-nbitq), 
to_sfixed(-1941.0/65536.0,1,-nbitq), 
to_sfixed(-3729.0/65536.0,1,-nbitq), 
to_sfixed(-764.0/65536.0,1,-nbitq), 
to_sfixed(-3698.0/65536.0,1,-nbitq), 
to_sfixed(3890.0/65536.0,1,-nbitq), 
to_sfixed(-2321.0/65536.0,1,-nbitq), 
to_sfixed(569.0/65536.0,1,-nbitq), 
to_sfixed(2980.0/65536.0,1,-nbitq), 
to_sfixed(2844.0/65536.0,1,-nbitq), 
to_sfixed(120.0/65536.0,1,-nbitq), 
to_sfixed(2403.0/65536.0,1,-nbitq), 
to_sfixed(2128.0/65536.0,1,-nbitq), 
to_sfixed(3569.0/65536.0,1,-nbitq), 
to_sfixed(3746.0/65536.0,1,-nbitq), 
to_sfixed(-2734.0/65536.0,1,-nbitq), 
to_sfixed(-3280.0/65536.0,1,-nbitq), 
to_sfixed(-3473.0/65536.0,1,-nbitq), 
to_sfixed(-2846.0/65536.0,1,-nbitq), 
to_sfixed(-6188.0/65536.0,1,-nbitq), 
to_sfixed(796.0/65536.0,1,-nbitq), 
to_sfixed(-2860.0/65536.0,1,-nbitq), 
to_sfixed(-780.0/65536.0,1,-nbitq), 
to_sfixed(-35.0/65536.0,1,-nbitq), 
to_sfixed(-2380.0/65536.0,1,-nbitq), 
to_sfixed(-2019.0/65536.0,1,-nbitq), 
to_sfixed(-4711.0/65536.0,1,-nbitq), 
to_sfixed(13107.0/65536.0,1,-nbitq), 
to_sfixed(-2813.0/65536.0,1,-nbitq), 
to_sfixed(4674.0/65536.0,1,-nbitq), 
to_sfixed(-6154.0/65536.0,1,-nbitq), 
to_sfixed(1864.0/65536.0,1,-nbitq), 
to_sfixed(-3930.0/65536.0,1,-nbitq), 
to_sfixed(923.0/65536.0,1,-nbitq), 
to_sfixed(-3260.0/65536.0,1,-nbitq), 
to_sfixed(1610.0/65536.0,1,-nbitq), 
to_sfixed(-1587.0/65536.0,1,-nbitq), 
to_sfixed(2052.0/65536.0,1,-nbitq), 
to_sfixed(2621.0/65536.0,1,-nbitq), 
to_sfixed(-4531.0/65536.0,1,-nbitq), 
to_sfixed(1657.0/65536.0,1,-nbitq), 
to_sfixed(5066.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-196.0/65536.0,1,-nbitq), 
to_sfixed(-2438.0/65536.0,1,-nbitq), 
to_sfixed(-5091.0/65536.0,1,-nbitq), 
to_sfixed(4832.0/65536.0,1,-nbitq), 
to_sfixed(6313.0/65536.0,1,-nbitq), 
to_sfixed(3660.0/65536.0,1,-nbitq), 
to_sfixed(-2243.0/65536.0,1,-nbitq), 
to_sfixed(1141.0/65536.0,1,-nbitq), 
to_sfixed(-263.0/65536.0,1,-nbitq), 
to_sfixed(1913.0/65536.0,1,-nbitq), 
to_sfixed(-3536.0/65536.0,1,-nbitq), 
to_sfixed(-110.0/65536.0,1,-nbitq), 
to_sfixed(-922.0/65536.0,1,-nbitq), 
to_sfixed(3416.0/65536.0,1,-nbitq), 
to_sfixed(1362.0/65536.0,1,-nbitq), 
to_sfixed(-2596.0/65536.0,1,-nbitq), 
to_sfixed(-2823.0/65536.0,1,-nbitq), 
to_sfixed(-9119.0/65536.0,1,-nbitq), 
to_sfixed(1056.0/65536.0,1,-nbitq), 
to_sfixed(940.0/65536.0,1,-nbitq), 
to_sfixed(-1610.0/65536.0,1,-nbitq), 
to_sfixed(4069.0/65536.0,1,-nbitq), 
to_sfixed(-5126.0/65536.0,1,-nbitq), 
to_sfixed(4801.0/65536.0,1,-nbitq), 
to_sfixed(-5818.0/65536.0,1,-nbitq), 
to_sfixed(2085.0/65536.0,1,-nbitq), 
to_sfixed(8759.0/65536.0,1,-nbitq), 
to_sfixed(-6559.0/65536.0,1,-nbitq), 
to_sfixed(-3157.0/65536.0,1,-nbitq), 
to_sfixed(799.0/65536.0,1,-nbitq), 
to_sfixed(-2702.0/65536.0,1,-nbitq), 
to_sfixed(3570.0/65536.0,1,-nbitq), 
to_sfixed(-5967.0/65536.0,1,-nbitq), 
to_sfixed(2655.0/65536.0,1,-nbitq), 
to_sfixed(-625.0/65536.0,1,-nbitq), 
to_sfixed(186.0/65536.0,1,-nbitq), 
to_sfixed(-1670.0/65536.0,1,-nbitq), 
to_sfixed(-4860.0/65536.0,1,-nbitq), 
to_sfixed(3317.0/65536.0,1,-nbitq), 
to_sfixed(391.0/65536.0,1,-nbitq), 
to_sfixed(1660.0/65536.0,1,-nbitq), 
to_sfixed(-1301.0/65536.0,1,-nbitq), 
to_sfixed(-5048.0/65536.0,1,-nbitq), 
to_sfixed(3915.0/65536.0,1,-nbitq), 
to_sfixed(-2362.0/65536.0,1,-nbitq), 
to_sfixed(191.0/65536.0,1,-nbitq), 
to_sfixed(40.0/65536.0,1,-nbitq), 
to_sfixed(1681.0/65536.0,1,-nbitq), 
to_sfixed(895.0/65536.0,1,-nbitq), 
to_sfixed(4512.0/65536.0,1,-nbitq), 
to_sfixed(1874.0/65536.0,1,-nbitq), 
to_sfixed(6341.0/65536.0,1,-nbitq), 
to_sfixed(5620.0/65536.0,1,-nbitq), 
to_sfixed(-10457.0/65536.0,1,-nbitq), 
to_sfixed(-1259.0/65536.0,1,-nbitq), 
to_sfixed(-4211.0/65536.0,1,-nbitq), 
to_sfixed(-2154.0/65536.0,1,-nbitq), 
to_sfixed(-5026.0/65536.0,1,-nbitq), 
to_sfixed(2699.0/65536.0,1,-nbitq), 
to_sfixed(-3685.0/65536.0,1,-nbitq), 
to_sfixed(2027.0/65536.0,1,-nbitq), 
to_sfixed(92.0/65536.0,1,-nbitq), 
to_sfixed(2090.0/65536.0,1,-nbitq), 
to_sfixed(-694.0/65536.0,1,-nbitq), 
to_sfixed(3278.0/65536.0,1,-nbitq), 
to_sfixed(10129.0/65536.0,1,-nbitq), 
to_sfixed(-345.0/65536.0,1,-nbitq), 
to_sfixed(3947.0/65536.0,1,-nbitq), 
to_sfixed(-4619.0/65536.0,1,-nbitq), 
to_sfixed(-2426.0/65536.0,1,-nbitq), 
to_sfixed(-2378.0/65536.0,1,-nbitq), 
to_sfixed(3209.0/65536.0,1,-nbitq), 
to_sfixed(-332.0/65536.0,1,-nbitq), 
to_sfixed(-2279.0/65536.0,1,-nbitq), 
to_sfixed(1356.0/65536.0,1,-nbitq), 
to_sfixed(2412.0/65536.0,1,-nbitq), 
to_sfixed(7204.0/65536.0,1,-nbitq), 
to_sfixed(-3299.0/65536.0,1,-nbitq), 
to_sfixed(2121.0/65536.0,1,-nbitq), 
to_sfixed(9116.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3522.0/65536.0,1,-nbitq), 
to_sfixed(-2823.0/65536.0,1,-nbitq), 
to_sfixed(-1885.0/65536.0,1,-nbitq), 
to_sfixed(770.0/65536.0,1,-nbitq), 
to_sfixed(4929.0/65536.0,1,-nbitq), 
to_sfixed(-3259.0/65536.0,1,-nbitq), 
to_sfixed(-3638.0/65536.0,1,-nbitq), 
to_sfixed(3723.0/65536.0,1,-nbitq), 
to_sfixed(1037.0/65536.0,1,-nbitq), 
to_sfixed(-3109.0/65536.0,1,-nbitq), 
to_sfixed(-3121.0/65536.0,1,-nbitq), 
to_sfixed(-124.0/65536.0,1,-nbitq), 
to_sfixed(2024.0/65536.0,1,-nbitq), 
to_sfixed(2616.0/65536.0,1,-nbitq), 
to_sfixed(-3126.0/65536.0,1,-nbitq), 
to_sfixed(-2122.0/65536.0,1,-nbitq), 
to_sfixed(-2723.0/65536.0,1,-nbitq), 
to_sfixed(-4137.0/65536.0,1,-nbitq), 
to_sfixed(1492.0/65536.0,1,-nbitq), 
to_sfixed(-1205.0/65536.0,1,-nbitq), 
to_sfixed(-5046.0/65536.0,1,-nbitq), 
to_sfixed(5503.0/65536.0,1,-nbitq), 
to_sfixed(-5760.0/65536.0,1,-nbitq), 
to_sfixed(6271.0/65536.0,1,-nbitq), 
to_sfixed(-5720.0/65536.0,1,-nbitq), 
to_sfixed(2229.0/65536.0,1,-nbitq), 
to_sfixed(3611.0/65536.0,1,-nbitq), 
to_sfixed(-5651.0/65536.0,1,-nbitq), 
to_sfixed(-8756.0/65536.0,1,-nbitq), 
to_sfixed(2486.0/65536.0,1,-nbitq), 
to_sfixed(-3960.0/65536.0,1,-nbitq), 
to_sfixed(2942.0/65536.0,1,-nbitq), 
to_sfixed(-864.0/65536.0,1,-nbitq), 
to_sfixed(6260.0/65536.0,1,-nbitq), 
to_sfixed(557.0/65536.0,1,-nbitq), 
to_sfixed(-1363.0/65536.0,1,-nbitq), 
to_sfixed(24.0/65536.0,1,-nbitq), 
to_sfixed(-1084.0/65536.0,1,-nbitq), 
to_sfixed(7221.0/65536.0,1,-nbitq), 
to_sfixed(-1562.0/65536.0,1,-nbitq), 
to_sfixed(7941.0/65536.0,1,-nbitq), 
to_sfixed(-344.0/65536.0,1,-nbitq), 
to_sfixed(-3043.0/65536.0,1,-nbitq), 
to_sfixed(-1019.0/65536.0,1,-nbitq), 
to_sfixed(54.0/65536.0,1,-nbitq), 
to_sfixed(-2359.0/65536.0,1,-nbitq), 
to_sfixed(3048.0/65536.0,1,-nbitq), 
to_sfixed(1129.0/65536.0,1,-nbitq), 
to_sfixed(172.0/65536.0,1,-nbitq), 
to_sfixed(-827.0/65536.0,1,-nbitq), 
to_sfixed(-2039.0/65536.0,1,-nbitq), 
to_sfixed(6818.0/65536.0,1,-nbitq), 
to_sfixed(-639.0/65536.0,1,-nbitq), 
to_sfixed(-6032.0/65536.0,1,-nbitq), 
to_sfixed(-1909.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(-886.0/65536.0,1,-nbitq), 
to_sfixed(-3718.0/65536.0,1,-nbitq), 
to_sfixed(768.0/65536.0,1,-nbitq), 
to_sfixed(4326.0/65536.0,1,-nbitq), 
to_sfixed(4073.0/65536.0,1,-nbitq), 
to_sfixed(-1742.0/65536.0,1,-nbitq), 
to_sfixed(1930.0/65536.0,1,-nbitq), 
to_sfixed(-1309.0/65536.0,1,-nbitq), 
to_sfixed(8279.0/65536.0,1,-nbitq), 
to_sfixed(9203.0/65536.0,1,-nbitq), 
to_sfixed(1196.0/65536.0,1,-nbitq), 
to_sfixed(1617.0/65536.0,1,-nbitq), 
to_sfixed(-8911.0/65536.0,1,-nbitq), 
to_sfixed(-10269.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(-908.0/65536.0,1,-nbitq), 
to_sfixed(1563.0/65536.0,1,-nbitq), 
to_sfixed(2275.0/65536.0,1,-nbitq), 
to_sfixed(-1083.0/65536.0,1,-nbitq), 
to_sfixed(-1218.0/65536.0,1,-nbitq), 
to_sfixed(3397.0/65536.0,1,-nbitq), 
to_sfixed(-4307.0/65536.0,1,-nbitq), 
to_sfixed(-175.0/65536.0,1,-nbitq), 
to_sfixed(5949.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1541.0/65536.0,1,-nbitq), 
to_sfixed(-603.0/65536.0,1,-nbitq), 
to_sfixed(5431.0/65536.0,1,-nbitq), 
to_sfixed(1123.0/65536.0,1,-nbitq), 
to_sfixed(4459.0/65536.0,1,-nbitq), 
to_sfixed(-3173.0/65536.0,1,-nbitq), 
to_sfixed(-1607.0/65536.0,1,-nbitq), 
to_sfixed(3918.0/65536.0,1,-nbitq), 
to_sfixed(1819.0/65536.0,1,-nbitq), 
to_sfixed(2152.0/65536.0,1,-nbitq), 
to_sfixed(-3718.0/65536.0,1,-nbitq), 
to_sfixed(-894.0/65536.0,1,-nbitq), 
to_sfixed(2529.0/65536.0,1,-nbitq), 
to_sfixed(-1157.0/65536.0,1,-nbitq), 
to_sfixed(-246.0/65536.0,1,-nbitq), 
to_sfixed(-1898.0/65536.0,1,-nbitq), 
to_sfixed(-347.0/65536.0,1,-nbitq), 
to_sfixed(-3179.0/65536.0,1,-nbitq), 
to_sfixed(2350.0/65536.0,1,-nbitq), 
to_sfixed(146.0/65536.0,1,-nbitq), 
to_sfixed(-3625.0/65536.0,1,-nbitq), 
to_sfixed(2784.0/65536.0,1,-nbitq), 
to_sfixed(497.0/65536.0,1,-nbitq), 
to_sfixed(4875.0/65536.0,1,-nbitq), 
to_sfixed(-829.0/65536.0,1,-nbitq), 
to_sfixed(-1884.0/65536.0,1,-nbitq), 
to_sfixed(5081.0/65536.0,1,-nbitq), 
to_sfixed(-6240.0/65536.0,1,-nbitq), 
to_sfixed(-8348.0/65536.0,1,-nbitq), 
to_sfixed(2457.0/65536.0,1,-nbitq), 
to_sfixed(-3552.0/65536.0,1,-nbitq), 
to_sfixed(1847.0/65536.0,1,-nbitq), 
to_sfixed(1906.0/65536.0,1,-nbitq), 
to_sfixed(7491.0/65536.0,1,-nbitq), 
to_sfixed(-603.0/65536.0,1,-nbitq), 
to_sfixed(-969.0/65536.0,1,-nbitq), 
to_sfixed(785.0/65536.0,1,-nbitq), 
to_sfixed(-3349.0/65536.0,1,-nbitq), 
to_sfixed(4375.0/65536.0,1,-nbitq), 
to_sfixed(-2204.0/65536.0,1,-nbitq), 
to_sfixed(11256.0/65536.0,1,-nbitq), 
to_sfixed(686.0/65536.0,1,-nbitq), 
to_sfixed(-2216.0/65536.0,1,-nbitq), 
to_sfixed(2643.0/65536.0,1,-nbitq), 
to_sfixed(-1813.0/65536.0,1,-nbitq), 
to_sfixed(1740.0/65536.0,1,-nbitq), 
to_sfixed(2533.0/65536.0,1,-nbitq), 
to_sfixed(416.0/65536.0,1,-nbitq), 
to_sfixed(-853.0/65536.0,1,-nbitq), 
to_sfixed(-1123.0/65536.0,1,-nbitq), 
to_sfixed(-1832.0/65536.0,1,-nbitq), 
to_sfixed(-300.0/65536.0,1,-nbitq), 
to_sfixed(1420.0/65536.0,1,-nbitq), 
to_sfixed(-8586.0/65536.0,1,-nbitq), 
to_sfixed(-1108.0/65536.0,1,-nbitq), 
to_sfixed(3936.0/65536.0,1,-nbitq), 
to_sfixed(-1412.0/65536.0,1,-nbitq), 
to_sfixed(1259.0/65536.0,1,-nbitq), 
to_sfixed(-646.0/65536.0,1,-nbitq), 
to_sfixed(5449.0/65536.0,1,-nbitq), 
to_sfixed(1312.0/65536.0,1,-nbitq), 
to_sfixed(-603.0/65536.0,1,-nbitq), 
to_sfixed(-2134.0/65536.0,1,-nbitq), 
to_sfixed(2497.0/65536.0,1,-nbitq), 
to_sfixed(6298.0/65536.0,1,-nbitq), 
to_sfixed(3954.0/65536.0,1,-nbitq), 
to_sfixed(-1533.0/65536.0,1,-nbitq), 
to_sfixed(2433.0/65536.0,1,-nbitq), 
to_sfixed(-2122.0/65536.0,1,-nbitq), 
to_sfixed(-8820.0/65536.0,1,-nbitq), 
to_sfixed(599.0/65536.0,1,-nbitq), 
to_sfixed(-895.0/65536.0,1,-nbitq), 
to_sfixed(2062.0/65536.0,1,-nbitq), 
to_sfixed(-1474.0/65536.0,1,-nbitq), 
to_sfixed(-1471.0/65536.0,1,-nbitq), 
to_sfixed(-1933.0/65536.0,1,-nbitq), 
to_sfixed(5834.0/65536.0,1,-nbitq), 
to_sfixed(-3206.0/65536.0,1,-nbitq), 
to_sfixed(-1646.0/65536.0,1,-nbitq), 
to_sfixed(8088.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2758.0/65536.0,1,-nbitq), 
to_sfixed(-1005.0/65536.0,1,-nbitq), 
to_sfixed(6446.0/65536.0,1,-nbitq), 
to_sfixed(-125.0/65536.0,1,-nbitq), 
to_sfixed(-970.0/65536.0,1,-nbitq), 
to_sfixed(255.0/65536.0,1,-nbitq), 
to_sfixed(-150.0/65536.0,1,-nbitq), 
to_sfixed(4782.0/65536.0,1,-nbitq), 
to_sfixed(-1704.0/65536.0,1,-nbitq), 
to_sfixed(-2767.0/65536.0,1,-nbitq), 
to_sfixed(-863.0/65536.0,1,-nbitq), 
to_sfixed(-266.0/65536.0,1,-nbitq), 
to_sfixed(-753.0/65536.0,1,-nbitq), 
to_sfixed(2554.0/65536.0,1,-nbitq), 
to_sfixed(-4615.0/65536.0,1,-nbitq), 
to_sfixed(3279.0/65536.0,1,-nbitq), 
to_sfixed(1107.0/65536.0,1,-nbitq), 
to_sfixed(-2964.0/65536.0,1,-nbitq), 
to_sfixed(-837.0/65536.0,1,-nbitq), 
to_sfixed(-2658.0/65536.0,1,-nbitq), 
to_sfixed(-363.0/65536.0,1,-nbitq), 
to_sfixed(-2464.0/65536.0,1,-nbitq), 
to_sfixed(4363.0/65536.0,1,-nbitq), 
to_sfixed(1960.0/65536.0,1,-nbitq), 
to_sfixed(-3282.0/65536.0,1,-nbitq), 
to_sfixed(1926.0/65536.0,1,-nbitq), 
to_sfixed(219.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(-8871.0/65536.0,1,-nbitq), 
to_sfixed(1132.0/65536.0,1,-nbitq), 
to_sfixed(787.0/65536.0,1,-nbitq), 
to_sfixed(2011.0/65536.0,1,-nbitq), 
to_sfixed(334.0/65536.0,1,-nbitq), 
to_sfixed(5214.0/65536.0,1,-nbitq), 
to_sfixed(2487.0/65536.0,1,-nbitq), 
to_sfixed(2088.0/65536.0,1,-nbitq), 
to_sfixed(-2269.0/65536.0,1,-nbitq), 
to_sfixed(-1576.0/65536.0,1,-nbitq), 
to_sfixed(1599.0/65536.0,1,-nbitq), 
to_sfixed(2456.0/65536.0,1,-nbitq), 
to_sfixed(6754.0/65536.0,1,-nbitq), 
to_sfixed(-2885.0/65536.0,1,-nbitq), 
to_sfixed(-491.0/65536.0,1,-nbitq), 
to_sfixed(197.0/65536.0,1,-nbitq), 
to_sfixed(1883.0/65536.0,1,-nbitq), 
to_sfixed(2675.0/65536.0,1,-nbitq), 
to_sfixed(1659.0/65536.0,1,-nbitq), 
to_sfixed(-1832.0/65536.0,1,-nbitq), 
to_sfixed(2129.0/65536.0,1,-nbitq), 
to_sfixed(-1255.0/65536.0,1,-nbitq), 
to_sfixed(2410.0/65536.0,1,-nbitq), 
to_sfixed(-659.0/65536.0,1,-nbitq), 
to_sfixed(1951.0/65536.0,1,-nbitq), 
to_sfixed(-4840.0/65536.0,1,-nbitq), 
to_sfixed(630.0/65536.0,1,-nbitq), 
to_sfixed(1879.0/65536.0,1,-nbitq), 
to_sfixed(-2421.0/65536.0,1,-nbitq), 
to_sfixed(3265.0/65536.0,1,-nbitq), 
to_sfixed(872.0/65536.0,1,-nbitq), 
to_sfixed(4705.0/65536.0,1,-nbitq), 
to_sfixed(-1337.0/65536.0,1,-nbitq), 
to_sfixed(-930.0/65536.0,1,-nbitq), 
to_sfixed(-1546.0/65536.0,1,-nbitq), 
to_sfixed(-3208.0/65536.0,1,-nbitq), 
to_sfixed(333.0/65536.0,1,-nbitq), 
to_sfixed(3388.0/65536.0,1,-nbitq), 
to_sfixed(1278.0/65536.0,1,-nbitq), 
to_sfixed(5146.0/65536.0,1,-nbitq), 
to_sfixed(-2183.0/65536.0,1,-nbitq), 
to_sfixed(-6061.0/65536.0,1,-nbitq), 
to_sfixed(3448.0/65536.0,1,-nbitq), 
to_sfixed(-1584.0/65536.0,1,-nbitq), 
to_sfixed(-4159.0/65536.0,1,-nbitq), 
to_sfixed(-2466.0/65536.0,1,-nbitq), 
to_sfixed(837.0/65536.0,1,-nbitq), 
to_sfixed(2348.0/65536.0,1,-nbitq), 
to_sfixed(320.0/65536.0,1,-nbitq), 
to_sfixed(-150.0/65536.0,1,-nbitq), 
to_sfixed(631.0/65536.0,1,-nbitq), 
to_sfixed(6987.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2205.0/65536.0,1,-nbitq), 
to_sfixed(-3582.0/65536.0,1,-nbitq), 
to_sfixed(7460.0/65536.0,1,-nbitq), 
to_sfixed(2034.0/65536.0,1,-nbitq), 
to_sfixed(1871.0/65536.0,1,-nbitq), 
to_sfixed(-1505.0/65536.0,1,-nbitq), 
to_sfixed(2544.0/65536.0,1,-nbitq), 
to_sfixed(6189.0/65536.0,1,-nbitq), 
to_sfixed(2355.0/65536.0,1,-nbitq), 
to_sfixed(1240.0/65536.0,1,-nbitq), 
to_sfixed(2625.0/65536.0,1,-nbitq), 
to_sfixed(2411.0/65536.0,1,-nbitq), 
to_sfixed(-379.0/65536.0,1,-nbitq), 
to_sfixed(1521.0/65536.0,1,-nbitq), 
to_sfixed(-2407.0/65536.0,1,-nbitq), 
to_sfixed(2695.0/65536.0,1,-nbitq), 
to_sfixed(2840.0/65536.0,1,-nbitq), 
to_sfixed(456.0/65536.0,1,-nbitq), 
to_sfixed(-1538.0/65536.0,1,-nbitq), 
to_sfixed(-2413.0/65536.0,1,-nbitq), 
to_sfixed(-625.0/65536.0,1,-nbitq), 
to_sfixed(-3314.0/65536.0,1,-nbitq), 
to_sfixed(-1993.0/65536.0,1,-nbitq), 
to_sfixed(-2310.0/65536.0,1,-nbitq), 
to_sfixed(-3741.0/65536.0,1,-nbitq), 
to_sfixed(-1946.0/65536.0,1,-nbitq), 
to_sfixed(-2357.0/65536.0,1,-nbitq), 
to_sfixed(-1449.0/65536.0,1,-nbitq), 
to_sfixed(-1643.0/65536.0,1,-nbitq), 
to_sfixed(631.0/65536.0,1,-nbitq), 
to_sfixed(-1531.0/65536.0,1,-nbitq), 
to_sfixed(2039.0/65536.0,1,-nbitq), 
to_sfixed(-352.0/65536.0,1,-nbitq), 
to_sfixed(4894.0/65536.0,1,-nbitq), 
to_sfixed(542.0/65536.0,1,-nbitq), 
to_sfixed(-2768.0/65536.0,1,-nbitq), 
to_sfixed(-5501.0/65536.0,1,-nbitq), 
to_sfixed(3490.0/65536.0,1,-nbitq), 
to_sfixed(-2659.0/65536.0,1,-nbitq), 
to_sfixed(2051.0/65536.0,1,-nbitq), 
to_sfixed(2136.0/65536.0,1,-nbitq), 
to_sfixed(-3190.0/65536.0,1,-nbitq), 
to_sfixed(1452.0/65536.0,1,-nbitq), 
to_sfixed(3421.0/65536.0,1,-nbitq), 
to_sfixed(1910.0/65536.0,1,-nbitq), 
to_sfixed(-323.0/65536.0,1,-nbitq), 
to_sfixed(1073.0/65536.0,1,-nbitq), 
to_sfixed(965.0/65536.0,1,-nbitq), 
to_sfixed(-6.0/65536.0,1,-nbitq), 
to_sfixed(3500.0/65536.0,1,-nbitq), 
to_sfixed(804.0/65536.0,1,-nbitq), 
to_sfixed(670.0/65536.0,1,-nbitq), 
to_sfixed(484.0/65536.0,1,-nbitq), 
to_sfixed(501.0/65536.0,1,-nbitq), 
to_sfixed(-843.0/65536.0,1,-nbitq), 
to_sfixed(1466.0/65536.0,1,-nbitq), 
to_sfixed(-2052.0/65536.0,1,-nbitq), 
to_sfixed(1855.0/65536.0,1,-nbitq), 
to_sfixed(196.0/65536.0,1,-nbitq), 
to_sfixed(1086.0/65536.0,1,-nbitq), 
to_sfixed(225.0/65536.0,1,-nbitq), 
to_sfixed(-1207.0/65536.0,1,-nbitq), 
to_sfixed(2311.0/65536.0,1,-nbitq), 
to_sfixed(-3375.0/65536.0,1,-nbitq), 
to_sfixed(-3261.0/65536.0,1,-nbitq), 
to_sfixed(6207.0/65536.0,1,-nbitq), 
to_sfixed(-4413.0/65536.0,1,-nbitq), 
to_sfixed(2091.0/65536.0,1,-nbitq), 
to_sfixed(-2504.0/65536.0,1,-nbitq), 
to_sfixed(2072.0/65536.0,1,-nbitq), 
to_sfixed(2219.0/65536.0,1,-nbitq), 
to_sfixed(310.0/65536.0,1,-nbitq), 
to_sfixed(-7146.0/65536.0,1,-nbitq), 
to_sfixed(-1871.0/65536.0,1,-nbitq), 
to_sfixed(620.0/65536.0,1,-nbitq), 
to_sfixed(2219.0/65536.0,1,-nbitq), 
to_sfixed(3104.0/65536.0,1,-nbitq), 
to_sfixed(-1279.0/65536.0,1,-nbitq), 
to_sfixed(1714.0/65536.0,1,-nbitq), 
to_sfixed(881.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-851.0/65536.0,1,-nbitq), 
to_sfixed(1110.0/65536.0,1,-nbitq), 
to_sfixed(5161.0/65536.0,1,-nbitq), 
to_sfixed(-2572.0/65536.0,1,-nbitq), 
to_sfixed(1547.0/65536.0,1,-nbitq), 
to_sfixed(-2064.0/65536.0,1,-nbitq), 
to_sfixed(-472.0/65536.0,1,-nbitq), 
to_sfixed(2587.0/65536.0,1,-nbitq), 
to_sfixed(-536.0/65536.0,1,-nbitq), 
to_sfixed(681.0/65536.0,1,-nbitq), 
to_sfixed(4241.0/65536.0,1,-nbitq), 
to_sfixed(-1303.0/65536.0,1,-nbitq), 
to_sfixed(-1138.0/65536.0,1,-nbitq), 
to_sfixed(2830.0/65536.0,1,-nbitq), 
to_sfixed(1508.0/65536.0,1,-nbitq), 
to_sfixed(-808.0/65536.0,1,-nbitq), 
to_sfixed(-2528.0/65536.0,1,-nbitq), 
to_sfixed(287.0/65536.0,1,-nbitq), 
to_sfixed(-850.0/65536.0,1,-nbitq), 
to_sfixed(135.0/65536.0,1,-nbitq), 
to_sfixed(1209.0/65536.0,1,-nbitq), 
to_sfixed(-2207.0/65536.0,1,-nbitq), 
to_sfixed(-3739.0/65536.0,1,-nbitq), 
to_sfixed(-1420.0/65536.0,1,-nbitq), 
to_sfixed(-2918.0/65536.0,1,-nbitq), 
to_sfixed(-6163.0/65536.0,1,-nbitq), 
to_sfixed(-2014.0/65536.0,1,-nbitq), 
to_sfixed(-3451.0/65536.0,1,-nbitq), 
to_sfixed(2385.0/65536.0,1,-nbitq), 
to_sfixed(2644.0/65536.0,1,-nbitq), 
to_sfixed(-88.0/65536.0,1,-nbitq), 
to_sfixed(-216.0/65536.0,1,-nbitq), 
to_sfixed(512.0/65536.0,1,-nbitq), 
to_sfixed(4449.0/65536.0,1,-nbitq), 
to_sfixed(-1671.0/65536.0,1,-nbitq), 
to_sfixed(-1850.0/65536.0,1,-nbitq), 
to_sfixed(-1314.0/65536.0,1,-nbitq), 
to_sfixed(2551.0/65536.0,1,-nbitq), 
to_sfixed(-620.0/65536.0,1,-nbitq), 
to_sfixed(2939.0/65536.0,1,-nbitq), 
to_sfixed(159.0/65536.0,1,-nbitq), 
to_sfixed(2232.0/65536.0,1,-nbitq), 
to_sfixed(-658.0/65536.0,1,-nbitq), 
to_sfixed(5001.0/65536.0,1,-nbitq), 
to_sfixed(1569.0/65536.0,1,-nbitq), 
to_sfixed(-1387.0/65536.0,1,-nbitq), 
to_sfixed(-3243.0/65536.0,1,-nbitq), 
to_sfixed(628.0/65536.0,1,-nbitq), 
to_sfixed(-242.0/65536.0,1,-nbitq), 
to_sfixed(1951.0/65536.0,1,-nbitq), 
to_sfixed(542.0/65536.0,1,-nbitq), 
to_sfixed(-2037.0/65536.0,1,-nbitq), 
to_sfixed(2556.0/65536.0,1,-nbitq), 
to_sfixed(5954.0/65536.0,1,-nbitq), 
to_sfixed(-4110.0/65536.0,1,-nbitq), 
to_sfixed(-1413.0/65536.0,1,-nbitq), 
to_sfixed(1804.0/65536.0,1,-nbitq), 
to_sfixed(-1664.0/65536.0,1,-nbitq), 
to_sfixed(-1902.0/65536.0,1,-nbitq), 
to_sfixed(802.0/65536.0,1,-nbitq), 
to_sfixed(3665.0/65536.0,1,-nbitq), 
to_sfixed(462.0/65536.0,1,-nbitq), 
to_sfixed(-2760.0/65536.0,1,-nbitq), 
to_sfixed(-1539.0/65536.0,1,-nbitq), 
to_sfixed(-3431.0/65536.0,1,-nbitq), 
to_sfixed(2027.0/65536.0,1,-nbitq), 
to_sfixed(-6064.0/65536.0,1,-nbitq), 
to_sfixed(2895.0/65536.0,1,-nbitq), 
to_sfixed(2534.0/65536.0,1,-nbitq), 
to_sfixed(2592.0/65536.0,1,-nbitq), 
to_sfixed(2651.0/65536.0,1,-nbitq), 
to_sfixed(1256.0/65536.0,1,-nbitq), 
to_sfixed(-9129.0/65536.0,1,-nbitq), 
to_sfixed(-837.0/65536.0,1,-nbitq), 
to_sfixed(-3036.0/65536.0,1,-nbitq), 
to_sfixed(918.0/65536.0,1,-nbitq), 
to_sfixed(-1930.0/65536.0,1,-nbitq), 
to_sfixed(-4341.0/65536.0,1,-nbitq), 
to_sfixed(-2215.0/65536.0,1,-nbitq), 
to_sfixed(1871.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4176.0/65536.0,1,-nbitq), 
to_sfixed(-74.0/65536.0,1,-nbitq), 
to_sfixed(827.0/65536.0,1,-nbitq), 
to_sfixed(-731.0/65536.0,1,-nbitq), 
to_sfixed(-226.0/65536.0,1,-nbitq), 
to_sfixed(-4830.0/65536.0,1,-nbitq), 
to_sfixed(-2357.0/65536.0,1,-nbitq), 
to_sfixed(-278.0/65536.0,1,-nbitq), 
to_sfixed(-2802.0/65536.0,1,-nbitq), 
to_sfixed(133.0/65536.0,1,-nbitq), 
to_sfixed(1966.0/65536.0,1,-nbitq), 
to_sfixed(-69.0/65536.0,1,-nbitq), 
to_sfixed(-1509.0/65536.0,1,-nbitq), 
to_sfixed(-3908.0/65536.0,1,-nbitq), 
to_sfixed(498.0/65536.0,1,-nbitq), 
to_sfixed(-1180.0/65536.0,1,-nbitq), 
to_sfixed(823.0/65536.0,1,-nbitq), 
to_sfixed(-2345.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(1948.0/65536.0,1,-nbitq), 
to_sfixed(-1997.0/65536.0,1,-nbitq), 
to_sfixed(400.0/65536.0,1,-nbitq), 
to_sfixed(-2423.0/65536.0,1,-nbitq), 
to_sfixed(848.0/65536.0,1,-nbitq), 
to_sfixed(474.0/65536.0,1,-nbitq), 
to_sfixed(-4924.0/65536.0,1,-nbitq), 
to_sfixed(-471.0/65536.0,1,-nbitq), 
to_sfixed(-3703.0/65536.0,1,-nbitq), 
to_sfixed(-1273.0/65536.0,1,-nbitq), 
to_sfixed(2752.0/65536.0,1,-nbitq), 
to_sfixed(-452.0/65536.0,1,-nbitq), 
to_sfixed(2484.0/65536.0,1,-nbitq), 
to_sfixed(-1147.0/65536.0,1,-nbitq), 
to_sfixed(3261.0/65536.0,1,-nbitq), 
to_sfixed(-3070.0/65536.0,1,-nbitq), 
to_sfixed(9.0/65536.0,1,-nbitq), 
to_sfixed(172.0/65536.0,1,-nbitq), 
to_sfixed(373.0/65536.0,1,-nbitq), 
to_sfixed(4042.0/65536.0,1,-nbitq), 
to_sfixed(2526.0/65536.0,1,-nbitq), 
to_sfixed(-3732.0/65536.0,1,-nbitq), 
to_sfixed(673.0/65536.0,1,-nbitq), 
to_sfixed(-4338.0/65536.0,1,-nbitq), 
to_sfixed(1668.0/65536.0,1,-nbitq), 
to_sfixed(-1518.0/65536.0,1,-nbitq), 
to_sfixed(1315.0/65536.0,1,-nbitq), 
to_sfixed(1736.0/65536.0,1,-nbitq), 
to_sfixed(2249.0/65536.0,1,-nbitq), 
to_sfixed(496.0/65536.0,1,-nbitq), 
to_sfixed(3216.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(2907.0/65536.0,1,-nbitq), 
to_sfixed(5437.0/65536.0,1,-nbitq), 
to_sfixed(-2182.0/65536.0,1,-nbitq), 
to_sfixed(-2763.0/65536.0,1,-nbitq), 
to_sfixed(240.0/65536.0,1,-nbitq), 
to_sfixed(-1495.0/65536.0,1,-nbitq), 
to_sfixed(2279.0/65536.0,1,-nbitq), 
to_sfixed(-611.0/65536.0,1,-nbitq), 
to_sfixed(-1508.0/65536.0,1,-nbitq), 
to_sfixed(-191.0/65536.0,1,-nbitq), 
to_sfixed(2100.0/65536.0,1,-nbitq), 
to_sfixed(2874.0/65536.0,1,-nbitq), 
to_sfixed(-292.0/65536.0,1,-nbitq), 
to_sfixed(-2210.0/65536.0,1,-nbitq), 
to_sfixed(1770.0/65536.0,1,-nbitq), 
to_sfixed(-3691.0/65536.0,1,-nbitq), 
to_sfixed(-461.0/65536.0,1,-nbitq), 
to_sfixed(3771.0/65536.0,1,-nbitq), 
to_sfixed(606.0/65536.0,1,-nbitq), 
to_sfixed(511.0/65536.0,1,-nbitq), 
to_sfixed(3075.0/65536.0,1,-nbitq), 
to_sfixed(-2400.0/65536.0,1,-nbitq), 
to_sfixed(-3110.0/65536.0,1,-nbitq), 
to_sfixed(2546.0/65536.0,1,-nbitq), 
to_sfixed(-2098.0/65536.0,1,-nbitq), 
to_sfixed(-1166.0/65536.0,1,-nbitq), 
to_sfixed(-1427.0/65536.0,1,-nbitq), 
to_sfixed(2710.0/65536.0,1,-nbitq), 
to_sfixed(1884.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3593.0/65536.0,1,-nbitq), 
to_sfixed(-2736.0/65536.0,1,-nbitq), 
to_sfixed(-2417.0/65536.0,1,-nbitq), 
to_sfixed(-1730.0/65536.0,1,-nbitq), 
to_sfixed(-1812.0/65536.0,1,-nbitq), 
to_sfixed(-3121.0/65536.0,1,-nbitq), 
to_sfixed(-508.0/65536.0,1,-nbitq), 
to_sfixed(3495.0/65536.0,1,-nbitq), 
to_sfixed(-2376.0/65536.0,1,-nbitq), 
to_sfixed(-2823.0/65536.0,1,-nbitq), 
to_sfixed(-3066.0/65536.0,1,-nbitq), 
to_sfixed(-1848.0/65536.0,1,-nbitq), 
to_sfixed(2638.0/65536.0,1,-nbitq), 
to_sfixed(-386.0/65536.0,1,-nbitq), 
to_sfixed(-144.0/65536.0,1,-nbitq), 
to_sfixed(-732.0/65536.0,1,-nbitq), 
to_sfixed(-1335.0/65536.0,1,-nbitq), 
to_sfixed(2910.0/65536.0,1,-nbitq), 
to_sfixed(3728.0/65536.0,1,-nbitq), 
to_sfixed(-126.0/65536.0,1,-nbitq), 
to_sfixed(2053.0/65536.0,1,-nbitq), 
to_sfixed(-1863.0/65536.0,1,-nbitq), 
to_sfixed(-1940.0/65536.0,1,-nbitq), 
to_sfixed(-2979.0/65536.0,1,-nbitq), 
to_sfixed(-86.0/65536.0,1,-nbitq), 
to_sfixed(-2010.0/65536.0,1,-nbitq), 
to_sfixed(-6919.0/65536.0,1,-nbitq), 
to_sfixed(187.0/65536.0,1,-nbitq), 
to_sfixed(-3278.0/65536.0,1,-nbitq), 
to_sfixed(-1285.0/65536.0,1,-nbitq), 
to_sfixed(-487.0/65536.0,1,-nbitq), 
to_sfixed(248.0/65536.0,1,-nbitq), 
to_sfixed(-3688.0/65536.0,1,-nbitq), 
to_sfixed(3111.0/65536.0,1,-nbitq), 
to_sfixed(-2828.0/65536.0,1,-nbitq), 
to_sfixed(-330.0/65536.0,1,-nbitq), 
to_sfixed(2110.0/65536.0,1,-nbitq), 
to_sfixed(125.0/65536.0,1,-nbitq), 
to_sfixed(-1277.0/65536.0,1,-nbitq), 
to_sfixed(-1667.0/65536.0,1,-nbitq), 
to_sfixed(1939.0/65536.0,1,-nbitq), 
to_sfixed(-1540.0/65536.0,1,-nbitq), 
to_sfixed(-4649.0/65536.0,1,-nbitq), 
to_sfixed(4034.0/65536.0,1,-nbitq), 
to_sfixed(-2607.0/65536.0,1,-nbitq), 
to_sfixed(-4052.0/65536.0,1,-nbitq), 
to_sfixed(-1157.0/65536.0,1,-nbitq), 
to_sfixed(-3029.0/65536.0,1,-nbitq), 
to_sfixed(1742.0/65536.0,1,-nbitq), 
to_sfixed(2693.0/65536.0,1,-nbitq), 
to_sfixed(2407.0/65536.0,1,-nbitq), 
to_sfixed(511.0/65536.0,1,-nbitq), 
to_sfixed(1327.0/65536.0,1,-nbitq), 
to_sfixed(-631.0/65536.0,1,-nbitq), 
to_sfixed(719.0/65536.0,1,-nbitq), 
to_sfixed(-391.0/65536.0,1,-nbitq), 
to_sfixed(-512.0/65536.0,1,-nbitq), 
to_sfixed(1787.0/65536.0,1,-nbitq), 
to_sfixed(-1106.0/65536.0,1,-nbitq), 
to_sfixed(-2911.0/65536.0,1,-nbitq), 
to_sfixed(699.0/65536.0,1,-nbitq), 
to_sfixed(-1821.0/65536.0,1,-nbitq), 
to_sfixed(1035.0/65536.0,1,-nbitq), 
to_sfixed(1354.0/65536.0,1,-nbitq), 
to_sfixed(819.0/65536.0,1,-nbitq), 
to_sfixed(585.0/65536.0,1,-nbitq), 
to_sfixed(1298.0/65536.0,1,-nbitq), 
to_sfixed(-2698.0/65536.0,1,-nbitq), 
to_sfixed(5250.0/65536.0,1,-nbitq), 
to_sfixed(2712.0/65536.0,1,-nbitq), 
to_sfixed(-1918.0/65536.0,1,-nbitq), 
to_sfixed(1066.0/65536.0,1,-nbitq), 
to_sfixed(-3673.0/65536.0,1,-nbitq), 
to_sfixed(-90.0/65536.0,1,-nbitq), 
to_sfixed(1264.0/65536.0,1,-nbitq), 
to_sfixed(-96.0/65536.0,1,-nbitq), 
to_sfixed(-482.0/65536.0,1,-nbitq), 
to_sfixed(2713.0/65536.0,1,-nbitq), 
to_sfixed(-2163.0/65536.0,1,-nbitq), 
to_sfixed(-66.0/65536.0,1,-nbitq)  ), 
( to_sfixed(45.0/65536.0,1,-nbitq), 
to_sfixed(-603.0/65536.0,1,-nbitq), 
to_sfixed(-3535.0/65536.0,1,-nbitq), 
to_sfixed(985.0/65536.0,1,-nbitq), 
to_sfixed(-1478.0/65536.0,1,-nbitq), 
to_sfixed(6.0/65536.0,1,-nbitq), 
to_sfixed(1779.0/65536.0,1,-nbitq), 
to_sfixed(1462.0/65536.0,1,-nbitq), 
to_sfixed(-3665.0/65536.0,1,-nbitq), 
to_sfixed(253.0/65536.0,1,-nbitq), 
to_sfixed(890.0/65536.0,1,-nbitq), 
to_sfixed(-3488.0/65536.0,1,-nbitq), 
to_sfixed(883.0/65536.0,1,-nbitq), 
to_sfixed(1746.0/65536.0,1,-nbitq), 
to_sfixed(-1501.0/65536.0,1,-nbitq), 
to_sfixed(-31.0/65536.0,1,-nbitq), 
to_sfixed(2651.0/65536.0,1,-nbitq), 
to_sfixed(1968.0/65536.0,1,-nbitq), 
to_sfixed(3482.0/65536.0,1,-nbitq), 
to_sfixed(-90.0/65536.0,1,-nbitq), 
to_sfixed(-2147.0/65536.0,1,-nbitq), 
to_sfixed(-1159.0/65536.0,1,-nbitq), 
to_sfixed(976.0/65536.0,1,-nbitq), 
to_sfixed(-1788.0/65536.0,1,-nbitq), 
to_sfixed(-55.0/65536.0,1,-nbitq), 
to_sfixed(-2352.0/65536.0,1,-nbitq), 
to_sfixed(-6075.0/65536.0,1,-nbitq), 
to_sfixed(1593.0/65536.0,1,-nbitq), 
to_sfixed(276.0/65536.0,1,-nbitq), 
to_sfixed(-2478.0/65536.0,1,-nbitq), 
to_sfixed(4358.0/65536.0,1,-nbitq), 
to_sfixed(417.0/65536.0,1,-nbitq), 
to_sfixed(-1947.0/65536.0,1,-nbitq), 
to_sfixed(-660.0/65536.0,1,-nbitq), 
to_sfixed(710.0/65536.0,1,-nbitq), 
to_sfixed(524.0/65536.0,1,-nbitq), 
to_sfixed(-1946.0/65536.0,1,-nbitq), 
to_sfixed(-1944.0/65536.0,1,-nbitq), 
to_sfixed(2053.0/65536.0,1,-nbitq), 
to_sfixed(-288.0/65536.0,1,-nbitq), 
to_sfixed(-249.0/65536.0,1,-nbitq), 
to_sfixed(-3162.0/65536.0,1,-nbitq), 
to_sfixed(-2653.0/65536.0,1,-nbitq), 
to_sfixed(4973.0/65536.0,1,-nbitq), 
to_sfixed(-983.0/65536.0,1,-nbitq), 
to_sfixed(2060.0/65536.0,1,-nbitq), 
to_sfixed(-2437.0/65536.0,1,-nbitq), 
to_sfixed(769.0/65536.0,1,-nbitq), 
to_sfixed(2112.0/65536.0,1,-nbitq), 
to_sfixed(1994.0/65536.0,1,-nbitq), 
to_sfixed(-1561.0/65536.0,1,-nbitq), 
to_sfixed(2996.0/65536.0,1,-nbitq), 
to_sfixed(-8.0/65536.0,1,-nbitq), 
to_sfixed(-4473.0/65536.0,1,-nbitq), 
to_sfixed(610.0/65536.0,1,-nbitq), 
to_sfixed(-76.0/65536.0,1,-nbitq), 
to_sfixed(-9.0/65536.0,1,-nbitq), 
to_sfixed(1083.0/65536.0,1,-nbitq), 
to_sfixed(1166.0/65536.0,1,-nbitq), 
to_sfixed(781.0/65536.0,1,-nbitq), 
to_sfixed(512.0/65536.0,1,-nbitq), 
to_sfixed(-631.0/65536.0,1,-nbitq), 
to_sfixed(-2119.0/65536.0,1,-nbitq), 
to_sfixed(-1262.0/65536.0,1,-nbitq), 
to_sfixed(2304.0/65536.0,1,-nbitq), 
to_sfixed(-2930.0/65536.0,1,-nbitq), 
to_sfixed(888.0/65536.0,1,-nbitq), 
to_sfixed(-2160.0/65536.0,1,-nbitq), 
to_sfixed(5219.0/65536.0,1,-nbitq), 
to_sfixed(-280.0/65536.0,1,-nbitq), 
to_sfixed(-2533.0/65536.0,1,-nbitq), 
to_sfixed(46.0/65536.0,1,-nbitq), 
to_sfixed(-1074.0/65536.0,1,-nbitq), 
to_sfixed(-1259.0/65536.0,1,-nbitq), 
to_sfixed(-1168.0/65536.0,1,-nbitq), 
to_sfixed(-678.0/65536.0,1,-nbitq), 
to_sfixed(812.0/65536.0,1,-nbitq), 
to_sfixed(3578.0/65536.0,1,-nbitq), 
to_sfixed(2153.0/65536.0,1,-nbitq), 
to_sfixed(1793.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3002.0/65536.0,1,-nbitq), 
to_sfixed(2019.0/65536.0,1,-nbitq), 
to_sfixed(-1511.0/65536.0,1,-nbitq), 
to_sfixed(-2516.0/65536.0,1,-nbitq), 
to_sfixed(-2687.0/65536.0,1,-nbitq), 
to_sfixed(-2529.0/65536.0,1,-nbitq), 
to_sfixed(-2454.0/65536.0,1,-nbitq), 
to_sfixed(-718.0/65536.0,1,-nbitq), 
to_sfixed(-2478.0/65536.0,1,-nbitq), 
to_sfixed(-2823.0/65536.0,1,-nbitq), 
to_sfixed(-2894.0/65536.0,1,-nbitq), 
to_sfixed(-76.0/65536.0,1,-nbitq), 
to_sfixed(2516.0/65536.0,1,-nbitq), 
to_sfixed(-1977.0/65536.0,1,-nbitq), 
to_sfixed(318.0/65536.0,1,-nbitq), 
to_sfixed(3070.0/65536.0,1,-nbitq), 
to_sfixed(-153.0/65536.0,1,-nbitq), 
to_sfixed(47.0/65536.0,1,-nbitq), 
to_sfixed(1902.0/65536.0,1,-nbitq), 
to_sfixed(755.0/65536.0,1,-nbitq), 
to_sfixed(-3560.0/65536.0,1,-nbitq), 
to_sfixed(537.0/65536.0,1,-nbitq), 
to_sfixed(-1615.0/65536.0,1,-nbitq), 
to_sfixed(357.0/65536.0,1,-nbitq), 
to_sfixed(100.0/65536.0,1,-nbitq), 
to_sfixed(2793.0/65536.0,1,-nbitq), 
to_sfixed(-1429.0/65536.0,1,-nbitq), 
to_sfixed(-432.0/65536.0,1,-nbitq), 
to_sfixed(1298.0/65536.0,1,-nbitq), 
to_sfixed(909.0/65536.0,1,-nbitq), 
to_sfixed(2400.0/65536.0,1,-nbitq), 
to_sfixed(-654.0/65536.0,1,-nbitq), 
to_sfixed(-316.0/65536.0,1,-nbitq), 
to_sfixed(-2614.0/65536.0,1,-nbitq), 
to_sfixed(2397.0/65536.0,1,-nbitq), 
to_sfixed(-1493.0/65536.0,1,-nbitq), 
to_sfixed(-3662.0/65536.0,1,-nbitq), 
to_sfixed(-2315.0/65536.0,1,-nbitq), 
to_sfixed(-708.0/65536.0,1,-nbitq), 
to_sfixed(-132.0/65536.0,1,-nbitq), 
to_sfixed(-551.0/65536.0,1,-nbitq), 
to_sfixed(1255.0/65536.0,1,-nbitq), 
to_sfixed(-2749.0/65536.0,1,-nbitq), 
to_sfixed(3273.0/65536.0,1,-nbitq), 
to_sfixed(2933.0/65536.0,1,-nbitq), 
to_sfixed(3654.0/65536.0,1,-nbitq), 
to_sfixed(-2734.0/65536.0,1,-nbitq), 
to_sfixed(2309.0/65536.0,1,-nbitq), 
to_sfixed(2855.0/65536.0,1,-nbitq), 
to_sfixed(2613.0/65536.0,1,-nbitq), 
to_sfixed(-2483.0/65536.0,1,-nbitq), 
to_sfixed(3319.0/65536.0,1,-nbitq), 
to_sfixed(1578.0/65536.0,1,-nbitq), 
to_sfixed(-2325.0/65536.0,1,-nbitq), 
to_sfixed(1146.0/65536.0,1,-nbitq), 
to_sfixed(-92.0/65536.0,1,-nbitq), 
to_sfixed(2912.0/65536.0,1,-nbitq), 
to_sfixed(2315.0/65536.0,1,-nbitq), 
to_sfixed(-310.0/65536.0,1,-nbitq), 
to_sfixed(4716.0/65536.0,1,-nbitq), 
to_sfixed(-1211.0/65536.0,1,-nbitq), 
to_sfixed(-2844.0/65536.0,1,-nbitq), 
to_sfixed(-995.0/65536.0,1,-nbitq), 
to_sfixed(-1475.0/65536.0,1,-nbitq), 
to_sfixed(2028.0/65536.0,1,-nbitq), 
to_sfixed(182.0/65536.0,1,-nbitq), 
to_sfixed(3493.0/65536.0,1,-nbitq), 
to_sfixed(-2103.0/65536.0,1,-nbitq), 
to_sfixed(5057.0/65536.0,1,-nbitq), 
to_sfixed(-2189.0/65536.0,1,-nbitq), 
to_sfixed(63.0/65536.0,1,-nbitq), 
to_sfixed(3942.0/65536.0,1,-nbitq), 
to_sfixed(2007.0/65536.0,1,-nbitq), 
to_sfixed(2118.0/65536.0,1,-nbitq), 
to_sfixed(-2835.0/65536.0,1,-nbitq), 
to_sfixed(-2138.0/65536.0,1,-nbitq), 
to_sfixed(-3213.0/65536.0,1,-nbitq), 
to_sfixed(1174.0/65536.0,1,-nbitq), 
to_sfixed(-719.0/65536.0,1,-nbitq), 
to_sfixed(126.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-714.0/65536.0,1,-nbitq), 
to_sfixed(-1472.0/65536.0,1,-nbitq), 
to_sfixed(2534.0/65536.0,1,-nbitq), 
to_sfixed(34.0/65536.0,1,-nbitq), 
to_sfixed(-3003.0/65536.0,1,-nbitq), 
to_sfixed(-3602.0/65536.0,1,-nbitq), 
to_sfixed(-3454.0/65536.0,1,-nbitq), 
to_sfixed(-1214.0/65536.0,1,-nbitq), 
to_sfixed(-1046.0/65536.0,1,-nbitq), 
to_sfixed(787.0/65536.0,1,-nbitq), 
to_sfixed(-3637.0/65536.0,1,-nbitq), 
to_sfixed(-3104.0/65536.0,1,-nbitq), 
to_sfixed(-1225.0/65536.0,1,-nbitq), 
to_sfixed(-3196.0/65536.0,1,-nbitq), 
to_sfixed(-282.0/65536.0,1,-nbitq), 
to_sfixed(-1146.0/65536.0,1,-nbitq), 
to_sfixed(675.0/65536.0,1,-nbitq), 
to_sfixed(-463.0/65536.0,1,-nbitq), 
to_sfixed(2310.0/65536.0,1,-nbitq), 
to_sfixed(-1370.0/65536.0,1,-nbitq), 
to_sfixed(-3836.0/65536.0,1,-nbitq), 
to_sfixed(2323.0/65536.0,1,-nbitq), 
to_sfixed(402.0/65536.0,1,-nbitq), 
to_sfixed(1528.0/65536.0,1,-nbitq), 
to_sfixed(-2497.0/65536.0,1,-nbitq), 
to_sfixed(1369.0/65536.0,1,-nbitq), 
to_sfixed(-3954.0/65536.0,1,-nbitq), 
to_sfixed(-1576.0/65536.0,1,-nbitq), 
to_sfixed(-3873.0/65536.0,1,-nbitq), 
to_sfixed(-2279.0/65536.0,1,-nbitq), 
to_sfixed(843.0/65536.0,1,-nbitq), 
to_sfixed(2863.0/65536.0,1,-nbitq), 
to_sfixed(-557.0/65536.0,1,-nbitq), 
to_sfixed(-966.0/65536.0,1,-nbitq), 
to_sfixed(-2504.0/65536.0,1,-nbitq), 
to_sfixed(-696.0/65536.0,1,-nbitq), 
to_sfixed(-1843.0/65536.0,1,-nbitq), 
to_sfixed(-863.0/65536.0,1,-nbitq), 
to_sfixed(1502.0/65536.0,1,-nbitq), 
to_sfixed(-1592.0/65536.0,1,-nbitq), 
to_sfixed(-2757.0/65536.0,1,-nbitq), 
to_sfixed(1533.0/65536.0,1,-nbitq), 
to_sfixed(-5071.0/65536.0,1,-nbitq), 
to_sfixed(5214.0/65536.0,1,-nbitq), 
to_sfixed(2164.0/65536.0,1,-nbitq), 
to_sfixed(5243.0/65536.0,1,-nbitq), 
to_sfixed(1779.0/65536.0,1,-nbitq), 
to_sfixed(275.0/65536.0,1,-nbitq), 
to_sfixed(3473.0/65536.0,1,-nbitq), 
to_sfixed(2145.0/65536.0,1,-nbitq), 
to_sfixed(388.0/65536.0,1,-nbitq), 
to_sfixed(-1147.0/65536.0,1,-nbitq), 
to_sfixed(155.0/65536.0,1,-nbitq), 
to_sfixed(-1243.0/65536.0,1,-nbitq), 
to_sfixed(2610.0/65536.0,1,-nbitq), 
to_sfixed(2838.0/65536.0,1,-nbitq), 
to_sfixed(-814.0/65536.0,1,-nbitq), 
to_sfixed(-1661.0/65536.0,1,-nbitq), 
to_sfixed(-1101.0/65536.0,1,-nbitq), 
to_sfixed(574.0/65536.0,1,-nbitq), 
to_sfixed(-444.0/65536.0,1,-nbitq), 
to_sfixed(-917.0/65536.0,1,-nbitq), 
to_sfixed(2514.0/65536.0,1,-nbitq), 
to_sfixed(-841.0/65536.0,1,-nbitq), 
to_sfixed(3455.0/65536.0,1,-nbitq), 
to_sfixed(-843.0/65536.0,1,-nbitq), 
to_sfixed(3040.0/65536.0,1,-nbitq), 
to_sfixed(429.0/65536.0,1,-nbitq), 
to_sfixed(684.0/65536.0,1,-nbitq), 
to_sfixed(338.0/65536.0,1,-nbitq), 
to_sfixed(-2407.0/65536.0,1,-nbitq), 
to_sfixed(-147.0/65536.0,1,-nbitq), 
to_sfixed(2029.0/65536.0,1,-nbitq), 
to_sfixed(-180.0/65536.0,1,-nbitq), 
to_sfixed(2297.0/65536.0,1,-nbitq), 
to_sfixed(985.0/65536.0,1,-nbitq), 
to_sfixed(-292.0/65536.0,1,-nbitq), 
to_sfixed(3824.0/65536.0,1,-nbitq), 
to_sfixed(-2657.0/65536.0,1,-nbitq), 
to_sfixed(-605.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1127.0/65536.0,1,-nbitq), 
to_sfixed(-1284.0/65536.0,1,-nbitq), 
to_sfixed(-1106.0/65536.0,1,-nbitq), 
to_sfixed(1897.0/65536.0,1,-nbitq), 
to_sfixed(-3411.0/65536.0,1,-nbitq), 
to_sfixed(-4117.0/65536.0,1,-nbitq), 
to_sfixed(-30.0/65536.0,1,-nbitq), 
to_sfixed(-335.0/65536.0,1,-nbitq), 
to_sfixed(-3463.0/65536.0,1,-nbitq), 
to_sfixed(-2549.0/65536.0,1,-nbitq), 
to_sfixed(-2563.0/65536.0,1,-nbitq), 
to_sfixed(-3394.0/65536.0,1,-nbitq), 
to_sfixed(626.0/65536.0,1,-nbitq), 
to_sfixed(-954.0/65536.0,1,-nbitq), 
to_sfixed(-1954.0/65536.0,1,-nbitq), 
to_sfixed(-198.0/65536.0,1,-nbitq), 
to_sfixed(2343.0/65536.0,1,-nbitq), 
to_sfixed(1503.0/65536.0,1,-nbitq), 
to_sfixed(2667.0/65536.0,1,-nbitq), 
to_sfixed(3385.0/65536.0,1,-nbitq), 
to_sfixed(-742.0/65536.0,1,-nbitq), 
to_sfixed(-137.0/65536.0,1,-nbitq), 
to_sfixed(50.0/65536.0,1,-nbitq), 
to_sfixed(2214.0/65536.0,1,-nbitq), 
to_sfixed(1505.0/65536.0,1,-nbitq), 
to_sfixed(1599.0/65536.0,1,-nbitq), 
to_sfixed(158.0/65536.0,1,-nbitq), 
to_sfixed(-185.0/65536.0,1,-nbitq), 
to_sfixed(121.0/65536.0,1,-nbitq), 
to_sfixed(-2688.0/65536.0,1,-nbitq), 
to_sfixed(2206.0/65536.0,1,-nbitq), 
to_sfixed(-1632.0/65536.0,1,-nbitq), 
to_sfixed(-3670.0/65536.0,1,-nbitq), 
to_sfixed(-3824.0/65536.0,1,-nbitq), 
to_sfixed(2819.0/65536.0,1,-nbitq), 
to_sfixed(-2105.0/65536.0,1,-nbitq), 
to_sfixed(-3006.0/65536.0,1,-nbitq), 
to_sfixed(-8.0/65536.0,1,-nbitq), 
to_sfixed(-3828.0/65536.0,1,-nbitq), 
to_sfixed(-1741.0/65536.0,1,-nbitq), 
to_sfixed(-217.0/65536.0,1,-nbitq), 
to_sfixed(991.0/65536.0,1,-nbitq), 
to_sfixed(241.0/65536.0,1,-nbitq), 
to_sfixed(1784.0/65536.0,1,-nbitq), 
to_sfixed(2526.0/65536.0,1,-nbitq), 
to_sfixed(3861.0/65536.0,1,-nbitq), 
to_sfixed(1834.0/65536.0,1,-nbitq), 
to_sfixed(571.0/65536.0,1,-nbitq), 
to_sfixed(-2373.0/65536.0,1,-nbitq), 
to_sfixed(-97.0/65536.0,1,-nbitq), 
to_sfixed(41.0/65536.0,1,-nbitq), 
to_sfixed(722.0/65536.0,1,-nbitq), 
to_sfixed(-340.0/65536.0,1,-nbitq), 
to_sfixed(45.0/65536.0,1,-nbitq), 
to_sfixed(1692.0/65536.0,1,-nbitq), 
to_sfixed(1837.0/65536.0,1,-nbitq), 
to_sfixed(-1785.0/65536.0,1,-nbitq), 
to_sfixed(392.0/65536.0,1,-nbitq), 
to_sfixed(-876.0/65536.0,1,-nbitq), 
to_sfixed(5628.0/65536.0,1,-nbitq), 
to_sfixed(1452.0/65536.0,1,-nbitq), 
to_sfixed(2097.0/65536.0,1,-nbitq), 
to_sfixed(-176.0/65536.0,1,-nbitq), 
to_sfixed(1129.0/65536.0,1,-nbitq), 
to_sfixed(3085.0/65536.0,1,-nbitq), 
to_sfixed(232.0/65536.0,1,-nbitq), 
to_sfixed(-1824.0/65536.0,1,-nbitq), 
to_sfixed(-1133.0/65536.0,1,-nbitq), 
to_sfixed(-270.0/65536.0,1,-nbitq), 
to_sfixed(2312.0/65536.0,1,-nbitq), 
to_sfixed(-1605.0/65536.0,1,-nbitq), 
to_sfixed(-1298.0/65536.0,1,-nbitq), 
to_sfixed(1524.0/65536.0,1,-nbitq), 
to_sfixed(-2777.0/65536.0,1,-nbitq), 
to_sfixed(-1730.0/65536.0,1,-nbitq), 
to_sfixed(1938.0/65536.0,1,-nbitq), 
to_sfixed(-2559.0/65536.0,1,-nbitq), 
to_sfixed(3113.0/65536.0,1,-nbitq), 
to_sfixed(2163.0/65536.0,1,-nbitq), 
to_sfixed(2213.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1573.0/65536.0,1,-nbitq), 
to_sfixed(1414.0/65536.0,1,-nbitq), 
to_sfixed(4429.0/65536.0,1,-nbitq), 
to_sfixed(218.0/65536.0,1,-nbitq), 
to_sfixed(-964.0/65536.0,1,-nbitq), 
to_sfixed(-1960.0/65536.0,1,-nbitq), 
to_sfixed(-2313.0/65536.0,1,-nbitq), 
to_sfixed(-345.0/65536.0,1,-nbitq), 
to_sfixed(-945.0/65536.0,1,-nbitq), 
to_sfixed(2234.0/65536.0,1,-nbitq), 
to_sfixed(281.0/65536.0,1,-nbitq), 
to_sfixed(-478.0/65536.0,1,-nbitq), 
to_sfixed(-2545.0/65536.0,1,-nbitq), 
to_sfixed(-3136.0/65536.0,1,-nbitq), 
to_sfixed(901.0/65536.0,1,-nbitq), 
to_sfixed(-38.0/65536.0,1,-nbitq), 
to_sfixed(143.0/65536.0,1,-nbitq), 
to_sfixed(-1984.0/65536.0,1,-nbitq), 
to_sfixed(1624.0/65536.0,1,-nbitq), 
to_sfixed(1256.0/65536.0,1,-nbitq), 
to_sfixed(-1333.0/65536.0,1,-nbitq), 
to_sfixed(-2095.0/65536.0,1,-nbitq), 
to_sfixed(1406.0/65536.0,1,-nbitq), 
to_sfixed(3317.0/65536.0,1,-nbitq), 
to_sfixed(-1369.0/65536.0,1,-nbitq), 
to_sfixed(952.0/65536.0,1,-nbitq), 
to_sfixed(-2912.0/65536.0,1,-nbitq), 
to_sfixed(-1662.0/65536.0,1,-nbitq), 
to_sfixed(1026.0/65536.0,1,-nbitq), 
to_sfixed(-3345.0/65536.0,1,-nbitq), 
to_sfixed(-1880.0/65536.0,1,-nbitq), 
to_sfixed(2845.0/65536.0,1,-nbitq), 
to_sfixed(-2403.0/65536.0,1,-nbitq), 
to_sfixed(-2136.0/65536.0,1,-nbitq), 
to_sfixed(2713.0/65536.0,1,-nbitq), 
to_sfixed(-2626.0/65536.0,1,-nbitq), 
to_sfixed(1885.0/65536.0,1,-nbitq), 
to_sfixed(1152.0/65536.0,1,-nbitq), 
to_sfixed(-2851.0/65536.0,1,-nbitq), 
to_sfixed(-1851.0/65536.0,1,-nbitq), 
to_sfixed(114.0/65536.0,1,-nbitq), 
to_sfixed(-2230.0/65536.0,1,-nbitq), 
to_sfixed(-4467.0/65536.0,1,-nbitq), 
to_sfixed(264.0/65536.0,1,-nbitq), 
to_sfixed(-231.0/65536.0,1,-nbitq), 
to_sfixed(343.0/65536.0,1,-nbitq), 
to_sfixed(1221.0/65536.0,1,-nbitq), 
to_sfixed(699.0/65536.0,1,-nbitq), 
to_sfixed(3472.0/65536.0,1,-nbitq), 
to_sfixed(-11.0/65536.0,1,-nbitq), 
to_sfixed(2887.0/65536.0,1,-nbitq), 
to_sfixed(1416.0/65536.0,1,-nbitq), 
to_sfixed(1849.0/65536.0,1,-nbitq), 
to_sfixed(-1708.0/65536.0,1,-nbitq), 
to_sfixed(1023.0/65536.0,1,-nbitq), 
to_sfixed(-2054.0/65536.0,1,-nbitq), 
to_sfixed(2438.0/65536.0,1,-nbitq), 
to_sfixed(-50.0/65536.0,1,-nbitq), 
to_sfixed(836.0/65536.0,1,-nbitq), 
to_sfixed(4134.0/65536.0,1,-nbitq), 
to_sfixed(-2456.0/65536.0,1,-nbitq), 
to_sfixed(346.0/65536.0,1,-nbitq), 
to_sfixed(-617.0/65536.0,1,-nbitq), 
to_sfixed(1397.0/65536.0,1,-nbitq), 
to_sfixed(-1644.0/65536.0,1,-nbitq), 
to_sfixed(3952.0/65536.0,1,-nbitq), 
to_sfixed(2017.0/65536.0,1,-nbitq), 
to_sfixed(-4367.0/65536.0,1,-nbitq), 
to_sfixed(3120.0/65536.0,1,-nbitq), 
to_sfixed(2410.0/65536.0,1,-nbitq), 
to_sfixed(1485.0/65536.0,1,-nbitq), 
to_sfixed(2789.0/65536.0,1,-nbitq), 
to_sfixed(1130.0/65536.0,1,-nbitq), 
to_sfixed(-1068.0/65536.0,1,-nbitq), 
to_sfixed(-2676.0/65536.0,1,-nbitq), 
to_sfixed(4184.0/65536.0,1,-nbitq), 
to_sfixed(2101.0/65536.0,1,-nbitq), 
to_sfixed(-525.0/65536.0,1,-nbitq), 
to_sfixed(903.0/65536.0,1,-nbitq), 
to_sfixed(3245.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1019.0/65536.0,1,-nbitq), 
to_sfixed(-516.0/65536.0,1,-nbitq), 
to_sfixed(1587.0/65536.0,1,-nbitq), 
to_sfixed(-982.0/65536.0,1,-nbitq), 
to_sfixed(-3723.0/65536.0,1,-nbitq), 
to_sfixed(-2229.0/65536.0,1,-nbitq), 
to_sfixed(-3263.0/65536.0,1,-nbitq), 
to_sfixed(-2859.0/65536.0,1,-nbitq), 
to_sfixed(-462.0/65536.0,1,-nbitq), 
to_sfixed(737.0/65536.0,1,-nbitq), 
to_sfixed(453.0/65536.0,1,-nbitq), 
to_sfixed(-3432.0/65536.0,1,-nbitq), 
to_sfixed(1257.0/65536.0,1,-nbitq), 
to_sfixed(105.0/65536.0,1,-nbitq), 
to_sfixed(445.0/65536.0,1,-nbitq), 
to_sfixed(2598.0/65536.0,1,-nbitq), 
to_sfixed(1583.0/65536.0,1,-nbitq), 
to_sfixed(-244.0/65536.0,1,-nbitq), 
to_sfixed(2156.0/65536.0,1,-nbitq), 
to_sfixed(1449.0/65536.0,1,-nbitq), 
to_sfixed(2059.0/65536.0,1,-nbitq), 
to_sfixed(-2462.0/65536.0,1,-nbitq), 
to_sfixed(1981.0/65536.0,1,-nbitq), 
to_sfixed(1836.0/65536.0,1,-nbitq), 
to_sfixed(-2498.0/65536.0,1,-nbitq), 
to_sfixed(3508.0/65536.0,1,-nbitq), 
to_sfixed(560.0/65536.0,1,-nbitq), 
to_sfixed(-2423.0/65536.0,1,-nbitq), 
to_sfixed(-2805.0/65536.0,1,-nbitq), 
to_sfixed(-1503.0/65536.0,1,-nbitq), 
to_sfixed(764.0/65536.0,1,-nbitq), 
to_sfixed(2809.0/65536.0,1,-nbitq), 
to_sfixed(-3301.0/65536.0,1,-nbitq), 
to_sfixed(-537.0/65536.0,1,-nbitq), 
to_sfixed(2873.0/65536.0,1,-nbitq), 
to_sfixed(-641.0/65536.0,1,-nbitq), 
to_sfixed(697.0/65536.0,1,-nbitq), 
to_sfixed(1160.0/65536.0,1,-nbitq), 
to_sfixed(1171.0/65536.0,1,-nbitq), 
to_sfixed(-1750.0/65536.0,1,-nbitq), 
to_sfixed(-2375.0/65536.0,1,-nbitq), 
to_sfixed(450.0/65536.0,1,-nbitq), 
to_sfixed(-450.0/65536.0,1,-nbitq), 
to_sfixed(163.0/65536.0,1,-nbitq), 
to_sfixed(-443.0/65536.0,1,-nbitq), 
to_sfixed(1704.0/65536.0,1,-nbitq), 
to_sfixed(-65.0/65536.0,1,-nbitq), 
to_sfixed(-1314.0/65536.0,1,-nbitq), 
to_sfixed(2057.0/65536.0,1,-nbitq), 
to_sfixed(-1030.0/65536.0,1,-nbitq), 
to_sfixed(2723.0/65536.0,1,-nbitq), 
to_sfixed(-1916.0/65536.0,1,-nbitq), 
to_sfixed(2503.0/65536.0,1,-nbitq), 
to_sfixed(398.0/65536.0,1,-nbitq), 
to_sfixed(855.0/65536.0,1,-nbitq), 
to_sfixed(913.0/65536.0,1,-nbitq), 
to_sfixed(-715.0/65536.0,1,-nbitq), 
to_sfixed(1610.0/65536.0,1,-nbitq), 
to_sfixed(265.0/65536.0,1,-nbitq), 
to_sfixed(3569.0/65536.0,1,-nbitq), 
to_sfixed(673.0/65536.0,1,-nbitq), 
to_sfixed(-462.0/65536.0,1,-nbitq), 
to_sfixed(2479.0/65536.0,1,-nbitq), 
to_sfixed(-445.0/65536.0,1,-nbitq), 
to_sfixed(2277.0/65536.0,1,-nbitq), 
to_sfixed(942.0/65536.0,1,-nbitq), 
to_sfixed(1602.0/65536.0,1,-nbitq), 
to_sfixed(-1230.0/65536.0,1,-nbitq), 
to_sfixed(2854.0/65536.0,1,-nbitq), 
to_sfixed(-60.0/65536.0,1,-nbitq), 
to_sfixed(2876.0/65536.0,1,-nbitq), 
to_sfixed(-1886.0/65536.0,1,-nbitq), 
to_sfixed(4427.0/65536.0,1,-nbitq), 
to_sfixed(1048.0/65536.0,1,-nbitq), 
to_sfixed(159.0/65536.0,1,-nbitq), 
to_sfixed(-761.0/65536.0,1,-nbitq), 
to_sfixed(2016.0/65536.0,1,-nbitq), 
to_sfixed(3512.0/65536.0,1,-nbitq), 
to_sfixed(-681.0/65536.0,1,-nbitq), 
to_sfixed(1104.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1682.0/65536.0,1,-nbitq), 
to_sfixed(799.0/65536.0,1,-nbitq), 
to_sfixed(4552.0/65536.0,1,-nbitq), 
to_sfixed(1021.0/65536.0,1,-nbitq), 
to_sfixed(-777.0/65536.0,1,-nbitq), 
to_sfixed(-2507.0/65536.0,1,-nbitq), 
to_sfixed(-523.0/65536.0,1,-nbitq), 
to_sfixed(-2584.0/65536.0,1,-nbitq), 
to_sfixed(2086.0/65536.0,1,-nbitq), 
to_sfixed(1702.0/65536.0,1,-nbitq), 
to_sfixed(-1632.0/65536.0,1,-nbitq), 
to_sfixed(-3566.0/65536.0,1,-nbitq), 
to_sfixed(21.0/65536.0,1,-nbitq), 
to_sfixed(-3148.0/65536.0,1,-nbitq), 
to_sfixed(-1591.0/65536.0,1,-nbitq), 
to_sfixed(-441.0/65536.0,1,-nbitq), 
to_sfixed(-1499.0/65536.0,1,-nbitq), 
to_sfixed(-5151.0/65536.0,1,-nbitq), 
to_sfixed(437.0/65536.0,1,-nbitq), 
to_sfixed(3093.0/65536.0,1,-nbitq), 
to_sfixed(-1591.0/65536.0,1,-nbitq), 
to_sfixed(2336.0/65536.0,1,-nbitq), 
to_sfixed(1304.0/65536.0,1,-nbitq), 
to_sfixed(-2372.0/65536.0,1,-nbitq), 
to_sfixed(1099.0/65536.0,1,-nbitq), 
to_sfixed(1143.0/65536.0,1,-nbitq), 
to_sfixed(-3684.0/65536.0,1,-nbitq), 
to_sfixed(89.0/65536.0,1,-nbitq), 
to_sfixed(-5732.0/65536.0,1,-nbitq), 
to_sfixed(-3373.0/65536.0,1,-nbitq), 
to_sfixed(1996.0/65536.0,1,-nbitq), 
to_sfixed(-2807.0/65536.0,1,-nbitq), 
to_sfixed(-1438.0/65536.0,1,-nbitq), 
to_sfixed(1378.0/65536.0,1,-nbitq), 
to_sfixed(1769.0/65536.0,1,-nbitq), 
to_sfixed(1056.0/65536.0,1,-nbitq), 
to_sfixed(4705.0/65536.0,1,-nbitq), 
to_sfixed(-2277.0/65536.0,1,-nbitq), 
to_sfixed(3159.0/65536.0,1,-nbitq), 
to_sfixed(1489.0/65536.0,1,-nbitq), 
to_sfixed(786.0/65536.0,1,-nbitq), 
to_sfixed(2424.0/65536.0,1,-nbitq), 
to_sfixed(-4417.0/65536.0,1,-nbitq), 
to_sfixed(5502.0/65536.0,1,-nbitq), 
to_sfixed(-1699.0/65536.0,1,-nbitq), 
to_sfixed(4715.0/65536.0,1,-nbitq), 
to_sfixed(3008.0/65536.0,1,-nbitq), 
to_sfixed(-1481.0/65536.0,1,-nbitq), 
to_sfixed(-2052.0/65536.0,1,-nbitq), 
to_sfixed(-503.0/65536.0,1,-nbitq), 
to_sfixed(704.0/65536.0,1,-nbitq), 
to_sfixed(3119.0/65536.0,1,-nbitq), 
to_sfixed(2822.0/65536.0,1,-nbitq), 
to_sfixed(-4781.0/65536.0,1,-nbitq), 
to_sfixed(168.0/65536.0,1,-nbitq), 
to_sfixed(1957.0/65536.0,1,-nbitq), 
to_sfixed(919.0/65536.0,1,-nbitq), 
to_sfixed(-1280.0/65536.0,1,-nbitq), 
to_sfixed(-106.0/65536.0,1,-nbitq), 
to_sfixed(4145.0/65536.0,1,-nbitq), 
to_sfixed(-2753.0/65536.0,1,-nbitq), 
to_sfixed(1655.0/65536.0,1,-nbitq), 
to_sfixed(-1767.0/65536.0,1,-nbitq), 
to_sfixed(-2857.0/65536.0,1,-nbitq), 
to_sfixed(1304.0/65536.0,1,-nbitq), 
to_sfixed(-3785.0/65536.0,1,-nbitq), 
to_sfixed(3213.0/65536.0,1,-nbitq), 
to_sfixed(-1698.0/65536.0,1,-nbitq), 
to_sfixed(-906.0/65536.0,1,-nbitq), 
to_sfixed(2730.0/65536.0,1,-nbitq), 
to_sfixed(3085.0/65536.0,1,-nbitq), 
to_sfixed(-1931.0/65536.0,1,-nbitq), 
to_sfixed(-1326.0/65536.0,1,-nbitq), 
to_sfixed(-1155.0/65536.0,1,-nbitq), 
to_sfixed(1185.0/65536.0,1,-nbitq), 
to_sfixed(820.0/65536.0,1,-nbitq), 
to_sfixed(-867.0/65536.0,1,-nbitq), 
to_sfixed(3511.0/65536.0,1,-nbitq), 
to_sfixed(-3194.0/65536.0,1,-nbitq), 
to_sfixed(3442.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2834.0/65536.0,1,-nbitq), 
to_sfixed(958.0/65536.0,1,-nbitq), 
to_sfixed(2789.0/65536.0,1,-nbitq), 
to_sfixed(462.0/65536.0,1,-nbitq), 
to_sfixed(204.0/65536.0,1,-nbitq), 
to_sfixed(-2756.0/65536.0,1,-nbitq), 
to_sfixed(482.0/65536.0,1,-nbitq), 
to_sfixed(-1517.0/65536.0,1,-nbitq), 
to_sfixed(16.0/65536.0,1,-nbitq), 
to_sfixed(1101.0/65536.0,1,-nbitq), 
to_sfixed(-2952.0/65536.0,1,-nbitq), 
to_sfixed(-3875.0/65536.0,1,-nbitq), 
to_sfixed(1930.0/65536.0,1,-nbitq), 
to_sfixed(-3475.0/65536.0,1,-nbitq), 
to_sfixed(-741.0/65536.0,1,-nbitq), 
to_sfixed(1355.0/65536.0,1,-nbitq), 
to_sfixed(-1791.0/65536.0,1,-nbitq), 
to_sfixed(-1681.0/65536.0,1,-nbitq), 
to_sfixed(-4654.0/65536.0,1,-nbitq), 
to_sfixed(368.0/65536.0,1,-nbitq), 
to_sfixed(-521.0/65536.0,1,-nbitq), 
to_sfixed(-2297.0/65536.0,1,-nbitq), 
to_sfixed(-1950.0/65536.0,1,-nbitq), 
to_sfixed(435.0/65536.0,1,-nbitq), 
to_sfixed(-2006.0/65536.0,1,-nbitq), 
to_sfixed(236.0/65536.0,1,-nbitq), 
to_sfixed(-1759.0/65536.0,1,-nbitq), 
to_sfixed(1515.0/65536.0,1,-nbitq), 
to_sfixed(-1648.0/65536.0,1,-nbitq), 
to_sfixed(199.0/65536.0,1,-nbitq), 
to_sfixed(441.0/65536.0,1,-nbitq), 
to_sfixed(-3868.0/65536.0,1,-nbitq), 
to_sfixed(-1503.0/65536.0,1,-nbitq), 
to_sfixed(-539.0/65536.0,1,-nbitq), 
to_sfixed(-265.0/65536.0,1,-nbitq), 
to_sfixed(742.0/65536.0,1,-nbitq), 
to_sfixed(2821.0/65536.0,1,-nbitq), 
to_sfixed(598.0/65536.0,1,-nbitq), 
to_sfixed(3733.0/65536.0,1,-nbitq), 
to_sfixed(3401.0/65536.0,1,-nbitq), 
to_sfixed(1539.0/65536.0,1,-nbitq), 
to_sfixed(-2779.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(772.0/65536.0,1,-nbitq), 
to_sfixed(1806.0/65536.0,1,-nbitq), 
to_sfixed(3793.0/65536.0,1,-nbitq), 
to_sfixed(2046.0/65536.0,1,-nbitq), 
to_sfixed(441.0/65536.0,1,-nbitq), 
to_sfixed(-623.0/65536.0,1,-nbitq), 
to_sfixed(2210.0/65536.0,1,-nbitq), 
to_sfixed(306.0/65536.0,1,-nbitq), 
to_sfixed(1344.0/65536.0,1,-nbitq), 
to_sfixed(1927.0/65536.0,1,-nbitq), 
to_sfixed(-4341.0/65536.0,1,-nbitq), 
to_sfixed(-1734.0/65536.0,1,-nbitq), 
to_sfixed(-2627.0/65536.0,1,-nbitq), 
to_sfixed(2408.0/65536.0,1,-nbitq), 
to_sfixed(2749.0/65536.0,1,-nbitq), 
to_sfixed(-367.0/65536.0,1,-nbitq), 
to_sfixed(562.0/65536.0,1,-nbitq), 
to_sfixed(864.0/65536.0,1,-nbitq), 
to_sfixed(-2348.0/65536.0,1,-nbitq), 
to_sfixed(684.0/65536.0,1,-nbitq), 
to_sfixed(-2252.0/65536.0,1,-nbitq), 
to_sfixed(2119.0/65536.0,1,-nbitq), 
to_sfixed(-5257.0/65536.0,1,-nbitq), 
to_sfixed(3417.0/65536.0,1,-nbitq), 
to_sfixed(-4161.0/65536.0,1,-nbitq), 
to_sfixed(46.0/65536.0,1,-nbitq), 
to_sfixed(4608.0/65536.0,1,-nbitq), 
to_sfixed(417.0/65536.0,1,-nbitq), 
to_sfixed(-867.0/65536.0,1,-nbitq), 
to_sfixed(1868.0/65536.0,1,-nbitq), 
to_sfixed(-937.0/65536.0,1,-nbitq), 
to_sfixed(-1891.0/65536.0,1,-nbitq), 
to_sfixed(-579.0/65536.0,1,-nbitq), 
to_sfixed(-5061.0/65536.0,1,-nbitq), 
to_sfixed(-1336.0/65536.0,1,-nbitq), 
to_sfixed(-1171.0/65536.0,1,-nbitq), 
to_sfixed(3145.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-225.0/65536.0,1,-nbitq), 
to_sfixed(-841.0/65536.0,1,-nbitq), 
to_sfixed(2172.0/65536.0,1,-nbitq), 
to_sfixed(1156.0/65536.0,1,-nbitq), 
to_sfixed(4952.0/65536.0,1,-nbitq), 
to_sfixed(-484.0/65536.0,1,-nbitq), 
to_sfixed(1065.0/65536.0,1,-nbitq), 
to_sfixed(105.0/65536.0,1,-nbitq), 
to_sfixed(-1485.0/65536.0,1,-nbitq), 
to_sfixed(2339.0/65536.0,1,-nbitq), 
to_sfixed(488.0/65536.0,1,-nbitq), 
to_sfixed(-11320.0/65536.0,1,-nbitq), 
to_sfixed(-1906.0/65536.0,1,-nbitq), 
to_sfixed(-3249.0/65536.0,1,-nbitq), 
to_sfixed(-1756.0/65536.0,1,-nbitq), 
to_sfixed(349.0/65536.0,1,-nbitq), 
to_sfixed(-2332.0/65536.0,1,-nbitq), 
to_sfixed(-5081.0/65536.0,1,-nbitq), 
to_sfixed(-3703.0/65536.0,1,-nbitq), 
to_sfixed(3228.0/65536.0,1,-nbitq), 
to_sfixed(1568.0/65536.0,1,-nbitq), 
to_sfixed(-3190.0/65536.0,1,-nbitq), 
to_sfixed(-3265.0/65536.0,1,-nbitq), 
to_sfixed(-7145.0/65536.0,1,-nbitq), 
to_sfixed(891.0/65536.0,1,-nbitq), 
to_sfixed(-3231.0/65536.0,1,-nbitq), 
to_sfixed(-267.0/65536.0,1,-nbitq), 
to_sfixed(-350.0/65536.0,1,-nbitq), 
to_sfixed(6428.0/65536.0,1,-nbitq), 
to_sfixed(-4672.0/65536.0,1,-nbitq), 
to_sfixed(-464.0/65536.0,1,-nbitq), 
to_sfixed(-2866.0/65536.0,1,-nbitq), 
to_sfixed(-2124.0/65536.0,1,-nbitq), 
to_sfixed(-421.0/65536.0,1,-nbitq), 
to_sfixed(-1707.0/65536.0,1,-nbitq), 
to_sfixed(1316.0/65536.0,1,-nbitq), 
to_sfixed(4787.0/65536.0,1,-nbitq), 
to_sfixed(-281.0/65536.0,1,-nbitq), 
to_sfixed(4657.0/65536.0,1,-nbitq), 
to_sfixed(-2613.0/65536.0,1,-nbitq), 
to_sfixed(2305.0/65536.0,1,-nbitq), 
to_sfixed(-1086.0/65536.0,1,-nbitq), 
to_sfixed(2276.0/65536.0,1,-nbitq), 
to_sfixed(1742.0/65536.0,1,-nbitq), 
to_sfixed(-1432.0/65536.0,1,-nbitq), 
to_sfixed(2289.0/65536.0,1,-nbitq), 
to_sfixed(378.0/65536.0,1,-nbitq), 
to_sfixed(1824.0/65536.0,1,-nbitq), 
to_sfixed(2370.0/65536.0,1,-nbitq), 
to_sfixed(-376.0/65536.0,1,-nbitq), 
to_sfixed(3051.0/65536.0,1,-nbitq), 
to_sfixed(-915.0/65536.0,1,-nbitq), 
to_sfixed(1054.0/65536.0,1,-nbitq), 
to_sfixed(2359.0/65536.0,1,-nbitq), 
to_sfixed(-2550.0/65536.0,1,-nbitq), 
to_sfixed(-2991.0/65536.0,1,-nbitq), 
to_sfixed(-873.0/65536.0,1,-nbitq), 
to_sfixed(1229.0/65536.0,1,-nbitq), 
to_sfixed(1351.0/65536.0,1,-nbitq), 
to_sfixed(-4599.0/65536.0,1,-nbitq), 
to_sfixed(-2034.0/65536.0,1,-nbitq), 
to_sfixed(2463.0/65536.0,1,-nbitq), 
to_sfixed(2199.0/65536.0,1,-nbitq), 
to_sfixed(1532.0/65536.0,1,-nbitq), 
to_sfixed(3942.0/65536.0,1,-nbitq), 
to_sfixed(-4316.0/65536.0,1,-nbitq), 
to_sfixed(2923.0/65536.0,1,-nbitq), 
to_sfixed(-2712.0/65536.0,1,-nbitq), 
to_sfixed(4642.0/65536.0,1,-nbitq), 
to_sfixed(3769.0/65536.0,1,-nbitq), 
to_sfixed(-1437.0/65536.0,1,-nbitq), 
to_sfixed(-425.0/65536.0,1,-nbitq), 
to_sfixed(-1657.0/65536.0,1,-nbitq), 
to_sfixed(-1642.0/65536.0,1,-nbitq), 
to_sfixed(1844.0/65536.0,1,-nbitq), 
to_sfixed(3523.0/65536.0,1,-nbitq), 
to_sfixed(-4780.0/65536.0,1,-nbitq), 
to_sfixed(5052.0/65536.0,1,-nbitq), 
to_sfixed(-3017.0/65536.0,1,-nbitq), 
to_sfixed(3654.0/65536.0,1,-nbitq)  ), 
( to_sfixed(360.0/65536.0,1,-nbitq), 
to_sfixed(6246.0/65536.0,1,-nbitq), 
to_sfixed(6704.0/65536.0,1,-nbitq), 
to_sfixed(357.0/65536.0,1,-nbitq), 
to_sfixed(3481.0/65536.0,1,-nbitq), 
to_sfixed(-7066.0/65536.0,1,-nbitq), 
to_sfixed(1608.0/65536.0,1,-nbitq), 
to_sfixed(-3173.0/65536.0,1,-nbitq), 
to_sfixed(-2222.0/65536.0,1,-nbitq), 
to_sfixed(2471.0/65536.0,1,-nbitq), 
to_sfixed(654.0/65536.0,1,-nbitq), 
to_sfixed(-5194.0/65536.0,1,-nbitq), 
to_sfixed(2128.0/65536.0,1,-nbitq), 
to_sfixed(344.0/65536.0,1,-nbitq), 
to_sfixed(-1663.0/65536.0,1,-nbitq), 
to_sfixed(1767.0/65536.0,1,-nbitq), 
to_sfixed(-663.0/65536.0,1,-nbitq), 
to_sfixed(-3000.0/65536.0,1,-nbitq), 
to_sfixed(-5385.0/65536.0,1,-nbitq), 
to_sfixed(3192.0/65536.0,1,-nbitq), 
to_sfixed(3116.0/65536.0,1,-nbitq), 
to_sfixed(-832.0/65536.0,1,-nbitq), 
to_sfixed(-504.0/65536.0,1,-nbitq), 
to_sfixed(-11590.0/65536.0,1,-nbitq), 
to_sfixed(-3931.0/65536.0,1,-nbitq), 
to_sfixed(-10553.0/65536.0,1,-nbitq), 
to_sfixed(-2507.0/65536.0,1,-nbitq), 
to_sfixed(1302.0/65536.0,1,-nbitq), 
to_sfixed(5100.0/65536.0,1,-nbitq), 
to_sfixed(129.0/65536.0,1,-nbitq), 
to_sfixed(3559.0/65536.0,1,-nbitq), 
to_sfixed(1699.0/65536.0,1,-nbitq), 
to_sfixed(4902.0/65536.0,1,-nbitq), 
to_sfixed(5089.0/65536.0,1,-nbitq), 
to_sfixed(-2131.0/65536.0,1,-nbitq), 
to_sfixed(-499.0/65536.0,1,-nbitq), 
to_sfixed(3680.0/65536.0,1,-nbitq), 
to_sfixed(91.0/65536.0,1,-nbitq), 
to_sfixed(4064.0/65536.0,1,-nbitq), 
to_sfixed(-3397.0/65536.0,1,-nbitq), 
to_sfixed(2489.0/65536.0,1,-nbitq), 
to_sfixed(512.0/65536.0,1,-nbitq), 
to_sfixed(6900.0/65536.0,1,-nbitq), 
to_sfixed(-3411.0/65536.0,1,-nbitq), 
to_sfixed(2138.0/65536.0,1,-nbitq), 
to_sfixed(3147.0/65536.0,1,-nbitq), 
to_sfixed(-1025.0/65536.0,1,-nbitq), 
to_sfixed(5351.0/65536.0,1,-nbitq), 
to_sfixed(940.0/65536.0,1,-nbitq), 
to_sfixed(2570.0/65536.0,1,-nbitq), 
to_sfixed(1536.0/65536.0,1,-nbitq), 
to_sfixed(2565.0/65536.0,1,-nbitq), 
to_sfixed(407.0/65536.0,1,-nbitq), 
to_sfixed(6335.0/65536.0,1,-nbitq), 
to_sfixed(-858.0/65536.0,1,-nbitq), 
to_sfixed(238.0/65536.0,1,-nbitq), 
to_sfixed(-2034.0/65536.0,1,-nbitq), 
to_sfixed(4017.0/65536.0,1,-nbitq), 
to_sfixed(-2633.0/65536.0,1,-nbitq), 
to_sfixed(-4151.0/65536.0,1,-nbitq), 
to_sfixed(-1767.0/65536.0,1,-nbitq), 
to_sfixed(436.0/65536.0,1,-nbitq), 
to_sfixed(-537.0/65536.0,1,-nbitq), 
to_sfixed(-962.0/65536.0,1,-nbitq), 
to_sfixed(-3734.0/65536.0,1,-nbitq), 
to_sfixed(-3687.0/65536.0,1,-nbitq), 
to_sfixed(4754.0/65536.0,1,-nbitq), 
to_sfixed(-3269.0/65536.0,1,-nbitq), 
to_sfixed(5841.0/65536.0,1,-nbitq), 
to_sfixed(4235.0/65536.0,1,-nbitq), 
to_sfixed(1634.0/65536.0,1,-nbitq), 
to_sfixed(931.0/65536.0,1,-nbitq), 
to_sfixed(-1046.0/65536.0,1,-nbitq), 
to_sfixed(-2714.0/65536.0,1,-nbitq), 
to_sfixed(1840.0/65536.0,1,-nbitq), 
to_sfixed(1361.0/65536.0,1,-nbitq), 
to_sfixed(-2258.0/65536.0,1,-nbitq), 
to_sfixed(2818.0/65536.0,1,-nbitq), 
to_sfixed(-1117.0/65536.0,1,-nbitq), 
to_sfixed(-1869.0/65536.0,1,-nbitq)  ), 
( to_sfixed(773.0/65536.0,1,-nbitq), 
to_sfixed(3820.0/65536.0,1,-nbitq), 
to_sfixed(2886.0/65536.0,1,-nbitq), 
to_sfixed(1562.0/65536.0,1,-nbitq), 
to_sfixed(-2896.0/65536.0,1,-nbitq), 
to_sfixed(-8919.0/65536.0,1,-nbitq), 
to_sfixed(1210.0/65536.0,1,-nbitq), 
to_sfixed(-2247.0/65536.0,1,-nbitq), 
to_sfixed(-3303.0/65536.0,1,-nbitq), 
to_sfixed(3058.0/65536.0,1,-nbitq), 
to_sfixed(3965.0/65536.0,1,-nbitq), 
to_sfixed(-7366.0/65536.0,1,-nbitq), 
to_sfixed(-1019.0/65536.0,1,-nbitq), 
to_sfixed(-4274.0/65536.0,1,-nbitq), 
to_sfixed(-3866.0/65536.0,1,-nbitq), 
to_sfixed(1072.0/65536.0,1,-nbitq), 
to_sfixed(1915.0/65536.0,1,-nbitq), 
to_sfixed(5717.0/65536.0,1,-nbitq), 
to_sfixed(-10150.0/65536.0,1,-nbitq), 
to_sfixed(-879.0/65536.0,1,-nbitq), 
to_sfixed(7537.0/65536.0,1,-nbitq), 
to_sfixed(423.0/65536.0,1,-nbitq), 
to_sfixed(-1011.0/65536.0,1,-nbitq), 
to_sfixed(-10209.0/65536.0,1,-nbitq), 
to_sfixed(3472.0/65536.0,1,-nbitq), 
to_sfixed(-15549.0/65536.0,1,-nbitq), 
to_sfixed(-2598.0/65536.0,1,-nbitq), 
to_sfixed(-1859.0/65536.0,1,-nbitq), 
to_sfixed(-4314.0/65536.0,1,-nbitq), 
to_sfixed(109.0/65536.0,1,-nbitq), 
to_sfixed(-444.0/65536.0,1,-nbitq), 
to_sfixed(-2873.0/65536.0,1,-nbitq), 
to_sfixed(8324.0/65536.0,1,-nbitq), 
to_sfixed(5215.0/65536.0,1,-nbitq), 
to_sfixed(345.0/65536.0,1,-nbitq), 
to_sfixed(2154.0/65536.0,1,-nbitq), 
to_sfixed(5476.0/65536.0,1,-nbitq), 
to_sfixed(3374.0/65536.0,1,-nbitq), 
to_sfixed(5153.0/65536.0,1,-nbitq), 
to_sfixed(-1655.0/65536.0,1,-nbitq), 
to_sfixed(1900.0/65536.0,1,-nbitq), 
to_sfixed(-988.0/65536.0,1,-nbitq), 
to_sfixed(8004.0/65536.0,1,-nbitq), 
to_sfixed(-719.0/65536.0,1,-nbitq), 
to_sfixed(2662.0/65536.0,1,-nbitq), 
to_sfixed(-4227.0/65536.0,1,-nbitq), 
to_sfixed(-2816.0/65536.0,1,-nbitq), 
to_sfixed(3869.0/65536.0,1,-nbitq), 
to_sfixed(-3082.0/65536.0,1,-nbitq), 
to_sfixed(81.0/65536.0,1,-nbitq), 
to_sfixed(-2411.0/65536.0,1,-nbitq), 
to_sfixed(1372.0/65536.0,1,-nbitq), 
to_sfixed(-833.0/65536.0,1,-nbitq), 
to_sfixed(3732.0/65536.0,1,-nbitq), 
to_sfixed(2316.0/65536.0,1,-nbitq), 
to_sfixed(-1552.0/65536.0,1,-nbitq), 
to_sfixed(-224.0/65536.0,1,-nbitq), 
to_sfixed(-448.0/65536.0,1,-nbitq), 
to_sfixed(364.0/65536.0,1,-nbitq), 
to_sfixed(-5174.0/65536.0,1,-nbitq), 
to_sfixed(5872.0/65536.0,1,-nbitq), 
to_sfixed(2179.0/65536.0,1,-nbitq), 
to_sfixed(2421.0/65536.0,1,-nbitq), 
to_sfixed(-432.0/65536.0,1,-nbitq), 
to_sfixed(-6840.0/65536.0,1,-nbitq), 
to_sfixed(-5271.0/65536.0,1,-nbitq), 
to_sfixed(3378.0/65536.0,1,-nbitq), 
to_sfixed(-1847.0/65536.0,1,-nbitq), 
to_sfixed(-831.0/65536.0,1,-nbitq), 
to_sfixed(4928.0/65536.0,1,-nbitq), 
to_sfixed(-1611.0/65536.0,1,-nbitq), 
to_sfixed(-408.0/65536.0,1,-nbitq), 
to_sfixed(-479.0/65536.0,1,-nbitq), 
to_sfixed(-716.0/65536.0,1,-nbitq), 
to_sfixed(-2848.0/65536.0,1,-nbitq), 
to_sfixed(-1617.0/65536.0,1,-nbitq), 
to_sfixed(-1063.0/65536.0,1,-nbitq), 
to_sfixed(1720.0/65536.0,1,-nbitq), 
to_sfixed(1352.0/65536.0,1,-nbitq), 
to_sfixed(-5219.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1529.0/65536.0,1,-nbitq), 
to_sfixed(-1064.0/65536.0,1,-nbitq), 
to_sfixed(2106.0/65536.0,1,-nbitq), 
to_sfixed(-1229.0/65536.0,1,-nbitq), 
to_sfixed(3941.0/65536.0,1,-nbitq), 
to_sfixed(-4635.0/65536.0,1,-nbitq), 
to_sfixed(-3769.0/65536.0,1,-nbitq), 
to_sfixed(-1333.0/65536.0,1,-nbitq), 
to_sfixed(436.0/65536.0,1,-nbitq), 
to_sfixed(-1099.0/65536.0,1,-nbitq), 
to_sfixed(4576.0/65536.0,1,-nbitq), 
to_sfixed(-10643.0/65536.0,1,-nbitq), 
to_sfixed(1154.0/65536.0,1,-nbitq), 
to_sfixed(-4705.0/65536.0,1,-nbitq), 
to_sfixed(-2583.0/65536.0,1,-nbitq), 
to_sfixed(189.0/65536.0,1,-nbitq), 
to_sfixed(1210.0/65536.0,1,-nbitq), 
to_sfixed(4883.0/65536.0,1,-nbitq), 
to_sfixed(-8130.0/65536.0,1,-nbitq), 
to_sfixed(910.0/65536.0,1,-nbitq), 
to_sfixed(9511.0/65536.0,1,-nbitq), 
to_sfixed(-2445.0/65536.0,1,-nbitq), 
to_sfixed(-2981.0/65536.0,1,-nbitq), 
to_sfixed(-16917.0/65536.0,1,-nbitq), 
to_sfixed(-23.0/65536.0,1,-nbitq), 
to_sfixed(-13978.0/65536.0,1,-nbitq), 
to_sfixed(6018.0/65536.0,1,-nbitq), 
to_sfixed(-50.0/65536.0,1,-nbitq), 
to_sfixed(-3097.0/65536.0,1,-nbitq), 
to_sfixed(-2946.0/65536.0,1,-nbitq), 
to_sfixed(3044.0/65536.0,1,-nbitq), 
to_sfixed(251.0/65536.0,1,-nbitq), 
to_sfixed(3212.0/65536.0,1,-nbitq), 
to_sfixed(3844.0/65536.0,1,-nbitq), 
to_sfixed(1748.0/65536.0,1,-nbitq), 
to_sfixed(-991.0/65536.0,1,-nbitq), 
to_sfixed(3967.0/65536.0,1,-nbitq), 
to_sfixed(3999.0/65536.0,1,-nbitq), 
to_sfixed(7618.0/65536.0,1,-nbitq), 
to_sfixed(-2720.0/65536.0,1,-nbitq), 
to_sfixed(-378.0/65536.0,1,-nbitq), 
to_sfixed(1304.0/65536.0,1,-nbitq), 
to_sfixed(5754.0/65536.0,1,-nbitq), 
to_sfixed(-483.0/65536.0,1,-nbitq), 
to_sfixed(1076.0/65536.0,1,-nbitq), 
to_sfixed(-3974.0/65536.0,1,-nbitq), 
to_sfixed(-781.0/65536.0,1,-nbitq), 
to_sfixed(-556.0/65536.0,1,-nbitq), 
to_sfixed(2187.0/65536.0,1,-nbitq), 
to_sfixed(2384.0/65536.0,1,-nbitq), 
to_sfixed(814.0/65536.0,1,-nbitq), 
to_sfixed(1550.0/65536.0,1,-nbitq), 
to_sfixed(6608.0/65536.0,1,-nbitq), 
to_sfixed(-4413.0/65536.0,1,-nbitq), 
to_sfixed(3164.0/65536.0,1,-nbitq), 
to_sfixed(994.0/65536.0,1,-nbitq), 
to_sfixed(252.0/65536.0,1,-nbitq), 
to_sfixed(1777.0/65536.0,1,-nbitq), 
to_sfixed(1979.0/65536.0,1,-nbitq), 
to_sfixed(-6840.0/65536.0,1,-nbitq), 
to_sfixed(6477.0/65536.0,1,-nbitq), 
to_sfixed(-1987.0/65536.0,1,-nbitq), 
to_sfixed(1862.0/65536.0,1,-nbitq), 
to_sfixed(-2105.0/65536.0,1,-nbitq), 
to_sfixed(-4799.0/65536.0,1,-nbitq), 
to_sfixed(6327.0/65536.0,1,-nbitq), 
to_sfixed(3558.0/65536.0,1,-nbitq), 
to_sfixed(-3800.0/65536.0,1,-nbitq), 
to_sfixed(-1888.0/65536.0,1,-nbitq), 
to_sfixed(-121.0/65536.0,1,-nbitq), 
to_sfixed(2845.0/65536.0,1,-nbitq), 
to_sfixed(-6798.0/65536.0,1,-nbitq), 
to_sfixed(-2326.0/65536.0,1,-nbitq), 
to_sfixed(-2046.0/65536.0,1,-nbitq), 
to_sfixed(2095.0/65536.0,1,-nbitq), 
to_sfixed(2331.0/65536.0,1,-nbitq), 
to_sfixed(3021.0/65536.0,1,-nbitq), 
to_sfixed(3645.0/65536.0,1,-nbitq), 
to_sfixed(-2408.0/65536.0,1,-nbitq), 
to_sfixed(-5707.0/65536.0,1,-nbitq)  ), 
( to_sfixed(806.0/65536.0,1,-nbitq), 
to_sfixed(3726.0/65536.0,1,-nbitq), 
to_sfixed(11812.0/65536.0,1,-nbitq), 
to_sfixed(-4821.0/65536.0,1,-nbitq), 
to_sfixed(-60.0/65536.0,1,-nbitq), 
to_sfixed(2264.0/65536.0,1,-nbitq), 
to_sfixed(-7125.0/65536.0,1,-nbitq), 
to_sfixed(2873.0/65536.0,1,-nbitq), 
to_sfixed(359.0/65536.0,1,-nbitq), 
to_sfixed(2052.0/65536.0,1,-nbitq), 
to_sfixed(-690.0/65536.0,1,-nbitq), 
to_sfixed(-5777.0/65536.0,1,-nbitq), 
to_sfixed(1177.0/65536.0,1,-nbitq), 
to_sfixed(-2228.0/65536.0,1,-nbitq), 
to_sfixed(1392.0/65536.0,1,-nbitq), 
to_sfixed(-1136.0/65536.0,1,-nbitq), 
to_sfixed(-2130.0/65536.0,1,-nbitq), 
to_sfixed(3056.0/65536.0,1,-nbitq), 
to_sfixed(363.0/65536.0,1,-nbitq), 
to_sfixed(1164.0/65536.0,1,-nbitq), 
to_sfixed(5144.0/65536.0,1,-nbitq), 
to_sfixed(6624.0/65536.0,1,-nbitq), 
to_sfixed(-556.0/65536.0,1,-nbitq), 
to_sfixed(-17296.0/65536.0,1,-nbitq), 
to_sfixed(-1508.0/65536.0,1,-nbitq), 
to_sfixed(-11842.0/65536.0,1,-nbitq), 
to_sfixed(9662.0/65536.0,1,-nbitq), 
to_sfixed(-1537.0/65536.0,1,-nbitq), 
to_sfixed(-56.0/65536.0,1,-nbitq), 
to_sfixed(606.0/65536.0,1,-nbitq), 
to_sfixed(-1776.0/65536.0,1,-nbitq), 
to_sfixed(-3612.0/65536.0,1,-nbitq), 
to_sfixed(6255.0/65536.0,1,-nbitq), 
to_sfixed(-1764.0/65536.0,1,-nbitq), 
to_sfixed(-893.0/65536.0,1,-nbitq), 
to_sfixed(-903.0/65536.0,1,-nbitq), 
to_sfixed(6285.0/65536.0,1,-nbitq), 
to_sfixed(-159.0/65536.0,1,-nbitq), 
to_sfixed(6932.0/65536.0,1,-nbitq), 
to_sfixed(-312.0/65536.0,1,-nbitq), 
to_sfixed(-1183.0/65536.0,1,-nbitq), 
to_sfixed(837.0/65536.0,1,-nbitq), 
to_sfixed(4840.0/65536.0,1,-nbitq), 
to_sfixed(-225.0/65536.0,1,-nbitq), 
to_sfixed(-1339.0/65536.0,1,-nbitq), 
to_sfixed(-4232.0/65536.0,1,-nbitq), 
to_sfixed(-788.0/65536.0,1,-nbitq), 
to_sfixed(4489.0/65536.0,1,-nbitq), 
to_sfixed(-194.0/65536.0,1,-nbitq), 
to_sfixed(3312.0/65536.0,1,-nbitq), 
to_sfixed(-591.0/65536.0,1,-nbitq), 
to_sfixed(825.0/65536.0,1,-nbitq), 
to_sfixed(3380.0/65536.0,1,-nbitq), 
to_sfixed(-4668.0/65536.0,1,-nbitq), 
to_sfixed(-1215.0/65536.0,1,-nbitq), 
to_sfixed(-2357.0/65536.0,1,-nbitq), 
to_sfixed(-339.0/65536.0,1,-nbitq), 
to_sfixed(801.0/65536.0,1,-nbitq), 
to_sfixed(-3011.0/65536.0,1,-nbitq), 
to_sfixed(-6580.0/65536.0,1,-nbitq), 
to_sfixed(3951.0/65536.0,1,-nbitq), 
to_sfixed(-1326.0/65536.0,1,-nbitq), 
to_sfixed(-272.0/65536.0,1,-nbitq), 
to_sfixed(-2832.0/65536.0,1,-nbitq), 
to_sfixed(-4511.0/65536.0,1,-nbitq), 
to_sfixed(4882.0/65536.0,1,-nbitq), 
to_sfixed(1838.0/65536.0,1,-nbitq), 
to_sfixed(-844.0/65536.0,1,-nbitq), 
to_sfixed(-5357.0/65536.0,1,-nbitq), 
to_sfixed(3905.0/65536.0,1,-nbitq), 
to_sfixed(146.0/65536.0,1,-nbitq), 
to_sfixed(-2888.0/65536.0,1,-nbitq), 
to_sfixed(-3390.0/65536.0,1,-nbitq), 
to_sfixed(2292.0/65536.0,1,-nbitq), 
to_sfixed(1137.0/65536.0,1,-nbitq), 
to_sfixed(1025.0/65536.0,1,-nbitq), 
to_sfixed(3842.0/65536.0,1,-nbitq), 
to_sfixed(707.0/65536.0,1,-nbitq), 
to_sfixed(575.0/65536.0,1,-nbitq), 
to_sfixed(-1217.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-791.0/65536.0,1,-nbitq), 
to_sfixed(-2125.0/65536.0,1,-nbitq), 
to_sfixed(4616.0/65536.0,1,-nbitq), 
to_sfixed(-5052.0/65536.0,1,-nbitq), 
to_sfixed(3856.0/65536.0,1,-nbitq), 
to_sfixed(-7092.0/65536.0,1,-nbitq), 
to_sfixed(-9423.0/65536.0,1,-nbitq), 
to_sfixed(-2999.0/65536.0,1,-nbitq), 
to_sfixed(5131.0/65536.0,1,-nbitq), 
to_sfixed(2489.0/65536.0,1,-nbitq), 
to_sfixed(-1555.0/65536.0,1,-nbitq), 
to_sfixed(-11495.0/65536.0,1,-nbitq), 
to_sfixed(-2037.0/65536.0,1,-nbitq), 
to_sfixed(5766.0/65536.0,1,-nbitq), 
to_sfixed(-4097.0/65536.0,1,-nbitq), 
to_sfixed(566.0/65536.0,1,-nbitq), 
to_sfixed(-1722.0/65536.0,1,-nbitq), 
to_sfixed(801.0/65536.0,1,-nbitq), 
to_sfixed(2202.0/65536.0,1,-nbitq), 
to_sfixed(199.0/65536.0,1,-nbitq), 
to_sfixed(-554.0/65536.0,1,-nbitq), 
to_sfixed(5519.0/65536.0,1,-nbitq), 
to_sfixed(4864.0/65536.0,1,-nbitq), 
to_sfixed(-3846.0/65536.0,1,-nbitq), 
to_sfixed(-1487.0/65536.0,1,-nbitq), 
to_sfixed(-13508.0/65536.0,1,-nbitq), 
to_sfixed(3937.0/65536.0,1,-nbitq), 
to_sfixed(-3176.0/65536.0,1,-nbitq), 
to_sfixed(-6093.0/65536.0,1,-nbitq), 
to_sfixed(7767.0/65536.0,1,-nbitq), 
to_sfixed(1863.0/65536.0,1,-nbitq), 
to_sfixed(-1785.0/65536.0,1,-nbitq), 
to_sfixed(1839.0/65536.0,1,-nbitq), 
to_sfixed(-3753.0/65536.0,1,-nbitq), 
to_sfixed(1678.0/65536.0,1,-nbitq), 
to_sfixed(2814.0/65536.0,1,-nbitq), 
to_sfixed(9616.0/65536.0,1,-nbitq), 
to_sfixed(-2510.0/65536.0,1,-nbitq), 
to_sfixed(2661.0/65536.0,1,-nbitq), 
to_sfixed(2042.0/65536.0,1,-nbitq), 
to_sfixed(-1641.0/65536.0,1,-nbitq), 
to_sfixed(-355.0/65536.0,1,-nbitq), 
to_sfixed(-6920.0/65536.0,1,-nbitq), 
to_sfixed(-2013.0/65536.0,1,-nbitq), 
to_sfixed(2759.0/65536.0,1,-nbitq), 
to_sfixed(-10980.0/65536.0,1,-nbitq), 
to_sfixed(-1754.0/65536.0,1,-nbitq), 
to_sfixed(4182.0/65536.0,1,-nbitq), 
to_sfixed(-1908.0/65536.0,1,-nbitq), 
to_sfixed(109.0/65536.0,1,-nbitq), 
to_sfixed(1645.0/65536.0,1,-nbitq), 
to_sfixed(566.0/65536.0,1,-nbitq), 
to_sfixed(-1561.0/65536.0,1,-nbitq), 
to_sfixed(-8127.0/65536.0,1,-nbitq), 
to_sfixed(-2295.0/65536.0,1,-nbitq), 
to_sfixed(-2685.0/65536.0,1,-nbitq), 
to_sfixed(-1009.0/65536.0,1,-nbitq), 
to_sfixed(426.0/65536.0,1,-nbitq), 
to_sfixed(1750.0/65536.0,1,-nbitq), 
to_sfixed(-1133.0/65536.0,1,-nbitq), 
to_sfixed(-1785.0/65536.0,1,-nbitq), 
to_sfixed(321.0/65536.0,1,-nbitq), 
to_sfixed(-1022.0/65536.0,1,-nbitq), 
to_sfixed(-1866.0/65536.0,1,-nbitq), 
to_sfixed(-1843.0/65536.0,1,-nbitq), 
to_sfixed(1410.0/65536.0,1,-nbitq), 
to_sfixed(2659.0/65536.0,1,-nbitq), 
to_sfixed(-879.0/65536.0,1,-nbitq), 
to_sfixed(-9809.0/65536.0,1,-nbitq), 
to_sfixed(-2792.0/65536.0,1,-nbitq), 
to_sfixed(597.0/65536.0,1,-nbitq), 
to_sfixed(-5098.0/65536.0,1,-nbitq), 
to_sfixed(-3341.0/65536.0,1,-nbitq), 
to_sfixed(2557.0/65536.0,1,-nbitq), 
to_sfixed(1530.0/65536.0,1,-nbitq), 
to_sfixed(-4524.0/65536.0,1,-nbitq), 
to_sfixed(8961.0/65536.0,1,-nbitq), 
to_sfixed(285.0/65536.0,1,-nbitq), 
to_sfixed(814.0/65536.0,1,-nbitq), 
to_sfixed(-2632.0/65536.0,1,-nbitq)  ), 
( to_sfixed(997.0/65536.0,1,-nbitq), 
to_sfixed(-374.0/65536.0,1,-nbitq), 
to_sfixed(-7044.0/65536.0,1,-nbitq), 
to_sfixed(-6420.0/65536.0,1,-nbitq), 
to_sfixed(3496.0/65536.0,1,-nbitq), 
to_sfixed(-4829.0/65536.0,1,-nbitq), 
to_sfixed(-8707.0/65536.0,1,-nbitq), 
to_sfixed(1583.0/65536.0,1,-nbitq), 
to_sfixed(1279.0/65536.0,1,-nbitq), 
to_sfixed(2089.0/65536.0,1,-nbitq), 
to_sfixed(579.0/65536.0,1,-nbitq), 
to_sfixed(-5969.0/65536.0,1,-nbitq), 
to_sfixed(2791.0/65536.0,1,-nbitq), 
to_sfixed(8112.0/65536.0,1,-nbitq), 
to_sfixed(-4131.0/65536.0,1,-nbitq), 
to_sfixed(1500.0/65536.0,1,-nbitq), 
to_sfixed(2738.0/65536.0,1,-nbitq), 
to_sfixed(-6559.0/65536.0,1,-nbitq), 
to_sfixed(3044.0/65536.0,1,-nbitq), 
to_sfixed(-681.0/65536.0,1,-nbitq), 
to_sfixed(-3510.0/65536.0,1,-nbitq), 
to_sfixed(688.0/65536.0,1,-nbitq), 
to_sfixed(-1329.0/65536.0,1,-nbitq), 
to_sfixed(2912.0/65536.0,1,-nbitq), 
to_sfixed(-2932.0/65536.0,1,-nbitq), 
to_sfixed(-6856.0/65536.0,1,-nbitq), 
to_sfixed(683.0/65536.0,1,-nbitq), 
to_sfixed(-4023.0/65536.0,1,-nbitq), 
to_sfixed(-8661.0/65536.0,1,-nbitq), 
to_sfixed(10133.0/65536.0,1,-nbitq), 
to_sfixed(5492.0/65536.0,1,-nbitq), 
to_sfixed(2286.0/65536.0,1,-nbitq), 
to_sfixed(-3944.0/65536.0,1,-nbitq), 
to_sfixed(-4241.0/65536.0,1,-nbitq), 
to_sfixed(3106.0/65536.0,1,-nbitq), 
to_sfixed(-2069.0/65536.0,1,-nbitq), 
to_sfixed(9611.0/65536.0,1,-nbitq), 
to_sfixed(-1373.0/65536.0,1,-nbitq), 
to_sfixed(1673.0/65536.0,1,-nbitq), 
to_sfixed(649.0/65536.0,1,-nbitq), 
to_sfixed(-8509.0/65536.0,1,-nbitq), 
to_sfixed(-1232.0/65536.0,1,-nbitq), 
to_sfixed(-11578.0/65536.0,1,-nbitq), 
to_sfixed(7048.0/65536.0,1,-nbitq), 
to_sfixed(2298.0/65536.0,1,-nbitq), 
to_sfixed(-3911.0/65536.0,1,-nbitq), 
to_sfixed(2089.0/65536.0,1,-nbitq), 
to_sfixed(7182.0/65536.0,1,-nbitq), 
to_sfixed(2495.0/65536.0,1,-nbitq), 
to_sfixed(1448.0/65536.0,1,-nbitq), 
to_sfixed(1756.0/65536.0,1,-nbitq), 
to_sfixed(826.0/65536.0,1,-nbitq), 
to_sfixed(-3029.0/65536.0,1,-nbitq), 
to_sfixed(-7019.0/65536.0,1,-nbitq), 
to_sfixed(81.0/65536.0,1,-nbitq), 
to_sfixed(-3357.0/65536.0,1,-nbitq), 
to_sfixed(1299.0/65536.0,1,-nbitq), 
to_sfixed(36.0/65536.0,1,-nbitq), 
to_sfixed(2032.0/65536.0,1,-nbitq), 
to_sfixed(-2405.0/65536.0,1,-nbitq), 
to_sfixed(-2806.0/65536.0,1,-nbitq), 
to_sfixed(623.0/65536.0,1,-nbitq), 
to_sfixed(-2157.0/65536.0,1,-nbitq), 
to_sfixed(1458.0/65536.0,1,-nbitq), 
to_sfixed(1381.0/65536.0,1,-nbitq), 
to_sfixed(-1581.0/65536.0,1,-nbitq), 
to_sfixed(651.0/65536.0,1,-nbitq), 
to_sfixed(2081.0/65536.0,1,-nbitq), 
to_sfixed(-10170.0/65536.0,1,-nbitq), 
to_sfixed(-1470.0/65536.0,1,-nbitq), 
to_sfixed(69.0/65536.0,1,-nbitq), 
to_sfixed(-4524.0/65536.0,1,-nbitq), 
to_sfixed(-2521.0/65536.0,1,-nbitq), 
to_sfixed(1472.0/65536.0,1,-nbitq), 
to_sfixed(-2404.0/65536.0,1,-nbitq), 
to_sfixed(-4804.0/65536.0,1,-nbitq), 
to_sfixed(9194.0/65536.0,1,-nbitq), 
to_sfixed(-1171.0/65536.0,1,-nbitq), 
to_sfixed(-1310.0/65536.0,1,-nbitq), 
to_sfixed(-4847.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1379.0/65536.0,1,-nbitq), 
to_sfixed(-4148.0/65536.0,1,-nbitq), 
to_sfixed(-10887.0/65536.0,1,-nbitq), 
to_sfixed(-2985.0/65536.0,1,-nbitq), 
to_sfixed(-601.0/65536.0,1,-nbitq), 
to_sfixed(3719.0/65536.0,1,-nbitq), 
to_sfixed(-5743.0/65536.0,1,-nbitq), 
to_sfixed(5374.0/65536.0,1,-nbitq), 
to_sfixed(-4488.0/65536.0,1,-nbitq), 
to_sfixed(2487.0/65536.0,1,-nbitq), 
to_sfixed(-2705.0/65536.0,1,-nbitq), 
to_sfixed(2258.0/65536.0,1,-nbitq), 
to_sfixed(1395.0/65536.0,1,-nbitq), 
to_sfixed(7609.0/65536.0,1,-nbitq), 
to_sfixed(-2521.0/65536.0,1,-nbitq), 
to_sfixed(458.0/65536.0,1,-nbitq), 
to_sfixed(3010.0/65536.0,1,-nbitq), 
to_sfixed(-10092.0/65536.0,1,-nbitq), 
to_sfixed(-549.0/65536.0,1,-nbitq), 
to_sfixed(-2484.0/65536.0,1,-nbitq), 
to_sfixed(-5517.0/65536.0,1,-nbitq), 
to_sfixed(161.0/65536.0,1,-nbitq), 
to_sfixed(-4837.0/65536.0,1,-nbitq), 
to_sfixed(-2282.0/65536.0,1,-nbitq), 
to_sfixed(-1446.0/65536.0,1,-nbitq), 
to_sfixed(-2280.0/65536.0,1,-nbitq), 
to_sfixed(8402.0/65536.0,1,-nbitq), 
to_sfixed(-4799.0/65536.0,1,-nbitq), 
to_sfixed(92.0/65536.0,1,-nbitq), 
to_sfixed(4875.0/65536.0,1,-nbitq), 
to_sfixed(1747.0/65536.0,1,-nbitq), 
to_sfixed(5280.0/65536.0,1,-nbitq), 
to_sfixed(-4082.0/65536.0,1,-nbitq), 
to_sfixed(-4800.0/65536.0,1,-nbitq), 
to_sfixed(-1591.0/65536.0,1,-nbitq), 
to_sfixed(-2361.0/65536.0,1,-nbitq), 
to_sfixed(-3000.0/65536.0,1,-nbitq), 
to_sfixed(-1784.0/65536.0,1,-nbitq), 
to_sfixed(4257.0/65536.0,1,-nbitq), 
to_sfixed(339.0/65536.0,1,-nbitq), 
to_sfixed(-8284.0/65536.0,1,-nbitq), 
to_sfixed(2527.0/65536.0,1,-nbitq), 
to_sfixed(-3419.0/65536.0,1,-nbitq), 
to_sfixed(1538.0/65536.0,1,-nbitq), 
to_sfixed(559.0/65536.0,1,-nbitq), 
to_sfixed(-2059.0/65536.0,1,-nbitq), 
to_sfixed(-697.0/65536.0,1,-nbitq), 
to_sfixed(7668.0/65536.0,1,-nbitq), 
to_sfixed(359.0/65536.0,1,-nbitq), 
to_sfixed(1103.0/65536.0,1,-nbitq), 
to_sfixed(-1152.0/65536.0,1,-nbitq), 
to_sfixed(2085.0/65536.0,1,-nbitq), 
to_sfixed(-283.0/65536.0,1,-nbitq), 
to_sfixed(-6855.0/65536.0,1,-nbitq), 
to_sfixed(-1542.0/65536.0,1,-nbitq), 
to_sfixed(-4044.0/65536.0,1,-nbitq), 
to_sfixed(-459.0/65536.0,1,-nbitq), 
to_sfixed(1855.0/65536.0,1,-nbitq), 
to_sfixed(2337.0/65536.0,1,-nbitq), 
to_sfixed(-1772.0/65536.0,1,-nbitq), 
to_sfixed(1230.0/65536.0,1,-nbitq), 
to_sfixed(-2492.0/65536.0,1,-nbitq), 
to_sfixed(708.0/65536.0,1,-nbitq), 
to_sfixed(2116.0/65536.0,1,-nbitq), 
to_sfixed(1039.0/65536.0,1,-nbitq), 
to_sfixed(5808.0/65536.0,1,-nbitq), 
to_sfixed(-2837.0/65536.0,1,-nbitq), 
to_sfixed(10163.0/65536.0,1,-nbitq), 
to_sfixed(-8593.0/65536.0,1,-nbitq), 
to_sfixed(449.0/65536.0,1,-nbitq), 
to_sfixed(-1973.0/65536.0,1,-nbitq), 
to_sfixed(1526.0/65536.0,1,-nbitq), 
to_sfixed(-3923.0/65536.0,1,-nbitq), 
to_sfixed(1223.0/65536.0,1,-nbitq), 
to_sfixed(708.0/65536.0,1,-nbitq), 
to_sfixed(-3067.0/65536.0,1,-nbitq), 
to_sfixed(6379.0/65536.0,1,-nbitq), 
to_sfixed(-2753.0/65536.0,1,-nbitq), 
to_sfixed(1051.0/65536.0,1,-nbitq), 
to_sfixed(-2968.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1394.0/65536.0,1,-nbitq), 
to_sfixed(-4424.0/65536.0,1,-nbitq), 
to_sfixed(-3025.0/65536.0,1,-nbitq), 
to_sfixed(705.0/65536.0,1,-nbitq), 
to_sfixed(-5627.0/65536.0,1,-nbitq), 
to_sfixed(-3000.0/65536.0,1,-nbitq), 
to_sfixed(-951.0/65536.0,1,-nbitq), 
to_sfixed(4058.0/65536.0,1,-nbitq), 
to_sfixed(-7.0/65536.0,1,-nbitq), 
to_sfixed(2565.0/65536.0,1,-nbitq), 
to_sfixed(-2354.0/65536.0,1,-nbitq), 
to_sfixed(-1324.0/65536.0,1,-nbitq), 
to_sfixed(3322.0/65536.0,1,-nbitq), 
to_sfixed(5708.0/65536.0,1,-nbitq), 
to_sfixed(827.0/65536.0,1,-nbitq), 
to_sfixed(1056.0/65536.0,1,-nbitq), 
to_sfixed(1867.0/65536.0,1,-nbitq), 
to_sfixed(-10283.0/65536.0,1,-nbitq), 
to_sfixed(2765.0/65536.0,1,-nbitq), 
to_sfixed(-2126.0/65536.0,1,-nbitq), 
to_sfixed(-7334.0/65536.0,1,-nbitq), 
to_sfixed(5608.0/65536.0,1,-nbitq), 
to_sfixed(3214.0/65536.0,1,-nbitq), 
to_sfixed(-1684.0/65536.0,1,-nbitq), 
to_sfixed(-3098.0/65536.0,1,-nbitq), 
to_sfixed(-1357.0/65536.0,1,-nbitq), 
to_sfixed(4354.0/65536.0,1,-nbitq), 
to_sfixed(-2646.0/65536.0,1,-nbitq), 
to_sfixed(-5481.0/65536.0,1,-nbitq), 
to_sfixed(4533.0/65536.0,1,-nbitq), 
to_sfixed(1689.0/65536.0,1,-nbitq), 
to_sfixed(3990.0/65536.0,1,-nbitq), 
to_sfixed(-6553.0/65536.0,1,-nbitq), 
to_sfixed(5885.0/65536.0,1,-nbitq), 
to_sfixed(-388.0/65536.0,1,-nbitq), 
to_sfixed(3108.0/65536.0,1,-nbitq), 
to_sfixed(-3069.0/65536.0,1,-nbitq), 
to_sfixed(1246.0/65536.0,1,-nbitq), 
to_sfixed(5278.0/65536.0,1,-nbitq), 
to_sfixed(2910.0/65536.0,1,-nbitq), 
to_sfixed(-1615.0/65536.0,1,-nbitq), 
to_sfixed(-2348.0/65536.0,1,-nbitq), 
to_sfixed(-1400.0/65536.0,1,-nbitq), 
to_sfixed(5848.0/65536.0,1,-nbitq), 
to_sfixed(410.0/65536.0,1,-nbitq), 
to_sfixed(5252.0/65536.0,1,-nbitq), 
to_sfixed(-112.0/65536.0,1,-nbitq), 
to_sfixed(3769.0/65536.0,1,-nbitq), 
to_sfixed(-681.0/65536.0,1,-nbitq), 
to_sfixed(419.0/65536.0,1,-nbitq), 
to_sfixed(558.0/65536.0,1,-nbitq), 
to_sfixed(1948.0/65536.0,1,-nbitq), 
to_sfixed(1791.0/65536.0,1,-nbitq), 
to_sfixed(-383.0/65536.0,1,-nbitq), 
to_sfixed(-102.0/65536.0,1,-nbitq), 
to_sfixed(-4313.0/65536.0,1,-nbitq), 
to_sfixed(-1303.0/65536.0,1,-nbitq), 
to_sfixed(-4718.0/65536.0,1,-nbitq), 
to_sfixed(-867.0/65536.0,1,-nbitq), 
to_sfixed(-4821.0/65536.0,1,-nbitq), 
to_sfixed(3828.0/65536.0,1,-nbitq), 
to_sfixed(558.0/65536.0,1,-nbitq), 
to_sfixed(-1383.0/65536.0,1,-nbitq), 
to_sfixed(-2686.0/65536.0,1,-nbitq), 
to_sfixed(2349.0/65536.0,1,-nbitq), 
to_sfixed(6818.0/65536.0,1,-nbitq), 
to_sfixed(-3654.0/65536.0,1,-nbitq), 
to_sfixed(703.0/65536.0,1,-nbitq), 
to_sfixed(-11845.0/65536.0,1,-nbitq), 
to_sfixed(1882.0/65536.0,1,-nbitq), 
to_sfixed(-1699.0/65536.0,1,-nbitq), 
to_sfixed(4330.0/65536.0,1,-nbitq), 
to_sfixed(627.0/65536.0,1,-nbitq), 
to_sfixed(-747.0/65536.0,1,-nbitq), 
to_sfixed(109.0/65536.0,1,-nbitq), 
to_sfixed(-3144.0/65536.0,1,-nbitq), 
to_sfixed(5168.0/65536.0,1,-nbitq), 
to_sfixed(-4189.0/65536.0,1,-nbitq), 
to_sfixed(148.0/65536.0,1,-nbitq), 
to_sfixed(963.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-37.0/65536.0,1,-nbitq), 
to_sfixed(-6958.0/65536.0,1,-nbitq), 
to_sfixed(3373.0/65536.0,1,-nbitq), 
to_sfixed(-2335.0/65536.0,1,-nbitq), 
to_sfixed(-6331.0/65536.0,1,-nbitq), 
to_sfixed(-2468.0/65536.0,1,-nbitq), 
to_sfixed(4355.0/65536.0,1,-nbitq), 
to_sfixed(4018.0/65536.0,1,-nbitq), 
to_sfixed(58.0/65536.0,1,-nbitq), 
to_sfixed(-2701.0/65536.0,1,-nbitq), 
to_sfixed(-1757.0/65536.0,1,-nbitq), 
to_sfixed(670.0/65536.0,1,-nbitq), 
to_sfixed(-1214.0/65536.0,1,-nbitq), 
to_sfixed(675.0/65536.0,1,-nbitq), 
to_sfixed(-2367.0/65536.0,1,-nbitq), 
to_sfixed(-471.0/65536.0,1,-nbitq), 
to_sfixed(1256.0/65536.0,1,-nbitq), 
to_sfixed(-10180.0/65536.0,1,-nbitq), 
to_sfixed(643.0/65536.0,1,-nbitq), 
to_sfixed(818.0/65536.0,1,-nbitq), 
to_sfixed(287.0/65536.0,1,-nbitq), 
to_sfixed(9203.0/65536.0,1,-nbitq), 
to_sfixed(2367.0/65536.0,1,-nbitq), 
to_sfixed(1604.0/65536.0,1,-nbitq), 
to_sfixed(-3287.0/65536.0,1,-nbitq), 
to_sfixed(-1753.0/65536.0,1,-nbitq), 
to_sfixed(6591.0/65536.0,1,-nbitq), 
to_sfixed(-1905.0/65536.0,1,-nbitq), 
to_sfixed(-6106.0/65536.0,1,-nbitq), 
to_sfixed(2954.0/65536.0,1,-nbitq), 
to_sfixed(1622.0/65536.0,1,-nbitq), 
to_sfixed(2280.0/65536.0,1,-nbitq), 
to_sfixed(-2197.0/65536.0,1,-nbitq), 
to_sfixed(8433.0/65536.0,1,-nbitq), 
to_sfixed(857.0/65536.0,1,-nbitq), 
to_sfixed(-879.0/65536.0,1,-nbitq), 
to_sfixed(-3765.0/65536.0,1,-nbitq), 
to_sfixed(1988.0/65536.0,1,-nbitq), 
to_sfixed(3647.0/65536.0,1,-nbitq), 
to_sfixed(-779.0/65536.0,1,-nbitq), 
to_sfixed(3787.0/65536.0,1,-nbitq), 
to_sfixed(-1760.0/65536.0,1,-nbitq), 
to_sfixed(2081.0/65536.0,1,-nbitq), 
to_sfixed(7908.0/65536.0,1,-nbitq), 
to_sfixed(-551.0/65536.0,1,-nbitq), 
to_sfixed(2617.0/65536.0,1,-nbitq), 
to_sfixed(-1072.0/65536.0,1,-nbitq), 
to_sfixed(6975.0/65536.0,1,-nbitq), 
to_sfixed(2864.0/65536.0,1,-nbitq), 
to_sfixed(2187.0/65536.0,1,-nbitq), 
to_sfixed(-1028.0/65536.0,1,-nbitq), 
to_sfixed(225.0/65536.0,1,-nbitq), 
to_sfixed(1556.0/65536.0,1,-nbitq), 
to_sfixed(261.0/65536.0,1,-nbitq), 
to_sfixed(258.0/65536.0,1,-nbitq), 
to_sfixed(-4793.0/65536.0,1,-nbitq), 
to_sfixed(135.0/65536.0,1,-nbitq), 
to_sfixed(-5209.0/65536.0,1,-nbitq), 
to_sfixed(2330.0/65536.0,1,-nbitq), 
to_sfixed(-7246.0/65536.0,1,-nbitq), 
to_sfixed(-1187.0/65536.0,1,-nbitq), 
to_sfixed(-2685.0/65536.0,1,-nbitq), 
to_sfixed(-842.0/65536.0,1,-nbitq), 
to_sfixed(75.0/65536.0,1,-nbitq), 
to_sfixed(3135.0/65536.0,1,-nbitq), 
to_sfixed(6416.0/65536.0,1,-nbitq), 
to_sfixed(-4226.0/65536.0,1,-nbitq), 
to_sfixed(1441.0/65536.0,1,-nbitq), 
to_sfixed(-8977.0/65536.0,1,-nbitq), 
to_sfixed(-888.0/65536.0,1,-nbitq), 
to_sfixed(-3626.0/65536.0,1,-nbitq), 
to_sfixed(2618.0/65536.0,1,-nbitq), 
to_sfixed(-491.0/65536.0,1,-nbitq), 
to_sfixed(-1470.0/65536.0,1,-nbitq), 
to_sfixed(-524.0/65536.0,1,-nbitq), 
to_sfixed(-203.0/65536.0,1,-nbitq), 
to_sfixed(7820.0/65536.0,1,-nbitq), 
to_sfixed(-404.0/65536.0,1,-nbitq), 
to_sfixed(-2570.0/65536.0,1,-nbitq), 
to_sfixed(1633.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2271.0/65536.0,1,-nbitq), 
to_sfixed(-4132.0/65536.0,1,-nbitq), 
to_sfixed(421.0/65536.0,1,-nbitq), 
to_sfixed(1968.0/65536.0,1,-nbitq), 
to_sfixed(-4679.0/65536.0,1,-nbitq), 
to_sfixed(-4094.0/65536.0,1,-nbitq), 
to_sfixed(455.0/65536.0,1,-nbitq), 
to_sfixed(-1.0/65536.0,1,-nbitq), 
to_sfixed(2319.0/65536.0,1,-nbitq), 
to_sfixed(-2179.0/65536.0,1,-nbitq), 
to_sfixed(-1537.0/65536.0,1,-nbitq), 
to_sfixed(2271.0/65536.0,1,-nbitq), 
to_sfixed(4299.0/65536.0,1,-nbitq), 
to_sfixed(445.0/65536.0,1,-nbitq), 
to_sfixed(-1481.0/65536.0,1,-nbitq), 
to_sfixed(2750.0/65536.0,1,-nbitq), 
to_sfixed(-441.0/65536.0,1,-nbitq), 
to_sfixed(-7957.0/65536.0,1,-nbitq), 
to_sfixed(-2548.0/65536.0,1,-nbitq), 
to_sfixed(1045.0/65536.0,1,-nbitq), 
to_sfixed(3117.0/65536.0,1,-nbitq), 
to_sfixed(11499.0/65536.0,1,-nbitq), 
to_sfixed(-616.0/65536.0,1,-nbitq), 
to_sfixed(9001.0/65536.0,1,-nbitq), 
to_sfixed(-2547.0/65536.0,1,-nbitq), 
to_sfixed(648.0/65536.0,1,-nbitq), 
to_sfixed(6936.0/65536.0,1,-nbitq), 
to_sfixed(-5652.0/65536.0,1,-nbitq), 
to_sfixed(-2150.0/65536.0,1,-nbitq), 
to_sfixed(387.0/65536.0,1,-nbitq), 
to_sfixed(-7017.0/65536.0,1,-nbitq), 
to_sfixed(442.0/65536.0,1,-nbitq), 
to_sfixed(-3474.0/65536.0,1,-nbitq), 
to_sfixed(4397.0/65536.0,1,-nbitq), 
to_sfixed(2270.0/65536.0,1,-nbitq), 
to_sfixed(1746.0/65536.0,1,-nbitq), 
to_sfixed(-1631.0/65536.0,1,-nbitq), 
to_sfixed(-1411.0/65536.0,1,-nbitq), 
to_sfixed(6466.0/65536.0,1,-nbitq), 
to_sfixed(2640.0/65536.0,1,-nbitq), 
to_sfixed(9031.0/65536.0,1,-nbitq), 
to_sfixed(1906.0/65536.0,1,-nbitq), 
to_sfixed(-2214.0/65536.0,1,-nbitq), 
to_sfixed(9866.0/65536.0,1,-nbitq), 
to_sfixed(-666.0/65536.0,1,-nbitq), 
to_sfixed(2023.0/65536.0,1,-nbitq), 
to_sfixed(-704.0/65536.0,1,-nbitq), 
to_sfixed(3272.0/65536.0,1,-nbitq), 
to_sfixed(3384.0/65536.0,1,-nbitq), 
to_sfixed(1275.0/65536.0,1,-nbitq), 
to_sfixed(1442.0/65536.0,1,-nbitq), 
to_sfixed(5115.0/65536.0,1,-nbitq), 
to_sfixed(-1731.0/65536.0,1,-nbitq), 
to_sfixed(-7250.0/65536.0,1,-nbitq), 
to_sfixed(-139.0/65536.0,1,-nbitq), 
to_sfixed(2869.0/65536.0,1,-nbitq), 
to_sfixed(2614.0/65536.0,1,-nbitq), 
to_sfixed(-99.0/65536.0,1,-nbitq), 
to_sfixed(-1930.0/65536.0,1,-nbitq), 
to_sfixed(-1500.0/65536.0,1,-nbitq), 
to_sfixed(-4904.0/65536.0,1,-nbitq), 
to_sfixed(1252.0/65536.0,1,-nbitq), 
to_sfixed(2971.0/65536.0,1,-nbitq), 
to_sfixed(1112.0/65536.0,1,-nbitq), 
to_sfixed(5864.0/65536.0,1,-nbitq), 
to_sfixed(5689.0/65536.0,1,-nbitq), 
to_sfixed(-1936.0/65536.0,1,-nbitq), 
to_sfixed(2313.0/65536.0,1,-nbitq), 
to_sfixed(-9244.0/65536.0,1,-nbitq), 
to_sfixed(-994.0/65536.0,1,-nbitq), 
to_sfixed(1344.0/65536.0,1,-nbitq), 
to_sfixed(-3486.0/65536.0,1,-nbitq), 
to_sfixed(-2690.0/65536.0,1,-nbitq), 
to_sfixed(751.0/65536.0,1,-nbitq), 
to_sfixed(477.0/65536.0,1,-nbitq), 
to_sfixed(1430.0/65536.0,1,-nbitq), 
to_sfixed(6477.0/65536.0,1,-nbitq), 
to_sfixed(-3527.0/65536.0,1,-nbitq), 
to_sfixed(-1452.0/65536.0,1,-nbitq), 
to_sfixed(4989.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-588.0/65536.0,1,-nbitq), 
to_sfixed(-1509.0/65536.0,1,-nbitq), 
to_sfixed(2368.0/65536.0,1,-nbitq), 
to_sfixed(3914.0/65536.0,1,-nbitq), 
to_sfixed(-897.0/65536.0,1,-nbitq), 
to_sfixed(-1629.0/65536.0,1,-nbitq), 
to_sfixed(3562.0/65536.0,1,-nbitq), 
to_sfixed(-3698.0/65536.0,1,-nbitq), 
to_sfixed(2920.0/65536.0,1,-nbitq), 
to_sfixed(1877.0/65536.0,1,-nbitq), 
to_sfixed(-2835.0/65536.0,1,-nbitq), 
to_sfixed(-348.0/65536.0,1,-nbitq), 
to_sfixed(-676.0/65536.0,1,-nbitq), 
to_sfixed(-3037.0/65536.0,1,-nbitq), 
to_sfixed(-3928.0/65536.0,1,-nbitq), 
to_sfixed(-653.0/65536.0,1,-nbitq), 
to_sfixed(-648.0/65536.0,1,-nbitq), 
to_sfixed(-4634.0/65536.0,1,-nbitq), 
to_sfixed(-1548.0/65536.0,1,-nbitq), 
to_sfixed(1273.0/65536.0,1,-nbitq), 
to_sfixed(2617.0/65536.0,1,-nbitq), 
to_sfixed(3385.0/65536.0,1,-nbitq), 
to_sfixed(-1007.0/65536.0,1,-nbitq), 
to_sfixed(7642.0/65536.0,1,-nbitq), 
to_sfixed(1120.0/65536.0,1,-nbitq), 
to_sfixed(5311.0/65536.0,1,-nbitq), 
to_sfixed(6521.0/65536.0,1,-nbitq), 
to_sfixed(-4985.0/65536.0,1,-nbitq), 
to_sfixed(-5408.0/65536.0,1,-nbitq), 
to_sfixed(1625.0/65536.0,1,-nbitq), 
to_sfixed(-10054.0/65536.0,1,-nbitq), 
to_sfixed(3630.0/65536.0,1,-nbitq), 
to_sfixed(-1835.0/65536.0,1,-nbitq), 
to_sfixed(-431.0/65536.0,1,-nbitq), 
to_sfixed(-362.0/65536.0,1,-nbitq), 
to_sfixed(2531.0/65536.0,1,-nbitq), 
to_sfixed(-7691.0/65536.0,1,-nbitq), 
to_sfixed(-2712.0/65536.0,1,-nbitq), 
to_sfixed(4589.0/65536.0,1,-nbitq), 
to_sfixed(1886.0/65536.0,1,-nbitq), 
to_sfixed(13140.0/65536.0,1,-nbitq), 
to_sfixed(-1149.0/65536.0,1,-nbitq), 
to_sfixed(-2435.0/65536.0,1,-nbitq), 
to_sfixed(8173.0/65536.0,1,-nbitq), 
to_sfixed(1418.0/65536.0,1,-nbitq), 
to_sfixed(1099.0/65536.0,1,-nbitq), 
to_sfixed(-1951.0/65536.0,1,-nbitq), 
to_sfixed(1285.0/65536.0,1,-nbitq), 
to_sfixed(-2037.0/65536.0,1,-nbitq), 
to_sfixed(1836.0/65536.0,1,-nbitq), 
to_sfixed(2129.0/65536.0,1,-nbitq), 
to_sfixed(5033.0/65536.0,1,-nbitq), 
to_sfixed(-6872.0/65536.0,1,-nbitq), 
to_sfixed(-9691.0/65536.0,1,-nbitq), 
to_sfixed(-1274.0/65536.0,1,-nbitq), 
to_sfixed(2645.0/65536.0,1,-nbitq), 
to_sfixed(1580.0/65536.0,1,-nbitq), 
to_sfixed(-2233.0/65536.0,1,-nbitq), 
to_sfixed(-422.0/65536.0,1,-nbitq), 
to_sfixed(-753.0/65536.0,1,-nbitq), 
to_sfixed(-4057.0/65536.0,1,-nbitq), 
to_sfixed(-111.0/65536.0,1,-nbitq), 
to_sfixed(-1080.0/65536.0,1,-nbitq), 
to_sfixed(-1178.0/65536.0,1,-nbitq), 
to_sfixed(4758.0/65536.0,1,-nbitq), 
to_sfixed(1518.0/65536.0,1,-nbitq), 
to_sfixed(936.0/65536.0,1,-nbitq), 
to_sfixed(2598.0/65536.0,1,-nbitq), 
to_sfixed(-8226.0/65536.0,1,-nbitq), 
to_sfixed(-5045.0/65536.0,1,-nbitq), 
to_sfixed(283.0/65536.0,1,-nbitq), 
to_sfixed(-2701.0/65536.0,1,-nbitq), 
to_sfixed(1065.0/65536.0,1,-nbitq), 
to_sfixed(574.0/65536.0,1,-nbitq), 
to_sfixed(-944.0/65536.0,1,-nbitq), 
to_sfixed(3905.0/65536.0,1,-nbitq), 
to_sfixed(5561.0/65536.0,1,-nbitq), 
to_sfixed(-3252.0/65536.0,1,-nbitq), 
to_sfixed(1459.0/65536.0,1,-nbitq), 
to_sfixed(7768.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2192.0/65536.0,1,-nbitq), 
to_sfixed(-1444.0/65536.0,1,-nbitq), 
to_sfixed(4750.0/65536.0,1,-nbitq), 
to_sfixed(951.0/65536.0,1,-nbitq), 
to_sfixed(230.0/65536.0,1,-nbitq), 
to_sfixed(-193.0/65536.0,1,-nbitq), 
to_sfixed(-449.0/65536.0,1,-nbitq), 
to_sfixed(1234.0/65536.0,1,-nbitq), 
to_sfixed(1597.0/65536.0,1,-nbitq), 
to_sfixed(2143.0/65536.0,1,-nbitq), 
to_sfixed(483.0/65536.0,1,-nbitq), 
to_sfixed(3194.0/65536.0,1,-nbitq), 
to_sfixed(3565.0/65536.0,1,-nbitq), 
to_sfixed(1244.0/65536.0,1,-nbitq), 
to_sfixed(850.0/65536.0,1,-nbitq), 
to_sfixed(-103.0/65536.0,1,-nbitq), 
to_sfixed(2078.0/65536.0,1,-nbitq), 
to_sfixed(-228.0/65536.0,1,-nbitq), 
to_sfixed(-708.0/65536.0,1,-nbitq), 
to_sfixed(-2033.0/65536.0,1,-nbitq), 
to_sfixed(3460.0/65536.0,1,-nbitq), 
to_sfixed(2681.0/65536.0,1,-nbitq), 
to_sfixed(4408.0/65536.0,1,-nbitq), 
to_sfixed(2867.0/65536.0,1,-nbitq), 
to_sfixed(-1270.0/65536.0,1,-nbitq), 
to_sfixed(4454.0/65536.0,1,-nbitq), 
to_sfixed(3114.0/65536.0,1,-nbitq), 
to_sfixed(-1731.0/65536.0,1,-nbitq), 
to_sfixed(-8091.0/65536.0,1,-nbitq), 
to_sfixed(166.0/65536.0,1,-nbitq), 
to_sfixed(-6020.0/65536.0,1,-nbitq), 
to_sfixed(4085.0/65536.0,1,-nbitq), 
to_sfixed(3625.0/65536.0,1,-nbitq), 
to_sfixed(748.0/65536.0,1,-nbitq), 
to_sfixed(2013.0/65536.0,1,-nbitq), 
to_sfixed(-1619.0/65536.0,1,-nbitq), 
to_sfixed(-4010.0/65536.0,1,-nbitq), 
to_sfixed(805.0/65536.0,1,-nbitq), 
to_sfixed(-473.0/65536.0,1,-nbitq), 
to_sfixed(1380.0/65536.0,1,-nbitq), 
to_sfixed(11641.0/65536.0,1,-nbitq), 
to_sfixed(-1503.0/65536.0,1,-nbitq), 
to_sfixed(3327.0/65536.0,1,-nbitq), 
to_sfixed(10316.0/65536.0,1,-nbitq), 
to_sfixed(59.0/65536.0,1,-nbitq), 
to_sfixed(-1631.0/65536.0,1,-nbitq), 
to_sfixed(-5.0/65536.0,1,-nbitq), 
to_sfixed(-821.0/65536.0,1,-nbitq), 
to_sfixed(-1363.0/65536.0,1,-nbitq), 
to_sfixed(-1454.0/65536.0,1,-nbitq), 
to_sfixed(-1917.0/65536.0,1,-nbitq), 
to_sfixed(2695.0/65536.0,1,-nbitq), 
to_sfixed(235.0/65536.0,1,-nbitq), 
to_sfixed(-5042.0/65536.0,1,-nbitq), 
to_sfixed(-3200.0/65536.0,1,-nbitq), 
to_sfixed(4864.0/65536.0,1,-nbitq), 
to_sfixed(-114.0/65536.0,1,-nbitq), 
to_sfixed(1347.0/65536.0,1,-nbitq), 
to_sfixed(1953.0/65536.0,1,-nbitq), 
to_sfixed(1794.0/65536.0,1,-nbitq), 
to_sfixed(-3723.0/65536.0,1,-nbitq), 
to_sfixed(-2134.0/65536.0,1,-nbitq), 
to_sfixed(1267.0/65536.0,1,-nbitq), 
to_sfixed(-36.0/65536.0,1,-nbitq), 
to_sfixed(434.0/65536.0,1,-nbitq), 
to_sfixed(-2664.0/65536.0,1,-nbitq), 
to_sfixed(-653.0/65536.0,1,-nbitq), 
to_sfixed(4961.0/65536.0,1,-nbitq), 
to_sfixed(-278.0/65536.0,1,-nbitq), 
to_sfixed(-2312.0/65536.0,1,-nbitq), 
to_sfixed(485.0/65536.0,1,-nbitq), 
to_sfixed(-5182.0/65536.0,1,-nbitq), 
to_sfixed(1349.0/65536.0,1,-nbitq), 
to_sfixed(-521.0/65536.0,1,-nbitq), 
to_sfixed(-1914.0/65536.0,1,-nbitq), 
to_sfixed(-298.0/65536.0,1,-nbitq), 
to_sfixed(6333.0/65536.0,1,-nbitq), 
to_sfixed(-402.0/65536.0,1,-nbitq), 
to_sfixed(1907.0/65536.0,1,-nbitq), 
to_sfixed(4222.0/65536.0,1,-nbitq)  ), 
( to_sfixed(548.0/65536.0,1,-nbitq), 
to_sfixed(874.0/65536.0,1,-nbitq), 
to_sfixed(6875.0/65536.0,1,-nbitq), 
to_sfixed(1198.0/65536.0,1,-nbitq), 
to_sfixed(-6506.0/65536.0,1,-nbitq), 
to_sfixed(-6353.0/65536.0,1,-nbitq), 
to_sfixed(2981.0/65536.0,1,-nbitq), 
to_sfixed(3583.0/65536.0,1,-nbitq), 
to_sfixed(-1124.0/65536.0,1,-nbitq), 
to_sfixed(-1357.0/65536.0,1,-nbitq), 
to_sfixed(78.0/65536.0,1,-nbitq), 
to_sfixed(1211.0/65536.0,1,-nbitq), 
to_sfixed(709.0/65536.0,1,-nbitq), 
to_sfixed(2501.0/65536.0,1,-nbitq), 
to_sfixed(1842.0/65536.0,1,-nbitq), 
to_sfixed(-3012.0/65536.0,1,-nbitq), 
to_sfixed(-1939.0/65536.0,1,-nbitq), 
to_sfixed(-1730.0/65536.0,1,-nbitq), 
to_sfixed(-1489.0/65536.0,1,-nbitq), 
to_sfixed(2782.0/65536.0,1,-nbitq), 
to_sfixed(3757.0/65536.0,1,-nbitq), 
to_sfixed(-996.0/65536.0,1,-nbitq), 
to_sfixed(1505.0/65536.0,1,-nbitq), 
to_sfixed(803.0/65536.0,1,-nbitq), 
to_sfixed(1741.0/65536.0,1,-nbitq), 
to_sfixed(2224.0/65536.0,1,-nbitq), 
to_sfixed(-2993.0/65536.0,1,-nbitq), 
to_sfixed(-3527.0/65536.0,1,-nbitq), 
to_sfixed(-5661.0/65536.0,1,-nbitq), 
to_sfixed(554.0/65536.0,1,-nbitq), 
to_sfixed(-2599.0/65536.0,1,-nbitq), 
to_sfixed(3923.0/65536.0,1,-nbitq), 
to_sfixed(3683.0/65536.0,1,-nbitq), 
to_sfixed(-2279.0/65536.0,1,-nbitq), 
to_sfixed(4421.0/65536.0,1,-nbitq), 
to_sfixed(1166.0/65536.0,1,-nbitq), 
to_sfixed(-4947.0/65536.0,1,-nbitq), 
to_sfixed(474.0/65536.0,1,-nbitq), 
to_sfixed(1565.0/65536.0,1,-nbitq), 
to_sfixed(-83.0/65536.0,1,-nbitq), 
to_sfixed(8813.0/65536.0,1,-nbitq), 
to_sfixed(2129.0/65536.0,1,-nbitq), 
to_sfixed(6047.0/65536.0,1,-nbitq), 
to_sfixed(12.0/65536.0,1,-nbitq), 
to_sfixed(-564.0/65536.0,1,-nbitq), 
to_sfixed(3115.0/65536.0,1,-nbitq), 
to_sfixed(142.0/65536.0,1,-nbitq), 
to_sfixed(-3089.0/65536.0,1,-nbitq), 
to_sfixed(-837.0/65536.0,1,-nbitq), 
to_sfixed(2325.0/65536.0,1,-nbitq), 
to_sfixed(-1064.0/65536.0,1,-nbitq), 
to_sfixed(-2794.0/65536.0,1,-nbitq), 
to_sfixed(3014.0/65536.0,1,-nbitq), 
to_sfixed(-2136.0/65536.0,1,-nbitq), 
to_sfixed(-4517.0/65536.0,1,-nbitq), 
to_sfixed(6614.0/65536.0,1,-nbitq), 
to_sfixed(1301.0/65536.0,1,-nbitq), 
to_sfixed(468.0/65536.0,1,-nbitq), 
to_sfixed(-284.0/65536.0,1,-nbitq), 
to_sfixed(3517.0/65536.0,1,-nbitq), 
to_sfixed(270.0/65536.0,1,-nbitq), 
to_sfixed(1757.0/65536.0,1,-nbitq), 
to_sfixed(2049.0/65536.0,1,-nbitq), 
to_sfixed(-428.0/65536.0,1,-nbitq), 
to_sfixed(3576.0/65536.0,1,-nbitq), 
to_sfixed(-4082.0/65536.0,1,-nbitq), 
to_sfixed(-12.0/65536.0,1,-nbitq), 
to_sfixed(-602.0/65536.0,1,-nbitq), 
to_sfixed(-1401.0/65536.0,1,-nbitq), 
to_sfixed(-757.0/65536.0,1,-nbitq), 
to_sfixed(478.0/65536.0,1,-nbitq), 
to_sfixed(-4143.0/65536.0,1,-nbitq), 
to_sfixed(-1528.0/65536.0,1,-nbitq), 
to_sfixed(-331.0/65536.0,1,-nbitq), 
to_sfixed(1360.0/65536.0,1,-nbitq), 
to_sfixed(-672.0/65536.0,1,-nbitq), 
to_sfixed(4216.0/65536.0,1,-nbitq), 
to_sfixed(-1276.0/65536.0,1,-nbitq), 
to_sfixed(-841.0/65536.0,1,-nbitq), 
to_sfixed(2763.0/65536.0,1,-nbitq)  ), 
( to_sfixed(568.0/65536.0,1,-nbitq), 
to_sfixed(-985.0/65536.0,1,-nbitq), 
to_sfixed(5128.0/65536.0,1,-nbitq), 
to_sfixed(-1768.0/65536.0,1,-nbitq), 
to_sfixed(-2215.0/65536.0,1,-nbitq), 
to_sfixed(412.0/65536.0,1,-nbitq), 
to_sfixed(1937.0/65536.0,1,-nbitq), 
to_sfixed(2402.0/65536.0,1,-nbitq), 
to_sfixed(1392.0/65536.0,1,-nbitq), 
to_sfixed(-860.0/65536.0,1,-nbitq), 
to_sfixed(3455.0/65536.0,1,-nbitq), 
to_sfixed(2715.0/65536.0,1,-nbitq), 
to_sfixed(2335.0/65536.0,1,-nbitq), 
to_sfixed(784.0/65536.0,1,-nbitq), 
to_sfixed(-746.0/65536.0,1,-nbitq), 
to_sfixed(1973.0/65536.0,1,-nbitq), 
to_sfixed(2368.0/65536.0,1,-nbitq), 
to_sfixed(-2123.0/65536.0,1,-nbitq), 
to_sfixed(49.0/65536.0,1,-nbitq), 
to_sfixed(-1161.0/65536.0,1,-nbitq), 
to_sfixed(4671.0/65536.0,1,-nbitq), 
to_sfixed(-4628.0/65536.0,1,-nbitq), 
to_sfixed(225.0/65536.0,1,-nbitq), 
to_sfixed(1335.0/65536.0,1,-nbitq), 
to_sfixed(1898.0/65536.0,1,-nbitq), 
to_sfixed(-1504.0/65536.0,1,-nbitq), 
to_sfixed(-6476.0/65536.0,1,-nbitq), 
to_sfixed(-2641.0/65536.0,1,-nbitq), 
to_sfixed(2490.0/65536.0,1,-nbitq), 
to_sfixed(4735.0/65536.0,1,-nbitq), 
to_sfixed(-1211.0/65536.0,1,-nbitq), 
to_sfixed(5830.0/65536.0,1,-nbitq), 
to_sfixed(4928.0/65536.0,1,-nbitq), 
to_sfixed(780.0/65536.0,1,-nbitq), 
to_sfixed(2525.0/65536.0,1,-nbitq), 
to_sfixed(-560.0/65536.0,1,-nbitq), 
to_sfixed(-5414.0/65536.0,1,-nbitq), 
to_sfixed(-2962.0/65536.0,1,-nbitq), 
to_sfixed(1492.0/65536.0,1,-nbitq), 
to_sfixed(-680.0/65536.0,1,-nbitq), 
to_sfixed(4637.0/65536.0,1,-nbitq), 
to_sfixed(2712.0/65536.0,1,-nbitq), 
to_sfixed(2447.0/65536.0,1,-nbitq), 
to_sfixed(-1226.0/65536.0,1,-nbitq), 
to_sfixed(-2309.0/65536.0,1,-nbitq), 
to_sfixed(1438.0/65536.0,1,-nbitq), 
to_sfixed(67.0/65536.0,1,-nbitq), 
to_sfixed(41.0/65536.0,1,-nbitq), 
to_sfixed(2490.0/65536.0,1,-nbitq), 
to_sfixed(2048.0/65536.0,1,-nbitq), 
to_sfixed(1252.0/65536.0,1,-nbitq), 
to_sfixed(889.0/65536.0,1,-nbitq), 
to_sfixed(3230.0/65536.0,1,-nbitq), 
to_sfixed(5.0/65536.0,1,-nbitq), 
to_sfixed(-3168.0/65536.0,1,-nbitq), 
to_sfixed(2390.0/65536.0,1,-nbitq), 
to_sfixed(-1828.0/65536.0,1,-nbitq), 
to_sfixed(-653.0/65536.0,1,-nbitq), 
to_sfixed(2476.0/65536.0,1,-nbitq), 
to_sfixed(-2086.0/65536.0,1,-nbitq), 
to_sfixed(5522.0/65536.0,1,-nbitq), 
to_sfixed(1002.0/65536.0,1,-nbitq), 
to_sfixed(-2818.0/65536.0,1,-nbitq), 
to_sfixed(-3356.0/65536.0,1,-nbitq), 
to_sfixed(1162.0/65536.0,1,-nbitq), 
to_sfixed(-4321.0/65536.0,1,-nbitq), 
to_sfixed(-620.0/65536.0,1,-nbitq), 
to_sfixed(1467.0/65536.0,1,-nbitq), 
to_sfixed(1509.0/65536.0,1,-nbitq), 
to_sfixed(1070.0/65536.0,1,-nbitq), 
to_sfixed(4463.0/65536.0,1,-nbitq), 
to_sfixed(3530.0/65536.0,1,-nbitq), 
to_sfixed(-4110.0/65536.0,1,-nbitq), 
to_sfixed(2413.0/65536.0,1,-nbitq), 
to_sfixed(631.0/65536.0,1,-nbitq), 
to_sfixed(4228.0/65536.0,1,-nbitq), 
to_sfixed(2394.0/65536.0,1,-nbitq), 
to_sfixed(-1901.0/65536.0,1,-nbitq), 
to_sfixed(2359.0/65536.0,1,-nbitq), 
to_sfixed(1576.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-810.0/65536.0,1,-nbitq), 
to_sfixed(-127.0/65536.0,1,-nbitq), 
to_sfixed(1762.0/65536.0,1,-nbitq), 
to_sfixed(-515.0/65536.0,1,-nbitq), 
to_sfixed(-944.0/65536.0,1,-nbitq), 
to_sfixed(-6316.0/65536.0,1,-nbitq), 
to_sfixed(3653.0/65536.0,1,-nbitq), 
to_sfixed(2388.0/65536.0,1,-nbitq), 
to_sfixed(2115.0/65536.0,1,-nbitq), 
to_sfixed(-434.0/65536.0,1,-nbitq), 
to_sfixed(3049.0/65536.0,1,-nbitq), 
to_sfixed(4784.0/65536.0,1,-nbitq), 
to_sfixed(-89.0/65536.0,1,-nbitq), 
to_sfixed(1380.0/65536.0,1,-nbitq), 
to_sfixed(-1974.0/65536.0,1,-nbitq), 
to_sfixed(-1972.0/65536.0,1,-nbitq), 
to_sfixed(-153.0/65536.0,1,-nbitq), 
to_sfixed(-886.0/65536.0,1,-nbitq), 
to_sfixed(-2779.0/65536.0,1,-nbitq), 
to_sfixed(1057.0/65536.0,1,-nbitq), 
to_sfixed(3131.0/65536.0,1,-nbitq), 
to_sfixed(-2433.0/65536.0,1,-nbitq), 
to_sfixed(-353.0/65536.0,1,-nbitq), 
to_sfixed(-767.0/65536.0,1,-nbitq), 
to_sfixed(-1746.0/65536.0,1,-nbitq), 
to_sfixed(844.0/65536.0,1,-nbitq), 
to_sfixed(-5890.0/65536.0,1,-nbitq), 
to_sfixed(42.0/65536.0,1,-nbitq), 
to_sfixed(1258.0/65536.0,1,-nbitq), 
to_sfixed(22.0/65536.0,1,-nbitq), 
to_sfixed(-4825.0/65536.0,1,-nbitq), 
to_sfixed(795.0/65536.0,1,-nbitq), 
to_sfixed(2299.0/65536.0,1,-nbitq), 
to_sfixed(170.0/65536.0,1,-nbitq), 
to_sfixed(-281.0/65536.0,1,-nbitq), 
to_sfixed(-599.0/65536.0,1,-nbitq), 
to_sfixed(-194.0/65536.0,1,-nbitq), 
to_sfixed(2751.0/65536.0,1,-nbitq), 
to_sfixed(1212.0/65536.0,1,-nbitq), 
to_sfixed(1767.0/65536.0,1,-nbitq), 
to_sfixed(201.0/65536.0,1,-nbitq), 
to_sfixed(2713.0/65536.0,1,-nbitq), 
to_sfixed(33.0/65536.0,1,-nbitq), 
to_sfixed(2695.0/65536.0,1,-nbitq), 
to_sfixed(-976.0/65536.0,1,-nbitq), 
to_sfixed(889.0/65536.0,1,-nbitq), 
to_sfixed(-2060.0/65536.0,1,-nbitq), 
to_sfixed(-1208.0/65536.0,1,-nbitq), 
to_sfixed(566.0/65536.0,1,-nbitq), 
to_sfixed(2901.0/65536.0,1,-nbitq), 
to_sfixed(3044.0/65536.0,1,-nbitq), 
to_sfixed(2081.0/65536.0,1,-nbitq), 
to_sfixed(2107.0/65536.0,1,-nbitq), 
to_sfixed(713.0/65536.0,1,-nbitq), 
to_sfixed(-8075.0/65536.0,1,-nbitq), 
to_sfixed(2561.0/65536.0,1,-nbitq), 
to_sfixed(1245.0/65536.0,1,-nbitq), 
to_sfixed(4868.0/65536.0,1,-nbitq), 
to_sfixed(972.0/65536.0,1,-nbitq), 
to_sfixed(1991.0/65536.0,1,-nbitq), 
to_sfixed(1263.0/65536.0,1,-nbitq), 
to_sfixed(876.0/65536.0,1,-nbitq), 
to_sfixed(-966.0/65536.0,1,-nbitq), 
to_sfixed(-3248.0/65536.0,1,-nbitq), 
to_sfixed(1887.0/65536.0,1,-nbitq), 
to_sfixed(-4089.0/65536.0,1,-nbitq), 
to_sfixed(-4618.0/65536.0,1,-nbitq), 
to_sfixed(416.0/65536.0,1,-nbitq), 
to_sfixed(5144.0/65536.0,1,-nbitq), 
to_sfixed(-39.0/65536.0,1,-nbitq), 
to_sfixed(-2466.0/65536.0,1,-nbitq), 
to_sfixed(-1277.0/65536.0,1,-nbitq), 
to_sfixed(-5983.0/65536.0,1,-nbitq), 
to_sfixed(-284.0/65536.0,1,-nbitq), 
to_sfixed(-755.0/65536.0,1,-nbitq), 
to_sfixed(720.0/65536.0,1,-nbitq), 
to_sfixed(-933.0/65536.0,1,-nbitq), 
to_sfixed(260.0/65536.0,1,-nbitq), 
to_sfixed(-1637.0/65536.0,1,-nbitq), 
to_sfixed(5154.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-572.0/65536.0,1,-nbitq), 
to_sfixed(-760.0/65536.0,1,-nbitq), 
to_sfixed(88.0/65536.0,1,-nbitq), 
to_sfixed(-2942.0/65536.0,1,-nbitq), 
to_sfixed(-3134.0/65536.0,1,-nbitq), 
to_sfixed(-5181.0/65536.0,1,-nbitq), 
to_sfixed(-85.0/65536.0,1,-nbitq), 
to_sfixed(2729.0/65536.0,1,-nbitq), 
to_sfixed(-917.0/65536.0,1,-nbitq), 
to_sfixed(-1766.0/65536.0,1,-nbitq), 
to_sfixed(2139.0/65536.0,1,-nbitq), 
to_sfixed(6297.0/65536.0,1,-nbitq), 
to_sfixed(-1910.0/65536.0,1,-nbitq), 
to_sfixed(-411.0/65536.0,1,-nbitq), 
to_sfixed(-3383.0/65536.0,1,-nbitq), 
to_sfixed(-425.0/65536.0,1,-nbitq), 
to_sfixed(-1070.0/65536.0,1,-nbitq), 
to_sfixed(415.0/65536.0,1,-nbitq), 
to_sfixed(-178.0/65536.0,1,-nbitq), 
to_sfixed(-1945.0/65536.0,1,-nbitq), 
to_sfixed(2217.0/65536.0,1,-nbitq), 
to_sfixed(-3216.0/65536.0,1,-nbitq), 
to_sfixed(-3694.0/65536.0,1,-nbitq), 
to_sfixed(-3884.0/65536.0,1,-nbitq), 
to_sfixed(-36.0/65536.0,1,-nbitq), 
to_sfixed(-2738.0/65536.0,1,-nbitq), 
to_sfixed(-4595.0/65536.0,1,-nbitq), 
to_sfixed(-3511.0/65536.0,1,-nbitq), 
to_sfixed(3527.0/65536.0,1,-nbitq), 
to_sfixed(1481.0/65536.0,1,-nbitq), 
to_sfixed(-4278.0/65536.0,1,-nbitq), 
to_sfixed(-721.0/65536.0,1,-nbitq), 
to_sfixed(-1595.0/65536.0,1,-nbitq), 
to_sfixed(1320.0/65536.0,1,-nbitq), 
to_sfixed(1006.0/65536.0,1,-nbitq), 
to_sfixed(3394.0/65536.0,1,-nbitq), 
to_sfixed(2697.0/65536.0,1,-nbitq), 
to_sfixed(4596.0/65536.0,1,-nbitq), 
to_sfixed(518.0/65536.0,1,-nbitq), 
to_sfixed(-2197.0/65536.0,1,-nbitq), 
to_sfixed(-2894.0/65536.0,1,-nbitq), 
to_sfixed(-1280.0/65536.0,1,-nbitq), 
to_sfixed(1510.0/65536.0,1,-nbitq), 
to_sfixed(668.0/65536.0,1,-nbitq), 
to_sfixed(-492.0/65536.0,1,-nbitq), 
to_sfixed(1579.0/65536.0,1,-nbitq), 
to_sfixed(1312.0/65536.0,1,-nbitq), 
to_sfixed(-3734.0/65536.0,1,-nbitq), 
to_sfixed(2046.0/65536.0,1,-nbitq), 
to_sfixed(-1358.0/65536.0,1,-nbitq), 
to_sfixed(-920.0/65536.0,1,-nbitq), 
to_sfixed(-1442.0/65536.0,1,-nbitq), 
to_sfixed(2424.0/65536.0,1,-nbitq), 
to_sfixed(1218.0/65536.0,1,-nbitq), 
to_sfixed(-4477.0/65536.0,1,-nbitq), 
to_sfixed(4097.0/65536.0,1,-nbitq), 
to_sfixed(-2182.0/65536.0,1,-nbitq), 
to_sfixed(3971.0/65536.0,1,-nbitq), 
to_sfixed(385.0/65536.0,1,-nbitq), 
to_sfixed(-4377.0/65536.0,1,-nbitq), 
to_sfixed(242.0/65536.0,1,-nbitq), 
to_sfixed(-1594.0/65536.0,1,-nbitq), 
to_sfixed(-2633.0/65536.0,1,-nbitq), 
to_sfixed(778.0/65536.0,1,-nbitq), 
to_sfixed(-2003.0/65536.0,1,-nbitq), 
to_sfixed(-1138.0/65536.0,1,-nbitq), 
to_sfixed(1120.0/65536.0,1,-nbitq), 
to_sfixed(-3106.0/65536.0,1,-nbitq), 
to_sfixed(8496.0/65536.0,1,-nbitq), 
to_sfixed(-3553.0/65536.0,1,-nbitq), 
to_sfixed(604.0/65536.0,1,-nbitq), 
to_sfixed(-1730.0/65536.0,1,-nbitq), 
to_sfixed(-3947.0/65536.0,1,-nbitq), 
to_sfixed(-1039.0/65536.0,1,-nbitq), 
to_sfixed(-947.0/65536.0,1,-nbitq), 
to_sfixed(-2865.0/65536.0,1,-nbitq), 
to_sfixed(-529.0/65536.0,1,-nbitq), 
to_sfixed(-187.0/65536.0,1,-nbitq), 
to_sfixed(1515.0/65536.0,1,-nbitq), 
to_sfixed(3193.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3071.0/65536.0,1,-nbitq), 
to_sfixed(-2133.0/65536.0,1,-nbitq), 
to_sfixed(-2442.0/65536.0,1,-nbitq), 
to_sfixed(723.0/65536.0,1,-nbitq), 
to_sfixed(-3420.0/65536.0,1,-nbitq), 
to_sfixed(-3429.0/65536.0,1,-nbitq), 
to_sfixed(-2941.0/65536.0,1,-nbitq), 
to_sfixed(-743.0/65536.0,1,-nbitq), 
to_sfixed(-689.0/65536.0,1,-nbitq), 
to_sfixed(1839.0/65536.0,1,-nbitq), 
to_sfixed(1248.0/65536.0,1,-nbitq), 
to_sfixed(4912.0/65536.0,1,-nbitq), 
to_sfixed(705.0/65536.0,1,-nbitq), 
to_sfixed(-4162.0/65536.0,1,-nbitq), 
to_sfixed(-4487.0/65536.0,1,-nbitq), 
to_sfixed(1711.0/65536.0,1,-nbitq), 
to_sfixed(1435.0/65536.0,1,-nbitq), 
to_sfixed(1577.0/65536.0,1,-nbitq), 
to_sfixed(2516.0/65536.0,1,-nbitq), 
to_sfixed(-1306.0/65536.0,1,-nbitq), 
to_sfixed(1714.0/65536.0,1,-nbitq), 
to_sfixed(2389.0/65536.0,1,-nbitq), 
to_sfixed(-2836.0/65536.0,1,-nbitq), 
to_sfixed(-4645.0/65536.0,1,-nbitq), 
to_sfixed(551.0/65536.0,1,-nbitq), 
to_sfixed(-1095.0/65536.0,1,-nbitq), 
to_sfixed(-2548.0/65536.0,1,-nbitq), 
to_sfixed(1924.0/65536.0,1,-nbitq), 
to_sfixed(-819.0/65536.0,1,-nbitq), 
to_sfixed(-71.0/65536.0,1,-nbitq), 
to_sfixed(-1790.0/65536.0,1,-nbitq), 
to_sfixed(-2379.0/65536.0,1,-nbitq), 
to_sfixed(-2463.0/65536.0,1,-nbitq), 
to_sfixed(-537.0/65536.0,1,-nbitq), 
to_sfixed(-502.0/65536.0,1,-nbitq), 
to_sfixed(542.0/65536.0,1,-nbitq), 
to_sfixed(2016.0/65536.0,1,-nbitq), 
to_sfixed(433.0/65536.0,1,-nbitq), 
to_sfixed(1290.0/65536.0,1,-nbitq), 
to_sfixed(282.0/65536.0,1,-nbitq), 
to_sfixed(-2051.0/65536.0,1,-nbitq), 
to_sfixed(-1760.0/65536.0,1,-nbitq), 
to_sfixed(694.0/65536.0,1,-nbitq), 
to_sfixed(121.0/65536.0,1,-nbitq), 
to_sfixed(2108.0/65536.0,1,-nbitq), 
to_sfixed(-65.0/65536.0,1,-nbitq), 
to_sfixed(-1396.0/65536.0,1,-nbitq), 
to_sfixed(52.0/65536.0,1,-nbitq), 
to_sfixed(-2386.0/65536.0,1,-nbitq), 
to_sfixed(-1038.0/65536.0,1,-nbitq), 
to_sfixed(2835.0/65536.0,1,-nbitq), 
to_sfixed(2313.0/65536.0,1,-nbitq), 
to_sfixed(2425.0/65536.0,1,-nbitq), 
to_sfixed(2998.0/65536.0,1,-nbitq), 
to_sfixed(-1217.0/65536.0,1,-nbitq), 
to_sfixed(1215.0/65536.0,1,-nbitq), 
to_sfixed(1347.0/65536.0,1,-nbitq), 
to_sfixed(-947.0/65536.0,1,-nbitq), 
to_sfixed(-368.0/65536.0,1,-nbitq), 
to_sfixed(1491.0/65536.0,1,-nbitq), 
to_sfixed(-1955.0/65536.0,1,-nbitq), 
to_sfixed(134.0/65536.0,1,-nbitq), 
to_sfixed(-240.0/65536.0,1,-nbitq), 
to_sfixed(-3018.0/65536.0,1,-nbitq), 
to_sfixed(-376.0/65536.0,1,-nbitq), 
to_sfixed(52.0/65536.0,1,-nbitq), 
to_sfixed(3462.0/65536.0,1,-nbitq), 
to_sfixed(1388.0/65536.0,1,-nbitq), 
to_sfixed(8477.0/65536.0,1,-nbitq), 
to_sfixed(81.0/65536.0,1,-nbitq), 
to_sfixed(577.0/65536.0,1,-nbitq), 
to_sfixed(4812.0/65536.0,1,-nbitq), 
to_sfixed(-414.0/65536.0,1,-nbitq), 
to_sfixed(-159.0/65536.0,1,-nbitq), 
to_sfixed(727.0/65536.0,1,-nbitq), 
to_sfixed(-1803.0/65536.0,1,-nbitq), 
to_sfixed(-3451.0/65536.0,1,-nbitq), 
to_sfixed(-1243.0/65536.0,1,-nbitq), 
to_sfixed(-621.0/65536.0,1,-nbitq), 
to_sfixed(-1621.0/65536.0,1,-nbitq)  ), 
( to_sfixed(556.0/65536.0,1,-nbitq), 
to_sfixed(-2973.0/65536.0,1,-nbitq), 
to_sfixed(-1170.0/65536.0,1,-nbitq), 
to_sfixed(-19.0/65536.0,1,-nbitq), 
to_sfixed(-592.0/65536.0,1,-nbitq), 
to_sfixed(-1715.0/65536.0,1,-nbitq), 
to_sfixed(-2788.0/65536.0,1,-nbitq), 
to_sfixed(-249.0/65536.0,1,-nbitq), 
to_sfixed(-4241.0/65536.0,1,-nbitq), 
to_sfixed(1436.0/65536.0,1,-nbitq), 
to_sfixed(-2804.0/65536.0,1,-nbitq), 
to_sfixed(2158.0/65536.0,1,-nbitq), 
to_sfixed(-291.0/65536.0,1,-nbitq), 
to_sfixed(-2079.0/65536.0,1,-nbitq), 
to_sfixed(-1935.0/65536.0,1,-nbitq), 
to_sfixed(-2270.0/65536.0,1,-nbitq), 
to_sfixed(-916.0/65536.0,1,-nbitq), 
to_sfixed(583.0/65536.0,1,-nbitq), 
to_sfixed(1095.0/65536.0,1,-nbitq), 
to_sfixed(2274.0/65536.0,1,-nbitq), 
to_sfixed(140.0/65536.0,1,-nbitq), 
to_sfixed(2170.0/65536.0,1,-nbitq), 
to_sfixed(-1228.0/65536.0,1,-nbitq), 
to_sfixed(1749.0/65536.0,1,-nbitq), 
to_sfixed(-281.0/65536.0,1,-nbitq), 
to_sfixed(-1701.0/65536.0,1,-nbitq), 
to_sfixed(-2024.0/65536.0,1,-nbitq), 
to_sfixed(247.0/65536.0,1,-nbitq), 
to_sfixed(986.0/65536.0,1,-nbitq), 
to_sfixed(-1707.0/65536.0,1,-nbitq), 
to_sfixed(317.0/65536.0,1,-nbitq), 
to_sfixed(-2415.0/65536.0,1,-nbitq), 
to_sfixed(-3172.0/65536.0,1,-nbitq), 
to_sfixed(-3980.0/65536.0,1,-nbitq), 
to_sfixed(2585.0/65536.0,1,-nbitq), 
to_sfixed(800.0/65536.0,1,-nbitq), 
to_sfixed(1637.0/65536.0,1,-nbitq), 
to_sfixed(-1427.0/65536.0,1,-nbitq), 
to_sfixed(-1563.0/65536.0,1,-nbitq), 
to_sfixed(450.0/65536.0,1,-nbitq), 
to_sfixed(307.0/65536.0,1,-nbitq), 
to_sfixed(-251.0/65536.0,1,-nbitq), 
to_sfixed(-1419.0/65536.0,1,-nbitq), 
to_sfixed(-988.0/65536.0,1,-nbitq), 
to_sfixed(1928.0/65536.0,1,-nbitq), 
to_sfixed(2999.0/65536.0,1,-nbitq), 
to_sfixed(-800.0/65536.0,1,-nbitq), 
to_sfixed(-1296.0/65536.0,1,-nbitq), 
to_sfixed(-797.0/65536.0,1,-nbitq), 
to_sfixed(-405.0/65536.0,1,-nbitq), 
to_sfixed(-571.0/65536.0,1,-nbitq), 
to_sfixed(2386.0/65536.0,1,-nbitq), 
to_sfixed(-742.0/65536.0,1,-nbitq), 
to_sfixed(-2855.0/65536.0,1,-nbitq), 
to_sfixed(626.0/65536.0,1,-nbitq), 
to_sfixed(-2929.0/65536.0,1,-nbitq), 
to_sfixed(-361.0/65536.0,1,-nbitq), 
to_sfixed(-2358.0/65536.0,1,-nbitq), 
to_sfixed(1198.0/65536.0,1,-nbitq), 
to_sfixed(1561.0/65536.0,1,-nbitq), 
to_sfixed(-30.0/65536.0,1,-nbitq), 
to_sfixed(709.0/65536.0,1,-nbitq), 
to_sfixed(1092.0/65536.0,1,-nbitq), 
to_sfixed(848.0/65536.0,1,-nbitq), 
to_sfixed(-822.0/65536.0,1,-nbitq), 
to_sfixed(-2714.0/65536.0,1,-nbitq), 
to_sfixed(2833.0/65536.0,1,-nbitq), 
to_sfixed(-2121.0/65536.0,1,-nbitq), 
to_sfixed(4816.0/65536.0,1,-nbitq), 
to_sfixed(-539.0/65536.0,1,-nbitq), 
to_sfixed(1193.0/65536.0,1,-nbitq), 
to_sfixed(1325.0/65536.0,1,-nbitq), 
to_sfixed(789.0/65536.0,1,-nbitq), 
to_sfixed(250.0/65536.0,1,-nbitq), 
to_sfixed(2242.0/65536.0,1,-nbitq), 
to_sfixed(-2910.0/65536.0,1,-nbitq), 
to_sfixed(2240.0/65536.0,1,-nbitq), 
to_sfixed(3507.0/65536.0,1,-nbitq), 
to_sfixed(-3117.0/65536.0,1,-nbitq), 
to_sfixed(3838.0/65536.0,1,-nbitq)  ), 
( to_sfixed(739.0/65536.0,1,-nbitq), 
to_sfixed(-23.0/65536.0,1,-nbitq), 
to_sfixed(331.0/65536.0,1,-nbitq), 
to_sfixed(-1398.0/65536.0,1,-nbitq), 
to_sfixed(-2613.0/65536.0,1,-nbitq), 
to_sfixed(-1706.0/65536.0,1,-nbitq), 
to_sfixed(439.0/65536.0,1,-nbitq), 
to_sfixed(1207.0/65536.0,1,-nbitq), 
to_sfixed(-1316.0/65536.0,1,-nbitq), 
to_sfixed(2666.0/65536.0,1,-nbitq), 
to_sfixed(-2529.0/65536.0,1,-nbitq), 
to_sfixed(3605.0/65536.0,1,-nbitq), 
to_sfixed(-2892.0/65536.0,1,-nbitq), 
to_sfixed(-1171.0/65536.0,1,-nbitq), 
to_sfixed(997.0/65536.0,1,-nbitq), 
to_sfixed(1442.0/65536.0,1,-nbitq), 
to_sfixed(-75.0/65536.0,1,-nbitq), 
to_sfixed(1888.0/65536.0,1,-nbitq), 
to_sfixed(2875.0/65536.0,1,-nbitq), 
to_sfixed(2299.0/65536.0,1,-nbitq), 
to_sfixed(-2310.0/65536.0,1,-nbitq), 
to_sfixed(365.0/65536.0,1,-nbitq), 
to_sfixed(1565.0/65536.0,1,-nbitq), 
to_sfixed(1756.0/65536.0,1,-nbitq), 
to_sfixed(-295.0/65536.0,1,-nbitq), 
to_sfixed(2557.0/65536.0,1,-nbitq), 
to_sfixed(-393.0/65536.0,1,-nbitq), 
to_sfixed(-1889.0/65536.0,1,-nbitq), 
to_sfixed(-593.0/65536.0,1,-nbitq), 
to_sfixed(-3123.0/65536.0,1,-nbitq), 
to_sfixed(-442.0/65536.0,1,-nbitq), 
to_sfixed(2321.0/65536.0,1,-nbitq), 
to_sfixed(-5065.0/65536.0,1,-nbitq), 
to_sfixed(942.0/65536.0,1,-nbitq), 
to_sfixed(-1908.0/65536.0,1,-nbitq), 
to_sfixed(-957.0/65536.0,1,-nbitq), 
to_sfixed(-2515.0/65536.0,1,-nbitq), 
to_sfixed(-3924.0/65536.0,1,-nbitq), 
to_sfixed(-1880.0/65536.0,1,-nbitq), 
to_sfixed(-1323.0/65536.0,1,-nbitq), 
to_sfixed(-3222.0/65536.0,1,-nbitq), 
to_sfixed(-295.0/65536.0,1,-nbitq), 
to_sfixed(-3708.0/65536.0,1,-nbitq), 
to_sfixed(341.0/65536.0,1,-nbitq), 
to_sfixed(702.0/65536.0,1,-nbitq), 
to_sfixed(3181.0/65536.0,1,-nbitq), 
to_sfixed(-62.0/65536.0,1,-nbitq), 
to_sfixed(-260.0/65536.0,1,-nbitq), 
to_sfixed(-136.0/65536.0,1,-nbitq), 
to_sfixed(382.0/65536.0,1,-nbitq), 
to_sfixed(-1486.0/65536.0,1,-nbitq), 
to_sfixed(-1941.0/65536.0,1,-nbitq), 
to_sfixed(-2435.0/65536.0,1,-nbitq), 
to_sfixed(862.0/65536.0,1,-nbitq), 
to_sfixed(1460.0/65536.0,1,-nbitq), 
to_sfixed(1293.0/65536.0,1,-nbitq), 
to_sfixed(1758.0/65536.0,1,-nbitq), 
to_sfixed(-1402.0/65536.0,1,-nbitq), 
to_sfixed(-2022.0/65536.0,1,-nbitq), 
to_sfixed(963.0/65536.0,1,-nbitq), 
to_sfixed(-1103.0/65536.0,1,-nbitq), 
to_sfixed(983.0/65536.0,1,-nbitq), 
to_sfixed(3055.0/65536.0,1,-nbitq), 
to_sfixed(-88.0/65536.0,1,-nbitq), 
to_sfixed(-2253.0/65536.0,1,-nbitq), 
to_sfixed(1300.0/65536.0,1,-nbitq), 
to_sfixed(-745.0/65536.0,1,-nbitq), 
to_sfixed(-1252.0/65536.0,1,-nbitq), 
to_sfixed(568.0/65536.0,1,-nbitq), 
to_sfixed(-1716.0/65536.0,1,-nbitq), 
to_sfixed(-302.0/65536.0,1,-nbitq), 
to_sfixed(3156.0/65536.0,1,-nbitq), 
to_sfixed(4146.0/65536.0,1,-nbitq), 
to_sfixed(842.0/65536.0,1,-nbitq), 
to_sfixed(2636.0/65536.0,1,-nbitq), 
to_sfixed(-1811.0/65536.0,1,-nbitq), 
to_sfixed(520.0/65536.0,1,-nbitq), 
to_sfixed(1377.0/65536.0,1,-nbitq), 
to_sfixed(215.0/65536.0,1,-nbitq), 
to_sfixed(79.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1133.0/65536.0,1,-nbitq), 
to_sfixed(-1421.0/65536.0,1,-nbitq), 
to_sfixed(1192.0/65536.0,1,-nbitq), 
to_sfixed(-1380.0/65536.0,1,-nbitq), 
to_sfixed(-2014.0/65536.0,1,-nbitq), 
to_sfixed(-1540.0/65536.0,1,-nbitq), 
to_sfixed(1362.0/65536.0,1,-nbitq), 
to_sfixed(-947.0/65536.0,1,-nbitq), 
to_sfixed(-681.0/65536.0,1,-nbitq), 
to_sfixed(-2147.0/65536.0,1,-nbitq), 
to_sfixed(-1218.0/65536.0,1,-nbitq), 
to_sfixed(183.0/65536.0,1,-nbitq), 
to_sfixed(-1027.0/65536.0,1,-nbitq), 
to_sfixed(1350.0/65536.0,1,-nbitq), 
to_sfixed(-504.0/65536.0,1,-nbitq), 
to_sfixed(-59.0/65536.0,1,-nbitq), 
to_sfixed(-1756.0/65536.0,1,-nbitq), 
to_sfixed(2707.0/65536.0,1,-nbitq), 
to_sfixed(-78.0/65536.0,1,-nbitq), 
to_sfixed(622.0/65536.0,1,-nbitq), 
to_sfixed(-1103.0/65536.0,1,-nbitq), 
to_sfixed(1972.0/65536.0,1,-nbitq), 
to_sfixed(2476.0/65536.0,1,-nbitq), 
to_sfixed(-577.0/65536.0,1,-nbitq), 
to_sfixed(2499.0/65536.0,1,-nbitq), 
to_sfixed(1790.0/65536.0,1,-nbitq), 
to_sfixed(-3702.0/65536.0,1,-nbitq), 
to_sfixed(-1386.0/65536.0,1,-nbitq), 
to_sfixed(-1603.0/65536.0,1,-nbitq), 
to_sfixed(-537.0/65536.0,1,-nbitq), 
to_sfixed(1520.0/65536.0,1,-nbitq), 
to_sfixed(2454.0/65536.0,1,-nbitq), 
to_sfixed(-2047.0/65536.0,1,-nbitq), 
to_sfixed(60.0/65536.0,1,-nbitq), 
to_sfixed(1573.0/65536.0,1,-nbitq), 
to_sfixed(-41.0/65536.0,1,-nbitq), 
to_sfixed(2190.0/65536.0,1,-nbitq), 
to_sfixed(-141.0/65536.0,1,-nbitq), 
to_sfixed(-3629.0/65536.0,1,-nbitq), 
to_sfixed(1744.0/65536.0,1,-nbitq), 
to_sfixed(-150.0/65536.0,1,-nbitq), 
to_sfixed(-907.0/65536.0,1,-nbitq), 
to_sfixed(-63.0/65536.0,1,-nbitq), 
to_sfixed(-1600.0/65536.0,1,-nbitq), 
to_sfixed(-2069.0/65536.0,1,-nbitq), 
to_sfixed(6178.0/65536.0,1,-nbitq), 
to_sfixed(-146.0/65536.0,1,-nbitq), 
to_sfixed(624.0/65536.0,1,-nbitq), 
to_sfixed(2976.0/65536.0,1,-nbitq), 
to_sfixed(741.0/65536.0,1,-nbitq), 
to_sfixed(1380.0/65536.0,1,-nbitq), 
to_sfixed(1778.0/65536.0,1,-nbitq), 
to_sfixed(-1149.0/65536.0,1,-nbitq), 
to_sfixed(-441.0/65536.0,1,-nbitq), 
to_sfixed(969.0/65536.0,1,-nbitq), 
to_sfixed(1184.0/65536.0,1,-nbitq), 
to_sfixed(447.0/65536.0,1,-nbitq), 
to_sfixed(134.0/65536.0,1,-nbitq), 
to_sfixed(-1449.0/65536.0,1,-nbitq), 
to_sfixed(5910.0/65536.0,1,-nbitq), 
to_sfixed(1823.0/65536.0,1,-nbitq), 
to_sfixed(1590.0/65536.0,1,-nbitq), 
to_sfixed(3005.0/65536.0,1,-nbitq), 
to_sfixed(-254.0/65536.0,1,-nbitq), 
to_sfixed(-1718.0/65536.0,1,-nbitq), 
to_sfixed(1926.0/65536.0,1,-nbitq), 
to_sfixed(-1399.0/65536.0,1,-nbitq), 
to_sfixed(-103.0/65536.0,1,-nbitq), 
to_sfixed(3256.0/65536.0,1,-nbitq), 
to_sfixed(-2156.0/65536.0,1,-nbitq), 
to_sfixed(-648.0/65536.0,1,-nbitq), 
to_sfixed(3121.0/65536.0,1,-nbitq), 
to_sfixed(1111.0/65536.0,1,-nbitq), 
to_sfixed(-349.0/65536.0,1,-nbitq), 
to_sfixed(-2993.0/65536.0,1,-nbitq), 
to_sfixed(837.0/65536.0,1,-nbitq), 
to_sfixed(269.0/65536.0,1,-nbitq), 
to_sfixed(3912.0/65536.0,1,-nbitq), 
to_sfixed(-2709.0/65536.0,1,-nbitq), 
to_sfixed(4182.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2425.0/65536.0,1,-nbitq), 
to_sfixed(709.0/65536.0,1,-nbitq), 
to_sfixed(4425.0/65536.0,1,-nbitq), 
to_sfixed(2293.0/65536.0,1,-nbitq), 
to_sfixed(605.0/65536.0,1,-nbitq), 
to_sfixed(-2716.0/65536.0,1,-nbitq), 
to_sfixed(1297.0/65536.0,1,-nbitq), 
to_sfixed(-1772.0/65536.0,1,-nbitq), 
to_sfixed(-269.0/65536.0,1,-nbitq), 
to_sfixed(1022.0/65536.0,1,-nbitq), 
to_sfixed(-3374.0/65536.0,1,-nbitq), 
to_sfixed(-780.0/65536.0,1,-nbitq), 
to_sfixed(2700.0/65536.0,1,-nbitq), 
to_sfixed(1043.0/65536.0,1,-nbitq), 
to_sfixed(1980.0/65536.0,1,-nbitq), 
to_sfixed(1441.0/65536.0,1,-nbitq), 
to_sfixed(-1701.0/65536.0,1,-nbitq), 
to_sfixed(-3841.0/65536.0,1,-nbitq), 
to_sfixed(871.0/65536.0,1,-nbitq), 
to_sfixed(-1843.0/65536.0,1,-nbitq), 
to_sfixed(-2703.0/65536.0,1,-nbitq), 
to_sfixed(-509.0/65536.0,1,-nbitq), 
to_sfixed(874.0/65536.0,1,-nbitq), 
to_sfixed(4222.0/65536.0,1,-nbitq), 
to_sfixed(-1378.0/65536.0,1,-nbitq), 
to_sfixed(1176.0/65536.0,1,-nbitq), 
to_sfixed(1205.0/65536.0,1,-nbitq), 
to_sfixed(-2257.0/65536.0,1,-nbitq), 
to_sfixed(943.0/65536.0,1,-nbitq), 
to_sfixed(-2968.0/65536.0,1,-nbitq), 
to_sfixed(2296.0/65536.0,1,-nbitq), 
to_sfixed(72.0/65536.0,1,-nbitq), 
to_sfixed(-20.0/65536.0,1,-nbitq), 
to_sfixed(-1351.0/65536.0,1,-nbitq), 
to_sfixed(1344.0/65536.0,1,-nbitq), 
to_sfixed(-2962.0/65536.0,1,-nbitq), 
to_sfixed(-2278.0/65536.0,1,-nbitq), 
to_sfixed(-3023.0/65536.0,1,-nbitq), 
to_sfixed(-1684.0/65536.0,1,-nbitq), 
to_sfixed(1667.0/65536.0,1,-nbitq), 
to_sfixed(2169.0/65536.0,1,-nbitq), 
to_sfixed(-1238.0/65536.0,1,-nbitq), 
to_sfixed(-4074.0/65536.0,1,-nbitq), 
to_sfixed(1379.0/65536.0,1,-nbitq), 
to_sfixed(2331.0/65536.0,1,-nbitq), 
to_sfixed(3863.0/65536.0,1,-nbitq), 
to_sfixed(-2093.0/65536.0,1,-nbitq), 
to_sfixed(-457.0/65536.0,1,-nbitq), 
to_sfixed(1698.0/65536.0,1,-nbitq), 
to_sfixed(1811.0/65536.0,1,-nbitq), 
to_sfixed(3246.0/65536.0,1,-nbitq), 
to_sfixed(-608.0/65536.0,1,-nbitq), 
to_sfixed(3116.0/65536.0,1,-nbitq), 
to_sfixed(-1764.0/65536.0,1,-nbitq), 
to_sfixed(-1019.0/65536.0,1,-nbitq), 
to_sfixed(-2255.0/65536.0,1,-nbitq), 
to_sfixed(1576.0/65536.0,1,-nbitq), 
to_sfixed(-1268.0/65536.0,1,-nbitq), 
to_sfixed(-1083.0/65536.0,1,-nbitq), 
to_sfixed(1567.0/65536.0,1,-nbitq), 
to_sfixed(-2344.0/65536.0,1,-nbitq), 
to_sfixed(-1611.0/65536.0,1,-nbitq), 
to_sfixed(-55.0/65536.0,1,-nbitq), 
to_sfixed(2566.0/65536.0,1,-nbitq), 
to_sfixed(2897.0/65536.0,1,-nbitq), 
to_sfixed(2924.0/65536.0,1,-nbitq), 
to_sfixed(-1484.0/65536.0,1,-nbitq), 
to_sfixed(494.0/65536.0,1,-nbitq), 
to_sfixed(2342.0/65536.0,1,-nbitq), 
to_sfixed(2517.0/65536.0,1,-nbitq), 
to_sfixed(895.0/65536.0,1,-nbitq), 
to_sfixed(-1893.0/65536.0,1,-nbitq), 
to_sfixed(1063.0/65536.0,1,-nbitq), 
to_sfixed(614.0/65536.0,1,-nbitq), 
to_sfixed(-2854.0/65536.0,1,-nbitq), 
to_sfixed(-1960.0/65536.0,1,-nbitq), 
to_sfixed(-1710.0/65536.0,1,-nbitq), 
to_sfixed(5045.0/65536.0,1,-nbitq), 
to_sfixed(-70.0/65536.0,1,-nbitq), 
to_sfixed(4632.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1287.0/65536.0,1,-nbitq), 
to_sfixed(2831.0/65536.0,1,-nbitq), 
to_sfixed(3365.0/65536.0,1,-nbitq), 
to_sfixed(1736.0/65536.0,1,-nbitq), 
to_sfixed(-5349.0/65536.0,1,-nbitq), 
to_sfixed(-3302.0/65536.0,1,-nbitq), 
to_sfixed(1325.0/65536.0,1,-nbitq), 
to_sfixed(-1130.0/65536.0,1,-nbitq), 
to_sfixed(-6960.0/65536.0,1,-nbitq), 
to_sfixed(-593.0/65536.0,1,-nbitq), 
to_sfixed(-2078.0/65536.0,1,-nbitq), 
to_sfixed(-3734.0/65536.0,1,-nbitq), 
to_sfixed(-1916.0/65536.0,1,-nbitq), 
to_sfixed(-2857.0/65536.0,1,-nbitq), 
to_sfixed(982.0/65536.0,1,-nbitq), 
to_sfixed(778.0/65536.0,1,-nbitq), 
to_sfixed(-2152.0/65536.0,1,-nbitq), 
to_sfixed(-51.0/65536.0,1,-nbitq), 
to_sfixed(-2619.0/65536.0,1,-nbitq), 
to_sfixed(-1332.0/65536.0,1,-nbitq), 
to_sfixed(-710.0/65536.0,1,-nbitq), 
to_sfixed(2175.0/65536.0,1,-nbitq), 
to_sfixed(-2119.0/65536.0,1,-nbitq), 
to_sfixed(3908.0/65536.0,1,-nbitq), 
to_sfixed(-470.0/65536.0,1,-nbitq), 
to_sfixed(-1713.0/65536.0,1,-nbitq), 
to_sfixed(-1457.0/65536.0,1,-nbitq), 
to_sfixed(-1631.0/65536.0,1,-nbitq), 
to_sfixed(857.0/65536.0,1,-nbitq), 
to_sfixed(1949.0/65536.0,1,-nbitq), 
to_sfixed(1126.0/65536.0,1,-nbitq), 
to_sfixed(-56.0/65536.0,1,-nbitq), 
to_sfixed(-5381.0/65536.0,1,-nbitq), 
to_sfixed(-5219.0/65536.0,1,-nbitq), 
to_sfixed(231.0/65536.0,1,-nbitq), 
to_sfixed(-2921.0/65536.0,1,-nbitq), 
to_sfixed(-1403.0/65536.0,1,-nbitq), 
to_sfixed(-1023.0/65536.0,1,-nbitq), 
to_sfixed(-25.0/65536.0,1,-nbitq), 
to_sfixed(-1563.0/65536.0,1,-nbitq), 
to_sfixed(1392.0/65536.0,1,-nbitq), 
to_sfixed(139.0/65536.0,1,-nbitq), 
to_sfixed(-1650.0/65536.0,1,-nbitq), 
to_sfixed(2885.0/65536.0,1,-nbitq), 
to_sfixed(1120.0/65536.0,1,-nbitq), 
to_sfixed(1823.0/65536.0,1,-nbitq), 
to_sfixed(190.0/65536.0,1,-nbitq), 
to_sfixed(2503.0/65536.0,1,-nbitq), 
to_sfixed(3602.0/65536.0,1,-nbitq), 
to_sfixed(3733.0/65536.0,1,-nbitq), 
to_sfixed(-482.0/65536.0,1,-nbitq), 
to_sfixed(2303.0/65536.0,1,-nbitq), 
to_sfixed(3504.0/65536.0,1,-nbitq), 
to_sfixed(-1186.0/65536.0,1,-nbitq), 
to_sfixed(1053.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(724.0/65536.0,1,-nbitq), 
to_sfixed(-1600.0/65536.0,1,-nbitq), 
to_sfixed(2421.0/65536.0,1,-nbitq), 
to_sfixed(2246.0/65536.0,1,-nbitq), 
to_sfixed(1673.0/65536.0,1,-nbitq), 
to_sfixed(827.0/65536.0,1,-nbitq), 
to_sfixed(1413.0/65536.0,1,-nbitq), 
to_sfixed(2383.0/65536.0,1,-nbitq), 
to_sfixed(6733.0/65536.0,1,-nbitq), 
to_sfixed(2324.0/65536.0,1,-nbitq), 
to_sfixed(-1527.0/65536.0,1,-nbitq), 
to_sfixed(-1388.0/65536.0,1,-nbitq), 
to_sfixed(1278.0/65536.0,1,-nbitq), 
to_sfixed(-842.0/65536.0,1,-nbitq), 
to_sfixed(411.0/65536.0,1,-nbitq), 
to_sfixed(3300.0/65536.0,1,-nbitq), 
to_sfixed(1578.0/65536.0,1,-nbitq), 
to_sfixed(-1733.0/65536.0,1,-nbitq), 
to_sfixed(-1079.0/65536.0,1,-nbitq), 
to_sfixed(-1489.0/65536.0,1,-nbitq), 
to_sfixed(-1313.0/65536.0,1,-nbitq), 
to_sfixed(640.0/65536.0,1,-nbitq), 
to_sfixed(1865.0/65536.0,1,-nbitq), 
to_sfixed(1570.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3617.0/65536.0,1,-nbitq), 
to_sfixed(-943.0/65536.0,1,-nbitq), 
to_sfixed(6444.0/65536.0,1,-nbitq), 
to_sfixed(-1772.0/65536.0,1,-nbitq), 
to_sfixed(-905.0/65536.0,1,-nbitq), 
to_sfixed(-1251.0/65536.0,1,-nbitq), 
to_sfixed(-2676.0/65536.0,1,-nbitq), 
to_sfixed(-913.0/65536.0,1,-nbitq), 
to_sfixed(-4987.0/65536.0,1,-nbitq), 
to_sfixed(1274.0/65536.0,1,-nbitq), 
to_sfixed(448.0/65536.0,1,-nbitq), 
to_sfixed(-4667.0/65536.0,1,-nbitq), 
to_sfixed(-1770.0/65536.0,1,-nbitq), 
to_sfixed(-2814.0/65536.0,1,-nbitq), 
to_sfixed(-531.0/65536.0,1,-nbitq), 
to_sfixed(1038.0/65536.0,1,-nbitq), 
to_sfixed(1734.0/65536.0,1,-nbitq), 
to_sfixed(-2266.0/65536.0,1,-nbitq), 
to_sfixed(-1727.0/65536.0,1,-nbitq), 
to_sfixed(-1775.0/65536.0,1,-nbitq), 
to_sfixed(-1749.0/65536.0,1,-nbitq), 
to_sfixed(1569.0/65536.0,1,-nbitq), 
to_sfixed(-2383.0/65536.0,1,-nbitq), 
to_sfixed(1177.0/65536.0,1,-nbitq), 
to_sfixed(2919.0/65536.0,1,-nbitq), 
to_sfixed(4767.0/65536.0,1,-nbitq), 
to_sfixed(-1692.0/65536.0,1,-nbitq), 
to_sfixed(1497.0/65536.0,1,-nbitq), 
to_sfixed(435.0/65536.0,1,-nbitq), 
to_sfixed(326.0/65536.0,1,-nbitq), 
to_sfixed(1187.0/65536.0,1,-nbitq), 
to_sfixed(-932.0/65536.0,1,-nbitq), 
to_sfixed(-2254.0/65536.0,1,-nbitq), 
to_sfixed(-3795.0/65536.0,1,-nbitq), 
to_sfixed(1933.0/65536.0,1,-nbitq), 
to_sfixed(-2912.0/65536.0,1,-nbitq), 
to_sfixed(-1886.0/65536.0,1,-nbitq), 
to_sfixed(1495.0/65536.0,1,-nbitq), 
to_sfixed(3843.0/65536.0,1,-nbitq), 
to_sfixed(1439.0/65536.0,1,-nbitq), 
to_sfixed(1442.0/65536.0,1,-nbitq), 
to_sfixed(1589.0/65536.0,1,-nbitq), 
to_sfixed(-2514.0/65536.0,1,-nbitq), 
to_sfixed(2181.0/65536.0,1,-nbitq), 
to_sfixed(-2475.0/65536.0,1,-nbitq), 
to_sfixed(3075.0/65536.0,1,-nbitq), 
to_sfixed(377.0/65536.0,1,-nbitq), 
to_sfixed(2444.0/65536.0,1,-nbitq), 
to_sfixed(-1202.0/65536.0,1,-nbitq), 
to_sfixed(3730.0/65536.0,1,-nbitq), 
to_sfixed(3244.0/65536.0,1,-nbitq), 
to_sfixed(99.0/65536.0,1,-nbitq), 
to_sfixed(1839.0/65536.0,1,-nbitq), 
to_sfixed(-2594.0/65536.0,1,-nbitq), 
to_sfixed(687.0/65536.0,1,-nbitq), 
to_sfixed(-564.0/65536.0,1,-nbitq), 
to_sfixed(-835.0/65536.0,1,-nbitq), 
to_sfixed(-3497.0/65536.0,1,-nbitq), 
to_sfixed(-1102.0/65536.0,1,-nbitq), 
to_sfixed(1462.0/65536.0,1,-nbitq), 
to_sfixed(-1021.0/65536.0,1,-nbitq), 
to_sfixed(957.0/65536.0,1,-nbitq), 
to_sfixed(-2033.0/65536.0,1,-nbitq), 
to_sfixed(1573.0/65536.0,1,-nbitq), 
to_sfixed(7209.0/65536.0,1,-nbitq), 
to_sfixed(2440.0/65536.0,1,-nbitq), 
to_sfixed(28.0/65536.0,1,-nbitq), 
to_sfixed(-2306.0/65536.0,1,-nbitq), 
to_sfixed(1697.0/65536.0,1,-nbitq), 
to_sfixed(-150.0/65536.0,1,-nbitq), 
to_sfixed(-2548.0/65536.0,1,-nbitq), 
to_sfixed(4111.0/65536.0,1,-nbitq), 
to_sfixed(-1543.0/65536.0,1,-nbitq), 
to_sfixed(-451.0/65536.0,1,-nbitq), 
to_sfixed(-888.0/65536.0,1,-nbitq), 
to_sfixed(798.0/65536.0,1,-nbitq), 
to_sfixed(2306.0/65536.0,1,-nbitq), 
to_sfixed(4211.0/65536.0,1,-nbitq), 
to_sfixed(-3099.0/65536.0,1,-nbitq), 
to_sfixed(4067.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-778.0/65536.0,1,-nbitq), 
to_sfixed(-20.0/65536.0,1,-nbitq), 
to_sfixed(4698.0/65536.0,1,-nbitq), 
to_sfixed(2048.0/65536.0,1,-nbitq), 
to_sfixed(3639.0/65536.0,1,-nbitq), 
to_sfixed(-3651.0/65536.0,1,-nbitq), 
to_sfixed(2377.0/65536.0,1,-nbitq), 
to_sfixed(-3306.0/65536.0,1,-nbitq), 
to_sfixed(-3969.0/65536.0,1,-nbitq), 
to_sfixed(1937.0/65536.0,1,-nbitq), 
to_sfixed(-1562.0/65536.0,1,-nbitq), 
to_sfixed(-5407.0/65536.0,1,-nbitq), 
to_sfixed(-2171.0/65536.0,1,-nbitq), 
to_sfixed(1307.0/65536.0,1,-nbitq), 
to_sfixed(1399.0/65536.0,1,-nbitq), 
to_sfixed(-1016.0/65536.0,1,-nbitq), 
to_sfixed(-1183.0/65536.0,1,-nbitq), 
to_sfixed(-2199.0/65536.0,1,-nbitq), 
to_sfixed(1913.0/65536.0,1,-nbitq), 
to_sfixed(1526.0/65536.0,1,-nbitq), 
to_sfixed(-734.0/65536.0,1,-nbitq), 
to_sfixed(-2299.0/65536.0,1,-nbitq), 
to_sfixed(-650.0/65536.0,1,-nbitq), 
to_sfixed(-933.0/65536.0,1,-nbitq), 
to_sfixed(-1860.0/65536.0,1,-nbitq), 
to_sfixed(309.0/65536.0,1,-nbitq), 
to_sfixed(315.0/65536.0,1,-nbitq), 
to_sfixed(1713.0/65536.0,1,-nbitq), 
to_sfixed(3355.0/65536.0,1,-nbitq), 
to_sfixed(-2752.0/65536.0,1,-nbitq), 
to_sfixed(-1527.0/65536.0,1,-nbitq), 
to_sfixed(118.0/65536.0,1,-nbitq), 
to_sfixed(-2844.0/65536.0,1,-nbitq), 
to_sfixed(-4893.0/65536.0,1,-nbitq), 
to_sfixed(2360.0/65536.0,1,-nbitq), 
to_sfixed(1825.0/65536.0,1,-nbitq), 
to_sfixed(-650.0/65536.0,1,-nbitq), 
to_sfixed(584.0/65536.0,1,-nbitq), 
to_sfixed(987.0/65536.0,1,-nbitq), 
to_sfixed(-4.0/65536.0,1,-nbitq), 
to_sfixed(139.0/65536.0,1,-nbitq), 
to_sfixed(-3180.0/65536.0,1,-nbitq), 
to_sfixed(1592.0/65536.0,1,-nbitq), 
to_sfixed(1893.0/65536.0,1,-nbitq), 
to_sfixed(-1253.0/65536.0,1,-nbitq), 
to_sfixed(1996.0/65536.0,1,-nbitq), 
to_sfixed(1925.0/65536.0,1,-nbitq), 
to_sfixed(-1079.0/65536.0,1,-nbitq), 
to_sfixed(-1248.0/65536.0,1,-nbitq), 
to_sfixed(1983.0/65536.0,1,-nbitq), 
to_sfixed(2050.0/65536.0,1,-nbitq), 
to_sfixed(2922.0/65536.0,1,-nbitq), 
to_sfixed(2007.0/65536.0,1,-nbitq), 
to_sfixed(-1469.0/65536.0,1,-nbitq), 
to_sfixed(289.0/65536.0,1,-nbitq), 
to_sfixed(-1825.0/65536.0,1,-nbitq), 
to_sfixed(-2820.0/65536.0,1,-nbitq), 
to_sfixed(152.0/65536.0,1,-nbitq), 
to_sfixed(-2486.0/65536.0,1,-nbitq), 
to_sfixed(82.0/65536.0,1,-nbitq), 
to_sfixed(-2604.0/65536.0,1,-nbitq), 
to_sfixed(-189.0/65536.0,1,-nbitq), 
to_sfixed(-2756.0/65536.0,1,-nbitq), 
to_sfixed(-581.0/65536.0,1,-nbitq), 
to_sfixed(2299.0/65536.0,1,-nbitq), 
to_sfixed(-853.0/65536.0,1,-nbitq), 
to_sfixed(-1501.0/65536.0,1,-nbitq), 
to_sfixed(-3172.0/65536.0,1,-nbitq), 
to_sfixed(5864.0/65536.0,1,-nbitq), 
to_sfixed(-257.0/65536.0,1,-nbitq), 
to_sfixed(-1635.0/65536.0,1,-nbitq), 
to_sfixed(-1044.0/65536.0,1,-nbitq), 
to_sfixed(330.0/65536.0,1,-nbitq), 
to_sfixed(-863.0/65536.0,1,-nbitq), 
to_sfixed(-2518.0/65536.0,1,-nbitq), 
to_sfixed(509.0/65536.0,1,-nbitq), 
to_sfixed(-2460.0/65536.0,1,-nbitq), 
to_sfixed(1414.0/65536.0,1,-nbitq), 
to_sfixed(-1098.0/65536.0,1,-nbitq), 
to_sfixed(2657.0/65536.0,1,-nbitq)  ), 
( to_sfixed(344.0/65536.0,1,-nbitq), 
to_sfixed(-470.0/65536.0,1,-nbitq), 
to_sfixed(-1409.0/65536.0,1,-nbitq), 
to_sfixed(3268.0/65536.0,1,-nbitq), 
to_sfixed(2981.0/65536.0,1,-nbitq), 
to_sfixed(-584.0/65536.0,1,-nbitq), 
to_sfixed(3574.0/65536.0,1,-nbitq), 
to_sfixed(-4919.0/65536.0,1,-nbitq), 
to_sfixed(-3083.0/65536.0,1,-nbitq), 
to_sfixed(-1041.0/65536.0,1,-nbitq), 
to_sfixed(-144.0/65536.0,1,-nbitq), 
to_sfixed(-4702.0/65536.0,1,-nbitq), 
to_sfixed(-116.0/65536.0,1,-nbitq), 
to_sfixed(-4141.0/65536.0,1,-nbitq), 
to_sfixed(517.0/65536.0,1,-nbitq), 
to_sfixed(-151.0/65536.0,1,-nbitq), 
to_sfixed(41.0/65536.0,1,-nbitq), 
to_sfixed(-3959.0/65536.0,1,-nbitq), 
to_sfixed(-2462.0/65536.0,1,-nbitq), 
to_sfixed(-51.0/65536.0,1,-nbitq), 
to_sfixed(1384.0/65536.0,1,-nbitq), 
to_sfixed(-1658.0/65536.0,1,-nbitq), 
to_sfixed(-1812.0/65536.0,1,-nbitq), 
to_sfixed(-4395.0/65536.0,1,-nbitq), 
to_sfixed(2083.0/65536.0,1,-nbitq), 
to_sfixed(1207.0/65536.0,1,-nbitq), 
to_sfixed(-2807.0/65536.0,1,-nbitq), 
to_sfixed(694.0/65536.0,1,-nbitq), 
to_sfixed(2970.0/65536.0,1,-nbitq), 
to_sfixed(-5534.0/65536.0,1,-nbitq), 
to_sfixed(-2107.0/65536.0,1,-nbitq), 
to_sfixed(-3880.0/65536.0,1,-nbitq), 
to_sfixed(-543.0/65536.0,1,-nbitq), 
to_sfixed(3150.0/65536.0,1,-nbitq), 
to_sfixed(620.0/65536.0,1,-nbitq), 
to_sfixed(2479.0/65536.0,1,-nbitq), 
to_sfixed(-2278.0/65536.0,1,-nbitq), 
to_sfixed(-346.0/65536.0,1,-nbitq), 
to_sfixed(5535.0/65536.0,1,-nbitq), 
to_sfixed(-2869.0/65536.0,1,-nbitq), 
to_sfixed(1039.0/65536.0,1,-nbitq), 
to_sfixed(1250.0/65536.0,1,-nbitq), 
to_sfixed(3772.0/65536.0,1,-nbitq), 
to_sfixed(-625.0/65536.0,1,-nbitq), 
to_sfixed(444.0/65536.0,1,-nbitq), 
to_sfixed(3401.0/65536.0,1,-nbitq), 
to_sfixed(1630.0/65536.0,1,-nbitq), 
to_sfixed(-770.0/65536.0,1,-nbitq), 
to_sfixed(1954.0/65536.0,1,-nbitq), 
to_sfixed(3001.0/65536.0,1,-nbitq), 
to_sfixed(3186.0/65536.0,1,-nbitq), 
to_sfixed(4328.0/65536.0,1,-nbitq), 
to_sfixed(2329.0/65536.0,1,-nbitq), 
to_sfixed(-5655.0/65536.0,1,-nbitq), 
to_sfixed(-2729.0/65536.0,1,-nbitq), 
to_sfixed(352.0/65536.0,1,-nbitq), 
to_sfixed(-1728.0/65536.0,1,-nbitq), 
to_sfixed(-3815.0/65536.0,1,-nbitq), 
to_sfixed(1222.0/65536.0,1,-nbitq), 
to_sfixed(-718.0/65536.0,1,-nbitq), 
to_sfixed(-1923.0/65536.0,1,-nbitq), 
to_sfixed(194.0/65536.0,1,-nbitq), 
to_sfixed(2331.0/65536.0,1,-nbitq), 
to_sfixed(464.0/65536.0,1,-nbitq), 
to_sfixed(2417.0/65536.0,1,-nbitq), 
to_sfixed(-1271.0/65536.0,1,-nbitq), 
to_sfixed(-542.0/65536.0,1,-nbitq), 
to_sfixed(-5162.0/65536.0,1,-nbitq), 
to_sfixed(2453.0/65536.0,1,-nbitq), 
to_sfixed(1604.0/65536.0,1,-nbitq), 
to_sfixed(2099.0/65536.0,1,-nbitq), 
to_sfixed(2140.0/65536.0,1,-nbitq), 
to_sfixed(2975.0/65536.0,1,-nbitq), 
to_sfixed(-996.0/65536.0,1,-nbitq), 
to_sfixed(-2182.0/65536.0,1,-nbitq), 
to_sfixed(2185.0/65536.0,1,-nbitq), 
to_sfixed(-4447.0/65536.0,1,-nbitq), 
to_sfixed(534.0/65536.0,1,-nbitq), 
to_sfixed(-2206.0/65536.0,1,-nbitq), 
to_sfixed(3029.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2493.0/65536.0,1,-nbitq), 
to_sfixed(442.0/65536.0,1,-nbitq), 
to_sfixed(5524.0/65536.0,1,-nbitq), 
to_sfixed(1766.0/65536.0,1,-nbitq), 
to_sfixed(2081.0/65536.0,1,-nbitq), 
to_sfixed(-3996.0/65536.0,1,-nbitq), 
to_sfixed(992.0/65536.0,1,-nbitq), 
to_sfixed(-2761.0/65536.0,1,-nbitq), 
to_sfixed(-5653.0/65536.0,1,-nbitq), 
to_sfixed(808.0/65536.0,1,-nbitq), 
to_sfixed(-2661.0/65536.0,1,-nbitq), 
to_sfixed(-3066.0/65536.0,1,-nbitq), 
to_sfixed(-326.0/65536.0,1,-nbitq), 
to_sfixed(2526.0/65536.0,1,-nbitq), 
to_sfixed(-2216.0/65536.0,1,-nbitq), 
to_sfixed(-291.0/65536.0,1,-nbitq), 
to_sfixed(852.0/65536.0,1,-nbitq), 
to_sfixed(-5042.0/65536.0,1,-nbitq), 
to_sfixed(-7978.0/65536.0,1,-nbitq), 
to_sfixed(-2082.0/65536.0,1,-nbitq), 
to_sfixed(3946.0/65536.0,1,-nbitq), 
to_sfixed(1873.0/65536.0,1,-nbitq), 
to_sfixed(-611.0/65536.0,1,-nbitq), 
to_sfixed(-8872.0/65536.0,1,-nbitq), 
to_sfixed(4202.0/65536.0,1,-nbitq), 
to_sfixed(-7026.0/65536.0,1,-nbitq), 
to_sfixed(-55.0/65536.0,1,-nbitq), 
to_sfixed(-603.0/65536.0,1,-nbitq), 
to_sfixed(874.0/65536.0,1,-nbitq), 
to_sfixed(-6016.0/65536.0,1,-nbitq), 
to_sfixed(2883.0/65536.0,1,-nbitq), 
to_sfixed(764.0/65536.0,1,-nbitq), 
to_sfixed(121.0/65536.0,1,-nbitq), 
to_sfixed(8148.0/65536.0,1,-nbitq), 
to_sfixed(1313.0/65536.0,1,-nbitq), 
to_sfixed(-1197.0/65536.0,1,-nbitq), 
to_sfixed(2302.0/65536.0,1,-nbitq), 
to_sfixed(-158.0/65536.0,1,-nbitq), 
to_sfixed(2964.0/65536.0,1,-nbitq), 
to_sfixed(-4293.0/65536.0,1,-nbitq), 
to_sfixed(4048.0/65536.0,1,-nbitq), 
to_sfixed(2289.0/65536.0,1,-nbitq), 
to_sfixed(7010.0/65536.0,1,-nbitq), 
to_sfixed(-3890.0/65536.0,1,-nbitq), 
to_sfixed(-2635.0/65536.0,1,-nbitq), 
to_sfixed(-2897.0/65536.0,1,-nbitq), 
to_sfixed(3224.0/65536.0,1,-nbitq), 
to_sfixed(-71.0/65536.0,1,-nbitq), 
to_sfixed(-2011.0/65536.0,1,-nbitq), 
to_sfixed(4403.0/65536.0,1,-nbitq), 
to_sfixed(-1832.0/65536.0,1,-nbitq), 
to_sfixed(1312.0/65536.0,1,-nbitq), 
to_sfixed(-2202.0/65536.0,1,-nbitq), 
to_sfixed(798.0/65536.0,1,-nbitq), 
to_sfixed(-3693.0/65536.0,1,-nbitq), 
to_sfixed(-2798.0/65536.0,1,-nbitq), 
to_sfixed(-1156.0/65536.0,1,-nbitq), 
to_sfixed(-2652.0/65536.0,1,-nbitq), 
to_sfixed(2153.0/65536.0,1,-nbitq), 
to_sfixed(-6118.0/65536.0,1,-nbitq), 
to_sfixed(110.0/65536.0,1,-nbitq), 
to_sfixed(-1045.0/65536.0,1,-nbitq), 
to_sfixed(1223.0/65536.0,1,-nbitq), 
to_sfixed(2365.0/65536.0,1,-nbitq), 
to_sfixed(-3824.0/65536.0,1,-nbitq), 
to_sfixed(-2030.0/65536.0,1,-nbitq), 
to_sfixed(1583.0/65536.0,1,-nbitq), 
to_sfixed(-7207.0/65536.0,1,-nbitq), 
to_sfixed(5629.0/65536.0,1,-nbitq), 
to_sfixed(755.0/65536.0,1,-nbitq), 
to_sfixed(1676.0/65536.0,1,-nbitq), 
to_sfixed(822.0/65536.0,1,-nbitq), 
to_sfixed(-680.0/65536.0,1,-nbitq), 
to_sfixed(562.0/65536.0,1,-nbitq), 
to_sfixed(720.0/65536.0,1,-nbitq), 
to_sfixed(1935.0/65536.0,1,-nbitq), 
to_sfixed(-981.0/65536.0,1,-nbitq), 
to_sfixed(-1232.0/65536.0,1,-nbitq), 
to_sfixed(-363.0/65536.0,1,-nbitq), 
to_sfixed(-1362.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2722.0/65536.0,1,-nbitq), 
to_sfixed(3622.0/65536.0,1,-nbitq), 
to_sfixed(3875.0/65536.0,1,-nbitq), 
to_sfixed(2605.0/65536.0,1,-nbitq), 
to_sfixed(3792.0/65536.0,1,-nbitq), 
to_sfixed(-5991.0/65536.0,1,-nbitq), 
to_sfixed(-1307.0/65536.0,1,-nbitq), 
to_sfixed(-392.0/65536.0,1,-nbitq), 
to_sfixed(-276.0/65536.0,1,-nbitq), 
to_sfixed(-2215.0/65536.0,1,-nbitq), 
to_sfixed(-1494.0/65536.0,1,-nbitq), 
to_sfixed(-8492.0/65536.0,1,-nbitq), 
to_sfixed(1405.0/65536.0,1,-nbitq), 
to_sfixed(786.0/65536.0,1,-nbitq), 
to_sfixed(-3002.0/65536.0,1,-nbitq), 
to_sfixed(-344.0/65536.0,1,-nbitq), 
to_sfixed(-898.0/65536.0,1,-nbitq), 
to_sfixed(-1043.0/65536.0,1,-nbitq), 
to_sfixed(-8565.0/65536.0,1,-nbitq), 
to_sfixed(1003.0/65536.0,1,-nbitq), 
to_sfixed(6420.0/65536.0,1,-nbitq), 
to_sfixed(1766.0/65536.0,1,-nbitq), 
to_sfixed(176.0/65536.0,1,-nbitq), 
to_sfixed(-12090.0/65536.0,1,-nbitq), 
to_sfixed(347.0/65536.0,1,-nbitq), 
to_sfixed(-14610.0/65536.0,1,-nbitq), 
to_sfixed(-6171.0/65536.0,1,-nbitq), 
to_sfixed(-2003.0/65536.0,1,-nbitq), 
to_sfixed(-1092.0/65536.0,1,-nbitq), 
to_sfixed(-2800.0/65536.0,1,-nbitq), 
to_sfixed(2394.0/65536.0,1,-nbitq), 
to_sfixed(216.0/65536.0,1,-nbitq), 
to_sfixed(671.0/65536.0,1,-nbitq), 
to_sfixed(3656.0/65536.0,1,-nbitq), 
to_sfixed(-1840.0/65536.0,1,-nbitq), 
to_sfixed(-201.0/65536.0,1,-nbitq), 
to_sfixed(791.0/65536.0,1,-nbitq), 
to_sfixed(2497.0/65536.0,1,-nbitq), 
to_sfixed(3698.0/65536.0,1,-nbitq), 
to_sfixed(-2170.0/65536.0,1,-nbitq), 
to_sfixed(5770.0/65536.0,1,-nbitq), 
to_sfixed(-1946.0/65536.0,1,-nbitq), 
to_sfixed(1658.0/65536.0,1,-nbitq), 
to_sfixed(-3297.0/65536.0,1,-nbitq), 
to_sfixed(-1414.0/65536.0,1,-nbitq), 
to_sfixed(-2105.0/65536.0,1,-nbitq), 
to_sfixed(3635.0/65536.0,1,-nbitq), 
to_sfixed(-1966.0/65536.0,1,-nbitq), 
to_sfixed(-2684.0/65536.0,1,-nbitq), 
to_sfixed(4148.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(294.0/65536.0,1,-nbitq), 
to_sfixed(-2061.0/65536.0,1,-nbitq), 
to_sfixed(5405.0/65536.0,1,-nbitq), 
to_sfixed(-3140.0/65536.0,1,-nbitq), 
to_sfixed(-3411.0/65536.0,1,-nbitq), 
to_sfixed(-558.0/65536.0,1,-nbitq), 
to_sfixed(-3147.0/65536.0,1,-nbitq), 
to_sfixed(320.0/65536.0,1,-nbitq), 
to_sfixed(-3516.0/65536.0,1,-nbitq), 
to_sfixed(-3513.0/65536.0,1,-nbitq), 
to_sfixed(-1125.0/65536.0,1,-nbitq), 
to_sfixed(-1243.0/65536.0,1,-nbitq), 
to_sfixed(2206.0/65536.0,1,-nbitq), 
to_sfixed(-475.0/65536.0,1,-nbitq), 
to_sfixed(-485.0/65536.0,1,-nbitq), 
to_sfixed(4662.0/65536.0,1,-nbitq), 
to_sfixed(-2692.0/65536.0,1,-nbitq), 
to_sfixed(7259.0/65536.0,1,-nbitq), 
to_sfixed(-747.0/65536.0,1,-nbitq), 
to_sfixed(1400.0/65536.0,1,-nbitq), 
to_sfixed(607.0/65536.0,1,-nbitq), 
to_sfixed(-2232.0/65536.0,1,-nbitq), 
to_sfixed(1981.0/65536.0,1,-nbitq), 
to_sfixed(-1559.0/65536.0,1,-nbitq), 
to_sfixed(-1691.0/65536.0,1,-nbitq), 
to_sfixed(223.0/65536.0,1,-nbitq), 
to_sfixed(962.0/65536.0,1,-nbitq), 
to_sfixed(2218.0/65536.0,1,-nbitq), 
to_sfixed(-3110.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1905.0/65536.0,1,-nbitq), 
to_sfixed(-2018.0/65536.0,1,-nbitq), 
to_sfixed(-1540.0/65536.0,1,-nbitq), 
to_sfixed(-838.0/65536.0,1,-nbitq), 
to_sfixed(-582.0/65536.0,1,-nbitq), 
to_sfixed(-1420.0/65536.0,1,-nbitq), 
to_sfixed(-3262.0/65536.0,1,-nbitq), 
to_sfixed(2642.0/65536.0,1,-nbitq), 
to_sfixed(-6634.0/65536.0,1,-nbitq), 
to_sfixed(-2089.0/65536.0,1,-nbitq), 
to_sfixed(-1424.0/65536.0,1,-nbitq), 
to_sfixed(-13556.0/65536.0,1,-nbitq), 
to_sfixed(979.0/65536.0,1,-nbitq), 
to_sfixed(-2703.0/65536.0,1,-nbitq), 
to_sfixed(-2897.0/65536.0,1,-nbitq), 
to_sfixed(-2798.0/65536.0,1,-nbitq), 
to_sfixed(1499.0/65536.0,1,-nbitq), 
to_sfixed(6986.0/65536.0,1,-nbitq), 
to_sfixed(-7404.0/65536.0,1,-nbitq), 
to_sfixed(1594.0/65536.0,1,-nbitq), 
to_sfixed(7079.0/65536.0,1,-nbitq), 
to_sfixed(-1838.0/65536.0,1,-nbitq), 
to_sfixed(-4036.0/65536.0,1,-nbitq), 
to_sfixed(-14621.0/65536.0,1,-nbitq), 
to_sfixed(1895.0/65536.0,1,-nbitq), 
to_sfixed(-16146.0/65536.0,1,-nbitq), 
to_sfixed(-3547.0/65536.0,1,-nbitq), 
to_sfixed(-2720.0/65536.0,1,-nbitq), 
to_sfixed(-3915.0/65536.0,1,-nbitq), 
to_sfixed(-3786.0/65536.0,1,-nbitq), 
to_sfixed(-4195.0/65536.0,1,-nbitq), 
to_sfixed(-637.0/65536.0,1,-nbitq), 
to_sfixed(4121.0/65536.0,1,-nbitq), 
to_sfixed(652.0/65536.0,1,-nbitq), 
to_sfixed(230.0/65536.0,1,-nbitq), 
to_sfixed(-1035.0/65536.0,1,-nbitq), 
to_sfixed(4828.0/65536.0,1,-nbitq), 
to_sfixed(3232.0/65536.0,1,-nbitq), 
to_sfixed(3428.0/65536.0,1,-nbitq), 
to_sfixed(-1110.0/65536.0,1,-nbitq), 
to_sfixed(3862.0/65536.0,1,-nbitq), 
to_sfixed(-866.0/65536.0,1,-nbitq), 
to_sfixed(9737.0/65536.0,1,-nbitq), 
to_sfixed(453.0/65536.0,1,-nbitq), 
to_sfixed(1545.0/65536.0,1,-nbitq), 
to_sfixed(-7660.0/65536.0,1,-nbitq), 
to_sfixed(-2371.0/65536.0,1,-nbitq), 
to_sfixed(-3123.0/65536.0,1,-nbitq), 
to_sfixed(160.0/65536.0,1,-nbitq), 
to_sfixed(5126.0/65536.0,1,-nbitq), 
to_sfixed(-639.0/65536.0,1,-nbitq), 
to_sfixed(-933.0/65536.0,1,-nbitq), 
to_sfixed(-3385.0/65536.0,1,-nbitq), 
to_sfixed(-846.0/65536.0,1,-nbitq), 
to_sfixed(251.0/65536.0,1,-nbitq), 
to_sfixed(-490.0/65536.0,1,-nbitq), 
to_sfixed(2754.0/65536.0,1,-nbitq), 
to_sfixed(-5534.0/65536.0,1,-nbitq), 
to_sfixed(946.0/65536.0,1,-nbitq), 
to_sfixed(-8743.0/65536.0,1,-nbitq), 
to_sfixed(1568.0/65536.0,1,-nbitq), 
to_sfixed(-2941.0/65536.0,1,-nbitq), 
to_sfixed(2113.0/65536.0,1,-nbitq), 
to_sfixed(2022.0/65536.0,1,-nbitq), 
to_sfixed(-893.0/65536.0,1,-nbitq), 
to_sfixed(8513.0/65536.0,1,-nbitq), 
to_sfixed(4004.0/65536.0,1,-nbitq), 
to_sfixed(-2277.0/65536.0,1,-nbitq), 
to_sfixed(3382.0/65536.0,1,-nbitq), 
to_sfixed(-2936.0/65536.0,1,-nbitq), 
to_sfixed(-3222.0/65536.0,1,-nbitq), 
to_sfixed(-2274.0/65536.0,1,-nbitq), 
to_sfixed(-2423.0/65536.0,1,-nbitq), 
to_sfixed(-1940.0/65536.0,1,-nbitq), 
to_sfixed(-1029.0/65536.0,1,-nbitq), 
to_sfixed(-178.0/65536.0,1,-nbitq), 
to_sfixed(3147.0/65536.0,1,-nbitq), 
to_sfixed(1135.0/65536.0,1,-nbitq), 
to_sfixed(448.0/65536.0,1,-nbitq), 
to_sfixed(-5611.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-38.0/65536.0,1,-nbitq), 
to_sfixed(-1055.0/65536.0,1,-nbitq), 
to_sfixed(1075.0/65536.0,1,-nbitq), 
to_sfixed(-947.0/65536.0,1,-nbitq), 
to_sfixed(2989.0/65536.0,1,-nbitq), 
to_sfixed(906.0/65536.0,1,-nbitq), 
to_sfixed(-5028.0/65536.0,1,-nbitq), 
to_sfixed(-468.0/65536.0,1,-nbitq), 
to_sfixed(3818.0/65536.0,1,-nbitq), 
to_sfixed(-1925.0/65536.0,1,-nbitq), 
to_sfixed(-502.0/65536.0,1,-nbitq), 
to_sfixed(-7473.0/65536.0,1,-nbitq), 
to_sfixed(-2638.0/65536.0,1,-nbitq), 
to_sfixed(-610.0/65536.0,1,-nbitq), 
to_sfixed(-94.0/65536.0,1,-nbitq), 
to_sfixed(2273.0/65536.0,1,-nbitq), 
to_sfixed(381.0/65536.0,1,-nbitq), 
to_sfixed(7031.0/65536.0,1,-nbitq), 
to_sfixed(-4808.0/65536.0,1,-nbitq), 
to_sfixed(2333.0/65536.0,1,-nbitq), 
to_sfixed(9268.0/65536.0,1,-nbitq), 
to_sfixed(2558.0/65536.0,1,-nbitq), 
to_sfixed(-170.0/65536.0,1,-nbitq), 
to_sfixed(-10301.0/65536.0,1,-nbitq), 
to_sfixed(960.0/65536.0,1,-nbitq), 
to_sfixed(-14946.0/65536.0,1,-nbitq), 
to_sfixed(5785.0/65536.0,1,-nbitq), 
to_sfixed(-2180.0/65536.0,1,-nbitq), 
to_sfixed(-76.0/65536.0,1,-nbitq), 
to_sfixed(1991.0/65536.0,1,-nbitq), 
to_sfixed(-4018.0/65536.0,1,-nbitq), 
to_sfixed(184.0/65536.0,1,-nbitq), 
to_sfixed(6052.0/65536.0,1,-nbitq), 
to_sfixed(3635.0/65536.0,1,-nbitq), 
to_sfixed(2823.0/65536.0,1,-nbitq), 
to_sfixed(-1320.0/65536.0,1,-nbitq), 
to_sfixed(631.0/65536.0,1,-nbitq), 
to_sfixed(-458.0/65536.0,1,-nbitq), 
to_sfixed(5646.0/65536.0,1,-nbitq), 
to_sfixed(807.0/65536.0,1,-nbitq), 
to_sfixed(354.0/65536.0,1,-nbitq), 
to_sfixed(-32.0/65536.0,1,-nbitq), 
to_sfixed(9519.0/65536.0,1,-nbitq), 
to_sfixed(-4622.0/65536.0,1,-nbitq), 
to_sfixed(-1417.0/65536.0,1,-nbitq), 
to_sfixed(-7156.0/65536.0,1,-nbitq), 
to_sfixed(-1631.0/65536.0,1,-nbitq), 
to_sfixed(1335.0/65536.0,1,-nbitq), 
to_sfixed(-884.0/65536.0,1,-nbitq), 
to_sfixed(5305.0/65536.0,1,-nbitq), 
to_sfixed(2105.0/65536.0,1,-nbitq), 
to_sfixed(-3036.0/65536.0,1,-nbitq), 
to_sfixed(-3674.0/65536.0,1,-nbitq), 
to_sfixed(-10394.0/65536.0,1,-nbitq), 
to_sfixed(-1012.0/65536.0,1,-nbitq), 
to_sfixed(-5892.0/65536.0,1,-nbitq), 
to_sfixed(2764.0/65536.0,1,-nbitq), 
to_sfixed(-2970.0/65536.0,1,-nbitq), 
to_sfixed(-2711.0/65536.0,1,-nbitq), 
to_sfixed(-6848.0/65536.0,1,-nbitq), 
to_sfixed(6339.0/65536.0,1,-nbitq), 
to_sfixed(-2991.0/65536.0,1,-nbitq), 
to_sfixed(-469.0/65536.0,1,-nbitq), 
to_sfixed(-5.0/65536.0,1,-nbitq), 
to_sfixed(-2525.0/65536.0,1,-nbitq), 
to_sfixed(7622.0/65536.0,1,-nbitq), 
to_sfixed(6464.0/65536.0,1,-nbitq), 
to_sfixed(-4211.0/65536.0,1,-nbitq), 
to_sfixed(-2964.0/65536.0,1,-nbitq), 
to_sfixed(647.0/65536.0,1,-nbitq), 
to_sfixed(-2196.0/65536.0,1,-nbitq), 
to_sfixed(-10267.0/65536.0,1,-nbitq), 
to_sfixed(-2032.0/65536.0,1,-nbitq), 
to_sfixed(-971.0/65536.0,1,-nbitq), 
to_sfixed(-1808.0/65536.0,1,-nbitq), 
to_sfixed(8257.0/65536.0,1,-nbitq), 
to_sfixed(6591.0/65536.0,1,-nbitq), 
to_sfixed(990.0/65536.0,1,-nbitq), 
to_sfixed(-259.0/65536.0,1,-nbitq), 
to_sfixed(-6473.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2330.0/65536.0,1,-nbitq), 
to_sfixed(1270.0/65536.0,1,-nbitq), 
to_sfixed(3019.0/65536.0,1,-nbitq), 
to_sfixed(-4672.0/65536.0,1,-nbitq), 
to_sfixed(1006.0/65536.0,1,-nbitq), 
to_sfixed(-5453.0/65536.0,1,-nbitq), 
to_sfixed(-9709.0/65536.0,1,-nbitq), 
to_sfixed(-5445.0/65536.0,1,-nbitq), 
to_sfixed(-2692.0/65536.0,1,-nbitq), 
to_sfixed(2795.0/65536.0,1,-nbitq), 
to_sfixed(3648.0/65536.0,1,-nbitq), 
to_sfixed(-14451.0/65536.0,1,-nbitq), 
to_sfixed(-952.0/65536.0,1,-nbitq), 
to_sfixed(-3344.0/65536.0,1,-nbitq), 
to_sfixed(-570.0/65536.0,1,-nbitq), 
to_sfixed(3545.0/65536.0,1,-nbitq), 
to_sfixed(-2598.0/65536.0,1,-nbitq), 
to_sfixed(4676.0/65536.0,1,-nbitq), 
to_sfixed(419.0/65536.0,1,-nbitq), 
to_sfixed(-1065.0/65536.0,1,-nbitq), 
to_sfixed(4595.0/65536.0,1,-nbitq), 
to_sfixed(6714.0/65536.0,1,-nbitq), 
to_sfixed(-1064.0/65536.0,1,-nbitq), 
to_sfixed(-11630.0/65536.0,1,-nbitq), 
to_sfixed(2139.0/65536.0,1,-nbitq), 
to_sfixed(-14308.0/65536.0,1,-nbitq), 
to_sfixed(52.0/65536.0,1,-nbitq), 
to_sfixed(-1367.0/65536.0,1,-nbitq), 
to_sfixed(-763.0/65536.0,1,-nbitq), 
to_sfixed(564.0/65536.0,1,-nbitq), 
to_sfixed(-837.0/65536.0,1,-nbitq), 
to_sfixed(-1680.0/65536.0,1,-nbitq), 
to_sfixed(6464.0/65536.0,1,-nbitq), 
to_sfixed(-261.0/65536.0,1,-nbitq), 
to_sfixed(-762.0/65536.0,1,-nbitq), 
to_sfixed(1292.0/65536.0,1,-nbitq), 
to_sfixed(2453.0/65536.0,1,-nbitq), 
to_sfixed(338.0/65536.0,1,-nbitq), 
to_sfixed(2562.0/65536.0,1,-nbitq), 
to_sfixed(-1484.0/65536.0,1,-nbitq), 
to_sfixed(-1084.0/65536.0,1,-nbitq), 
to_sfixed(-3123.0/65536.0,1,-nbitq), 
to_sfixed(-177.0/65536.0,1,-nbitq), 
to_sfixed(-3204.0/65536.0,1,-nbitq), 
to_sfixed(724.0/65536.0,1,-nbitq), 
to_sfixed(-4097.0/65536.0,1,-nbitq), 
to_sfixed(-59.0/65536.0,1,-nbitq), 
to_sfixed(1302.0/65536.0,1,-nbitq), 
to_sfixed(1201.0/65536.0,1,-nbitq), 
to_sfixed(-440.0/65536.0,1,-nbitq), 
to_sfixed(262.0/65536.0,1,-nbitq), 
to_sfixed(832.0/65536.0,1,-nbitq), 
to_sfixed(-4903.0/65536.0,1,-nbitq), 
to_sfixed(-14795.0/65536.0,1,-nbitq), 
to_sfixed(-4445.0/65536.0,1,-nbitq), 
to_sfixed(-1923.0/65536.0,1,-nbitq), 
to_sfixed(-1216.0/65536.0,1,-nbitq), 
to_sfixed(-59.0/65536.0,1,-nbitq), 
to_sfixed(-1298.0/65536.0,1,-nbitq), 
to_sfixed(-3982.0/65536.0,1,-nbitq), 
to_sfixed(9628.0/65536.0,1,-nbitq), 
to_sfixed(-1973.0/65536.0,1,-nbitq), 
to_sfixed(-2642.0/65536.0,1,-nbitq), 
to_sfixed(-1705.0/65536.0,1,-nbitq), 
to_sfixed(-827.0/65536.0,1,-nbitq), 
to_sfixed(5146.0/65536.0,1,-nbitq), 
to_sfixed(3214.0/65536.0,1,-nbitq), 
to_sfixed(1057.0/65536.0,1,-nbitq), 
to_sfixed(-401.0/65536.0,1,-nbitq), 
to_sfixed(-6478.0/65536.0,1,-nbitq), 
to_sfixed(-2466.0/65536.0,1,-nbitq), 
to_sfixed(-8888.0/65536.0,1,-nbitq), 
to_sfixed(-2312.0/65536.0,1,-nbitq), 
to_sfixed(1140.0/65536.0,1,-nbitq), 
to_sfixed(2281.0/65536.0,1,-nbitq), 
to_sfixed(-1939.0/65536.0,1,-nbitq), 
to_sfixed(9227.0/65536.0,1,-nbitq), 
to_sfixed(-64.0/65536.0,1,-nbitq), 
to_sfixed(1913.0/65536.0,1,-nbitq), 
to_sfixed(-7731.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-834.0/65536.0,1,-nbitq), 
to_sfixed(-2008.0/65536.0,1,-nbitq), 
to_sfixed(-7670.0/65536.0,1,-nbitq), 
to_sfixed(-10107.0/65536.0,1,-nbitq), 
to_sfixed(7695.0/65536.0,1,-nbitq), 
to_sfixed(-5421.0/65536.0,1,-nbitq), 
to_sfixed(-8693.0/65536.0,1,-nbitq), 
to_sfixed(-3615.0/65536.0,1,-nbitq), 
to_sfixed(-3303.0/65536.0,1,-nbitq), 
to_sfixed(-117.0/65536.0,1,-nbitq), 
to_sfixed(4439.0/65536.0,1,-nbitq), 
to_sfixed(-14015.0/65536.0,1,-nbitq), 
to_sfixed(3025.0/65536.0,1,-nbitq), 
to_sfixed(-2615.0/65536.0,1,-nbitq), 
to_sfixed(-2555.0/65536.0,1,-nbitq), 
to_sfixed(840.0/65536.0,1,-nbitq), 
to_sfixed(2095.0/65536.0,1,-nbitq), 
to_sfixed(-2234.0/65536.0,1,-nbitq), 
to_sfixed(4198.0/65536.0,1,-nbitq), 
to_sfixed(1219.0/65536.0,1,-nbitq), 
to_sfixed(637.0/65536.0,1,-nbitq), 
to_sfixed(9229.0/65536.0,1,-nbitq), 
to_sfixed(2038.0/65536.0,1,-nbitq), 
to_sfixed(-3914.0/65536.0,1,-nbitq), 
to_sfixed(-907.0/65536.0,1,-nbitq), 
to_sfixed(-9962.0/65536.0,1,-nbitq), 
to_sfixed(168.0/65536.0,1,-nbitq), 
to_sfixed(-1834.0/65536.0,1,-nbitq), 
to_sfixed(-10357.0/65536.0,1,-nbitq), 
to_sfixed(4264.0/65536.0,1,-nbitq), 
to_sfixed(1729.0/65536.0,1,-nbitq), 
to_sfixed(-1076.0/65536.0,1,-nbitq), 
to_sfixed(1745.0/65536.0,1,-nbitq), 
to_sfixed(-4384.0/65536.0,1,-nbitq), 
to_sfixed(-1831.0/65536.0,1,-nbitq), 
to_sfixed(2091.0/65536.0,1,-nbitq), 
to_sfixed(-428.0/65536.0,1,-nbitq), 
to_sfixed(-1483.0/65536.0,1,-nbitq), 
to_sfixed(6241.0/65536.0,1,-nbitq), 
to_sfixed(4037.0/65536.0,1,-nbitq), 
to_sfixed(2975.0/65536.0,1,-nbitq), 
to_sfixed(197.0/65536.0,1,-nbitq), 
to_sfixed(-11468.0/65536.0,1,-nbitq), 
to_sfixed(-3535.0/65536.0,1,-nbitq), 
to_sfixed(1337.0/65536.0,1,-nbitq), 
to_sfixed(-410.0/65536.0,1,-nbitq), 
to_sfixed(-1032.0/65536.0,1,-nbitq), 
to_sfixed(6555.0/65536.0,1,-nbitq), 
to_sfixed(-700.0/65536.0,1,-nbitq), 
to_sfixed(-235.0/65536.0,1,-nbitq), 
to_sfixed(-821.0/65536.0,1,-nbitq), 
to_sfixed(-1638.0/65536.0,1,-nbitq), 
to_sfixed(-2143.0/65536.0,1,-nbitq), 
to_sfixed(-10411.0/65536.0,1,-nbitq), 
to_sfixed(-3000.0/65536.0,1,-nbitq), 
to_sfixed(-4236.0/65536.0,1,-nbitq), 
to_sfixed(-1961.0/65536.0,1,-nbitq), 
to_sfixed(2380.0/65536.0,1,-nbitq), 
to_sfixed(-1320.0/65536.0,1,-nbitq), 
to_sfixed(3405.0/65536.0,1,-nbitq), 
to_sfixed(2440.0/65536.0,1,-nbitq), 
to_sfixed(757.0/65536.0,1,-nbitq), 
to_sfixed(-1685.0/65536.0,1,-nbitq), 
to_sfixed(-1083.0/65536.0,1,-nbitq), 
to_sfixed(3198.0/65536.0,1,-nbitq), 
to_sfixed(5679.0/65536.0,1,-nbitq), 
to_sfixed(4183.0/65536.0,1,-nbitq), 
to_sfixed(4322.0/65536.0,1,-nbitq), 
to_sfixed(-2188.0/65536.0,1,-nbitq), 
to_sfixed(-10362.0/65536.0,1,-nbitq), 
to_sfixed(-3597.0/65536.0,1,-nbitq), 
to_sfixed(-1112.0/65536.0,1,-nbitq), 
to_sfixed(-3851.0/65536.0,1,-nbitq), 
to_sfixed(-26.0/65536.0,1,-nbitq), 
to_sfixed(-1432.0/65536.0,1,-nbitq), 
to_sfixed(-2869.0/65536.0,1,-nbitq), 
to_sfixed(10991.0/65536.0,1,-nbitq), 
to_sfixed(2387.0/65536.0,1,-nbitq), 
to_sfixed(-304.0/65536.0,1,-nbitq), 
to_sfixed(-3773.0/65536.0,1,-nbitq)  ), 
( to_sfixed(366.0/65536.0,1,-nbitq), 
to_sfixed(902.0/65536.0,1,-nbitq), 
to_sfixed(-15905.0/65536.0,1,-nbitq), 
to_sfixed(-7474.0/65536.0,1,-nbitq), 
to_sfixed(-279.0/65536.0,1,-nbitq), 
to_sfixed(-4677.0/65536.0,1,-nbitq), 
to_sfixed(-2830.0/65536.0,1,-nbitq), 
to_sfixed(-1698.0/65536.0,1,-nbitq), 
to_sfixed(423.0/65536.0,1,-nbitq), 
to_sfixed(-1462.0/65536.0,1,-nbitq), 
to_sfixed(-1469.0/65536.0,1,-nbitq), 
to_sfixed(3100.0/65536.0,1,-nbitq), 
to_sfixed(403.0/65536.0,1,-nbitq), 
to_sfixed(4874.0/65536.0,1,-nbitq), 
to_sfixed(2562.0/65536.0,1,-nbitq), 
to_sfixed(2781.0/65536.0,1,-nbitq), 
to_sfixed(1576.0/65536.0,1,-nbitq), 
to_sfixed(-10861.0/65536.0,1,-nbitq), 
to_sfixed(5173.0/65536.0,1,-nbitq), 
to_sfixed(-502.0/65536.0,1,-nbitq), 
to_sfixed(-4747.0/65536.0,1,-nbitq), 
to_sfixed(6951.0/65536.0,1,-nbitq), 
to_sfixed(7152.0/65536.0,1,-nbitq), 
to_sfixed(-403.0/65536.0,1,-nbitq), 
to_sfixed(1837.0/65536.0,1,-nbitq), 
to_sfixed(-6769.0/65536.0,1,-nbitq), 
to_sfixed(5440.0/65536.0,1,-nbitq), 
to_sfixed(-1518.0/65536.0,1,-nbitq), 
to_sfixed(-12608.0/65536.0,1,-nbitq), 
to_sfixed(9776.0/65536.0,1,-nbitq), 
to_sfixed(4938.0/65536.0,1,-nbitq), 
to_sfixed(2602.0/65536.0,1,-nbitq), 
to_sfixed(-15.0/65536.0,1,-nbitq), 
to_sfixed(-6982.0/65536.0,1,-nbitq), 
to_sfixed(-2683.0/65536.0,1,-nbitq), 
to_sfixed(-1412.0/65536.0,1,-nbitq), 
to_sfixed(-1112.0/65536.0,1,-nbitq), 
to_sfixed(1771.0/65536.0,1,-nbitq), 
to_sfixed(3430.0/65536.0,1,-nbitq), 
to_sfixed(-871.0/65536.0,1,-nbitq), 
to_sfixed(-275.0/65536.0,1,-nbitq), 
to_sfixed(813.0/65536.0,1,-nbitq), 
to_sfixed(-7987.0/65536.0,1,-nbitq), 
to_sfixed(-3046.0/65536.0,1,-nbitq), 
to_sfixed(414.0/65536.0,1,-nbitq), 
to_sfixed(5018.0/65536.0,1,-nbitq), 
to_sfixed(1144.0/65536.0,1,-nbitq), 
to_sfixed(10378.0/65536.0,1,-nbitq), 
to_sfixed(2781.0/65536.0,1,-nbitq), 
to_sfixed(-524.0/65536.0,1,-nbitq), 
to_sfixed(887.0/65536.0,1,-nbitq), 
to_sfixed(-2219.0/65536.0,1,-nbitq), 
to_sfixed(-1508.0/65536.0,1,-nbitq), 
to_sfixed(512.0/65536.0,1,-nbitq), 
to_sfixed(1463.0/65536.0,1,-nbitq), 
to_sfixed(-5138.0/65536.0,1,-nbitq), 
to_sfixed(-1788.0/65536.0,1,-nbitq), 
to_sfixed(4291.0/65536.0,1,-nbitq), 
to_sfixed(2262.0/65536.0,1,-nbitq), 
to_sfixed(6409.0/65536.0,1,-nbitq), 
to_sfixed(74.0/65536.0,1,-nbitq), 
to_sfixed(-2096.0/65536.0,1,-nbitq), 
to_sfixed(-2787.0/65536.0,1,-nbitq), 
to_sfixed(2526.0/65536.0,1,-nbitq), 
to_sfixed(368.0/65536.0,1,-nbitq), 
to_sfixed(7851.0/65536.0,1,-nbitq), 
to_sfixed(2671.0/65536.0,1,-nbitq), 
to_sfixed(-881.0/65536.0,1,-nbitq), 
to_sfixed(-7413.0/65536.0,1,-nbitq), 
to_sfixed(-5152.0/65536.0,1,-nbitq), 
to_sfixed(-3728.0/65536.0,1,-nbitq), 
to_sfixed(-3067.0/65536.0,1,-nbitq), 
to_sfixed(-5888.0/65536.0,1,-nbitq), 
to_sfixed(1230.0/65536.0,1,-nbitq), 
to_sfixed(-2083.0/65536.0,1,-nbitq), 
to_sfixed(-2420.0/65536.0,1,-nbitq), 
to_sfixed(2087.0/65536.0,1,-nbitq), 
to_sfixed(2300.0/65536.0,1,-nbitq), 
to_sfixed(-2372.0/65536.0,1,-nbitq), 
to_sfixed(-3865.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1216.0/65536.0,1,-nbitq), 
to_sfixed(-1848.0/65536.0,1,-nbitq), 
to_sfixed(-13710.0/65536.0,1,-nbitq), 
to_sfixed(-8061.0/65536.0,1,-nbitq), 
to_sfixed(-365.0/65536.0,1,-nbitq), 
to_sfixed(-6434.0/65536.0,1,-nbitq), 
to_sfixed(-1346.0/65536.0,1,-nbitq), 
to_sfixed(-2344.0/65536.0,1,-nbitq), 
to_sfixed(338.0/65536.0,1,-nbitq), 
to_sfixed(2441.0/65536.0,1,-nbitq), 
to_sfixed(2846.0/65536.0,1,-nbitq), 
to_sfixed(-3882.0/65536.0,1,-nbitq), 
to_sfixed(2507.0/65536.0,1,-nbitq), 
to_sfixed(4771.0/65536.0,1,-nbitq), 
to_sfixed(-2545.0/65536.0,1,-nbitq), 
to_sfixed(939.0/65536.0,1,-nbitq), 
to_sfixed(2435.0/65536.0,1,-nbitq), 
to_sfixed(-9652.0/65536.0,1,-nbitq), 
to_sfixed(4336.0/65536.0,1,-nbitq), 
to_sfixed(-6.0/65536.0,1,-nbitq), 
to_sfixed(-5816.0/65536.0,1,-nbitq), 
to_sfixed(1967.0/65536.0,1,-nbitq), 
to_sfixed(7396.0/65536.0,1,-nbitq), 
to_sfixed(-1017.0/65536.0,1,-nbitq), 
to_sfixed(3294.0/65536.0,1,-nbitq), 
to_sfixed(-3349.0/65536.0,1,-nbitq), 
to_sfixed(185.0/65536.0,1,-nbitq), 
to_sfixed(-3174.0/65536.0,1,-nbitq), 
to_sfixed(-10056.0/65536.0,1,-nbitq), 
to_sfixed(9880.0/65536.0,1,-nbitq), 
to_sfixed(6459.0/65536.0,1,-nbitq), 
to_sfixed(3856.0/65536.0,1,-nbitq), 
to_sfixed(-8111.0/65536.0,1,-nbitq), 
to_sfixed(-2003.0/65536.0,1,-nbitq), 
to_sfixed(-2168.0/65536.0,1,-nbitq), 
to_sfixed(2919.0/65536.0,1,-nbitq), 
to_sfixed(521.0/65536.0,1,-nbitq), 
to_sfixed(4649.0/65536.0,1,-nbitq), 
to_sfixed(6697.0/65536.0,1,-nbitq), 
to_sfixed(434.0/65536.0,1,-nbitq), 
to_sfixed(-6919.0/65536.0,1,-nbitq), 
to_sfixed(389.0/65536.0,1,-nbitq), 
to_sfixed(-7858.0/65536.0,1,-nbitq), 
to_sfixed(2227.0/65536.0,1,-nbitq), 
to_sfixed(-1479.0/65536.0,1,-nbitq), 
to_sfixed(-4689.0/65536.0,1,-nbitq), 
to_sfixed(-1137.0/65536.0,1,-nbitq), 
to_sfixed(6309.0/65536.0,1,-nbitq), 
to_sfixed(-143.0/65536.0,1,-nbitq), 
to_sfixed(-816.0/65536.0,1,-nbitq), 
to_sfixed(-610.0/65536.0,1,-nbitq), 
to_sfixed(819.0/65536.0,1,-nbitq), 
to_sfixed(2550.0/65536.0,1,-nbitq), 
to_sfixed(6584.0/65536.0,1,-nbitq), 
to_sfixed(4901.0/65536.0,1,-nbitq), 
to_sfixed(-3935.0/65536.0,1,-nbitq), 
to_sfixed(-1432.0/65536.0,1,-nbitq), 
to_sfixed(-1607.0/65536.0,1,-nbitq), 
to_sfixed(2226.0/65536.0,1,-nbitq), 
to_sfixed(-873.0/65536.0,1,-nbitq), 
to_sfixed(-3888.0/65536.0,1,-nbitq), 
to_sfixed(-2537.0/65536.0,1,-nbitq), 
to_sfixed(853.0/65536.0,1,-nbitq), 
to_sfixed(-1562.0/65536.0,1,-nbitq), 
to_sfixed(3886.0/65536.0,1,-nbitq), 
to_sfixed(12758.0/65536.0,1,-nbitq), 
to_sfixed(-5748.0/65536.0,1,-nbitq), 
to_sfixed(4198.0/65536.0,1,-nbitq), 
to_sfixed(-8046.0/65536.0,1,-nbitq), 
to_sfixed(-5769.0/65536.0,1,-nbitq), 
to_sfixed(801.0/65536.0,1,-nbitq), 
to_sfixed(577.0/65536.0,1,-nbitq), 
to_sfixed(-5406.0/65536.0,1,-nbitq), 
to_sfixed(-1384.0/65536.0,1,-nbitq), 
to_sfixed(-1369.0/65536.0,1,-nbitq), 
to_sfixed(-5444.0/65536.0,1,-nbitq), 
to_sfixed(9168.0/65536.0,1,-nbitq), 
to_sfixed(74.0/65536.0,1,-nbitq), 
to_sfixed(1758.0/65536.0,1,-nbitq), 
to_sfixed(-5395.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2925.0/65536.0,1,-nbitq), 
to_sfixed(-2186.0/65536.0,1,-nbitq), 
to_sfixed(5083.0/65536.0,1,-nbitq), 
to_sfixed(-1534.0/65536.0,1,-nbitq), 
to_sfixed(-2811.0/65536.0,1,-nbitq), 
to_sfixed(-941.0/65536.0,1,-nbitq), 
to_sfixed(2821.0/65536.0,1,-nbitq), 
to_sfixed(-3037.0/65536.0,1,-nbitq), 
to_sfixed(-5983.0/65536.0,1,-nbitq), 
to_sfixed(2868.0/65536.0,1,-nbitq), 
to_sfixed(47.0/65536.0,1,-nbitq), 
to_sfixed(-1757.0/65536.0,1,-nbitq), 
to_sfixed(3002.0/65536.0,1,-nbitq), 
to_sfixed(2692.0/65536.0,1,-nbitq), 
to_sfixed(-2602.0/65536.0,1,-nbitq), 
to_sfixed(-522.0/65536.0,1,-nbitq), 
to_sfixed(1192.0/65536.0,1,-nbitq), 
to_sfixed(-12444.0/65536.0,1,-nbitq), 
to_sfixed(3999.0/65536.0,1,-nbitq), 
to_sfixed(-265.0/65536.0,1,-nbitq), 
to_sfixed(-3292.0/65536.0,1,-nbitq), 
to_sfixed(2933.0/65536.0,1,-nbitq), 
to_sfixed(5216.0/65536.0,1,-nbitq), 
to_sfixed(-3521.0/65536.0,1,-nbitq), 
to_sfixed(2595.0/65536.0,1,-nbitq), 
to_sfixed(-3017.0/65536.0,1,-nbitq), 
to_sfixed(3196.0/65536.0,1,-nbitq), 
to_sfixed(-4287.0/65536.0,1,-nbitq), 
to_sfixed(-281.0/65536.0,1,-nbitq), 
to_sfixed(7381.0/65536.0,1,-nbitq), 
to_sfixed(3597.0/65536.0,1,-nbitq), 
to_sfixed(9065.0/65536.0,1,-nbitq), 
to_sfixed(-10125.0/65536.0,1,-nbitq), 
to_sfixed(-827.0/65536.0,1,-nbitq), 
to_sfixed(1810.0/65536.0,1,-nbitq), 
to_sfixed(249.0/65536.0,1,-nbitq), 
to_sfixed(-871.0/65536.0,1,-nbitq), 
to_sfixed(3860.0/65536.0,1,-nbitq), 
to_sfixed(9237.0/65536.0,1,-nbitq), 
to_sfixed(-2426.0/65536.0,1,-nbitq), 
to_sfixed(-3658.0/65536.0,1,-nbitq), 
to_sfixed(-2144.0/65536.0,1,-nbitq), 
to_sfixed(4068.0/65536.0,1,-nbitq), 
to_sfixed(12425.0/65536.0,1,-nbitq), 
to_sfixed(1060.0/65536.0,1,-nbitq), 
to_sfixed(2428.0/65536.0,1,-nbitq), 
to_sfixed(-337.0/65536.0,1,-nbitq), 
to_sfixed(5420.0/65536.0,1,-nbitq), 
to_sfixed(-602.0/65536.0,1,-nbitq), 
to_sfixed(3533.0/65536.0,1,-nbitq), 
to_sfixed(1590.0/65536.0,1,-nbitq), 
to_sfixed(553.0/65536.0,1,-nbitq), 
to_sfixed(3397.0/65536.0,1,-nbitq), 
to_sfixed(5339.0/65536.0,1,-nbitq), 
to_sfixed(1676.0/65536.0,1,-nbitq), 
to_sfixed(-853.0/65536.0,1,-nbitq), 
to_sfixed(-1628.0/65536.0,1,-nbitq), 
to_sfixed(-4144.0/65536.0,1,-nbitq), 
to_sfixed(-2276.0/65536.0,1,-nbitq), 
to_sfixed(-3553.0/65536.0,1,-nbitq), 
to_sfixed(-6139.0/65536.0,1,-nbitq), 
to_sfixed(1636.0/65536.0,1,-nbitq), 
to_sfixed(-28.0/65536.0,1,-nbitq), 
to_sfixed(855.0/65536.0,1,-nbitq), 
to_sfixed(4145.0/65536.0,1,-nbitq), 
to_sfixed(2038.0/65536.0,1,-nbitq), 
to_sfixed(-4720.0/65536.0,1,-nbitq), 
to_sfixed(9069.0/65536.0,1,-nbitq), 
to_sfixed(-7554.0/65536.0,1,-nbitq), 
to_sfixed(-6165.0/65536.0,1,-nbitq), 
to_sfixed(162.0/65536.0,1,-nbitq), 
to_sfixed(3918.0/65536.0,1,-nbitq), 
to_sfixed(-543.0/65536.0,1,-nbitq), 
to_sfixed(-271.0/65536.0,1,-nbitq), 
to_sfixed(-2624.0/65536.0,1,-nbitq), 
to_sfixed(-8990.0/65536.0,1,-nbitq), 
to_sfixed(11731.0/65536.0,1,-nbitq), 
to_sfixed(712.0/65536.0,1,-nbitq), 
to_sfixed(1074.0/65536.0,1,-nbitq), 
to_sfixed(118.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2186.0/65536.0,1,-nbitq), 
to_sfixed(-5838.0/65536.0,1,-nbitq), 
to_sfixed(7714.0/65536.0,1,-nbitq), 
to_sfixed(199.0/65536.0,1,-nbitq), 
to_sfixed(1169.0/65536.0,1,-nbitq), 
to_sfixed(-7239.0/65536.0,1,-nbitq), 
to_sfixed(3528.0/65536.0,1,-nbitq), 
to_sfixed(-564.0/65536.0,1,-nbitq), 
to_sfixed(1748.0/65536.0,1,-nbitq), 
to_sfixed(-1698.0/65536.0,1,-nbitq), 
to_sfixed(-384.0/65536.0,1,-nbitq), 
to_sfixed(8863.0/65536.0,1,-nbitq), 
to_sfixed(1316.0/65536.0,1,-nbitq), 
to_sfixed(4115.0/65536.0,1,-nbitq), 
to_sfixed(171.0/65536.0,1,-nbitq), 
to_sfixed(-2861.0/65536.0,1,-nbitq), 
to_sfixed(-1550.0/65536.0,1,-nbitq), 
to_sfixed(-5307.0/65536.0,1,-nbitq), 
to_sfixed(1133.0/65536.0,1,-nbitq), 
to_sfixed(2849.0/65536.0,1,-nbitq), 
to_sfixed(-784.0/65536.0,1,-nbitq), 
to_sfixed(10676.0/65536.0,1,-nbitq), 
to_sfixed(8876.0/65536.0,1,-nbitq), 
to_sfixed(-1709.0/65536.0,1,-nbitq), 
to_sfixed(2478.0/65536.0,1,-nbitq), 
to_sfixed(-1202.0/65536.0,1,-nbitq), 
to_sfixed(3495.0/65536.0,1,-nbitq), 
to_sfixed(-3716.0/65536.0,1,-nbitq), 
to_sfixed(-5867.0/65536.0,1,-nbitq), 
to_sfixed(946.0/65536.0,1,-nbitq), 
to_sfixed(1744.0/65536.0,1,-nbitq), 
to_sfixed(5721.0/65536.0,1,-nbitq), 
to_sfixed(-7438.0/65536.0,1,-nbitq), 
to_sfixed(13144.0/65536.0,1,-nbitq), 
to_sfixed(-2288.0/65536.0,1,-nbitq), 
to_sfixed(2686.0/65536.0,1,-nbitq), 
to_sfixed(-8244.0/65536.0,1,-nbitq), 
to_sfixed(3345.0/65536.0,1,-nbitq), 
to_sfixed(2873.0/65536.0,1,-nbitq), 
to_sfixed(-105.0/65536.0,1,-nbitq), 
to_sfixed(1460.0/65536.0,1,-nbitq), 
to_sfixed(-505.0/65536.0,1,-nbitq), 
to_sfixed(1801.0/65536.0,1,-nbitq), 
to_sfixed(4447.0/65536.0,1,-nbitq), 
to_sfixed(53.0/65536.0,1,-nbitq), 
to_sfixed(1512.0/65536.0,1,-nbitq), 
to_sfixed(676.0/65536.0,1,-nbitq), 
to_sfixed(9154.0/65536.0,1,-nbitq), 
to_sfixed(527.0/65536.0,1,-nbitq), 
to_sfixed(1906.0/65536.0,1,-nbitq), 
to_sfixed(-752.0/65536.0,1,-nbitq), 
to_sfixed(1044.0/65536.0,1,-nbitq), 
to_sfixed(314.0/65536.0,1,-nbitq), 
to_sfixed(5848.0/65536.0,1,-nbitq), 
to_sfixed(2180.0/65536.0,1,-nbitq), 
to_sfixed(-993.0/65536.0,1,-nbitq), 
to_sfixed(2473.0/65536.0,1,-nbitq), 
to_sfixed(-7734.0/65536.0,1,-nbitq), 
to_sfixed(-304.0/65536.0,1,-nbitq), 
to_sfixed(-3275.0/65536.0,1,-nbitq), 
to_sfixed(-1985.0/65536.0,1,-nbitq), 
to_sfixed(719.0/65536.0,1,-nbitq), 
to_sfixed(-2818.0/65536.0,1,-nbitq), 
to_sfixed(1407.0/65536.0,1,-nbitq), 
to_sfixed(-984.0/65536.0,1,-nbitq), 
to_sfixed(-2477.0/65536.0,1,-nbitq), 
to_sfixed(-4966.0/65536.0,1,-nbitq), 
to_sfixed(555.0/65536.0,1,-nbitq), 
to_sfixed(-14228.0/65536.0,1,-nbitq), 
to_sfixed(2435.0/65536.0,1,-nbitq), 
to_sfixed(-844.0/65536.0,1,-nbitq), 
to_sfixed(364.0/65536.0,1,-nbitq), 
to_sfixed(-1977.0/65536.0,1,-nbitq), 
to_sfixed(-809.0/65536.0,1,-nbitq), 
to_sfixed(-747.0/65536.0,1,-nbitq), 
to_sfixed(1848.0/65536.0,1,-nbitq), 
to_sfixed(5899.0/65536.0,1,-nbitq), 
to_sfixed(-4837.0/65536.0,1,-nbitq), 
to_sfixed(1518.0/65536.0,1,-nbitq), 
to_sfixed(2903.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1503.0/65536.0,1,-nbitq), 
to_sfixed(-4775.0/65536.0,1,-nbitq), 
to_sfixed(5536.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(2347.0/65536.0,1,-nbitq), 
to_sfixed(-5750.0/65536.0,1,-nbitq), 
to_sfixed(8246.0/65536.0,1,-nbitq), 
to_sfixed(1410.0/65536.0,1,-nbitq), 
to_sfixed(3171.0/65536.0,1,-nbitq), 
to_sfixed(-2356.0/65536.0,1,-nbitq), 
to_sfixed(1482.0/65536.0,1,-nbitq), 
to_sfixed(9877.0/65536.0,1,-nbitq), 
to_sfixed(2330.0/65536.0,1,-nbitq), 
to_sfixed(379.0/65536.0,1,-nbitq), 
to_sfixed(-3986.0/65536.0,1,-nbitq), 
to_sfixed(2515.0/65536.0,1,-nbitq), 
to_sfixed(722.0/65536.0,1,-nbitq), 
to_sfixed(-3197.0/65536.0,1,-nbitq), 
to_sfixed(-3551.0/65536.0,1,-nbitq), 
to_sfixed(1109.0/65536.0,1,-nbitq), 
to_sfixed(-878.0/65536.0,1,-nbitq), 
to_sfixed(8491.0/65536.0,1,-nbitq), 
to_sfixed(7761.0/65536.0,1,-nbitq), 
to_sfixed(166.0/65536.0,1,-nbitq), 
to_sfixed(308.0/65536.0,1,-nbitq), 
to_sfixed(1031.0/65536.0,1,-nbitq), 
to_sfixed(3590.0/65536.0,1,-nbitq), 
to_sfixed(-2423.0/65536.0,1,-nbitq), 
to_sfixed(-5092.0/65536.0,1,-nbitq), 
to_sfixed(3785.0/65536.0,1,-nbitq), 
to_sfixed(-1354.0/65536.0,1,-nbitq), 
to_sfixed(5206.0/65536.0,1,-nbitq), 
to_sfixed(-2458.0/65536.0,1,-nbitq), 
to_sfixed(9790.0/65536.0,1,-nbitq), 
to_sfixed(-1418.0/65536.0,1,-nbitq), 
to_sfixed(-1799.0/65536.0,1,-nbitq), 
to_sfixed(-4632.0/65536.0,1,-nbitq), 
to_sfixed(-597.0/65536.0,1,-nbitq), 
to_sfixed(-2245.0/65536.0,1,-nbitq), 
to_sfixed(-1870.0/65536.0,1,-nbitq), 
to_sfixed(3804.0/65536.0,1,-nbitq), 
to_sfixed(-1055.0/65536.0,1,-nbitq), 
to_sfixed(-1689.0/65536.0,1,-nbitq), 
to_sfixed(4871.0/65536.0,1,-nbitq), 
to_sfixed(1313.0/65536.0,1,-nbitq), 
to_sfixed(-2716.0/65536.0,1,-nbitq), 
to_sfixed(1741.0/65536.0,1,-nbitq), 
to_sfixed(4441.0/65536.0,1,-nbitq), 
to_sfixed(-962.0/65536.0,1,-nbitq), 
to_sfixed(1487.0/65536.0,1,-nbitq), 
to_sfixed(-2424.0/65536.0,1,-nbitq), 
to_sfixed(8736.0/65536.0,1,-nbitq), 
to_sfixed(-357.0/65536.0,1,-nbitq), 
to_sfixed(-3405.0/65536.0,1,-nbitq), 
to_sfixed(-74.0/65536.0,1,-nbitq), 
to_sfixed(6348.0/65536.0,1,-nbitq), 
to_sfixed(1042.0/65536.0,1,-nbitq), 
to_sfixed(-3577.0/65536.0,1,-nbitq), 
to_sfixed(319.0/65536.0,1,-nbitq), 
to_sfixed(3339.0/65536.0,1,-nbitq), 
to_sfixed(-2926.0/65536.0,1,-nbitq), 
to_sfixed(1786.0/65536.0,1,-nbitq), 
to_sfixed(1195.0/65536.0,1,-nbitq), 
to_sfixed(2027.0/65536.0,1,-nbitq), 
to_sfixed(4006.0/65536.0,1,-nbitq), 
to_sfixed(-4378.0/65536.0,1,-nbitq), 
to_sfixed(-2616.0/65536.0,1,-nbitq), 
to_sfixed(-4512.0/65536.0,1,-nbitq), 
to_sfixed(-5509.0/65536.0,1,-nbitq), 
to_sfixed(703.0/65536.0,1,-nbitq), 
to_sfixed(445.0/65536.0,1,-nbitq), 
to_sfixed(-5553.0/65536.0,1,-nbitq), 
to_sfixed(-928.0/65536.0,1,-nbitq), 
to_sfixed(-55.0/65536.0,1,-nbitq), 
to_sfixed(-2582.0/65536.0,1,-nbitq), 
to_sfixed(7257.0/65536.0,1,-nbitq), 
to_sfixed(2359.0/65536.0,1,-nbitq), 
to_sfixed(-8894.0/65536.0,1,-nbitq), 
to_sfixed(-1347.0/65536.0,1,-nbitq), 
to_sfixed(3462.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2511.0/65536.0,1,-nbitq), 
to_sfixed(-6470.0/65536.0,1,-nbitq), 
to_sfixed(1701.0/65536.0,1,-nbitq), 
to_sfixed(-2499.0/65536.0,1,-nbitq), 
to_sfixed(2376.0/65536.0,1,-nbitq), 
to_sfixed(-6287.0/65536.0,1,-nbitq), 
to_sfixed(5634.0/65536.0,1,-nbitq), 
to_sfixed(684.0/65536.0,1,-nbitq), 
to_sfixed(2084.0/65536.0,1,-nbitq), 
to_sfixed(-2561.0/65536.0,1,-nbitq), 
to_sfixed(-1971.0/65536.0,1,-nbitq), 
to_sfixed(339.0/65536.0,1,-nbitq), 
to_sfixed(590.0/65536.0,1,-nbitq), 
to_sfixed(-5070.0/65536.0,1,-nbitq), 
to_sfixed(1735.0/65536.0,1,-nbitq), 
to_sfixed(-475.0/65536.0,1,-nbitq), 
to_sfixed(1553.0/65536.0,1,-nbitq), 
to_sfixed(-325.0/65536.0,1,-nbitq), 
to_sfixed(-458.0/65536.0,1,-nbitq), 
to_sfixed(2417.0/65536.0,1,-nbitq), 
to_sfixed(-918.0/65536.0,1,-nbitq), 
to_sfixed(5327.0/65536.0,1,-nbitq), 
to_sfixed(3797.0/65536.0,1,-nbitq), 
to_sfixed(-517.0/65536.0,1,-nbitq), 
to_sfixed(4649.0/65536.0,1,-nbitq), 
to_sfixed(-2307.0/65536.0,1,-nbitq), 
to_sfixed(5838.0/65536.0,1,-nbitq), 
to_sfixed(-2041.0/65536.0,1,-nbitq), 
to_sfixed(-6815.0/65536.0,1,-nbitq), 
to_sfixed(1107.0/65536.0,1,-nbitq), 
to_sfixed(-7756.0/65536.0,1,-nbitq), 
to_sfixed(3655.0/65536.0,1,-nbitq), 
to_sfixed(4753.0/65536.0,1,-nbitq), 
to_sfixed(1714.0/65536.0,1,-nbitq), 
to_sfixed(-2942.0/65536.0,1,-nbitq), 
to_sfixed(-42.0/65536.0,1,-nbitq), 
to_sfixed(-1883.0/65536.0,1,-nbitq), 
to_sfixed(-672.0/65536.0,1,-nbitq), 
to_sfixed(3020.0/65536.0,1,-nbitq), 
to_sfixed(685.0/65536.0,1,-nbitq), 
to_sfixed(9918.0/65536.0,1,-nbitq), 
to_sfixed(-1122.0/65536.0,1,-nbitq), 
to_sfixed(-2309.0/65536.0,1,-nbitq), 
to_sfixed(1467.0/65536.0,1,-nbitq), 
to_sfixed(1355.0/65536.0,1,-nbitq), 
to_sfixed(-3153.0/65536.0,1,-nbitq), 
to_sfixed(1805.0/65536.0,1,-nbitq), 
to_sfixed(-4407.0/65536.0,1,-nbitq), 
to_sfixed(2642.0/65536.0,1,-nbitq), 
to_sfixed(-2052.0/65536.0,1,-nbitq), 
to_sfixed(2469.0/65536.0,1,-nbitq), 
to_sfixed(6802.0/65536.0,1,-nbitq), 
to_sfixed(-5314.0/65536.0,1,-nbitq), 
to_sfixed(-10111.0/65536.0,1,-nbitq), 
to_sfixed(3715.0/65536.0,1,-nbitq), 
to_sfixed(6460.0/65536.0,1,-nbitq), 
to_sfixed(-3036.0/65536.0,1,-nbitq), 
to_sfixed(-7511.0/65536.0,1,-nbitq), 
to_sfixed(-1941.0/65536.0,1,-nbitq), 
to_sfixed(-1210.0/65536.0,1,-nbitq), 
to_sfixed(-4840.0/65536.0,1,-nbitq), 
to_sfixed(836.0/65536.0,1,-nbitq), 
to_sfixed(2391.0/65536.0,1,-nbitq), 
to_sfixed(-554.0/65536.0,1,-nbitq), 
to_sfixed(9466.0/65536.0,1,-nbitq), 
to_sfixed(-1834.0/65536.0,1,-nbitq), 
to_sfixed(1082.0/65536.0,1,-nbitq), 
to_sfixed(-1728.0/65536.0,1,-nbitq), 
to_sfixed(-5991.0/65536.0,1,-nbitq), 
to_sfixed(-2396.0/65536.0,1,-nbitq), 
to_sfixed(2181.0/65536.0,1,-nbitq), 
to_sfixed(-3287.0/65536.0,1,-nbitq), 
to_sfixed(-1778.0/65536.0,1,-nbitq), 
to_sfixed(-1069.0/65536.0,1,-nbitq), 
to_sfixed(1572.0/65536.0,1,-nbitq), 
to_sfixed(5426.0/65536.0,1,-nbitq), 
to_sfixed(8848.0/65536.0,1,-nbitq), 
to_sfixed(-4920.0/65536.0,1,-nbitq), 
to_sfixed(-136.0/65536.0,1,-nbitq), 
to_sfixed(-993.0/65536.0,1,-nbitq)  ), 
( to_sfixed(6837.0/65536.0,1,-nbitq), 
to_sfixed(141.0/65536.0,1,-nbitq), 
to_sfixed(-7677.0/65536.0,1,-nbitq), 
to_sfixed(1927.0/65536.0,1,-nbitq), 
to_sfixed(-4756.0/65536.0,1,-nbitq), 
to_sfixed(-7169.0/65536.0,1,-nbitq), 
to_sfixed(4380.0/65536.0,1,-nbitq), 
to_sfixed(-1559.0/65536.0,1,-nbitq), 
to_sfixed(-2022.0/65536.0,1,-nbitq), 
to_sfixed(1535.0/65536.0,1,-nbitq), 
to_sfixed(-756.0/65536.0,1,-nbitq), 
to_sfixed(-3212.0/65536.0,1,-nbitq), 
to_sfixed(931.0/65536.0,1,-nbitq), 
to_sfixed(-4591.0/65536.0,1,-nbitq), 
to_sfixed(-1951.0/65536.0,1,-nbitq), 
to_sfixed(241.0/65536.0,1,-nbitq), 
to_sfixed(-1441.0/65536.0,1,-nbitq), 
to_sfixed(-1306.0/65536.0,1,-nbitq), 
to_sfixed(-3410.0/65536.0,1,-nbitq), 
to_sfixed(604.0/65536.0,1,-nbitq), 
to_sfixed(-306.0/65536.0,1,-nbitq), 
to_sfixed(7213.0/65536.0,1,-nbitq), 
to_sfixed(1811.0/65536.0,1,-nbitq), 
to_sfixed(-2461.0/65536.0,1,-nbitq), 
to_sfixed(3186.0/65536.0,1,-nbitq), 
to_sfixed(-5629.0/65536.0,1,-nbitq), 
to_sfixed(1778.0/65536.0,1,-nbitq), 
to_sfixed(-4094.0/65536.0,1,-nbitq), 
to_sfixed(-7091.0/65536.0,1,-nbitq), 
to_sfixed(-3277.0/65536.0,1,-nbitq), 
to_sfixed(-11524.0/65536.0,1,-nbitq), 
to_sfixed(4506.0/65536.0,1,-nbitq), 
to_sfixed(3358.0/65536.0,1,-nbitq), 
to_sfixed(-5252.0/65536.0,1,-nbitq), 
to_sfixed(997.0/65536.0,1,-nbitq), 
to_sfixed(2348.0/65536.0,1,-nbitq), 
to_sfixed(-858.0/65536.0,1,-nbitq), 
to_sfixed(-1399.0/65536.0,1,-nbitq), 
to_sfixed(1974.0/65536.0,1,-nbitq), 
to_sfixed(-1159.0/65536.0,1,-nbitq), 
to_sfixed(11180.0/65536.0,1,-nbitq), 
to_sfixed(1650.0/65536.0,1,-nbitq), 
to_sfixed(1004.0/65536.0,1,-nbitq), 
to_sfixed(132.0/65536.0,1,-nbitq), 
to_sfixed(2505.0/65536.0,1,-nbitq), 
to_sfixed(-1263.0/65536.0,1,-nbitq), 
to_sfixed(2377.0/65536.0,1,-nbitq), 
to_sfixed(-3684.0/65536.0,1,-nbitq), 
to_sfixed(-1129.0/65536.0,1,-nbitq), 
to_sfixed(-2215.0/65536.0,1,-nbitq), 
to_sfixed(-1.0/65536.0,1,-nbitq), 
to_sfixed(3787.0/65536.0,1,-nbitq), 
to_sfixed(811.0/65536.0,1,-nbitq), 
to_sfixed(-3740.0/65536.0,1,-nbitq), 
to_sfixed(856.0/65536.0,1,-nbitq), 
to_sfixed(5006.0/65536.0,1,-nbitq), 
to_sfixed(2677.0/65536.0,1,-nbitq), 
to_sfixed(-3791.0/65536.0,1,-nbitq), 
to_sfixed(-744.0/65536.0,1,-nbitq), 
to_sfixed(-7452.0/65536.0,1,-nbitq), 
to_sfixed(-6121.0/65536.0,1,-nbitq), 
to_sfixed(-1905.0/65536.0,1,-nbitq), 
to_sfixed(-642.0/65536.0,1,-nbitq), 
to_sfixed(2340.0/65536.0,1,-nbitq), 
to_sfixed(2111.0/65536.0,1,-nbitq), 
to_sfixed(-5325.0/65536.0,1,-nbitq), 
to_sfixed(2671.0/65536.0,1,-nbitq), 
to_sfixed(232.0/65536.0,1,-nbitq), 
to_sfixed(-5838.0/65536.0,1,-nbitq), 
to_sfixed(-2919.0/65536.0,1,-nbitq), 
to_sfixed(1214.0/65536.0,1,-nbitq), 
to_sfixed(-5250.0/65536.0,1,-nbitq), 
to_sfixed(2320.0/65536.0,1,-nbitq), 
to_sfixed(-583.0/65536.0,1,-nbitq), 
to_sfixed(-419.0/65536.0,1,-nbitq), 
to_sfixed(2867.0/65536.0,1,-nbitq), 
to_sfixed(9188.0/65536.0,1,-nbitq), 
to_sfixed(-1624.0/65536.0,1,-nbitq), 
to_sfixed(2755.0/65536.0,1,-nbitq), 
to_sfixed(1504.0/65536.0,1,-nbitq)  ), 
( to_sfixed(6511.0/65536.0,1,-nbitq), 
to_sfixed(-2121.0/65536.0,1,-nbitq), 
to_sfixed(-2018.0/65536.0,1,-nbitq), 
to_sfixed(3439.0/65536.0,1,-nbitq), 
to_sfixed(-6772.0/65536.0,1,-nbitq), 
to_sfixed(-8071.0/65536.0,1,-nbitq), 
to_sfixed(4992.0/65536.0,1,-nbitq), 
to_sfixed(-1973.0/65536.0,1,-nbitq), 
to_sfixed(983.0/65536.0,1,-nbitq), 
to_sfixed(-2173.0/65536.0,1,-nbitq), 
to_sfixed(-2263.0/65536.0,1,-nbitq), 
to_sfixed(6035.0/65536.0,1,-nbitq), 
to_sfixed(2783.0/65536.0,1,-nbitq), 
to_sfixed(-1717.0/65536.0,1,-nbitq), 
to_sfixed(136.0/65536.0,1,-nbitq), 
to_sfixed(950.0/65536.0,1,-nbitq), 
to_sfixed(-602.0/65536.0,1,-nbitq), 
to_sfixed(588.0/65536.0,1,-nbitq), 
to_sfixed(1541.0/65536.0,1,-nbitq), 
to_sfixed(676.0/65536.0,1,-nbitq), 
to_sfixed(2386.0/65536.0,1,-nbitq), 
to_sfixed(841.0/65536.0,1,-nbitq), 
to_sfixed(1278.0/65536.0,1,-nbitq), 
to_sfixed(-1543.0/65536.0,1,-nbitq), 
to_sfixed(911.0/65536.0,1,-nbitq), 
to_sfixed(-663.0/65536.0,1,-nbitq), 
to_sfixed(1089.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(-7849.0/65536.0,1,-nbitq), 
to_sfixed(-1741.0/65536.0,1,-nbitq), 
to_sfixed(-5468.0/65536.0,1,-nbitq), 
to_sfixed(5579.0/65536.0,1,-nbitq), 
to_sfixed(3072.0/65536.0,1,-nbitq), 
to_sfixed(-2785.0/65536.0,1,-nbitq), 
to_sfixed(3336.0/65536.0,1,-nbitq), 
to_sfixed(-3038.0/65536.0,1,-nbitq), 
to_sfixed(-552.0/65536.0,1,-nbitq), 
to_sfixed(-6456.0/65536.0,1,-nbitq), 
to_sfixed(2685.0/65536.0,1,-nbitq), 
to_sfixed(-2533.0/65536.0,1,-nbitq), 
to_sfixed(7614.0/65536.0,1,-nbitq), 
to_sfixed(-2117.0/65536.0,1,-nbitq), 
to_sfixed(4228.0/65536.0,1,-nbitq), 
to_sfixed(-2472.0/65536.0,1,-nbitq), 
to_sfixed(448.0/65536.0,1,-nbitq), 
to_sfixed(3455.0/65536.0,1,-nbitq), 
to_sfixed(-1939.0/65536.0,1,-nbitq), 
to_sfixed(-2748.0/65536.0,1,-nbitq), 
to_sfixed(-75.0/65536.0,1,-nbitq), 
to_sfixed(-61.0/65536.0,1,-nbitq), 
to_sfixed(-1562.0/65536.0,1,-nbitq), 
to_sfixed(1252.0/65536.0,1,-nbitq), 
to_sfixed(1505.0/65536.0,1,-nbitq), 
to_sfixed(-1879.0/65536.0,1,-nbitq), 
to_sfixed(1271.0/65536.0,1,-nbitq), 
to_sfixed(7800.0/65536.0,1,-nbitq), 
to_sfixed(-133.0/65536.0,1,-nbitq), 
to_sfixed(2061.0/65536.0,1,-nbitq), 
to_sfixed(-1127.0/65536.0,1,-nbitq), 
to_sfixed(1126.0/65536.0,1,-nbitq), 
to_sfixed(-298.0/65536.0,1,-nbitq), 
to_sfixed(1563.0/65536.0,1,-nbitq), 
to_sfixed(-2552.0/65536.0,1,-nbitq), 
to_sfixed(212.0/65536.0,1,-nbitq), 
to_sfixed(592.0/65536.0,1,-nbitq), 
to_sfixed(-6866.0/65536.0,1,-nbitq), 
to_sfixed(-354.0/65536.0,1,-nbitq), 
to_sfixed(1878.0/65536.0,1,-nbitq), 
to_sfixed(-4870.0/65536.0,1,-nbitq), 
to_sfixed(-5250.0/65536.0,1,-nbitq), 
to_sfixed(2874.0/65536.0,1,-nbitq), 
to_sfixed(1669.0/65536.0,1,-nbitq), 
to_sfixed(1720.0/65536.0,1,-nbitq), 
to_sfixed(-2278.0/65536.0,1,-nbitq), 
to_sfixed(-1625.0/65536.0,1,-nbitq), 
to_sfixed(2968.0/65536.0,1,-nbitq), 
to_sfixed(2664.0/65536.0,1,-nbitq), 
to_sfixed(568.0/65536.0,1,-nbitq), 
to_sfixed(2407.0/65536.0,1,-nbitq), 
to_sfixed(-1145.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1196.0/65536.0,1,-nbitq), 
to_sfixed(-1462.0/65536.0,1,-nbitq), 
to_sfixed(6417.0/65536.0,1,-nbitq), 
to_sfixed(1183.0/65536.0,1,-nbitq), 
to_sfixed(-11563.0/65536.0,1,-nbitq), 
to_sfixed(-691.0/65536.0,1,-nbitq), 
to_sfixed(1533.0/65536.0,1,-nbitq), 
to_sfixed(-3730.0/65536.0,1,-nbitq), 
to_sfixed(-2346.0/65536.0,1,-nbitq), 
to_sfixed(2741.0/65536.0,1,-nbitq), 
to_sfixed(-882.0/65536.0,1,-nbitq), 
to_sfixed(2188.0/65536.0,1,-nbitq), 
to_sfixed(2104.0/65536.0,1,-nbitq), 
to_sfixed(-3967.0/65536.0,1,-nbitq), 
to_sfixed(4568.0/65536.0,1,-nbitq), 
to_sfixed(-1481.0/65536.0,1,-nbitq), 
to_sfixed(939.0/65536.0,1,-nbitq), 
to_sfixed(2337.0/65536.0,1,-nbitq), 
to_sfixed(261.0/65536.0,1,-nbitq), 
to_sfixed(2958.0/65536.0,1,-nbitq), 
to_sfixed(3639.0/65536.0,1,-nbitq), 
to_sfixed(-761.0/65536.0,1,-nbitq), 
to_sfixed(416.0/65536.0,1,-nbitq), 
to_sfixed(1792.0/65536.0,1,-nbitq), 
to_sfixed(2226.0/65536.0,1,-nbitq), 
to_sfixed(190.0/65536.0,1,-nbitq), 
to_sfixed(-700.0/65536.0,1,-nbitq), 
to_sfixed(1072.0/65536.0,1,-nbitq), 
to_sfixed(-4970.0/65536.0,1,-nbitq), 
to_sfixed(1945.0/65536.0,1,-nbitq), 
to_sfixed(-2096.0/65536.0,1,-nbitq), 
to_sfixed(6474.0/65536.0,1,-nbitq), 
to_sfixed(2769.0/65536.0,1,-nbitq), 
to_sfixed(-2063.0/65536.0,1,-nbitq), 
to_sfixed(3353.0/65536.0,1,-nbitq), 
to_sfixed(927.0/65536.0,1,-nbitq), 
to_sfixed(-1363.0/65536.0,1,-nbitq), 
to_sfixed(-2099.0/65536.0,1,-nbitq), 
to_sfixed(3312.0/65536.0,1,-nbitq), 
to_sfixed(229.0/65536.0,1,-nbitq), 
to_sfixed(4485.0/65536.0,1,-nbitq), 
to_sfixed(2722.0/65536.0,1,-nbitq), 
to_sfixed(3871.0/65536.0,1,-nbitq), 
to_sfixed(-2472.0/65536.0,1,-nbitq), 
to_sfixed(291.0/65536.0,1,-nbitq), 
to_sfixed(3545.0/65536.0,1,-nbitq), 
to_sfixed(-2736.0/65536.0,1,-nbitq), 
to_sfixed(470.0/65536.0,1,-nbitq), 
to_sfixed(-2608.0/65536.0,1,-nbitq), 
to_sfixed(366.0/65536.0,1,-nbitq), 
to_sfixed(-1504.0/65536.0,1,-nbitq), 
to_sfixed(2280.0/65536.0,1,-nbitq), 
to_sfixed(483.0/65536.0,1,-nbitq), 
to_sfixed(-1285.0/65536.0,1,-nbitq), 
to_sfixed(2174.0/65536.0,1,-nbitq), 
to_sfixed(5713.0/65536.0,1,-nbitq), 
to_sfixed(2330.0/65536.0,1,-nbitq), 
to_sfixed(2602.0/65536.0,1,-nbitq), 
to_sfixed(-1015.0/65536.0,1,-nbitq), 
to_sfixed(2646.0/65536.0,1,-nbitq), 
to_sfixed(2678.0/65536.0,1,-nbitq), 
to_sfixed(-1561.0/65536.0,1,-nbitq), 
to_sfixed(-1889.0/65536.0,1,-nbitq), 
to_sfixed(-3111.0/65536.0,1,-nbitq), 
to_sfixed(-3440.0/65536.0,1,-nbitq), 
to_sfixed(-1213.0/65536.0,1,-nbitq), 
to_sfixed(-4246.0/65536.0,1,-nbitq), 
to_sfixed(1179.0/65536.0,1,-nbitq), 
to_sfixed(-5502.0/65536.0,1,-nbitq), 
to_sfixed(719.0/65536.0,1,-nbitq), 
to_sfixed(1648.0/65536.0,1,-nbitq), 
to_sfixed(1583.0/65536.0,1,-nbitq), 
to_sfixed(-221.0/65536.0,1,-nbitq), 
to_sfixed(1708.0/65536.0,1,-nbitq), 
to_sfixed(-2572.0/65536.0,1,-nbitq), 
to_sfixed(-2522.0/65536.0,1,-nbitq), 
to_sfixed(1988.0/65536.0,1,-nbitq), 
to_sfixed(778.0/65536.0,1,-nbitq), 
to_sfixed(-1574.0/65536.0,1,-nbitq), 
to_sfixed(-62.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4689.0/65536.0,1,-nbitq), 
to_sfixed(1000.0/65536.0,1,-nbitq), 
to_sfixed(6760.0/65536.0,1,-nbitq), 
to_sfixed(2188.0/65536.0,1,-nbitq), 
to_sfixed(-8169.0/65536.0,1,-nbitq), 
to_sfixed(-4635.0/65536.0,1,-nbitq), 
to_sfixed(2012.0/65536.0,1,-nbitq), 
to_sfixed(900.0/65536.0,1,-nbitq), 
to_sfixed(-429.0/65536.0,1,-nbitq), 
to_sfixed(1570.0/65536.0,1,-nbitq), 
to_sfixed(-2803.0/65536.0,1,-nbitq), 
to_sfixed(-779.0/65536.0,1,-nbitq), 
to_sfixed(3392.0/65536.0,1,-nbitq), 
to_sfixed(-6904.0/65536.0,1,-nbitq), 
to_sfixed(-2701.0/65536.0,1,-nbitq), 
to_sfixed(-424.0/65536.0,1,-nbitq), 
to_sfixed(-2518.0/65536.0,1,-nbitq), 
to_sfixed(4421.0/65536.0,1,-nbitq), 
to_sfixed(-114.0/65536.0,1,-nbitq), 
to_sfixed(1216.0/65536.0,1,-nbitq), 
to_sfixed(1579.0/65536.0,1,-nbitq), 
to_sfixed(-1788.0/65536.0,1,-nbitq), 
to_sfixed(-2036.0/65536.0,1,-nbitq), 
to_sfixed(-4484.0/65536.0,1,-nbitq), 
to_sfixed(4404.0/65536.0,1,-nbitq), 
to_sfixed(-5210.0/65536.0,1,-nbitq), 
to_sfixed(-6662.0/65536.0,1,-nbitq), 
to_sfixed(1095.0/65536.0,1,-nbitq), 
to_sfixed(-788.0/65536.0,1,-nbitq), 
to_sfixed(3287.0/65536.0,1,-nbitq), 
to_sfixed(-3474.0/65536.0,1,-nbitq), 
to_sfixed(2424.0/65536.0,1,-nbitq), 
to_sfixed(5827.0/65536.0,1,-nbitq), 
to_sfixed(1992.0/65536.0,1,-nbitq), 
to_sfixed(2826.0/65536.0,1,-nbitq), 
to_sfixed(657.0/65536.0,1,-nbitq), 
to_sfixed(87.0/65536.0,1,-nbitq), 
to_sfixed(-3149.0/65536.0,1,-nbitq), 
to_sfixed(1135.0/65536.0,1,-nbitq), 
to_sfixed(-87.0/65536.0,1,-nbitq), 
to_sfixed(-519.0/65536.0,1,-nbitq), 
to_sfixed(296.0/65536.0,1,-nbitq), 
to_sfixed(-1648.0/65536.0,1,-nbitq), 
to_sfixed(-1891.0/65536.0,1,-nbitq), 
to_sfixed(1540.0/65536.0,1,-nbitq), 
to_sfixed(-1261.0/65536.0,1,-nbitq), 
to_sfixed(-143.0/65536.0,1,-nbitq), 
to_sfixed(2161.0/65536.0,1,-nbitq), 
to_sfixed(-1472.0/65536.0,1,-nbitq), 
to_sfixed(1315.0/65536.0,1,-nbitq), 
to_sfixed(-2282.0/65536.0,1,-nbitq), 
to_sfixed(3258.0/65536.0,1,-nbitq), 
to_sfixed(477.0/65536.0,1,-nbitq), 
to_sfixed(1135.0/65536.0,1,-nbitq), 
to_sfixed(-2988.0/65536.0,1,-nbitq), 
to_sfixed(5436.0/65536.0,1,-nbitq), 
to_sfixed(-2978.0/65536.0,1,-nbitq), 
to_sfixed(5698.0/65536.0,1,-nbitq), 
to_sfixed(1359.0/65536.0,1,-nbitq), 
to_sfixed(-419.0/65536.0,1,-nbitq), 
to_sfixed(6126.0/65536.0,1,-nbitq), 
to_sfixed(-2498.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(-40.0/65536.0,1,-nbitq), 
to_sfixed(-1180.0/65536.0,1,-nbitq), 
to_sfixed(-6930.0/65536.0,1,-nbitq), 
to_sfixed(-4869.0/65536.0,1,-nbitq), 
to_sfixed(-4339.0/65536.0,1,-nbitq), 
to_sfixed(4781.0/65536.0,1,-nbitq), 
to_sfixed(4832.0/65536.0,1,-nbitq), 
to_sfixed(-2016.0/65536.0,1,-nbitq), 
to_sfixed(3734.0/65536.0,1,-nbitq), 
to_sfixed(-5163.0/65536.0,1,-nbitq), 
to_sfixed(-165.0/65536.0,1,-nbitq), 
to_sfixed(1450.0/65536.0,1,-nbitq), 
to_sfixed(796.0/65536.0,1,-nbitq), 
to_sfixed(3529.0/65536.0,1,-nbitq), 
to_sfixed(1535.0/65536.0,1,-nbitq), 
to_sfixed(-1112.0/65536.0,1,-nbitq), 
to_sfixed(297.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-758.0/65536.0,1,-nbitq), 
to_sfixed(-1023.0/65536.0,1,-nbitq), 
to_sfixed(1517.0/65536.0,1,-nbitq), 
to_sfixed(511.0/65536.0,1,-nbitq), 
to_sfixed(-2799.0/65536.0,1,-nbitq), 
to_sfixed(-6284.0/65536.0,1,-nbitq), 
to_sfixed(3098.0/65536.0,1,-nbitq), 
to_sfixed(1770.0/65536.0,1,-nbitq), 
to_sfixed(-779.0/65536.0,1,-nbitq), 
to_sfixed(1293.0/65536.0,1,-nbitq), 
to_sfixed(-562.0/65536.0,1,-nbitq), 
to_sfixed(-71.0/65536.0,1,-nbitq), 
to_sfixed(-2205.0/65536.0,1,-nbitq), 
to_sfixed(-7456.0/65536.0,1,-nbitq), 
to_sfixed(766.0/65536.0,1,-nbitq), 
to_sfixed(-2143.0/65536.0,1,-nbitq), 
to_sfixed(-1612.0/65536.0,1,-nbitq), 
to_sfixed(2797.0/65536.0,1,-nbitq), 
to_sfixed(265.0/65536.0,1,-nbitq), 
to_sfixed(1302.0/65536.0,1,-nbitq), 
to_sfixed(-797.0/65536.0,1,-nbitq), 
to_sfixed(-2040.0/65536.0,1,-nbitq), 
to_sfixed(478.0/65536.0,1,-nbitq), 
to_sfixed(-4825.0/65536.0,1,-nbitq), 
to_sfixed(-1150.0/65536.0,1,-nbitq), 
to_sfixed(-1743.0/65536.0,1,-nbitq), 
to_sfixed(-3526.0/65536.0,1,-nbitq), 
to_sfixed(1689.0/65536.0,1,-nbitq), 
to_sfixed(-1457.0/65536.0,1,-nbitq), 
to_sfixed(1402.0/65536.0,1,-nbitq), 
to_sfixed(-4609.0/65536.0,1,-nbitq), 
to_sfixed(3579.0/65536.0,1,-nbitq), 
to_sfixed(60.0/65536.0,1,-nbitq), 
to_sfixed(3883.0/65536.0,1,-nbitq), 
to_sfixed(-2870.0/65536.0,1,-nbitq), 
to_sfixed(2399.0/65536.0,1,-nbitq), 
to_sfixed(5461.0/65536.0,1,-nbitq), 
to_sfixed(1051.0/65536.0,1,-nbitq), 
to_sfixed(1938.0/65536.0,1,-nbitq), 
to_sfixed(-531.0/65536.0,1,-nbitq), 
to_sfixed(-1704.0/65536.0,1,-nbitq), 
to_sfixed(1291.0/65536.0,1,-nbitq), 
to_sfixed(3771.0/65536.0,1,-nbitq), 
to_sfixed(-2242.0/65536.0,1,-nbitq), 
to_sfixed(-338.0/65536.0,1,-nbitq), 
to_sfixed(2229.0/65536.0,1,-nbitq), 
to_sfixed(1916.0/65536.0,1,-nbitq), 
to_sfixed(1582.0/65536.0,1,-nbitq), 
to_sfixed(1406.0/65536.0,1,-nbitq), 
to_sfixed(3142.0/65536.0,1,-nbitq), 
to_sfixed(736.0/65536.0,1,-nbitq), 
to_sfixed(-129.0/65536.0,1,-nbitq), 
to_sfixed(-4918.0/65536.0,1,-nbitq), 
to_sfixed(3386.0/65536.0,1,-nbitq), 
to_sfixed(-1802.0/65536.0,1,-nbitq), 
to_sfixed(5927.0/65536.0,1,-nbitq), 
to_sfixed(-809.0/65536.0,1,-nbitq), 
to_sfixed(2835.0/65536.0,1,-nbitq), 
to_sfixed(1302.0/65536.0,1,-nbitq), 
to_sfixed(-4805.0/65536.0,1,-nbitq), 
to_sfixed(125.0/65536.0,1,-nbitq), 
to_sfixed(-1322.0/65536.0,1,-nbitq), 
to_sfixed(-777.0/65536.0,1,-nbitq), 
to_sfixed(-2533.0/65536.0,1,-nbitq), 
to_sfixed(-1476.0/65536.0,1,-nbitq), 
to_sfixed(-1815.0/65536.0,1,-nbitq), 
to_sfixed(-1156.0/65536.0,1,-nbitq), 
to_sfixed(-3281.0/65536.0,1,-nbitq), 
to_sfixed(9188.0/65536.0,1,-nbitq), 
to_sfixed(1331.0/65536.0,1,-nbitq), 
to_sfixed(-557.0/65536.0,1,-nbitq), 
to_sfixed(978.0/65536.0,1,-nbitq), 
to_sfixed(-1396.0/65536.0,1,-nbitq), 
to_sfixed(-1305.0/65536.0,1,-nbitq), 
to_sfixed(-894.0/65536.0,1,-nbitq), 
to_sfixed(420.0/65536.0,1,-nbitq), 
to_sfixed(-1074.0/65536.0,1,-nbitq), 
to_sfixed(-1792.0/65536.0,1,-nbitq), 
to_sfixed(-1609.0/65536.0,1,-nbitq), 
to_sfixed(5025.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2799.0/65536.0,1,-nbitq), 
to_sfixed(3456.0/65536.0,1,-nbitq), 
to_sfixed(-2911.0/65536.0,1,-nbitq), 
to_sfixed(-2440.0/65536.0,1,-nbitq), 
to_sfixed(1245.0/65536.0,1,-nbitq), 
to_sfixed(-3359.0/65536.0,1,-nbitq), 
to_sfixed(-108.0/65536.0,1,-nbitq), 
to_sfixed(1736.0/65536.0,1,-nbitq), 
to_sfixed(-1754.0/65536.0,1,-nbitq), 
to_sfixed(1833.0/65536.0,1,-nbitq), 
to_sfixed(790.0/65536.0,1,-nbitq), 
to_sfixed(3420.0/65536.0,1,-nbitq), 
to_sfixed(-2055.0/65536.0,1,-nbitq), 
to_sfixed(-2401.0/65536.0,1,-nbitq), 
to_sfixed(1666.0/65536.0,1,-nbitq), 
to_sfixed(2940.0/65536.0,1,-nbitq), 
to_sfixed(1311.0/65536.0,1,-nbitq), 
to_sfixed(-1259.0/65536.0,1,-nbitq), 
to_sfixed(2731.0/65536.0,1,-nbitq), 
to_sfixed(-1791.0/65536.0,1,-nbitq), 
to_sfixed(2572.0/65536.0,1,-nbitq), 
to_sfixed(-3690.0/65536.0,1,-nbitq), 
to_sfixed(-2375.0/65536.0,1,-nbitq), 
to_sfixed(-8517.0/65536.0,1,-nbitq), 
to_sfixed(3614.0/65536.0,1,-nbitq), 
to_sfixed(-4881.0/65536.0,1,-nbitq), 
to_sfixed(-7508.0/65536.0,1,-nbitq), 
to_sfixed(-2089.0/65536.0,1,-nbitq), 
to_sfixed(3627.0/65536.0,1,-nbitq), 
to_sfixed(-2150.0/65536.0,1,-nbitq), 
to_sfixed(966.0/65536.0,1,-nbitq), 
to_sfixed(-2414.0/65536.0,1,-nbitq), 
to_sfixed(2043.0/65536.0,1,-nbitq), 
to_sfixed(2200.0/65536.0,1,-nbitq), 
to_sfixed(-1053.0/65536.0,1,-nbitq), 
to_sfixed(-2050.0/65536.0,1,-nbitq), 
to_sfixed(1629.0/65536.0,1,-nbitq), 
to_sfixed(-1003.0/65536.0,1,-nbitq), 
to_sfixed(611.0/65536.0,1,-nbitq), 
to_sfixed(31.0/65536.0,1,-nbitq), 
to_sfixed(685.0/65536.0,1,-nbitq), 
to_sfixed(2023.0/65536.0,1,-nbitq), 
to_sfixed(1045.0/65536.0,1,-nbitq), 
to_sfixed(2252.0/65536.0,1,-nbitq), 
to_sfixed(-91.0/65536.0,1,-nbitq), 
to_sfixed(2218.0/65536.0,1,-nbitq), 
to_sfixed(-2728.0/65536.0,1,-nbitq), 
to_sfixed(-1589.0/65536.0,1,-nbitq), 
to_sfixed(-166.0/65536.0,1,-nbitq), 
to_sfixed(809.0/65536.0,1,-nbitq), 
to_sfixed(-1021.0/65536.0,1,-nbitq), 
to_sfixed(-1730.0/65536.0,1,-nbitq), 
to_sfixed(-804.0/65536.0,1,-nbitq), 
to_sfixed(5195.0/65536.0,1,-nbitq), 
to_sfixed(-1788.0/65536.0,1,-nbitq), 
to_sfixed(-302.0/65536.0,1,-nbitq), 
to_sfixed(395.0/65536.0,1,-nbitq), 
to_sfixed(2978.0/65536.0,1,-nbitq), 
to_sfixed(-1533.0/65536.0,1,-nbitq), 
to_sfixed(-2474.0/65536.0,1,-nbitq), 
to_sfixed(2460.0/65536.0,1,-nbitq), 
to_sfixed(-1346.0/65536.0,1,-nbitq), 
to_sfixed(93.0/65536.0,1,-nbitq), 
to_sfixed(1363.0/65536.0,1,-nbitq), 
to_sfixed(-2135.0/65536.0,1,-nbitq), 
to_sfixed(-1077.0/65536.0,1,-nbitq), 
to_sfixed(3100.0/65536.0,1,-nbitq), 
to_sfixed(-1764.0/65536.0,1,-nbitq), 
to_sfixed(9107.0/65536.0,1,-nbitq), 
to_sfixed(1978.0/65536.0,1,-nbitq), 
to_sfixed(-732.0/65536.0,1,-nbitq), 
to_sfixed(-1613.0/65536.0,1,-nbitq), 
to_sfixed(-3114.0/65536.0,1,-nbitq), 
to_sfixed(-3108.0/65536.0,1,-nbitq), 
to_sfixed(-1173.0/65536.0,1,-nbitq), 
to_sfixed(2700.0/65536.0,1,-nbitq), 
to_sfixed(-1018.0/65536.0,1,-nbitq), 
to_sfixed(793.0/65536.0,1,-nbitq), 
to_sfixed(584.0/65536.0,1,-nbitq), 
to_sfixed(165.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1505.0/65536.0,1,-nbitq), 
to_sfixed(725.0/65536.0,1,-nbitq), 
to_sfixed(-1181.0/65536.0,1,-nbitq), 
to_sfixed(-258.0/65536.0,1,-nbitq), 
to_sfixed(-2557.0/65536.0,1,-nbitq), 
to_sfixed(-1780.0/65536.0,1,-nbitq), 
to_sfixed(2732.0/65536.0,1,-nbitq), 
to_sfixed(39.0/65536.0,1,-nbitq), 
to_sfixed(-3939.0/65536.0,1,-nbitq), 
to_sfixed(-1137.0/65536.0,1,-nbitq), 
to_sfixed(-1384.0/65536.0,1,-nbitq), 
to_sfixed(5149.0/65536.0,1,-nbitq), 
to_sfixed(-734.0/65536.0,1,-nbitq), 
to_sfixed(-3676.0/65536.0,1,-nbitq), 
to_sfixed(679.0/65536.0,1,-nbitq), 
to_sfixed(1485.0/65536.0,1,-nbitq), 
to_sfixed(1078.0/65536.0,1,-nbitq), 
to_sfixed(-1986.0/65536.0,1,-nbitq), 
to_sfixed(2838.0/65536.0,1,-nbitq), 
to_sfixed(-256.0/65536.0,1,-nbitq), 
to_sfixed(-469.0/65536.0,1,-nbitq), 
to_sfixed(3383.0/65536.0,1,-nbitq), 
to_sfixed(309.0/65536.0,1,-nbitq), 
to_sfixed(-745.0/65536.0,1,-nbitq), 
to_sfixed(348.0/65536.0,1,-nbitq), 
to_sfixed(1514.0/65536.0,1,-nbitq), 
to_sfixed(-3052.0/65536.0,1,-nbitq), 
to_sfixed(-460.0/65536.0,1,-nbitq), 
to_sfixed(3017.0/65536.0,1,-nbitq), 
to_sfixed(-2089.0/65536.0,1,-nbitq), 
to_sfixed(-2873.0/65536.0,1,-nbitq), 
to_sfixed(-1358.0/65536.0,1,-nbitq), 
to_sfixed(-756.0/65536.0,1,-nbitq), 
to_sfixed(-1753.0/65536.0,1,-nbitq), 
to_sfixed(56.0/65536.0,1,-nbitq), 
to_sfixed(2656.0/65536.0,1,-nbitq), 
to_sfixed(2029.0/65536.0,1,-nbitq), 
to_sfixed(-2420.0/65536.0,1,-nbitq), 
to_sfixed(309.0/65536.0,1,-nbitq), 
to_sfixed(-2547.0/65536.0,1,-nbitq), 
to_sfixed(1015.0/65536.0,1,-nbitq), 
to_sfixed(-1309.0/65536.0,1,-nbitq), 
to_sfixed(-2073.0/65536.0,1,-nbitq), 
to_sfixed(1582.0/65536.0,1,-nbitq), 
to_sfixed(-323.0/65536.0,1,-nbitq), 
to_sfixed(363.0/65536.0,1,-nbitq), 
to_sfixed(223.0/65536.0,1,-nbitq), 
to_sfixed(-2143.0/65536.0,1,-nbitq), 
to_sfixed(-1468.0/65536.0,1,-nbitq), 
to_sfixed(1034.0/65536.0,1,-nbitq), 
to_sfixed(-2459.0/65536.0,1,-nbitq), 
to_sfixed(-672.0/65536.0,1,-nbitq), 
to_sfixed(-2309.0/65536.0,1,-nbitq), 
to_sfixed(-911.0/65536.0,1,-nbitq), 
to_sfixed(-2900.0/65536.0,1,-nbitq), 
to_sfixed(-1840.0/65536.0,1,-nbitq), 
to_sfixed(808.0/65536.0,1,-nbitq), 
to_sfixed(-1006.0/65536.0,1,-nbitq), 
to_sfixed(307.0/65536.0,1,-nbitq), 
to_sfixed(1496.0/65536.0,1,-nbitq), 
to_sfixed(-1084.0/65536.0,1,-nbitq), 
to_sfixed(2670.0/65536.0,1,-nbitq), 
to_sfixed(-1966.0/65536.0,1,-nbitq), 
to_sfixed(1760.0/65536.0,1,-nbitq), 
to_sfixed(611.0/65536.0,1,-nbitq), 
to_sfixed(-559.0/65536.0,1,-nbitq), 
to_sfixed(-887.0/65536.0,1,-nbitq), 
to_sfixed(-599.0/65536.0,1,-nbitq), 
to_sfixed(5370.0/65536.0,1,-nbitq), 
to_sfixed(1591.0/65536.0,1,-nbitq), 
to_sfixed(230.0/65536.0,1,-nbitq), 
to_sfixed(1870.0/65536.0,1,-nbitq), 
to_sfixed(-1460.0/65536.0,1,-nbitq), 
to_sfixed(38.0/65536.0,1,-nbitq), 
to_sfixed(1542.0/65536.0,1,-nbitq), 
to_sfixed(847.0/65536.0,1,-nbitq), 
to_sfixed(-4720.0/65536.0,1,-nbitq), 
to_sfixed(1504.0/65536.0,1,-nbitq), 
to_sfixed(800.0/65536.0,1,-nbitq), 
to_sfixed(-775.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1783.0/65536.0,1,-nbitq), 
to_sfixed(-403.0/65536.0,1,-nbitq), 
to_sfixed(-752.0/65536.0,1,-nbitq), 
to_sfixed(-1730.0/65536.0,1,-nbitq), 
to_sfixed(483.0/65536.0,1,-nbitq), 
to_sfixed(-1450.0/65536.0,1,-nbitq), 
to_sfixed(-755.0/65536.0,1,-nbitq), 
to_sfixed(-616.0/65536.0,1,-nbitq), 
to_sfixed(-515.0/65536.0,1,-nbitq), 
to_sfixed(-2761.0/65536.0,1,-nbitq), 
to_sfixed(-1303.0/65536.0,1,-nbitq), 
to_sfixed(4505.0/65536.0,1,-nbitq), 
to_sfixed(-89.0/65536.0,1,-nbitq), 
to_sfixed(-2540.0/65536.0,1,-nbitq), 
to_sfixed(1237.0/65536.0,1,-nbitq), 
to_sfixed(-2016.0/65536.0,1,-nbitq), 
to_sfixed(-2736.0/65536.0,1,-nbitq), 
to_sfixed(443.0/65536.0,1,-nbitq), 
to_sfixed(811.0/65536.0,1,-nbitq), 
to_sfixed(1903.0/65536.0,1,-nbitq), 
to_sfixed(-222.0/65536.0,1,-nbitq), 
to_sfixed(508.0/65536.0,1,-nbitq), 
to_sfixed(-2812.0/65536.0,1,-nbitq), 
to_sfixed(-2616.0/65536.0,1,-nbitq), 
to_sfixed(-677.0/65536.0,1,-nbitq), 
to_sfixed(-434.0/65536.0,1,-nbitq), 
to_sfixed(603.0/65536.0,1,-nbitq), 
to_sfixed(2965.0/65536.0,1,-nbitq), 
to_sfixed(-1145.0/65536.0,1,-nbitq), 
to_sfixed(1620.0/65536.0,1,-nbitq), 
to_sfixed(289.0/65536.0,1,-nbitq), 
to_sfixed(211.0/65536.0,1,-nbitq), 
to_sfixed(-8.0/65536.0,1,-nbitq), 
to_sfixed(1215.0/65536.0,1,-nbitq), 
to_sfixed(268.0/65536.0,1,-nbitq), 
to_sfixed(-3092.0/65536.0,1,-nbitq), 
to_sfixed(-1089.0/65536.0,1,-nbitq), 
to_sfixed(-1441.0/65536.0,1,-nbitq), 
to_sfixed(-677.0/65536.0,1,-nbitq), 
to_sfixed(-1960.0/65536.0,1,-nbitq), 
to_sfixed(-361.0/65536.0,1,-nbitq), 
to_sfixed(-878.0/65536.0,1,-nbitq), 
to_sfixed(-4630.0/65536.0,1,-nbitq), 
to_sfixed(-1045.0/65536.0,1,-nbitq), 
to_sfixed(-299.0/65536.0,1,-nbitq), 
to_sfixed(2425.0/65536.0,1,-nbitq), 
to_sfixed(-727.0/65536.0,1,-nbitq), 
to_sfixed(2274.0/65536.0,1,-nbitq), 
to_sfixed(1192.0/65536.0,1,-nbitq), 
to_sfixed(-128.0/65536.0,1,-nbitq), 
to_sfixed(-1704.0/65536.0,1,-nbitq), 
to_sfixed(1866.0/65536.0,1,-nbitq), 
to_sfixed(1624.0/65536.0,1,-nbitq), 
to_sfixed(-1066.0/65536.0,1,-nbitq), 
to_sfixed(-1439.0/65536.0,1,-nbitq), 
to_sfixed(-726.0/65536.0,1,-nbitq), 
to_sfixed(-9.0/65536.0,1,-nbitq), 
to_sfixed(352.0/65536.0,1,-nbitq), 
to_sfixed(1844.0/65536.0,1,-nbitq), 
to_sfixed(6081.0/65536.0,1,-nbitq), 
to_sfixed(-1053.0/65536.0,1,-nbitq), 
to_sfixed(-2015.0/65536.0,1,-nbitq), 
to_sfixed(3144.0/65536.0,1,-nbitq), 
to_sfixed(694.0/65536.0,1,-nbitq), 
to_sfixed(2946.0/65536.0,1,-nbitq), 
to_sfixed(1016.0/65536.0,1,-nbitq), 
to_sfixed(1629.0/65536.0,1,-nbitq), 
to_sfixed(-1233.0/65536.0,1,-nbitq), 
to_sfixed(-1184.0/65536.0,1,-nbitq), 
to_sfixed(838.0/65536.0,1,-nbitq), 
to_sfixed(1968.0/65536.0,1,-nbitq), 
to_sfixed(2179.0/65536.0,1,-nbitq), 
to_sfixed(-1113.0/65536.0,1,-nbitq), 
to_sfixed(-2369.0/65536.0,1,-nbitq), 
to_sfixed(1350.0/65536.0,1,-nbitq), 
to_sfixed(337.0/65536.0,1,-nbitq), 
to_sfixed(-1477.0/65536.0,1,-nbitq), 
to_sfixed(452.0/65536.0,1,-nbitq), 
to_sfixed(-1986.0/65536.0,1,-nbitq), 
to_sfixed(4771.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1669.0/65536.0,1,-nbitq), 
to_sfixed(-2551.0/65536.0,1,-nbitq), 
to_sfixed(2563.0/65536.0,1,-nbitq), 
to_sfixed(-3728.0/65536.0,1,-nbitq), 
to_sfixed(-618.0/65536.0,1,-nbitq), 
to_sfixed(-2167.0/65536.0,1,-nbitq), 
to_sfixed(1038.0/65536.0,1,-nbitq), 
to_sfixed(-2606.0/65536.0,1,-nbitq), 
to_sfixed(-691.0/65536.0,1,-nbitq), 
to_sfixed(657.0/65536.0,1,-nbitq), 
to_sfixed(-3946.0/65536.0,1,-nbitq), 
to_sfixed(728.0/65536.0,1,-nbitq), 
to_sfixed(1578.0/65536.0,1,-nbitq), 
to_sfixed(-3535.0/65536.0,1,-nbitq), 
to_sfixed(1066.0/65536.0,1,-nbitq), 
to_sfixed(2218.0/65536.0,1,-nbitq), 
to_sfixed(-50.0/65536.0,1,-nbitq), 
to_sfixed(-2429.0/65536.0,1,-nbitq), 
to_sfixed(331.0/65536.0,1,-nbitq), 
to_sfixed(3334.0/65536.0,1,-nbitq), 
to_sfixed(-3434.0/65536.0,1,-nbitq), 
to_sfixed(2464.0/65536.0,1,-nbitq), 
to_sfixed(-884.0/65536.0,1,-nbitq), 
to_sfixed(-431.0/65536.0,1,-nbitq), 
to_sfixed(-45.0/65536.0,1,-nbitq), 
to_sfixed(-174.0/65536.0,1,-nbitq), 
to_sfixed(999.0/65536.0,1,-nbitq), 
to_sfixed(-329.0/65536.0,1,-nbitq), 
to_sfixed(-3066.0/65536.0,1,-nbitq), 
to_sfixed(-1728.0/65536.0,1,-nbitq), 
to_sfixed(-1936.0/65536.0,1,-nbitq), 
to_sfixed(2173.0/65536.0,1,-nbitq), 
to_sfixed(-1739.0/65536.0,1,-nbitq), 
to_sfixed(-630.0/65536.0,1,-nbitq), 
to_sfixed(1023.0/65536.0,1,-nbitq), 
to_sfixed(60.0/65536.0,1,-nbitq), 
to_sfixed(-1180.0/65536.0,1,-nbitq), 
to_sfixed(-3905.0/65536.0,1,-nbitq), 
to_sfixed(559.0/65536.0,1,-nbitq), 
to_sfixed(-821.0/65536.0,1,-nbitq), 
to_sfixed(-239.0/65536.0,1,-nbitq), 
to_sfixed(-477.0/65536.0,1,-nbitq), 
to_sfixed(-1133.0/65536.0,1,-nbitq), 
to_sfixed(-169.0/65536.0,1,-nbitq), 
to_sfixed(-938.0/65536.0,1,-nbitq), 
to_sfixed(4046.0/65536.0,1,-nbitq), 
to_sfixed(3219.0/65536.0,1,-nbitq), 
to_sfixed(-855.0/65536.0,1,-nbitq), 
to_sfixed(2691.0/65536.0,1,-nbitq), 
to_sfixed(4097.0/65536.0,1,-nbitq), 
to_sfixed(2409.0/65536.0,1,-nbitq), 
to_sfixed(1834.0/65536.0,1,-nbitq), 
to_sfixed(-466.0/65536.0,1,-nbitq), 
to_sfixed(2061.0/65536.0,1,-nbitq), 
to_sfixed(3646.0/65536.0,1,-nbitq), 
to_sfixed(2520.0/65536.0,1,-nbitq), 
to_sfixed(1861.0/65536.0,1,-nbitq), 
to_sfixed(-140.0/65536.0,1,-nbitq), 
to_sfixed(1977.0/65536.0,1,-nbitq), 
to_sfixed(5818.0/65536.0,1,-nbitq), 
to_sfixed(-3257.0/65536.0,1,-nbitq), 
to_sfixed(1139.0/65536.0,1,-nbitq), 
to_sfixed(-39.0/65536.0,1,-nbitq), 
to_sfixed(148.0/65536.0,1,-nbitq), 
to_sfixed(3884.0/65536.0,1,-nbitq), 
to_sfixed(2662.0/65536.0,1,-nbitq), 
to_sfixed(3229.0/65536.0,1,-nbitq), 
to_sfixed(-2037.0/65536.0,1,-nbitq), 
to_sfixed(-303.0/65536.0,1,-nbitq), 
to_sfixed(-666.0/65536.0,1,-nbitq), 
to_sfixed(-638.0/65536.0,1,-nbitq), 
to_sfixed(1471.0/65536.0,1,-nbitq), 
to_sfixed(72.0/65536.0,1,-nbitq), 
to_sfixed(2170.0/65536.0,1,-nbitq), 
to_sfixed(842.0/65536.0,1,-nbitq), 
to_sfixed(2393.0/65536.0,1,-nbitq), 
to_sfixed(-2253.0/65536.0,1,-nbitq), 
to_sfixed(-124.0/65536.0,1,-nbitq), 
to_sfixed(-2837.0/65536.0,1,-nbitq), 
to_sfixed(2930.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3.0/65536.0,1,-nbitq), 
to_sfixed(-236.0/65536.0,1,-nbitq), 
to_sfixed(-1038.0/65536.0,1,-nbitq), 
to_sfixed(-2648.0/65536.0,1,-nbitq), 
to_sfixed(-2214.0/65536.0,1,-nbitq), 
to_sfixed(149.0/65536.0,1,-nbitq), 
to_sfixed(1346.0/65536.0,1,-nbitq), 
to_sfixed(2596.0/65536.0,1,-nbitq), 
to_sfixed(-664.0/65536.0,1,-nbitq), 
to_sfixed(-178.0/65536.0,1,-nbitq), 
to_sfixed(-1933.0/65536.0,1,-nbitq), 
to_sfixed(-3614.0/65536.0,1,-nbitq), 
to_sfixed(333.0/65536.0,1,-nbitq), 
to_sfixed(-2713.0/65536.0,1,-nbitq), 
to_sfixed(-1937.0/65536.0,1,-nbitq), 
to_sfixed(1835.0/65536.0,1,-nbitq), 
to_sfixed(-400.0/65536.0,1,-nbitq), 
to_sfixed(204.0/65536.0,1,-nbitq), 
to_sfixed(-1302.0/65536.0,1,-nbitq), 
to_sfixed(104.0/65536.0,1,-nbitq), 
to_sfixed(-324.0/65536.0,1,-nbitq), 
to_sfixed(2080.0/65536.0,1,-nbitq), 
to_sfixed(2348.0/65536.0,1,-nbitq), 
to_sfixed(508.0/65536.0,1,-nbitq), 
to_sfixed(-818.0/65536.0,1,-nbitq), 
to_sfixed(-1429.0/65536.0,1,-nbitq), 
to_sfixed(-440.0/65536.0,1,-nbitq), 
to_sfixed(-1950.0/65536.0,1,-nbitq), 
to_sfixed(1408.0/65536.0,1,-nbitq), 
to_sfixed(-1283.0/65536.0,1,-nbitq), 
to_sfixed(-287.0/65536.0,1,-nbitq), 
to_sfixed(-2020.0/65536.0,1,-nbitq), 
to_sfixed(-5364.0/65536.0,1,-nbitq), 
to_sfixed(-1184.0/65536.0,1,-nbitq), 
to_sfixed(1824.0/65536.0,1,-nbitq), 
to_sfixed(-266.0/65536.0,1,-nbitq), 
to_sfixed(1697.0/65536.0,1,-nbitq), 
to_sfixed(-828.0/65536.0,1,-nbitq), 
to_sfixed(-1078.0/65536.0,1,-nbitq), 
to_sfixed(-2720.0/65536.0,1,-nbitq), 
to_sfixed(-2060.0/65536.0,1,-nbitq), 
to_sfixed(-1407.0/65536.0,1,-nbitq), 
to_sfixed(-472.0/65536.0,1,-nbitq), 
to_sfixed(2025.0/65536.0,1,-nbitq), 
to_sfixed(-1755.0/65536.0,1,-nbitq), 
to_sfixed(4594.0/65536.0,1,-nbitq), 
to_sfixed(-1938.0/65536.0,1,-nbitq), 
to_sfixed(1631.0/65536.0,1,-nbitq), 
to_sfixed(-1869.0/65536.0,1,-nbitq), 
to_sfixed(1083.0/65536.0,1,-nbitq), 
to_sfixed(2285.0/65536.0,1,-nbitq), 
to_sfixed(999.0/65536.0,1,-nbitq), 
to_sfixed(3595.0/65536.0,1,-nbitq), 
to_sfixed(-2104.0/65536.0,1,-nbitq), 
to_sfixed(1643.0/65536.0,1,-nbitq), 
to_sfixed(-1623.0/65536.0,1,-nbitq), 
to_sfixed(-488.0/65536.0,1,-nbitq), 
to_sfixed(2651.0/65536.0,1,-nbitq), 
to_sfixed(-1307.0/65536.0,1,-nbitq), 
to_sfixed(5165.0/65536.0,1,-nbitq), 
to_sfixed(49.0/65536.0,1,-nbitq), 
to_sfixed(-2959.0/65536.0,1,-nbitq), 
to_sfixed(53.0/65536.0,1,-nbitq), 
to_sfixed(676.0/65536.0,1,-nbitq), 
to_sfixed(3001.0/65536.0,1,-nbitq), 
to_sfixed(-1902.0/65536.0,1,-nbitq), 
to_sfixed(806.0/65536.0,1,-nbitq), 
to_sfixed(640.0/65536.0,1,-nbitq), 
to_sfixed(3565.0/65536.0,1,-nbitq), 
to_sfixed(3313.0/65536.0,1,-nbitq), 
to_sfixed(2304.0/65536.0,1,-nbitq), 
to_sfixed(1342.0/65536.0,1,-nbitq), 
to_sfixed(3613.0/65536.0,1,-nbitq), 
to_sfixed(1859.0/65536.0,1,-nbitq), 
to_sfixed(1360.0/65536.0,1,-nbitq), 
to_sfixed(-1074.0/65536.0,1,-nbitq), 
to_sfixed(-2992.0/65536.0,1,-nbitq), 
to_sfixed(2506.0/65536.0,1,-nbitq), 
to_sfixed(-2603.0/65536.0,1,-nbitq), 
to_sfixed(1897.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1707.0/65536.0,1,-nbitq), 
to_sfixed(-183.0/65536.0,1,-nbitq), 
to_sfixed(6182.0/65536.0,1,-nbitq), 
to_sfixed(1629.0/65536.0,1,-nbitq), 
to_sfixed(-352.0/65536.0,1,-nbitq), 
to_sfixed(-3019.0/65536.0,1,-nbitq), 
to_sfixed(-2650.0/65536.0,1,-nbitq), 
to_sfixed(1692.0/65536.0,1,-nbitq), 
to_sfixed(-2784.0/65536.0,1,-nbitq), 
to_sfixed(636.0/65536.0,1,-nbitq), 
to_sfixed(-2695.0/65536.0,1,-nbitq), 
to_sfixed(-2667.0/65536.0,1,-nbitq), 
to_sfixed(-2609.0/65536.0,1,-nbitq), 
to_sfixed(-1394.0/65536.0,1,-nbitq), 
to_sfixed(-1439.0/65536.0,1,-nbitq), 
to_sfixed(-848.0/65536.0,1,-nbitq), 
to_sfixed(2566.0/65536.0,1,-nbitq), 
to_sfixed(-646.0/65536.0,1,-nbitq), 
to_sfixed(-1324.0/65536.0,1,-nbitq), 
to_sfixed(-287.0/65536.0,1,-nbitq), 
to_sfixed(805.0/65536.0,1,-nbitq), 
to_sfixed(2153.0/65536.0,1,-nbitq), 
to_sfixed(-2967.0/65536.0,1,-nbitq), 
to_sfixed(-361.0/65536.0,1,-nbitq), 
to_sfixed(-2605.0/65536.0,1,-nbitq), 
to_sfixed(2493.0/65536.0,1,-nbitq), 
to_sfixed(-30.0/65536.0,1,-nbitq), 
to_sfixed(-1647.0/65536.0,1,-nbitq), 
to_sfixed(318.0/65536.0,1,-nbitq), 
to_sfixed(-2802.0/65536.0,1,-nbitq), 
to_sfixed(-727.0/65536.0,1,-nbitq), 
to_sfixed(2088.0/65536.0,1,-nbitq), 
to_sfixed(-1778.0/65536.0,1,-nbitq), 
to_sfixed(-2842.0/65536.0,1,-nbitq), 
to_sfixed(2151.0/65536.0,1,-nbitq), 
to_sfixed(-1240.0/65536.0,1,-nbitq), 
to_sfixed(803.0/65536.0,1,-nbitq), 
to_sfixed(-2816.0/65536.0,1,-nbitq), 
to_sfixed(4714.0/65536.0,1,-nbitq), 
to_sfixed(2157.0/65536.0,1,-nbitq), 
to_sfixed(2385.0/65536.0,1,-nbitq), 
to_sfixed(1152.0/65536.0,1,-nbitq), 
to_sfixed(-15.0/65536.0,1,-nbitq), 
to_sfixed(-388.0/65536.0,1,-nbitq), 
to_sfixed(-1863.0/65536.0,1,-nbitq), 
to_sfixed(808.0/65536.0,1,-nbitq), 
to_sfixed(1974.0/65536.0,1,-nbitq), 
to_sfixed(-2669.0/65536.0,1,-nbitq), 
to_sfixed(929.0/65536.0,1,-nbitq), 
to_sfixed(3583.0/65536.0,1,-nbitq), 
to_sfixed(3076.0/65536.0,1,-nbitq), 
to_sfixed(661.0/65536.0,1,-nbitq), 
to_sfixed(-1568.0/65536.0,1,-nbitq), 
to_sfixed(-1984.0/65536.0,1,-nbitq), 
to_sfixed(-676.0/65536.0,1,-nbitq), 
to_sfixed(-1003.0/65536.0,1,-nbitq), 
to_sfixed(2989.0/65536.0,1,-nbitq), 
to_sfixed(-2782.0/65536.0,1,-nbitq), 
to_sfixed(1290.0/65536.0,1,-nbitq), 
to_sfixed(1731.0/65536.0,1,-nbitq), 
to_sfixed(-1217.0/65536.0,1,-nbitq), 
to_sfixed(-2548.0/65536.0,1,-nbitq), 
to_sfixed(-2496.0/65536.0,1,-nbitq), 
to_sfixed(1798.0/65536.0,1,-nbitq), 
to_sfixed(1816.0/65536.0,1,-nbitq), 
to_sfixed(2619.0/65536.0,1,-nbitq), 
to_sfixed(-234.0/65536.0,1,-nbitq), 
to_sfixed(-3559.0/65536.0,1,-nbitq), 
to_sfixed(548.0/65536.0,1,-nbitq), 
to_sfixed(-2417.0/65536.0,1,-nbitq), 
to_sfixed(1647.0/65536.0,1,-nbitq), 
to_sfixed(307.0/65536.0,1,-nbitq), 
to_sfixed(2202.0/65536.0,1,-nbitq), 
to_sfixed(1310.0/65536.0,1,-nbitq), 
to_sfixed(851.0/65536.0,1,-nbitq), 
to_sfixed(388.0/65536.0,1,-nbitq), 
to_sfixed(1425.0/65536.0,1,-nbitq), 
to_sfixed(-202.0/65536.0,1,-nbitq), 
to_sfixed(-2993.0/65536.0,1,-nbitq), 
to_sfixed(1871.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2843.0/65536.0,1,-nbitq), 
to_sfixed(2162.0/65536.0,1,-nbitq), 
to_sfixed(450.0/65536.0,1,-nbitq), 
to_sfixed(-2951.0/65536.0,1,-nbitq), 
to_sfixed(-1551.0/65536.0,1,-nbitq), 
to_sfixed(-3234.0/65536.0,1,-nbitq), 
to_sfixed(1851.0/65536.0,1,-nbitq), 
to_sfixed(-2299.0/65536.0,1,-nbitq), 
to_sfixed(-2549.0/65536.0,1,-nbitq), 
to_sfixed(-1357.0/65536.0,1,-nbitq), 
to_sfixed(-375.0/65536.0,1,-nbitq), 
to_sfixed(-2827.0/65536.0,1,-nbitq), 
to_sfixed(3003.0/65536.0,1,-nbitq), 
to_sfixed(1032.0/65536.0,1,-nbitq), 
to_sfixed(1984.0/65536.0,1,-nbitq), 
to_sfixed(-2308.0/65536.0,1,-nbitq), 
to_sfixed(-649.0/65536.0,1,-nbitq), 
to_sfixed(-5909.0/65536.0,1,-nbitq), 
to_sfixed(847.0/65536.0,1,-nbitq), 
to_sfixed(1761.0/65536.0,1,-nbitq), 
to_sfixed(1159.0/65536.0,1,-nbitq), 
to_sfixed(-2865.0/65536.0,1,-nbitq), 
to_sfixed(1065.0/65536.0,1,-nbitq), 
to_sfixed(-902.0/65536.0,1,-nbitq), 
to_sfixed(-1142.0/65536.0,1,-nbitq), 
to_sfixed(3786.0/65536.0,1,-nbitq), 
to_sfixed(-4551.0/65536.0,1,-nbitq), 
to_sfixed(-1350.0/65536.0,1,-nbitq), 
to_sfixed(-1304.0/65536.0,1,-nbitq), 
to_sfixed(-423.0/65536.0,1,-nbitq), 
to_sfixed(-995.0/65536.0,1,-nbitq), 
to_sfixed(-733.0/65536.0,1,-nbitq), 
to_sfixed(-3371.0/65536.0,1,-nbitq), 
to_sfixed(-1624.0/65536.0,1,-nbitq), 
to_sfixed(1012.0/65536.0,1,-nbitq), 
to_sfixed(-1969.0/65536.0,1,-nbitq), 
to_sfixed(717.0/65536.0,1,-nbitq), 
to_sfixed(-3988.0/65536.0,1,-nbitq), 
to_sfixed(3777.0/65536.0,1,-nbitq), 
to_sfixed(-2404.0/65536.0,1,-nbitq), 
to_sfixed(-646.0/65536.0,1,-nbitq), 
to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(-3704.0/65536.0,1,-nbitq), 
to_sfixed(950.0/65536.0,1,-nbitq), 
to_sfixed(-1598.0/65536.0,1,-nbitq), 
to_sfixed(2813.0/65536.0,1,-nbitq), 
to_sfixed(-1666.0/65536.0,1,-nbitq), 
to_sfixed(-662.0/65536.0,1,-nbitq), 
to_sfixed(2875.0/65536.0,1,-nbitq), 
to_sfixed(-1962.0/65536.0,1,-nbitq), 
to_sfixed(1475.0/65536.0,1,-nbitq), 
to_sfixed(-8.0/65536.0,1,-nbitq), 
to_sfixed(2936.0/65536.0,1,-nbitq), 
to_sfixed(-3045.0/65536.0,1,-nbitq), 
to_sfixed(38.0/65536.0,1,-nbitq), 
to_sfixed(2635.0/65536.0,1,-nbitq), 
to_sfixed(2145.0/65536.0,1,-nbitq), 
to_sfixed(1923.0/65536.0,1,-nbitq), 
to_sfixed(2267.0/65536.0,1,-nbitq), 
to_sfixed(912.0/65536.0,1,-nbitq), 
to_sfixed(-1876.0/65536.0,1,-nbitq), 
to_sfixed(1033.0/65536.0,1,-nbitq), 
to_sfixed(919.0/65536.0,1,-nbitq), 
to_sfixed(1614.0/65536.0,1,-nbitq), 
to_sfixed(2341.0/65536.0,1,-nbitq), 
to_sfixed(-1180.0/65536.0,1,-nbitq), 
to_sfixed(-1698.0/65536.0,1,-nbitq), 
to_sfixed(-6001.0/65536.0,1,-nbitq), 
to_sfixed(4176.0/65536.0,1,-nbitq), 
to_sfixed(445.0/65536.0,1,-nbitq), 
to_sfixed(-2703.0/65536.0,1,-nbitq), 
to_sfixed(-719.0/65536.0,1,-nbitq), 
to_sfixed(-1142.0/65536.0,1,-nbitq), 
to_sfixed(-2860.0/65536.0,1,-nbitq), 
to_sfixed(289.0/65536.0,1,-nbitq), 
to_sfixed(-2529.0/65536.0,1,-nbitq), 
to_sfixed(725.0/65536.0,1,-nbitq), 
to_sfixed(-1273.0/65536.0,1,-nbitq), 
to_sfixed(-299.0/65536.0,1,-nbitq), 
to_sfixed(-160.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1127.0/65536.0,1,-nbitq), 
to_sfixed(3563.0/65536.0,1,-nbitq), 
to_sfixed(-1071.0/65536.0,1,-nbitq), 
to_sfixed(2986.0/65536.0,1,-nbitq), 
to_sfixed(1902.0/65536.0,1,-nbitq), 
to_sfixed(-3336.0/65536.0,1,-nbitq), 
to_sfixed(1999.0/65536.0,1,-nbitq), 
to_sfixed(900.0/65536.0,1,-nbitq), 
to_sfixed(-1447.0/65536.0,1,-nbitq), 
to_sfixed(-1707.0/65536.0,1,-nbitq), 
to_sfixed(-1261.0/65536.0,1,-nbitq), 
to_sfixed(-2684.0/65536.0,1,-nbitq), 
to_sfixed(-1308.0/65536.0,1,-nbitq), 
to_sfixed(2210.0/65536.0,1,-nbitq), 
to_sfixed(-5047.0/65536.0,1,-nbitq), 
to_sfixed(3077.0/65536.0,1,-nbitq), 
to_sfixed(2063.0/65536.0,1,-nbitq), 
to_sfixed(-2250.0/65536.0,1,-nbitq), 
to_sfixed(2051.0/65536.0,1,-nbitq), 
to_sfixed(-826.0/65536.0,1,-nbitq), 
to_sfixed(2812.0/65536.0,1,-nbitq), 
to_sfixed(-1710.0/65536.0,1,-nbitq), 
to_sfixed(-4393.0/65536.0,1,-nbitq), 
to_sfixed(-2048.0/65536.0,1,-nbitq), 
to_sfixed(-2427.0/65536.0,1,-nbitq), 
to_sfixed(2416.0/65536.0,1,-nbitq), 
to_sfixed(-1195.0/65536.0,1,-nbitq), 
to_sfixed(1115.0/65536.0,1,-nbitq), 
to_sfixed(-2117.0/65536.0,1,-nbitq), 
to_sfixed(154.0/65536.0,1,-nbitq), 
to_sfixed(-2577.0/65536.0,1,-nbitq), 
to_sfixed(-4065.0/65536.0,1,-nbitq), 
to_sfixed(-1605.0/65536.0,1,-nbitq), 
to_sfixed(-1995.0/65536.0,1,-nbitq), 
to_sfixed(-2067.0/65536.0,1,-nbitq), 
to_sfixed(2636.0/65536.0,1,-nbitq), 
to_sfixed(-4372.0/65536.0,1,-nbitq), 
to_sfixed(1916.0/65536.0,1,-nbitq), 
to_sfixed(2638.0/65536.0,1,-nbitq), 
to_sfixed(-986.0/65536.0,1,-nbitq), 
to_sfixed(-1829.0/65536.0,1,-nbitq), 
to_sfixed(2473.0/65536.0,1,-nbitq), 
to_sfixed(1410.0/65536.0,1,-nbitq), 
to_sfixed(-2745.0/65536.0,1,-nbitq), 
to_sfixed(-287.0/65536.0,1,-nbitq), 
to_sfixed(1108.0/65536.0,1,-nbitq), 
to_sfixed(1506.0/65536.0,1,-nbitq), 
to_sfixed(1912.0/65536.0,1,-nbitq), 
to_sfixed(3256.0/65536.0,1,-nbitq), 
to_sfixed(2049.0/65536.0,1,-nbitq), 
to_sfixed(1118.0/65536.0,1,-nbitq), 
to_sfixed(3881.0/65536.0,1,-nbitq), 
to_sfixed(-537.0/65536.0,1,-nbitq), 
to_sfixed(2145.0/65536.0,1,-nbitq), 
to_sfixed(1932.0/65536.0,1,-nbitq), 
to_sfixed(1102.0/65536.0,1,-nbitq), 
to_sfixed(-313.0/65536.0,1,-nbitq), 
to_sfixed(-2419.0/65536.0,1,-nbitq), 
to_sfixed(2225.0/65536.0,1,-nbitq), 
to_sfixed(1464.0/65536.0,1,-nbitq), 
to_sfixed(320.0/65536.0,1,-nbitq), 
to_sfixed(245.0/65536.0,1,-nbitq), 
to_sfixed(3161.0/65536.0,1,-nbitq), 
to_sfixed(-2435.0/65536.0,1,-nbitq), 
to_sfixed(2910.0/65536.0,1,-nbitq), 
to_sfixed(-3876.0/65536.0,1,-nbitq), 
to_sfixed(-2423.0/65536.0,1,-nbitq), 
to_sfixed(-1946.0/65536.0,1,-nbitq), 
to_sfixed(6365.0/65536.0,1,-nbitq), 
to_sfixed(7071.0/65536.0,1,-nbitq), 
to_sfixed(-3173.0/65536.0,1,-nbitq), 
to_sfixed(-3903.0/65536.0,1,-nbitq), 
to_sfixed(1774.0/65536.0,1,-nbitq), 
to_sfixed(1234.0/65536.0,1,-nbitq), 
to_sfixed(-2078.0/65536.0,1,-nbitq), 
to_sfixed(554.0/65536.0,1,-nbitq), 
to_sfixed(-5549.0/65536.0,1,-nbitq), 
to_sfixed(1176.0/65536.0,1,-nbitq), 
to_sfixed(-3009.0/65536.0,1,-nbitq), 
to_sfixed(-987.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2669.0/65536.0,1,-nbitq), 
to_sfixed(1134.0/65536.0,1,-nbitq), 
to_sfixed(1563.0/65536.0,1,-nbitq), 
to_sfixed(4330.0/65536.0,1,-nbitq), 
to_sfixed(-1658.0/65536.0,1,-nbitq), 
to_sfixed(933.0/65536.0,1,-nbitq), 
to_sfixed(2385.0/65536.0,1,-nbitq), 
to_sfixed(-2379.0/65536.0,1,-nbitq), 
to_sfixed(-3463.0/65536.0,1,-nbitq), 
to_sfixed(-2160.0/65536.0,1,-nbitq), 
to_sfixed(-1366.0/65536.0,1,-nbitq), 
to_sfixed(78.0/65536.0,1,-nbitq), 
to_sfixed(1018.0/65536.0,1,-nbitq), 
to_sfixed(-429.0/65536.0,1,-nbitq), 
to_sfixed(-3110.0/65536.0,1,-nbitq), 
to_sfixed(1956.0/65536.0,1,-nbitq), 
to_sfixed(-427.0/65536.0,1,-nbitq), 
to_sfixed(-2224.0/65536.0,1,-nbitq), 
to_sfixed(-5630.0/65536.0,1,-nbitq), 
to_sfixed(1179.0/65536.0,1,-nbitq), 
to_sfixed(5205.0/65536.0,1,-nbitq), 
to_sfixed(-668.0/65536.0,1,-nbitq), 
to_sfixed(-1965.0/65536.0,1,-nbitq), 
to_sfixed(-1990.0/65536.0,1,-nbitq), 
to_sfixed(1796.0/65536.0,1,-nbitq), 
to_sfixed(389.0/65536.0,1,-nbitq), 
to_sfixed(-268.0/65536.0,1,-nbitq), 
to_sfixed(2369.0/65536.0,1,-nbitq), 
to_sfixed(2691.0/65536.0,1,-nbitq), 
to_sfixed(-6015.0/65536.0,1,-nbitq), 
to_sfixed(2573.0/65536.0,1,-nbitq), 
to_sfixed(-653.0/65536.0,1,-nbitq), 
to_sfixed(1121.0/65536.0,1,-nbitq), 
to_sfixed(5848.0/65536.0,1,-nbitq), 
to_sfixed(-2340.0/65536.0,1,-nbitq), 
to_sfixed(-813.0/65536.0,1,-nbitq), 
to_sfixed(-2841.0/65536.0,1,-nbitq), 
to_sfixed(-943.0/65536.0,1,-nbitq), 
to_sfixed(-2154.0/65536.0,1,-nbitq), 
to_sfixed(-2266.0/65536.0,1,-nbitq), 
to_sfixed(3001.0/65536.0,1,-nbitq), 
to_sfixed(1398.0/65536.0,1,-nbitq), 
to_sfixed(2932.0/65536.0,1,-nbitq), 
to_sfixed(-2732.0/65536.0,1,-nbitq), 
to_sfixed(1534.0/65536.0,1,-nbitq), 
to_sfixed(2422.0/65536.0,1,-nbitq), 
to_sfixed(739.0/65536.0,1,-nbitq), 
to_sfixed(-173.0/65536.0,1,-nbitq), 
to_sfixed(3123.0/65536.0,1,-nbitq), 
to_sfixed(1844.0/65536.0,1,-nbitq), 
to_sfixed(2806.0/65536.0,1,-nbitq), 
to_sfixed(3263.0/65536.0,1,-nbitq), 
to_sfixed(-2796.0/65536.0,1,-nbitq), 
to_sfixed(1318.0/65536.0,1,-nbitq), 
to_sfixed(1911.0/65536.0,1,-nbitq), 
to_sfixed(-1045.0/65536.0,1,-nbitq), 
to_sfixed(1909.0/65536.0,1,-nbitq), 
to_sfixed(-2105.0/65536.0,1,-nbitq), 
to_sfixed(-2373.0/65536.0,1,-nbitq), 
to_sfixed(-801.0/65536.0,1,-nbitq), 
to_sfixed(-873.0/65536.0,1,-nbitq), 
to_sfixed(294.0/65536.0,1,-nbitq), 
to_sfixed(-1381.0/65536.0,1,-nbitq), 
to_sfixed(-1737.0/65536.0,1,-nbitq), 
to_sfixed(1002.0/65536.0,1,-nbitq), 
to_sfixed(-1015.0/65536.0,1,-nbitq), 
to_sfixed(-428.0/65536.0,1,-nbitq), 
to_sfixed(-2713.0/65536.0,1,-nbitq), 
to_sfixed(5511.0/65536.0,1,-nbitq), 
to_sfixed(4382.0/65536.0,1,-nbitq), 
to_sfixed(-557.0/65536.0,1,-nbitq), 
to_sfixed(-2476.0/65536.0,1,-nbitq), 
to_sfixed(-852.0/65536.0,1,-nbitq), 
to_sfixed(-276.0/65536.0,1,-nbitq), 
to_sfixed(93.0/65536.0,1,-nbitq), 
to_sfixed(-905.0/65536.0,1,-nbitq), 
to_sfixed(-9161.0/65536.0,1,-nbitq), 
to_sfixed(-1925.0/65536.0,1,-nbitq), 
to_sfixed(-672.0/65536.0,1,-nbitq), 
to_sfixed(-170.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1569.0/65536.0,1,-nbitq), 
to_sfixed(717.0/65536.0,1,-nbitq), 
to_sfixed(752.0/65536.0,1,-nbitq), 
to_sfixed(4738.0/65536.0,1,-nbitq), 
to_sfixed(2056.0/65536.0,1,-nbitq), 
to_sfixed(-3285.0/65536.0,1,-nbitq), 
to_sfixed(-1931.0/65536.0,1,-nbitq), 
to_sfixed(-4031.0/65536.0,1,-nbitq), 
to_sfixed(-4126.0/65536.0,1,-nbitq), 
to_sfixed(868.0/65536.0,1,-nbitq), 
to_sfixed(2437.0/65536.0,1,-nbitq), 
to_sfixed(-553.0/65536.0,1,-nbitq), 
to_sfixed(-860.0/65536.0,1,-nbitq), 
to_sfixed(1259.0/65536.0,1,-nbitq), 
to_sfixed(-2424.0/65536.0,1,-nbitq), 
to_sfixed(-1803.0/65536.0,1,-nbitq), 
to_sfixed(-3168.0/65536.0,1,-nbitq), 
to_sfixed(-4470.0/65536.0,1,-nbitq), 
to_sfixed(-7625.0/65536.0,1,-nbitq), 
to_sfixed(761.0/65536.0,1,-nbitq), 
to_sfixed(5816.0/65536.0,1,-nbitq), 
to_sfixed(389.0/65536.0,1,-nbitq), 
to_sfixed(-2008.0/65536.0,1,-nbitq), 
to_sfixed(-9599.0/65536.0,1,-nbitq), 
to_sfixed(2717.0/65536.0,1,-nbitq), 
to_sfixed(-10877.0/65536.0,1,-nbitq), 
to_sfixed(-680.0/65536.0,1,-nbitq), 
to_sfixed(-348.0/65536.0,1,-nbitq), 
to_sfixed(5747.0/65536.0,1,-nbitq), 
to_sfixed(-2458.0/65536.0,1,-nbitq), 
to_sfixed(3223.0/65536.0,1,-nbitq), 
to_sfixed(-906.0/65536.0,1,-nbitq), 
to_sfixed(2496.0/65536.0,1,-nbitq), 
to_sfixed(3791.0/65536.0,1,-nbitq), 
to_sfixed(1332.0/65536.0,1,-nbitq), 
to_sfixed(-1394.0/65536.0,1,-nbitq), 
to_sfixed(-839.0/65536.0,1,-nbitq), 
to_sfixed(2281.0/65536.0,1,-nbitq), 
to_sfixed(4759.0/65536.0,1,-nbitq), 
to_sfixed(-3741.0/65536.0,1,-nbitq), 
to_sfixed(4549.0/65536.0,1,-nbitq), 
to_sfixed(1144.0/65536.0,1,-nbitq), 
to_sfixed(9001.0/65536.0,1,-nbitq), 
to_sfixed(-1562.0/65536.0,1,-nbitq), 
to_sfixed(-2277.0/65536.0,1,-nbitq), 
to_sfixed(-1992.0/65536.0,1,-nbitq), 
to_sfixed(3773.0/65536.0,1,-nbitq), 
to_sfixed(-2522.0/65536.0,1,-nbitq), 
to_sfixed(1287.0/65536.0,1,-nbitq), 
to_sfixed(599.0/65536.0,1,-nbitq), 
to_sfixed(1409.0/65536.0,1,-nbitq), 
to_sfixed(-2608.0/65536.0,1,-nbitq), 
to_sfixed(-2674.0/65536.0,1,-nbitq), 
to_sfixed(1123.0/65536.0,1,-nbitq), 
to_sfixed(-802.0/65536.0,1,-nbitq), 
to_sfixed(-3186.0/65536.0,1,-nbitq), 
to_sfixed(-2387.0/65536.0,1,-nbitq), 
to_sfixed(443.0/65536.0,1,-nbitq), 
to_sfixed(-600.0/65536.0,1,-nbitq), 
to_sfixed(-9833.0/65536.0,1,-nbitq), 
to_sfixed(-2737.0/65536.0,1,-nbitq), 
to_sfixed(-1510.0/65536.0,1,-nbitq), 
to_sfixed(2259.0/65536.0,1,-nbitq), 
to_sfixed(2142.0/65536.0,1,-nbitq), 
to_sfixed(-3925.0/65536.0,1,-nbitq), 
to_sfixed(-821.0/65536.0,1,-nbitq), 
to_sfixed(369.0/65536.0,1,-nbitq), 
to_sfixed(179.0/65536.0,1,-nbitq), 
to_sfixed(10170.0/65536.0,1,-nbitq), 
to_sfixed(1066.0/65536.0,1,-nbitq), 
to_sfixed(-1294.0/65536.0,1,-nbitq), 
to_sfixed(-1074.0/65536.0,1,-nbitq), 
to_sfixed(375.0/65536.0,1,-nbitq), 
to_sfixed(518.0/65536.0,1,-nbitq), 
to_sfixed(2126.0/65536.0,1,-nbitq), 
to_sfixed(-3832.0/65536.0,1,-nbitq), 
to_sfixed(-258.0/65536.0,1,-nbitq), 
to_sfixed(-702.0/65536.0,1,-nbitq), 
to_sfixed(-1413.0/65536.0,1,-nbitq), 
to_sfixed(-2380.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1130.0/65536.0,1,-nbitq), 
to_sfixed(-4029.0/65536.0,1,-nbitq), 
to_sfixed(-2613.0/65536.0,1,-nbitq), 
to_sfixed(-1783.0/65536.0,1,-nbitq), 
to_sfixed(2835.0/65536.0,1,-nbitq), 
to_sfixed(-1491.0/65536.0,1,-nbitq), 
to_sfixed(-4498.0/65536.0,1,-nbitq), 
to_sfixed(3645.0/65536.0,1,-nbitq), 
to_sfixed(-5289.0/65536.0,1,-nbitq), 
to_sfixed(1514.0/65536.0,1,-nbitq), 
to_sfixed(-3344.0/65536.0,1,-nbitq), 
to_sfixed(-3842.0/65536.0,1,-nbitq), 
to_sfixed(-401.0/65536.0,1,-nbitq), 
to_sfixed(2698.0/65536.0,1,-nbitq), 
to_sfixed(-786.0/65536.0,1,-nbitq), 
to_sfixed(1310.0/65536.0,1,-nbitq), 
to_sfixed(1306.0/65536.0,1,-nbitq), 
to_sfixed(-859.0/65536.0,1,-nbitq), 
to_sfixed(-2345.0/65536.0,1,-nbitq), 
to_sfixed(2128.0/65536.0,1,-nbitq), 
to_sfixed(6316.0/65536.0,1,-nbitq), 
to_sfixed(-687.0/65536.0,1,-nbitq), 
to_sfixed(-3641.0/65536.0,1,-nbitq), 
to_sfixed(-13639.0/65536.0,1,-nbitq), 
to_sfixed(6728.0/65536.0,1,-nbitq), 
to_sfixed(-16206.0/65536.0,1,-nbitq), 
to_sfixed(-1597.0/65536.0,1,-nbitq), 
to_sfixed(1099.0/65536.0,1,-nbitq), 
to_sfixed(3448.0/65536.0,1,-nbitq), 
to_sfixed(-6198.0/65536.0,1,-nbitq), 
to_sfixed(2396.0/65536.0,1,-nbitq), 
to_sfixed(-1758.0/65536.0,1,-nbitq), 
to_sfixed(3741.0/65536.0,1,-nbitq), 
to_sfixed(-3351.0/65536.0,1,-nbitq), 
to_sfixed(2169.0/65536.0,1,-nbitq), 
to_sfixed(1536.0/65536.0,1,-nbitq), 
to_sfixed(1737.0/65536.0,1,-nbitq), 
to_sfixed(1050.0/65536.0,1,-nbitq), 
to_sfixed(4969.0/65536.0,1,-nbitq), 
to_sfixed(-2533.0/65536.0,1,-nbitq), 
to_sfixed(4638.0/65536.0,1,-nbitq), 
to_sfixed(-340.0/65536.0,1,-nbitq), 
to_sfixed(3854.0/65536.0,1,-nbitq), 
to_sfixed(-3249.0/65536.0,1,-nbitq), 
to_sfixed(-1189.0/65536.0,1,-nbitq), 
to_sfixed(-822.0/65536.0,1,-nbitq), 
to_sfixed(3791.0/65536.0,1,-nbitq), 
to_sfixed(-6961.0/65536.0,1,-nbitq), 
to_sfixed(-1359.0/65536.0,1,-nbitq), 
to_sfixed(1734.0/65536.0,1,-nbitq), 
to_sfixed(-2492.0/65536.0,1,-nbitq), 
to_sfixed(1721.0/65536.0,1,-nbitq), 
to_sfixed(-4364.0/65536.0,1,-nbitq), 
to_sfixed(3027.0/65536.0,1,-nbitq), 
to_sfixed(-4300.0/65536.0,1,-nbitq), 
to_sfixed(-5782.0/65536.0,1,-nbitq), 
to_sfixed(-271.0/65536.0,1,-nbitq), 
to_sfixed(2969.0/65536.0,1,-nbitq), 
to_sfixed(2174.0/65536.0,1,-nbitq), 
to_sfixed(-13693.0/65536.0,1,-nbitq), 
to_sfixed(2163.0/65536.0,1,-nbitq), 
to_sfixed(-2742.0/65536.0,1,-nbitq), 
to_sfixed(-2456.0/65536.0,1,-nbitq), 
to_sfixed(2056.0/65536.0,1,-nbitq), 
to_sfixed(377.0/65536.0,1,-nbitq), 
to_sfixed(1954.0/65536.0,1,-nbitq), 
to_sfixed(1215.0/65536.0,1,-nbitq), 
to_sfixed(699.0/65536.0,1,-nbitq), 
to_sfixed(9572.0/65536.0,1,-nbitq), 
to_sfixed(-2170.0/65536.0,1,-nbitq), 
to_sfixed(-551.0/65536.0,1,-nbitq), 
to_sfixed(-3767.0/65536.0,1,-nbitq), 
to_sfixed(-362.0/65536.0,1,-nbitq), 
to_sfixed(1110.0/65536.0,1,-nbitq), 
to_sfixed(50.0/65536.0,1,-nbitq), 
to_sfixed(-3729.0/65536.0,1,-nbitq), 
to_sfixed(6174.0/65536.0,1,-nbitq), 
to_sfixed(-190.0/65536.0,1,-nbitq), 
to_sfixed(-967.0/65536.0,1,-nbitq), 
to_sfixed(-7074.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3631.0/65536.0,1,-nbitq), 
to_sfixed(-4630.0/65536.0,1,-nbitq), 
to_sfixed(-669.0/65536.0,1,-nbitq), 
to_sfixed(-5331.0/65536.0,1,-nbitq), 
to_sfixed(2303.0/65536.0,1,-nbitq), 
to_sfixed(456.0/65536.0,1,-nbitq), 
to_sfixed(-6832.0/65536.0,1,-nbitq), 
to_sfixed(4179.0/65536.0,1,-nbitq), 
to_sfixed(5375.0/65536.0,1,-nbitq), 
to_sfixed(2479.0/65536.0,1,-nbitq), 
to_sfixed(-3063.0/65536.0,1,-nbitq), 
to_sfixed(-6665.0/65536.0,1,-nbitq), 
to_sfixed(-2337.0/65536.0,1,-nbitq), 
to_sfixed(-893.0/65536.0,1,-nbitq), 
to_sfixed(182.0/65536.0,1,-nbitq), 
to_sfixed(3078.0/65536.0,1,-nbitq), 
to_sfixed(635.0/65536.0,1,-nbitq), 
to_sfixed(7160.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(-2420.0/65536.0,1,-nbitq), 
to_sfixed(7569.0/65536.0,1,-nbitq), 
to_sfixed(1296.0/65536.0,1,-nbitq), 
to_sfixed(-6715.0/65536.0,1,-nbitq), 
to_sfixed(-13920.0/65536.0,1,-nbitq), 
to_sfixed(2496.0/65536.0,1,-nbitq), 
to_sfixed(-18163.0/65536.0,1,-nbitq), 
to_sfixed(4436.0/65536.0,1,-nbitq), 
to_sfixed(2362.0/65536.0,1,-nbitq), 
to_sfixed(-51.0/65536.0,1,-nbitq), 
to_sfixed(4045.0/65536.0,1,-nbitq), 
to_sfixed(-4598.0/65536.0,1,-nbitq), 
to_sfixed(-2527.0/65536.0,1,-nbitq), 
to_sfixed(1458.0/65536.0,1,-nbitq), 
to_sfixed(1393.0/65536.0,1,-nbitq), 
to_sfixed(1711.0/65536.0,1,-nbitq), 
to_sfixed(-2076.0/65536.0,1,-nbitq), 
to_sfixed(-2632.0/65536.0,1,-nbitq), 
to_sfixed(2151.0/65536.0,1,-nbitq), 
to_sfixed(-74.0/65536.0,1,-nbitq), 
to_sfixed(167.0/65536.0,1,-nbitq), 
to_sfixed(-130.0/65536.0,1,-nbitq), 
to_sfixed(2105.0/65536.0,1,-nbitq), 
to_sfixed(8381.0/65536.0,1,-nbitq), 
to_sfixed(-3548.0/65536.0,1,-nbitq), 
to_sfixed(-2192.0/65536.0,1,-nbitq), 
to_sfixed(-1559.0/65536.0,1,-nbitq), 
to_sfixed(320.0/65536.0,1,-nbitq), 
to_sfixed(-4629.0/65536.0,1,-nbitq), 
to_sfixed(2442.0/65536.0,1,-nbitq), 
to_sfixed(5494.0/65536.0,1,-nbitq), 
to_sfixed(2902.0/65536.0,1,-nbitq), 
to_sfixed(-2407.0/65536.0,1,-nbitq), 
to_sfixed(-2513.0/65536.0,1,-nbitq), 
to_sfixed(1029.0/65536.0,1,-nbitq), 
to_sfixed(-863.0/65536.0,1,-nbitq), 
to_sfixed(-4493.0/65536.0,1,-nbitq), 
to_sfixed(-2403.0/65536.0,1,-nbitq), 
to_sfixed(-95.0/65536.0,1,-nbitq), 
to_sfixed(521.0/65536.0,1,-nbitq), 
to_sfixed(-7046.0/65536.0,1,-nbitq), 
to_sfixed(8305.0/65536.0,1,-nbitq), 
to_sfixed(-341.0/65536.0,1,-nbitq), 
to_sfixed(2568.0/65536.0,1,-nbitq), 
to_sfixed(-2672.0/65536.0,1,-nbitq), 
to_sfixed(-4565.0/65536.0,1,-nbitq), 
to_sfixed(2670.0/65536.0,1,-nbitq), 
to_sfixed(3560.0/65536.0,1,-nbitq), 
to_sfixed(-2061.0/65536.0,1,-nbitq), 
to_sfixed(9321.0/65536.0,1,-nbitq), 
to_sfixed(2144.0/65536.0,1,-nbitq), 
to_sfixed(345.0/65536.0,1,-nbitq), 
to_sfixed(-5539.0/65536.0,1,-nbitq), 
to_sfixed(-323.0/65536.0,1,-nbitq), 
to_sfixed(-258.0/65536.0,1,-nbitq), 
to_sfixed(-2632.0/65536.0,1,-nbitq), 
to_sfixed(-1858.0/65536.0,1,-nbitq), 
to_sfixed(7789.0/65536.0,1,-nbitq), 
to_sfixed(663.0/65536.0,1,-nbitq), 
to_sfixed(-1892.0/65536.0,1,-nbitq), 
to_sfixed(-4894.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-986.0/65536.0,1,-nbitq), 
to_sfixed(-4841.0/65536.0,1,-nbitq), 
to_sfixed(3240.0/65536.0,1,-nbitq), 
to_sfixed(-6139.0/65536.0,1,-nbitq), 
to_sfixed(-3931.0/65536.0,1,-nbitq), 
to_sfixed(1914.0/65536.0,1,-nbitq), 
to_sfixed(-7325.0/65536.0,1,-nbitq), 
to_sfixed(296.0/65536.0,1,-nbitq), 
to_sfixed(4789.0/65536.0,1,-nbitq), 
to_sfixed(-1062.0/65536.0,1,-nbitq), 
to_sfixed(-2285.0/65536.0,1,-nbitq), 
to_sfixed(-4147.0/65536.0,1,-nbitq), 
to_sfixed(832.0/65536.0,1,-nbitq), 
to_sfixed(-3929.0/65536.0,1,-nbitq), 
to_sfixed(-274.0/65536.0,1,-nbitq), 
to_sfixed(2598.0/65536.0,1,-nbitq), 
to_sfixed(343.0/65536.0,1,-nbitq), 
to_sfixed(10070.0/65536.0,1,-nbitq), 
to_sfixed(1050.0/65536.0,1,-nbitq), 
to_sfixed(-2253.0/65536.0,1,-nbitq), 
to_sfixed(5056.0/65536.0,1,-nbitq), 
to_sfixed(10182.0/65536.0,1,-nbitq), 
to_sfixed(-1788.0/65536.0,1,-nbitq), 
to_sfixed(-12617.0/65536.0,1,-nbitq), 
to_sfixed(239.0/65536.0,1,-nbitq), 
to_sfixed(-15715.0/65536.0,1,-nbitq), 
to_sfixed(-974.0/65536.0,1,-nbitq), 
to_sfixed(4430.0/65536.0,1,-nbitq), 
to_sfixed(-2757.0/65536.0,1,-nbitq), 
to_sfixed(5284.0/65536.0,1,-nbitq), 
to_sfixed(-5850.0/65536.0,1,-nbitq), 
to_sfixed(-4215.0/65536.0,1,-nbitq), 
to_sfixed(4522.0/65536.0,1,-nbitq), 
to_sfixed(11300.0/65536.0,1,-nbitq), 
to_sfixed(2357.0/65536.0,1,-nbitq), 
to_sfixed(2232.0/65536.0,1,-nbitq), 
to_sfixed(-6222.0/65536.0,1,-nbitq), 
to_sfixed(1892.0/65536.0,1,-nbitq), 
to_sfixed(-3131.0/65536.0,1,-nbitq), 
to_sfixed(3967.0/65536.0,1,-nbitq), 
to_sfixed(1072.0/65536.0,1,-nbitq), 
to_sfixed(116.0/65536.0,1,-nbitq), 
to_sfixed(6224.0/65536.0,1,-nbitq), 
to_sfixed(-6008.0/65536.0,1,-nbitq), 
to_sfixed(-1336.0/65536.0,1,-nbitq), 
to_sfixed(-3564.0/65536.0,1,-nbitq), 
to_sfixed(-1986.0/65536.0,1,-nbitq), 
to_sfixed(-8981.0/65536.0,1,-nbitq), 
to_sfixed(-392.0/65536.0,1,-nbitq), 
to_sfixed(5209.0/65536.0,1,-nbitq), 
to_sfixed(-88.0/65536.0,1,-nbitq), 
to_sfixed(-3702.0/65536.0,1,-nbitq), 
to_sfixed(-5244.0/65536.0,1,-nbitq), 
to_sfixed(-12334.0/65536.0,1,-nbitq), 
to_sfixed(-2557.0/65536.0,1,-nbitq), 
to_sfixed(-7665.0/65536.0,1,-nbitq), 
to_sfixed(-2387.0/65536.0,1,-nbitq), 
to_sfixed(-2513.0/65536.0,1,-nbitq), 
to_sfixed(984.0/65536.0,1,-nbitq), 
to_sfixed(-463.0/65536.0,1,-nbitq), 
to_sfixed(12286.0/65536.0,1,-nbitq), 
to_sfixed(-2973.0/65536.0,1,-nbitq), 
to_sfixed(-877.0/65536.0,1,-nbitq), 
to_sfixed(-1080.0/65536.0,1,-nbitq), 
to_sfixed(-3186.0/65536.0,1,-nbitq), 
to_sfixed(-561.0/65536.0,1,-nbitq), 
to_sfixed(5975.0/65536.0,1,-nbitq), 
to_sfixed(-431.0/65536.0,1,-nbitq), 
to_sfixed(3202.0/65536.0,1,-nbitq), 
to_sfixed(-2363.0/65536.0,1,-nbitq), 
to_sfixed(-2248.0/65536.0,1,-nbitq), 
to_sfixed(-2710.0/65536.0,1,-nbitq), 
to_sfixed(-2045.0/65536.0,1,-nbitq), 
to_sfixed(705.0/65536.0,1,-nbitq), 
to_sfixed(1141.0/65536.0,1,-nbitq), 
to_sfixed(-621.0/65536.0,1,-nbitq), 
to_sfixed(7054.0/65536.0,1,-nbitq), 
to_sfixed(-3564.0/65536.0,1,-nbitq), 
to_sfixed(-1680.0/65536.0,1,-nbitq), 
to_sfixed(-5184.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4936.0/65536.0,1,-nbitq), 
to_sfixed(-4193.0/65536.0,1,-nbitq), 
to_sfixed(-2729.0/65536.0,1,-nbitq), 
to_sfixed(-5620.0/65536.0,1,-nbitq), 
to_sfixed(-1100.0/65536.0,1,-nbitq), 
to_sfixed(-9485.0/65536.0,1,-nbitq), 
to_sfixed(-9735.0/65536.0,1,-nbitq), 
to_sfixed(-5554.0/65536.0,1,-nbitq), 
to_sfixed(-3043.0/65536.0,1,-nbitq), 
to_sfixed(-2546.0/65536.0,1,-nbitq), 
to_sfixed(-1839.0/65536.0,1,-nbitq), 
to_sfixed(-15064.0/65536.0,1,-nbitq), 
to_sfixed(2158.0/65536.0,1,-nbitq), 
to_sfixed(-6503.0/65536.0,1,-nbitq), 
to_sfixed(715.0/65536.0,1,-nbitq), 
to_sfixed(-449.0/65536.0,1,-nbitq), 
to_sfixed(2970.0/65536.0,1,-nbitq), 
to_sfixed(5990.0/65536.0,1,-nbitq), 
to_sfixed(729.0/65536.0,1,-nbitq), 
to_sfixed(-1827.0/65536.0,1,-nbitq), 
to_sfixed(5646.0/65536.0,1,-nbitq), 
to_sfixed(5696.0/65536.0,1,-nbitq), 
to_sfixed(-2449.0/65536.0,1,-nbitq), 
to_sfixed(-9336.0/65536.0,1,-nbitq), 
to_sfixed(4237.0/65536.0,1,-nbitq), 
to_sfixed(-11982.0/65536.0,1,-nbitq), 
to_sfixed(-7951.0/65536.0,1,-nbitq), 
to_sfixed(2898.0/65536.0,1,-nbitq), 
to_sfixed(-1844.0/65536.0,1,-nbitq), 
to_sfixed(1358.0/65536.0,1,-nbitq), 
to_sfixed(-2641.0/65536.0,1,-nbitq), 
to_sfixed(-3304.0/65536.0,1,-nbitq), 
to_sfixed(2824.0/65536.0,1,-nbitq), 
to_sfixed(3168.0/65536.0,1,-nbitq), 
to_sfixed(-36.0/65536.0,1,-nbitq), 
to_sfixed(2913.0/65536.0,1,-nbitq), 
to_sfixed(-6123.0/65536.0,1,-nbitq), 
to_sfixed(2125.0/65536.0,1,-nbitq), 
to_sfixed(1160.0/65536.0,1,-nbitq), 
to_sfixed(279.0/65536.0,1,-nbitq), 
to_sfixed(4583.0/65536.0,1,-nbitq), 
to_sfixed(419.0/65536.0,1,-nbitq), 
to_sfixed(-3139.0/65536.0,1,-nbitq), 
to_sfixed(-1356.0/65536.0,1,-nbitq), 
to_sfixed(-1265.0/65536.0,1,-nbitq), 
to_sfixed(-6075.0/65536.0,1,-nbitq), 
to_sfixed(-2054.0/65536.0,1,-nbitq), 
to_sfixed(-4136.0/65536.0,1,-nbitq), 
to_sfixed(-264.0/65536.0,1,-nbitq), 
to_sfixed(3284.0/65536.0,1,-nbitq), 
to_sfixed(710.0/65536.0,1,-nbitq), 
to_sfixed(1485.0/65536.0,1,-nbitq), 
to_sfixed(-3867.0/65536.0,1,-nbitq), 
to_sfixed(-15729.0/65536.0,1,-nbitq), 
to_sfixed(-6435.0/65536.0,1,-nbitq), 
to_sfixed(-4811.0/65536.0,1,-nbitq), 
to_sfixed(-2771.0/65536.0,1,-nbitq), 
to_sfixed(2693.0/65536.0,1,-nbitq), 
to_sfixed(-1530.0/65536.0,1,-nbitq), 
to_sfixed(2566.0/65536.0,1,-nbitq), 
to_sfixed(10226.0/65536.0,1,-nbitq), 
to_sfixed(-2364.0/65536.0,1,-nbitq), 
to_sfixed(-1662.0/65536.0,1,-nbitq), 
to_sfixed(1435.0/65536.0,1,-nbitq), 
to_sfixed(7662.0/65536.0,1,-nbitq), 
to_sfixed(1368.0/65536.0,1,-nbitq), 
to_sfixed(1428.0/65536.0,1,-nbitq), 
to_sfixed(-2224.0/65536.0,1,-nbitq), 
to_sfixed(561.0/65536.0,1,-nbitq), 
to_sfixed(-7765.0/65536.0,1,-nbitq), 
to_sfixed(-840.0/65536.0,1,-nbitq), 
to_sfixed(-3519.0/65536.0,1,-nbitq), 
to_sfixed(-3388.0/65536.0,1,-nbitq), 
to_sfixed(-1711.0/65536.0,1,-nbitq), 
to_sfixed(-403.0/65536.0,1,-nbitq), 
to_sfixed(-560.0/65536.0,1,-nbitq), 
to_sfixed(7305.0/65536.0,1,-nbitq), 
to_sfixed(2831.0/65536.0,1,-nbitq), 
to_sfixed(1957.0/65536.0,1,-nbitq), 
to_sfixed(-4482.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2973.0/65536.0,1,-nbitq), 
to_sfixed(-1194.0/65536.0,1,-nbitq), 
to_sfixed(-15691.0/65536.0,1,-nbitq), 
to_sfixed(-4241.0/65536.0,1,-nbitq), 
to_sfixed(-807.0/65536.0,1,-nbitq), 
to_sfixed(-3679.0/65536.0,1,-nbitq), 
to_sfixed(-6948.0/65536.0,1,-nbitq), 
to_sfixed(-2677.0/65536.0,1,-nbitq), 
to_sfixed(-2057.0/65536.0,1,-nbitq), 
to_sfixed(652.0/65536.0,1,-nbitq), 
to_sfixed(-2868.0/65536.0,1,-nbitq), 
to_sfixed(-5823.0/65536.0,1,-nbitq), 
to_sfixed(-255.0/65536.0,1,-nbitq), 
to_sfixed(-6554.0/65536.0,1,-nbitq), 
to_sfixed(1533.0/65536.0,1,-nbitq), 
to_sfixed(-2466.0/65536.0,1,-nbitq), 
to_sfixed(1156.0/65536.0,1,-nbitq), 
to_sfixed(-2346.0/65536.0,1,-nbitq), 
to_sfixed(1924.0/65536.0,1,-nbitq), 
to_sfixed(789.0/65536.0,1,-nbitq), 
to_sfixed(-608.0/65536.0,1,-nbitq), 
to_sfixed(4964.0/65536.0,1,-nbitq), 
to_sfixed(-4713.0/65536.0,1,-nbitq), 
to_sfixed(-6799.0/65536.0,1,-nbitq), 
to_sfixed(5295.0/65536.0,1,-nbitq), 
to_sfixed(-11396.0/65536.0,1,-nbitq), 
to_sfixed(-2099.0/65536.0,1,-nbitq), 
to_sfixed(5956.0/65536.0,1,-nbitq), 
to_sfixed(-4815.0/65536.0,1,-nbitq), 
to_sfixed(5265.0/65536.0,1,-nbitq), 
to_sfixed(-2711.0/65536.0,1,-nbitq), 
to_sfixed(1140.0/65536.0,1,-nbitq), 
to_sfixed(3588.0/65536.0,1,-nbitq), 
to_sfixed(-3469.0/65536.0,1,-nbitq), 
to_sfixed(1132.0/65536.0,1,-nbitq), 
to_sfixed(1281.0/65536.0,1,-nbitq), 
to_sfixed(-11011.0/65536.0,1,-nbitq), 
to_sfixed(1815.0/65536.0,1,-nbitq), 
to_sfixed(4612.0/65536.0,1,-nbitq), 
to_sfixed(2544.0/65536.0,1,-nbitq), 
to_sfixed(4045.0/65536.0,1,-nbitq), 
to_sfixed(2188.0/65536.0,1,-nbitq), 
to_sfixed(-8835.0/65536.0,1,-nbitq), 
to_sfixed(-4169.0/65536.0,1,-nbitq), 
to_sfixed(-237.0/65536.0,1,-nbitq), 
to_sfixed(4170.0/65536.0,1,-nbitq), 
to_sfixed(-1266.0/65536.0,1,-nbitq), 
to_sfixed(1111.0/65536.0,1,-nbitq), 
to_sfixed(-518.0/65536.0,1,-nbitq), 
to_sfixed(3975.0/65536.0,1,-nbitq), 
to_sfixed(-966.0/65536.0,1,-nbitq), 
to_sfixed(379.0/65536.0,1,-nbitq), 
to_sfixed(-7213.0/65536.0,1,-nbitq), 
to_sfixed(-11350.0/65536.0,1,-nbitq), 
to_sfixed(-994.0/65536.0,1,-nbitq), 
to_sfixed(-8160.0/65536.0,1,-nbitq), 
to_sfixed(1571.0/65536.0,1,-nbitq), 
to_sfixed(344.0/65536.0,1,-nbitq), 
to_sfixed(2138.0/65536.0,1,-nbitq), 
to_sfixed(5241.0/65536.0,1,-nbitq), 
to_sfixed(1722.0/65536.0,1,-nbitq), 
to_sfixed(1059.0/65536.0,1,-nbitq), 
to_sfixed(2904.0/65536.0,1,-nbitq), 
to_sfixed(1999.0/65536.0,1,-nbitq), 
to_sfixed(-70.0/65536.0,1,-nbitq), 
to_sfixed(10710.0/65536.0,1,-nbitq), 
to_sfixed(2548.0/65536.0,1,-nbitq), 
to_sfixed(3015.0/65536.0,1,-nbitq), 
to_sfixed(-1179.0/65536.0,1,-nbitq), 
to_sfixed(-1848.0/65536.0,1,-nbitq), 
to_sfixed(-4838.0/65536.0,1,-nbitq), 
to_sfixed(-5486.0/65536.0,1,-nbitq), 
to_sfixed(-4227.0/65536.0,1,-nbitq), 
to_sfixed(1288.0/65536.0,1,-nbitq), 
to_sfixed(-1443.0/65536.0,1,-nbitq), 
to_sfixed(4326.0/65536.0,1,-nbitq), 
to_sfixed(4981.0/65536.0,1,-nbitq), 
to_sfixed(5815.0/65536.0,1,-nbitq), 
to_sfixed(2587.0/65536.0,1,-nbitq), 
to_sfixed(-10913.0/65536.0,1,-nbitq)  ), 
( to_sfixed(522.0/65536.0,1,-nbitq), 
to_sfixed(6247.0/65536.0,1,-nbitq), 
to_sfixed(-19539.0/65536.0,1,-nbitq), 
to_sfixed(-6036.0/65536.0,1,-nbitq), 
to_sfixed(-1214.0/65536.0,1,-nbitq), 
to_sfixed(-2345.0/65536.0,1,-nbitq), 
to_sfixed(-1725.0/65536.0,1,-nbitq), 
to_sfixed(-11400.0/65536.0,1,-nbitq), 
to_sfixed(-5513.0/65536.0,1,-nbitq), 
to_sfixed(-260.0/65536.0,1,-nbitq), 
to_sfixed(778.0/65536.0,1,-nbitq), 
to_sfixed(-4927.0/65536.0,1,-nbitq), 
to_sfixed(1610.0/65536.0,1,-nbitq), 
to_sfixed(1569.0/65536.0,1,-nbitq), 
to_sfixed(-1827.0/65536.0,1,-nbitq), 
to_sfixed(-2688.0/65536.0,1,-nbitq), 
to_sfixed(1933.0/65536.0,1,-nbitq), 
to_sfixed(-11407.0/65536.0,1,-nbitq), 
to_sfixed(2868.0/65536.0,1,-nbitq), 
to_sfixed(976.0/65536.0,1,-nbitq), 
to_sfixed(-2373.0/65536.0,1,-nbitq), 
to_sfixed(4632.0/65536.0,1,-nbitq), 
to_sfixed(-3261.0/65536.0,1,-nbitq), 
to_sfixed(-2495.0/65536.0,1,-nbitq), 
to_sfixed(6251.0/65536.0,1,-nbitq), 
to_sfixed(-4255.0/65536.0,1,-nbitq), 
to_sfixed(5106.0/65536.0,1,-nbitq), 
to_sfixed(-80.0/65536.0,1,-nbitq), 
to_sfixed(-2441.0/65536.0,1,-nbitq), 
to_sfixed(3479.0/65536.0,1,-nbitq), 
to_sfixed(-2025.0/65536.0,1,-nbitq), 
to_sfixed(2223.0/65536.0,1,-nbitq), 
to_sfixed(76.0/65536.0,1,-nbitq), 
to_sfixed(-3610.0/65536.0,1,-nbitq), 
to_sfixed(1250.0/65536.0,1,-nbitq), 
to_sfixed(-1160.0/65536.0,1,-nbitq), 
to_sfixed(-6123.0/65536.0,1,-nbitq), 
to_sfixed(5207.0/65536.0,1,-nbitq), 
to_sfixed(3829.0/65536.0,1,-nbitq), 
to_sfixed(3780.0/65536.0,1,-nbitq), 
to_sfixed(255.0/65536.0,1,-nbitq), 
to_sfixed(-1997.0/65536.0,1,-nbitq), 
to_sfixed(-6941.0/65536.0,1,-nbitq), 
to_sfixed(2242.0/65536.0,1,-nbitq), 
to_sfixed(-472.0/65536.0,1,-nbitq), 
to_sfixed(4149.0/65536.0,1,-nbitq), 
to_sfixed(-2818.0/65536.0,1,-nbitq), 
to_sfixed(3893.0/65536.0,1,-nbitq), 
to_sfixed(1319.0/65536.0,1,-nbitq), 
to_sfixed(-2158.0/65536.0,1,-nbitq), 
to_sfixed(-1898.0/65536.0,1,-nbitq), 
to_sfixed(-338.0/65536.0,1,-nbitq), 
to_sfixed(-1925.0/65536.0,1,-nbitq), 
to_sfixed(455.0/65536.0,1,-nbitq), 
to_sfixed(395.0/65536.0,1,-nbitq), 
to_sfixed(-9964.0/65536.0,1,-nbitq), 
to_sfixed(742.0/65536.0,1,-nbitq), 
to_sfixed(4544.0/65536.0,1,-nbitq), 
to_sfixed(3331.0/65536.0,1,-nbitq), 
to_sfixed(11519.0/65536.0,1,-nbitq), 
to_sfixed(-1956.0/65536.0,1,-nbitq), 
to_sfixed(-967.0/65536.0,1,-nbitq), 
to_sfixed(-1521.0/65536.0,1,-nbitq), 
to_sfixed(186.0/65536.0,1,-nbitq), 
to_sfixed(-3420.0/65536.0,1,-nbitq), 
to_sfixed(17355.0/65536.0,1,-nbitq), 
to_sfixed(1716.0/65536.0,1,-nbitq), 
to_sfixed(2066.0/65536.0,1,-nbitq), 
to_sfixed(-4509.0/65536.0,1,-nbitq), 
to_sfixed(-4356.0/65536.0,1,-nbitq), 
to_sfixed(-3357.0/65536.0,1,-nbitq), 
to_sfixed(-6698.0/65536.0,1,-nbitq), 
to_sfixed(-7753.0/65536.0,1,-nbitq), 
to_sfixed(912.0/65536.0,1,-nbitq), 
to_sfixed(-1160.0/65536.0,1,-nbitq), 
to_sfixed(754.0/65536.0,1,-nbitq), 
to_sfixed(2653.0/65536.0,1,-nbitq), 
to_sfixed(2010.0/65536.0,1,-nbitq), 
to_sfixed(1276.0/65536.0,1,-nbitq), 
to_sfixed(-7891.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2124.0/65536.0,1,-nbitq), 
to_sfixed(5140.0/65536.0,1,-nbitq), 
to_sfixed(-7311.0/65536.0,1,-nbitq), 
to_sfixed(-9510.0/65536.0,1,-nbitq), 
to_sfixed(-2391.0/65536.0,1,-nbitq), 
to_sfixed(-3243.0/65536.0,1,-nbitq), 
to_sfixed(1950.0/65536.0,1,-nbitq), 
to_sfixed(-8884.0/65536.0,1,-nbitq), 
to_sfixed(-4330.0/65536.0,1,-nbitq), 
to_sfixed(3604.0/65536.0,1,-nbitq), 
to_sfixed(-3695.0/65536.0,1,-nbitq), 
to_sfixed(-9752.0/65536.0,1,-nbitq), 
to_sfixed(357.0/65536.0,1,-nbitq), 
to_sfixed(765.0/65536.0,1,-nbitq), 
to_sfixed(-3073.0/65536.0,1,-nbitq), 
to_sfixed(-977.0/65536.0,1,-nbitq), 
to_sfixed(190.0/65536.0,1,-nbitq), 
to_sfixed(-12859.0/65536.0,1,-nbitq), 
to_sfixed(-1477.0/65536.0,1,-nbitq), 
to_sfixed(1538.0/65536.0,1,-nbitq), 
to_sfixed(-2958.0/65536.0,1,-nbitq), 
to_sfixed(2921.0/65536.0,1,-nbitq), 
to_sfixed(5520.0/65536.0,1,-nbitq), 
to_sfixed(-6145.0/65536.0,1,-nbitq), 
to_sfixed(6765.0/65536.0,1,-nbitq), 
to_sfixed(-2592.0/65536.0,1,-nbitq), 
to_sfixed(-10430.0/65536.0,1,-nbitq), 
to_sfixed(2515.0/65536.0,1,-nbitq), 
to_sfixed(-18506.0/65536.0,1,-nbitq), 
to_sfixed(3724.0/65536.0,1,-nbitq), 
to_sfixed(3362.0/65536.0,1,-nbitq), 
to_sfixed(5809.0/65536.0,1,-nbitq), 
to_sfixed(-8490.0/65536.0,1,-nbitq), 
to_sfixed(92.0/65536.0,1,-nbitq), 
to_sfixed(-3813.0/65536.0,1,-nbitq), 
to_sfixed(-750.0/65536.0,1,-nbitq), 
to_sfixed(-2955.0/65536.0,1,-nbitq), 
to_sfixed(8376.0/65536.0,1,-nbitq), 
to_sfixed(12527.0/65536.0,1,-nbitq), 
to_sfixed(-1293.0/65536.0,1,-nbitq), 
to_sfixed(2437.0/65536.0,1,-nbitq), 
to_sfixed(-1807.0/65536.0,1,-nbitq), 
to_sfixed(-10276.0/65536.0,1,-nbitq), 
to_sfixed(5712.0/65536.0,1,-nbitq), 
to_sfixed(2031.0/65536.0,1,-nbitq), 
to_sfixed(-7158.0/65536.0,1,-nbitq), 
to_sfixed(-2879.0/65536.0,1,-nbitq), 
to_sfixed(1354.0/65536.0,1,-nbitq), 
to_sfixed(2642.0/65536.0,1,-nbitq), 
to_sfixed(1237.0/65536.0,1,-nbitq), 
to_sfixed(3164.0/65536.0,1,-nbitq), 
to_sfixed(5439.0/65536.0,1,-nbitq), 
to_sfixed(1496.0/65536.0,1,-nbitq), 
to_sfixed(4418.0/65536.0,1,-nbitq), 
to_sfixed(2046.0/65536.0,1,-nbitq), 
to_sfixed(-7989.0/65536.0,1,-nbitq), 
to_sfixed(-1964.0/65536.0,1,-nbitq), 
to_sfixed(2049.0/65536.0,1,-nbitq), 
to_sfixed(-2421.0/65536.0,1,-nbitq), 
to_sfixed(4918.0/65536.0,1,-nbitq), 
to_sfixed(-13288.0/65536.0,1,-nbitq), 
to_sfixed(-1259.0/65536.0,1,-nbitq), 
to_sfixed(-132.0/65536.0,1,-nbitq), 
to_sfixed(-2587.0/65536.0,1,-nbitq), 
to_sfixed(4342.0/65536.0,1,-nbitq), 
to_sfixed(7775.0/65536.0,1,-nbitq), 
to_sfixed(-3441.0/65536.0,1,-nbitq), 
to_sfixed(4021.0/65536.0,1,-nbitq), 
to_sfixed(-2828.0/65536.0,1,-nbitq), 
to_sfixed(-9717.0/65536.0,1,-nbitq), 
to_sfixed(-162.0/65536.0,1,-nbitq), 
to_sfixed(1985.0/65536.0,1,-nbitq), 
to_sfixed(-7121.0/65536.0,1,-nbitq), 
to_sfixed(-2845.0/65536.0,1,-nbitq), 
to_sfixed(2301.0/65536.0,1,-nbitq), 
to_sfixed(-7679.0/65536.0,1,-nbitq), 
to_sfixed(7748.0/65536.0,1,-nbitq), 
to_sfixed(-3408.0/65536.0,1,-nbitq), 
to_sfixed(2387.0/65536.0,1,-nbitq), 
to_sfixed(141.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2277.0/65536.0,1,-nbitq), 
to_sfixed(828.0/65536.0,1,-nbitq), 
to_sfixed(-8679.0/65536.0,1,-nbitq), 
to_sfixed(-1339.0/65536.0,1,-nbitq), 
to_sfixed(10489.0/65536.0,1,-nbitq), 
to_sfixed(-2814.0/65536.0,1,-nbitq), 
to_sfixed(1471.0/65536.0,1,-nbitq), 
to_sfixed(-6587.0/65536.0,1,-nbitq), 
to_sfixed(-4263.0/65536.0,1,-nbitq), 
to_sfixed(3829.0/65536.0,1,-nbitq), 
to_sfixed(-2234.0/65536.0,1,-nbitq), 
to_sfixed(-764.0/65536.0,1,-nbitq), 
to_sfixed(259.0/65536.0,1,-nbitq), 
to_sfixed(-3470.0/65536.0,1,-nbitq), 
to_sfixed(-1629.0/65536.0,1,-nbitq), 
to_sfixed(2281.0/65536.0,1,-nbitq), 
to_sfixed(2273.0/65536.0,1,-nbitq), 
to_sfixed(-10256.0/65536.0,1,-nbitq), 
to_sfixed(2193.0/65536.0,1,-nbitq), 
to_sfixed(2278.0/65536.0,1,-nbitq), 
to_sfixed(-1495.0/65536.0,1,-nbitq), 
to_sfixed(5683.0/65536.0,1,-nbitq), 
to_sfixed(-1451.0/65536.0,1,-nbitq), 
to_sfixed(-901.0/65536.0,1,-nbitq), 
to_sfixed(6579.0/65536.0,1,-nbitq), 
to_sfixed(-7629.0/65536.0,1,-nbitq), 
to_sfixed(-3518.0/65536.0,1,-nbitq), 
to_sfixed(-2988.0/65536.0,1,-nbitq), 
to_sfixed(-7537.0/65536.0,1,-nbitq), 
to_sfixed(3293.0/65536.0,1,-nbitq), 
to_sfixed(4290.0/65536.0,1,-nbitq), 
to_sfixed(5027.0/65536.0,1,-nbitq), 
to_sfixed(-11961.0/65536.0,1,-nbitq), 
to_sfixed(497.0/65536.0,1,-nbitq), 
to_sfixed(318.0/65536.0,1,-nbitq), 
to_sfixed(-3168.0/65536.0,1,-nbitq), 
to_sfixed(-9080.0/65536.0,1,-nbitq), 
to_sfixed(7273.0/65536.0,1,-nbitq), 
to_sfixed(13213.0/65536.0,1,-nbitq), 
to_sfixed(-1384.0/65536.0,1,-nbitq), 
to_sfixed(3086.0/65536.0,1,-nbitq), 
to_sfixed(-2813.0/65536.0,1,-nbitq), 
to_sfixed(-5186.0/65536.0,1,-nbitq), 
to_sfixed(3002.0/65536.0,1,-nbitq), 
to_sfixed(1895.0/65536.0,1,-nbitq), 
to_sfixed(-474.0/65536.0,1,-nbitq), 
to_sfixed(-2097.0/65536.0,1,-nbitq), 
to_sfixed(5084.0/65536.0,1,-nbitq), 
to_sfixed(-1394.0/65536.0,1,-nbitq), 
to_sfixed(3180.0/65536.0,1,-nbitq), 
to_sfixed(-2541.0/65536.0,1,-nbitq), 
to_sfixed(3919.0/65536.0,1,-nbitq), 
to_sfixed(1999.0/65536.0,1,-nbitq), 
to_sfixed(5430.0/65536.0,1,-nbitq), 
to_sfixed(3267.0/65536.0,1,-nbitq), 
to_sfixed(-6431.0/65536.0,1,-nbitq), 
to_sfixed(2835.0/65536.0,1,-nbitq), 
to_sfixed(-2373.0/65536.0,1,-nbitq), 
to_sfixed(1513.0/65536.0,1,-nbitq), 
to_sfixed(4408.0/65536.0,1,-nbitq), 
to_sfixed(-6480.0/65536.0,1,-nbitq), 
to_sfixed(-1394.0/65536.0,1,-nbitq), 
to_sfixed(-2305.0/65536.0,1,-nbitq), 
to_sfixed(1043.0/65536.0,1,-nbitq), 
to_sfixed(535.0/65536.0,1,-nbitq), 
to_sfixed(-5711.0/65536.0,1,-nbitq), 
to_sfixed(-8608.0/65536.0,1,-nbitq), 
to_sfixed(3973.0/65536.0,1,-nbitq), 
to_sfixed(-3928.0/65536.0,1,-nbitq), 
to_sfixed(3329.0/65536.0,1,-nbitq), 
to_sfixed(-1696.0/65536.0,1,-nbitq), 
to_sfixed(11084.0/65536.0,1,-nbitq), 
to_sfixed(-4903.0/65536.0,1,-nbitq), 
to_sfixed(-658.0/65536.0,1,-nbitq), 
to_sfixed(391.0/65536.0,1,-nbitq), 
to_sfixed(-5640.0/65536.0,1,-nbitq), 
to_sfixed(9817.0/65536.0,1,-nbitq), 
to_sfixed(1170.0/65536.0,1,-nbitq), 
to_sfixed(1395.0/65536.0,1,-nbitq), 
to_sfixed(5645.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3290.0/65536.0,1,-nbitq), 
to_sfixed(-1169.0/65536.0,1,-nbitq), 
to_sfixed(10591.0/65536.0,1,-nbitq), 
to_sfixed(-3627.0/65536.0,1,-nbitq), 
to_sfixed(5986.0/65536.0,1,-nbitq), 
to_sfixed(-6417.0/65536.0,1,-nbitq), 
to_sfixed(3407.0/65536.0,1,-nbitq), 
to_sfixed(-9349.0/65536.0,1,-nbitq), 
to_sfixed(-1380.0/65536.0,1,-nbitq), 
to_sfixed(-910.0/65536.0,1,-nbitq), 
to_sfixed(-488.0/65536.0,1,-nbitq), 
to_sfixed(8240.0/65536.0,1,-nbitq), 
to_sfixed(876.0/65536.0,1,-nbitq), 
to_sfixed(-6402.0/65536.0,1,-nbitq), 
to_sfixed(-1966.0/65536.0,1,-nbitq), 
to_sfixed(1725.0/65536.0,1,-nbitq), 
to_sfixed(-208.0/65536.0,1,-nbitq), 
to_sfixed(-1815.0/65536.0,1,-nbitq), 
to_sfixed(-1457.0/65536.0,1,-nbitq), 
to_sfixed(2427.0/65536.0,1,-nbitq), 
to_sfixed(-769.0/65536.0,1,-nbitq), 
to_sfixed(11749.0/65536.0,1,-nbitq), 
to_sfixed(12163.0/65536.0,1,-nbitq), 
to_sfixed(-2653.0/65536.0,1,-nbitq), 
to_sfixed(7042.0/65536.0,1,-nbitq), 
to_sfixed(-8932.0/65536.0,1,-nbitq), 
to_sfixed(-239.0/65536.0,1,-nbitq), 
to_sfixed(1208.0/65536.0,1,-nbitq), 
to_sfixed(-6191.0/65536.0,1,-nbitq), 
to_sfixed(47.0/65536.0,1,-nbitq), 
to_sfixed(10867.0/65536.0,1,-nbitq), 
to_sfixed(9777.0/65536.0,1,-nbitq), 
to_sfixed(-3991.0/65536.0,1,-nbitq), 
to_sfixed(6005.0/65536.0,1,-nbitq), 
to_sfixed(-4364.0/65536.0,1,-nbitq), 
to_sfixed(-297.0/65536.0,1,-nbitq), 
to_sfixed(3558.0/65536.0,1,-nbitq), 
to_sfixed(6576.0/65536.0,1,-nbitq), 
to_sfixed(3791.0/65536.0,1,-nbitq), 
to_sfixed(-113.0/65536.0,1,-nbitq), 
to_sfixed(-2011.0/65536.0,1,-nbitq), 
to_sfixed(2608.0/65536.0,1,-nbitq), 
to_sfixed(4720.0/65536.0,1,-nbitq), 
to_sfixed(-6915.0/65536.0,1,-nbitq), 
to_sfixed(825.0/65536.0,1,-nbitq), 
to_sfixed(1284.0/65536.0,1,-nbitq), 
to_sfixed(-1051.0/65536.0,1,-nbitq), 
to_sfixed(4068.0/65536.0,1,-nbitq), 
to_sfixed(-365.0/65536.0,1,-nbitq), 
to_sfixed(-923.0/65536.0,1,-nbitq), 
to_sfixed(1043.0/65536.0,1,-nbitq), 
to_sfixed(-3176.0/65536.0,1,-nbitq), 
to_sfixed(-789.0/65536.0,1,-nbitq), 
to_sfixed(10632.0/65536.0,1,-nbitq), 
to_sfixed(6201.0/65536.0,1,-nbitq), 
to_sfixed(3919.0/65536.0,1,-nbitq), 
to_sfixed(428.0/65536.0,1,-nbitq), 
to_sfixed(-7946.0/65536.0,1,-nbitq), 
to_sfixed(-1829.0/65536.0,1,-nbitq), 
to_sfixed(-1599.0/65536.0,1,-nbitq), 
to_sfixed(-4358.0/65536.0,1,-nbitq), 
to_sfixed(-1668.0/65536.0,1,-nbitq), 
to_sfixed(2421.0/65536.0,1,-nbitq), 
to_sfixed(-2512.0/65536.0,1,-nbitq), 
to_sfixed(475.0/65536.0,1,-nbitq), 
to_sfixed(-9873.0/65536.0,1,-nbitq), 
to_sfixed(-4212.0/65536.0,1,-nbitq), 
to_sfixed(-3691.0/65536.0,1,-nbitq), 
to_sfixed(-5051.0/65536.0,1,-nbitq), 
to_sfixed(2360.0/65536.0,1,-nbitq), 
to_sfixed(2563.0/65536.0,1,-nbitq), 
to_sfixed(5603.0/65536.0,1,-nbitq), 
to_sfixed(-4591.0/65536.0,1,-nbitq), 
to_sfixed(-1937.0/65536.0,1,-nbitq), 
to_sfixed(476.0/65536.0,1,-nbitq), 
to_sfixed(2595.0/65536.0,1,-nbitq), 
to_sfixed(9210.0/65536.0,1,-nbitq), 
to_sfixed(1204.0/65536.0,1,-nbitq), 
to_sfixed(1996.0/65536.0,1,-nbitq), 
to_sfixed(4753.0/65536.0,1,-nbitq)  ), 
( to_sfixed(353.0/65536.0,1,-nbitq), 
to_sfixed(-1303.0/65536.0,1,-nbitq), 
to_sfixed(8730.0/65536.0,1,-nbitq), 
to_sfixed(1882.0/65536.0,1,-nbitq), 
to_sfixed(9458.0/65536.0,1,-nbitq), 
to_sfixed(-4896.0/65536.0,1,-nbitq), 
to_sfixed(7782.0/65536.0,1,-nbitq), 
to_sfixed(-5157.0/65536.0,1,-nbitq), 
to_sfixed(-1873.0/65536.0,1,-nbitq), 
to_sfixed(2907.0/65536.0,1,-nbitq), 
to_sfixed(-2356.0/65536.0,1,-nbitq), 
to_sfixed(4377.0/65536.0,1,-nbitq), 
to_sfixed(708.0/65536.0,1,-nbitq), 
to_sfixed(-2950.0/65536.0,1,-nbitq), 
to_sfixed(1962.0/65536.0,1,-nbitq), 
to_sfixed(-2264.0/65536.0,1,-nbitq), 
to_sfixed(1112.0/65536.0,1,-nbitq), 
to_sfixed(3589.0/65536.0,1,-nbitq), 
to_sfixed(-826.0/65536.0,1,-nbitq), 
to_sfixed(1862.0/65536.0,1,-nbitq), 
to_sfixed(-2258.0/65536.0,1,-nbitq), 
to_sfixed(8431.0/65536.0,1,-nbitq), 
to_sfixed(2285.0/65536.0,1,-nbitq), 
to_sfixed(2746.0/65536.0,1,-nbitq), 
to_sfixed(12706.0/65536.0,1,-nbitq), 
to_sfixed(-1458.0/65536.0,1,-nbitq), 
to_sfixed(-2254.0/65536.0,1,-nbitq), 
to_sfixed(5.0/65536.0,1,-nbitq), 
to_sfixed(685.0/65536.0,1,-nbitq), 
to_sfixed(-1893.0/65536.0,1,-nbitq), 
to_sfixed(2404.0/65536.0,1,-nbitq), 
to_sfixed(12253.0/65536.0,1,-nbitq), 
to_sfixed(-4615.0/65536.0,1,-nbitq), 
to_sfixed(4003.0/65536.0,1,-nbitq), 
to_sfixed(-3996.0/65536.0,1,-nbitq), 
to_sfixed(-256.0/65536.0,1,-nbitq), 
to_sfixed(3400.0/65536.0,1,-nbitq), 
to_sfixed(1647.0/65536.0,1,-nbitq), 
to_sfixed(-2751.0/65536.0,1,-nbitq), 
to_sfixed(-1765.0/65536.0,1,-nbitq), 
to_sfixed(4948.0/65536.0,1,-nbitq), 
to_sfixed(-940.0/65536.0,1,-nbitq), 
to_sfixed(-252.0/65536.0,1,-nbitq), 
to_sfixed(-11874.0/65536.0,1,-nbitq), 
to_sfixed(2115.0/65536.0,1,-nbitq), 
to_sfixed(-290.0/65536.0,1,-nbitq), 
to_sfixed(-155.0/65536.0,1,-nbitq), 
to_sfixed(-4261.0/65536.0,1,-nbitq), 
to_sfixed(117.0/65536.0,1,-nbitq), 
to_sfixed(3407.0/65536.0,1,-nbitq), 
to_sfixed(606.0/65536.0,1,-nbitq), 
to_sfixed(1584.0/65536.0,1,-nbitq), 
to_sfixed(-2091.0/65536.0,1,-nbitq), 
to_sfixed(-178.0/65536.0,1,-nbitq), 
to_sfixed(6060.0/65536.0,1,-nbitq), 
to_sfixed(5206.0/65536.0,1,-nbitq), 
to_sfixed(-573.0/65536.0,1,-nbitq), 
to_sfixed(-8255.0/65536.0,1,-nbitq), 
to_sfixed(-2562.0/65536.0,1,-nbitq), 
to_sfixed(2026.0/65536.0,1,-nbitq), 
to_sfixed(-1108.0/65536.0,1,-nbitq), 
to_sfixed(-2488.0/65536.0,1,-nbitq), 
to_sfixed(-1176.0/65536.0,1,-nbitq), 
to_sfixed(1517.0/65536.0,1,-nbitq), 
to_sfixed(1412.0/65536.0,1,-nbitq), 
to_sfixed(-4299.0/65536.0,1,-nbitq), 
to_sfixed(1414.0/65536.0,1,-nbitq), 
to_sfixed(-8766.0/65536.0,1,-nbitq), 
to_sfixed(-6570.0/65536.0,1,-nbitq), 
to_sfixed(-6348.0/65536.0,1,-nbitq), 
to_sfixed(610.0/65536.0,1,-nbitq), 
to_sfixed(1853.0/65536.0,1,-nbitq), 
to_sfixed(4724.0/65536.0,1,-nbitq), 
to_sfixed(901.0/65536.0,1,-nbitq), 
to_sfixed(-1682.0/65536.0,1,-nbitq), 
to_sfixed(9578.0/65536.0,1,-nbitq), 
to_sfixed(8671.0/65536.0,1,-nbitq), 
to_sfixed(396.0/65536.0,1,-nbitq), 
to_sfixed(1878.0/65536.0,1,-nbitq), 
to_sfixed(1342.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1164.0/65536.0,1,-nbitq), 
to_sfixed(-4468.0/65536.0,1,-nbitq), 
to_sfixed(6273.0/65536.0,1,-nbitq), 
to_sfixed(-1852.0/65536.0,1,-nbitq), 
to_sfixed(1671.0/65536.0,1,-nbitq), 
to_sfixed(-10858.0/65536.0,1,-nbitq), 
to_sfixed(5565.0/65536.0,1,-nbitq), 
to_sfixed(-1262.0/65536.0,1,-nbitq), 
to_sfixed(-583.0/65536.0,1,-nbitq), 
to_sfixed(-308.0/65536.0,1,-nbitq), 
to_sfixed(-5285.0/65536.0,1,-nbitq), 
to_sfixed(732.0/65536.0,1,-nbitq), 
to_sfixed(2415.0/65536.0,1,-nbitq), 
to_sfixed(-519.0/65536.0,1,-nbitq), 
to_sfixed(-2358.0/65536.0,1,-nbitq), 
to_sfixed(1917.0/65536.0,1,-nbitq), 
to_sfixed(1840.0/65536.0,1,-nbitq), 
to_sfixed(8379.0/65536.0,1,-nbitq), 
to_sfixed(-2433.0/65536.0,1,-nbitq), 
to_sfixed(-441.0/65536.0,1,-nbitq), 
to_sfixed(-1976.0/65536.0,1,-nbitq), 
to_sfixed(-1327.0/65536.0,1,-nbitq), 
to_sfixed(5498.0/65536.0,1,-nbitq), 
to_sfixed(6131.0/65536.0,1,-nbitq), 
to_sfixed(10265.0/65536.0,1,-nbitq), 
to_sfixed(3595.0/65536.0,1,-nbitq), 
to_sfixed(5838.0/65536.0,1,-nbitq), 
to_sfixed(1295.0/65536.0,1,-nbitq), 
to_sfixed(-8765.0/65536.0,1,-nbitq), 
to_sfixed(2911.0/65536.0,1,-nbitq), 
to_sfixed(-10422.0/65536.0,1,-nbitq), 
to_sfixed(7602.0/65536.0,1,-nbitq), 
to_sfixed(-551.0/65536.0,1,-nbitq), 
to_sfixed(-5675.0/65536.0,1,-nbitq), 
to_sfixed(-784.0/65536.0,1,-nbitq), 
to_sfixed(2052.0/65536.0,1,-nbitq), 
to_sfixed(-1822.0/65536.0,1,-nbitq), 
to_sfixed(-1963.0/65536.0,1,-nbitq), 
to_sfixed(-1590.0/65536.0,1,-nbitq), 
to_sfixed(1085.0/65536.0,1,-nbitq), 
to_sfixed(7546.0/65536.0,1,-nbitq), 
to_sfixed(2180.0/65536.0,1,-nbitq), 
to_sfixed(-3495.0/65536.0,1,-nbitq), 
to_sfixed(-9346.0/65536.0,1,-nbitq), 
to_sfixed(2213.0/65536.0,1,-nbitq), 
to_sfixed(-5267.0/65536.0,1,-nbitq), 
to_sfixed(1066.0/65536.0,1,-nbitq), 
to_sfixed(-7545.0/65536.0,1,-nbitq), 
to_sfixed(-1224.0/65536.0,1,-nbitq), 
to_sfixed(-632.0/65536.0,1,-nbitq), 
to_sfixed(2280.0/65536.0,1,-nbitq), 
to_sfixed(6757.0/65536.0,1,-nbitq), 
to_sfixed(1752.0/65536.0,1,-nbitq), 
to_sfixed(-9320.0/65536.0,1,-nbitq), 
to_sfixed(1454.0/65536.0,1,-nbitq), 
to_sfixed(8802.0/65536.0,1,-nbitq), 
to_sfixed(-1626.0/65536.0,1,-nbitq), 
to_sfixed(-5304.0/65536.0,1,-nbitq), 
to_sfixed(-1874.0/65536.0,1,-nbitq), 
to_sfixed(1793.0/65536.0,1,-nbitq), 
to_sfixed(-5309.0/65536.0,1,-nbitq), 
to_sfixed(-2117.0/65536.0,1,-nbitq), 
to_sfixed(-2544.0/65536.0,1,-nbitq), 
to_sfixed(921.0/65536.0,1,-nbitq), 
to_sfixed(-2361.0/65536.0,1,-nbitq), 
to_sfixed(-6822.0/65536.0,1,-nbitq), 
to_sfixed(769.0/65536.0,1,-nbitq), 
to_sfixed(-8229.0/65536.0,1,-nbitq), 
to_sfixed(-8008.0/65536.0,1,-nbitq), 
to_sfixed(-5690.0/65536.0,1,-nbitq), 
to_sfixed(414.0/65536.0,1,-nbitq), 
to_sfixed(216.0/65536.0,1,-nbitq), 
to_sfixed(1285.0/65536.0,1,-nbitq), 
to_sfixed(-1100.0/65536.0,1,-nbitq), 
to_sfixed(7.0/65536.0,1,-nbitq), 
to_sfixed(4304.0/65536.0,1,-nbitq), 
to_sfixed(13978.0/65536.0,1,-nbitq), 
to_sfixed(-5059.0/65536.0,1,-nbitq), 
to_sfixed(-2607.0/65536.0,1,-nbitq), 
to_sfixed(-2360.0/65536.0,1,-nbitq)  ), 
( to_sfixed(8018.0/65536.0,1,-nbitq), 
to_sfixed(-2893.0/65536.0,1,-nbitq), 
to_sfixed(1028.0/65536.0,1,-nbitq), 
to_sfixed(-1626.0/65536.0,1,-nbitq), 
to_sfixed(-7334.0/65536.0,1,-nbitq), 
to_sfixed(-4406.0/65536.0,1,-nbitq), 
to_sfixed(5572.0/65536.0,1,-nbitq), 
to_sfixed(-2562.0/65536.0,1,-nbitq), 
to_sfixed(-2989.0/65536.0,1,-nbitq), 
to_sfixed(1480.0/65536.0,1,-nbitq), 
to_sfixed(679.0/65536.0,1,-nbitq), 
to_sfixed(413.0/65536.0,1,-nbitq), 
to_sfixed(2228.0/65536.0,1,-nbitq), 
to_sfixed(-4473.0/65536.0,1,-nbitq), 
to_sfixed(1357.0/65536.0,1,-nbitq), 
to_sfixed(1479.0/65536.0,1,-nbitq), 
to_sfixed(147.0/65536.0,1,-nbitq), 
to_sfixed(6746.0/65536.0,1,-nbitq), 
to_sfixed(-5168.0/65536.0,1,-nbitq), 
to_sfixed(-1156.0/65536.0,1,-nbitq), 
to_sfixed(1643.0/65536.0,1,-nbitq), 
to_sfixed(2513.0/65536.0,1,-nbitq), 
to_sfixed(-1934.0/65536.0,1,-nbitq), 
to_sfixed(-3862.0/65536.0,1,-nbitq), 
to_sfixed(6968.0/65536.0,1,-nbitq), 
to_sfixed(-4510.0/65536.0,1,-nbitq), 
to_sfixed(7137.0/65536.0,1,-nbitq), 
to_sfixed(-867.0/65536.0,1,-nbitq), 
to_sfixed(-7452.0/65536.0,1,-nbitq), 
to_sfixed(3802.0/65536.0,1,-nbitq), 
to_sfixed(-12064.0/65536.0,1,-nbitq), 
to_sfixed(6579.0/65536.0,1,-nbitq), 
to_sfixed(-361.0/65536.0,1,-nbitq), 
to_sfixed(-12287.0/65536.0,1,-nbitq), 
to_sfixed(-958.0/65536.0,1,-nbitq), 
to_sfixed(1778.0/65536.0,1,-nbitq), 
to_sfixed(636.0/65536.0,1,-nbitq), 
to_sfixed(-3031.0/65536.0,1,-nbitq), 
to_sfixed(-5770.0/65536.0,1,-nbitq), 
to_sfixed(2737.0/65536.0,1,-nbitq), 
to_sfixed(7010.0/65536.0,1,-nbitq), 
to_sfixed(180.0/65536.0,1,-nbitq), 
to_sfixed(3121.0/65536.0,1,-nbitq), 
to_sfixed(-7294.0/65536.0,1,-nbitq), 
to_sfixed(620.0/65536.0,1,-nbitq), 
to_sfixed(749.0/65536.0,1,-nbitq), 
to_sfixed(1815.0/65536.0,1,-nbitq), 
to_sfixed(-7102.0/65536.0,1,-nbitq), 
to_sfixed(1378.0/65536.0,1,-nbitq), 
to_sfixed(-414.0/65536.0,1,-nbitq), 
to_sfixed(-2486.0/65536.0,1,-nbitq), 
to_sfixed(2999.0/65536.0,1,-nbitq), 
to_sfixed(6720.0/65536.0,1,-nbitq), 
to_sfixed(-7684.0/65536.0,1,-nbitq), 
to_sfixed(-797.0/65536.0,1,-nbitq), 
to_sfixed(5231.0/65536.0,1,-nbitq), 
to_sfixed(1051.0/65536.0,1,-nbitq), 
to_sfixed(-5839.0/65536.0,1,-nbitq), 
to_sfixed(2532.0/65536.0,1,-nbitq), 
to_sfixed(518.0/65536.0,1,-nbitq), 
to_sfixed(-3158.0/65536.0,1,-nbitq), 
to_sfixed(-1590.0/65536.0,1,-nbitq), 
to_sfixed(-894.0/65536.0,1,-nbitq), 
to_sfixed(-625.0/65536.0,1,-nbitq), 
to_sfixed(-6551.0/65536.0,1,-nbitq), 
to_sfixed(-2236.0/65536.0,1,-nbitq), 
to_sfixed(1945.0/65536.0,1,-nbitq), 
to_sfixed(274.0/65536.0,1,-nbitq), 
to_sfixed(-5580.0/65536.0,1,-nbitq), 
to_sfixed(-6914.0/65536.0,1,-nbitq), 
to_sfixed(2430.0/65536.0,1,-nbitq), 
to_sfixed(-6862.0/65536.0,1,-nbitq), 
to_sfixed(-537.0/65536.0,1,-nbitq), 
to_sfixed(-684.0/65536.0,1,-nbitq), 
to_sfixed(-2880.0/65536.0,1,-nbitq), 
to_sfixed(-1101.0/65536.0,1,-nbitq), 
to_sfixed(8237.0/65536.0,1,-nbitq), 
to_sfixed(-6390.0/65536.0,1,-nbitq), 
to_sfixed(-2735.0/65536.0,1,-nbitq), 
to_sfixed(3142.0/65536.0,1,-nbitq)  ), 
( to_sfixed(7601.0/65536.0,1,-nbitq), 
to_sfixed(180.0/65536.0,1,-nbitq), 
to_sfixed(4209.0/65536.0,1,-nbitq), 
to_sfixed(-2299.0/65536.0,1,-nbitq), 
to_sfixed(-1618.0/65536.0,1,-nbitq), 
to_sfixed(-3278.0/65536.0,1,-nbitq), 
to_sfixed(2184.0/65536.0,1,-nbitq), 
to_sfixed(-1104.0/65536.0,1,-nbitq), 
to_sfixed(-3211.0/65536.0,1,-nbitq), 
to_sfixed(-2345.0/65536.0,1,-nbitq), 
to_sfixed(-2878.0/65536.0,1,-nbitq), 
to_sfixed(-2707.0/65536.0,1,-nbitq), 
to_sfixed(-337.0/65536.0,1,-nbitq), 
to_sfixed(-5067.0/65536.0,1,-nbitq), 
to_sfixed(2295.0/65536.0,1,-nbitq), 
to_sfixed(2798.0/65536.0,1,-nbitq), 
to_sfixed(-1212.0/65536.0,1,-nbitq), 
to_sfixed(4606.0/65536.0,1,-nbitq), 
to_sfixed(-1917.0/65536.0,1,-nbitq), 
to_sfixed(-2267.0/65536.0,1,-nbitq), 
to_sfixed(2856.0/65536.0,1,-nbitq), 
to_sfixed(6059.0/65536.0,1,-nbitq), 
to_sfixed(-1084.0/65536.0,1,-nbitq), 
to_sfixed(-2302.0/65536.0,1,-nbitq), 
to_sfixed(6515.0/65536.0,1,-nbitq), 
to_sfixed(1014.0/65536.0,1,-nbitq), 
to_sfixed(7328.0/65536.0,1,-nbitq), 
to_sfixed(-3358.0/65536.0,1,-nbitq), 
to_sfixed(-12655.0/65536.0,1,-nbitq), 
to_sfixed(-986.0/65536.0,1,-nbitq), 
to_sfixed(-2544.0/65536.0,1,-nbitq), 
to_sfixed(6419.0/65536.0,1,-nbitq), 
to_sfixed(-2338.0/65536.0,1,-nbitq), 
to_sfixed(-6157.0/65536.0,1,-nbitq), 
to_sfixed(-983.0/65536.0,1,-nbitq), 
to_sfixed(2299.0/65536.0,1,-nbitq), 
to_sfixed(978.0/65536.0,1,-nbitq), 
to_sfixed(-4693.0/65536.0,1,-nbitq), 
to_sfixed(181.0/65536.0,1,-nbitq), 
to_sfixed(-1492.0/65536.0,1,-nbitq), 
to_sfixed(5969.0/65536.0,1,-nbitq), 
to_sfixed(2155.0/65536.0,1,-nbitq), 
to_sfixed(965.0/65536.0,1,-nbitq), 
to_sfixed(-5927.0/65536.0,1,-nbitq), 
to_sfixed(2416.0/65536.0,1,-nbitq), 
to_sfixed(5151.0/65536.0,1,-nbitq), 
to_sfixed(-1133.0/65536.0,1,-nbitq), 
to_sfixed(-3003.0/65536.0,1,-nbitq), 
to_sfixed(1676.0/65536.0,1,-nbitq), 
to_sfixed(-1302.0/65536.0,1,-nbitq), 
to_sfixed(1853.0/65536.0,1,-nbitq), 
to_sfixed(2971.0/65536.0,1,-nbitq), 
to_sfixed(-287.0/65536.0,1,-nbitq), 
to_sfixed(-1557.0/65536.0,1,-nbitq), 
to_sfixed(2020.0/65536.0,1,-nbitq), 
to_sfixed(4389.0/65536.0,1,-nbitq), 
to_sfixed(699.0/65536.0,1,-nbitq), 
to_sfixed(-2703.0/65536.0,1,-nbitq), 
to_sfixed(-2121.0/65536.0,1,-nbitq), 
to_sfixed(-1623.0/65536.0,1,-nbitq), 
to_sfixed(-2402.0/65536.0,1,-nbitq), 
to_sfixed(2317.0/65536.0,1,-nbitq), 
to_sfixed(2991.0/65536.0,1,-nbitq), 
to_sfixed(-420.0/65536.0,1,-nbitq), 
to_sfixed(-7833.0/65536.0,1,-nbitq), 
to_sfixed(-10079.0/65536.0,1,-nbitq), 
to_sfixed(484.0/65536.0,1,-nbitq), 
to_sfixed(-1322.0/65536.0,1,-nbitq), 
to_sfixed(-3195.0/65536.0,1,-nbitq), 
to_sfixed(-3442.0/65536.0,1,-nbitq), 
to_sfixed(-1946.0/65536.0,1,-nbitq), 
to_sfixed(-5069.0/65536.0,1,-nbitq), 
to_sfixed(2291.0/65536.0,1,-nbitq), 
to_sfixed(-2201.0/65536.0,1,-nbitq), 
to_sfixed(1314.0/65536.0,1,-nbitq), 
to_sfixed(-2070.0/65536.0,1,-nbitq), 
to_sfixed(1479.0/65536.0,1,-nbitq), 
to_sfixed(-3666.0/65536.0,1,-nbitq), 
to_sfixed(1187.0/65536.0,1,-nbitq), 
to_sfixed(-537.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4012.0/65536.0,1,-nbitq), 
to_sfixed(-4038.0/65536.0,1,-nbitq), 
to_sfixed(2775.0/65536.0,1,-nbitq), 
to_sfixed(-3343.0/65536.0,1,-nbitq), 
to_sfixed(-3114.0/65536.0,1,-nbitq), 
to_sfixed(-5698.0/65536.0,1,-nbitq), 
to_sfixed(415.0/65536.0,1,-nbitq), 
to_sfixed(-7416.0/65536.0,1,-nbitq), 
to_sfixed(-1272.0/65536.0,1,-nbitq), 
to_sfixed(-529.0/65536.0,1,-nbitq), 
to_sfixed(-3844.0/65536.0,1,-nbitq), 
to_sfixed(2877.0/65536.0,1,-nbitq), 
to_sfixed(3452.0/65536.0,1,-nbitq), 
to_sfixed(-3486.0/65536.0,1,-nbitq), 
to_sfixed(3886.0/65536.0,1,-nbitq), 
to_sfixed(1902.0/65536.0,1,-nbitq), 
to_sfixed(3031.0/65536.0,1,-nbitq), 
to_sfixed(1292.0/65536.0,1,-nbitq), 
to_sfixed(-3165.0/65536.0,1,-nbitq), 
to_sfixed(1808.0/65536.0,1,-nbitq), 
to_sfixed(4133.0/65536.0,1,-nbitq), 
to_sfixed(5405.0/65536.0,1,-nbitq), 
to_sfixed(-3627.0/65536.0,1,-nbitq), 
to_sfixed(622.0/65536.0,1,-nbitq), 
to_sfixed(4866.0/65536.0,1,-nbitq), 
to_sfixed(-2434.0/65536.0,1,-nbitq), 
to_sfixed(-1182.0/65536.0,1,-nbitq), 
to_sfixed(-482.0/65536.0,1,-nbitq), 
to_sfixed(-5745.0/65536.0,1,-nbitq), 
to_sfixed(2853.0/65536.0,1,-nbitq), 
to_sfixed(-2168.0/65536.0,1,-nbitq), 
to_sfixed(4726.0/65536.0,1,-nbitq), 
to_sfixed(3341.0/65536.0,1,-nbitq), 
to_sfixed(-2414.0/65536.0,1,-nbitq), 
to_sfixed(-1800.0/65536.0,1,-nbitq), 
to_sfixed(-1091.0/65536.0,1,-nbitq), 
to_sfixed(-3600.0/65536.0,1,-nbitq), 
to_sfixed(-4692.0/65536.0,1,-nbitq), 
to_sfixed(4218.0/65536.0,1,-nbitq), 
to_sfixed(1270.0/65536.0,1,-nbitq), 
to_sfixed(5533.0/65536.0,1,-nbitq), 
to_sfixed(-1939.0/65536.0,1,-nbitq), 
to_sfixed(3090.0/65536.0,1,-nbitq), 
to_sfixed(-7042.0/65536.0,1,-nbitq), 
to_sfixed(2324.0/65536.0,1,-nbitq), 
to_sfixed(5717.0/65536.0,1,-nbitq), 
to_sfixed(-1105.0/65536.0,1,-nbitq), 
to_sfixed(1122.0/65536.0,1,-nbitq), 
to_sfixed(-275.0/65536.0,1,-nbitq), 
to_sfixed(-281.0/65536.0,1,-nbitq), 
to_sfixed(1804.0/65536.0,1,-nbitq), 
to_sfixed(7678.0/65536.0,1,-nbitq), 
to_sfixed(874.0/65536.0,1,-nbitq), 
to_sfixed(-1944.0/65536.0,1,-nbitq), 
to_sfixed(-200.0/65536.0,1,-nbitq), 
to_sfixed(-498.0/65536.0,1,-nbitq), 
to_sfixed(2552.0/65536.0,1,-nbitq), 
to_sfixed(2942.0/65536.0,1,-nbitq), 
to_sfixed(138.0/65536.0,1,-nbitq), 
to_sfixed(-18.0/65536.0,1,-nbitq), 
to_sfixed(2338.0/65536.0,1,-nbitq), 
to_sfixed(2673.0/65536.0,1,-nbitq), 
to_sfixed(1378.0/65536.0,1,-nbitq), 
to_sfixed(-2687.0/65536.0,1,-nbitq), 
to_sfixed(-6936.0/65536.0,1,-nbitq), 
to_sfixed(-5286.0/65536.0,1,-nbitq), 
to_sfixed(-4447.0/65536.0,1,-nbitq), 
to_sfixed(-1503.0/65536.0,1,-nbitq), 
to_sfixed(-4126.0/65536.0,1,-nbitq), 
to_sfixed(863.0/65536.0,1,-nbitq), 
to_sfixed(-2416.0/65536.0,1,-nbitq), 
to_sfixed(2062.0/65536.0,1,-nbitq), 
to_sfixed(3001.0/65536.0,1,-nbitq), 
to_sfixed(-2888.0/65536.0,1,-nbitq), 
to_sfixed(-2246.0/65536.0,1,-nbitq), 
to_sfixed(55.0/65536.0,1,-nbitq), 
to_sfixed(-723.0/65536.0,1,-nbitq), 
to_sfixed(-148.0/65536.0,1,-nbitq), 
to_sfixed(1760.0/65536.0,1,-nbitq), 
to_sfixed(-139.0/65536.0,1,-nbitq)  ), 
( to_sfixed(667.0/65536.0,1,-nbitq), 
to_sfixed(93.0/65536.0,1,-nbitq), 
to_sfixed(6585.0/65536.0,1,-nbitq), 
to_sfixed(-3979.0/65536.0,1,-nbitq), 
to_sfixed(-4710.0/65536.0,1,-nbitq), 
to_sfixed(-5326.0/65536.0,1,-nbitq), 
to_sfixed(532.0/65536.0,1,-nbitq), 
to_sfixed(1088.0/65536.0,1,-nbitq), 
to_sfixed(-1334.0/65536.0,1,-nbitq), 
to_sfixed(-2682.0/65536.0,1,-nbitq), 
to_sfixed(-4388.0/65536.0,1,-nbitq), 
to_sfixed(1.0/65536.0,1,-nbitq), 
to_sfixed(3101.0/65536.0,1,-nbitq), 
to_sfixed(-6896.0/65536.0,1,-nbitq), 
to_sfixed(908.0/65536.0,1,-nbitq), 
to_sfixed(883.0/65536.0,1,-nbitq), 
to_sfixed(-2527.0/65536.0,1,-nbitq), 
to_sfixed(1628.0/65536.0,1,-nbitq), 
to_sfixed(-2865.0/65536.0,1,-nbitq), 
to_sfixed(-1206.0/65536.0,1,-nbitq), 
to_sfixed(-70.0/65536.0,1,-nbitq), 
to_sfixed(-126.0/65536.0,1,-nbitq), 
to_sfixed(-2696.0/65536.0,1,-nbitq), 
to_sfixed(-6418.0/65536.0,1,-nbitq), 
to_sfixed(6106.0/65536.0,1,-nbitq), 
to_sfixed(-6681.0/65536.0,1,-nbitq), 
to_sfixed(-5288.0/65536.0,1,-nbitq), 
to_sfixed(-2313.0/65536.0,1,-nbitq), 
to_sfixed(-916.0/65536.0,1,-nbitq), 
to_sfixed(3944.0/65536.0,1,-nbitq), 
to_sfixed(-6471.0/65536.0,1,-nbitq), 
to_sfixed(4931.0/65536.0,1,-nbitq), 
to_sfixed(-874.0/65536.0,1,-nbitq), 
to_sfixed(3765.0/65536.0,1,-nbitq), 
to_sfixed(3250.0/65536.0,1,-nbitq), 
to_sfixed(5.0/65536.0,1,-nbitq), 
to_sfixed(279.0/65536.0,1,-nbitq), 
to_sfixed(-4532.0/65536.0,1,-nbitq), 
to_sfixed(3676.0/65536.0,1,-nbitq), 
to_sfixed(2214.0/65536.0,1,-nbitq), 
to_sfixed(3420.0/65536.0,1,-nbitq), 
to_sfixed(-1122.0/65536.0,1,-nbitq), 
to_sfixed(491.0/65536.0,1,-nbitq), 
to_sfixed(-9068.0/65536.0,1,-nbitq), 
to_sfixed(-2071.0/65536.0,1,-nbitq), 
to_sfixed(843.0/65536.0,1,-nbitq), 
to_sfixed(-917.0/65536.0,1,-nbitq), 
to_sfixed(491.0/65536.0,1,-nbitq), 
to_sfixed(-799.0/65536.0,1,-nbitq), 
to_sfixed(3568.0/65536.0,1,-nbitq), 
to_sfixed(-1646.0/65536.0,1,-nbitq), 
to_sfixed(5703.0/65536.0,1,-nbitq), 
to_sfixed(-3931.0/65536.0,1,-nbitq), 
to_sfixed(3635.0/65536.0,1,-nbitq), 
to_sfixed(-1435.0/65536.0,1,-nbitq), 
to_sfixed(378.0/65536.0,1,-nbitq), 
to_sfixed(-1114.0/65536.0,1,-nbitq), 
to_sfixed(2921.0/65536.0,1,-nbitq), 
to_sfixed(-421.0/65536.0,1,-nbitq), 
to_sfixed(-3066.0/65536.0,1,-nbitq), 
to_sfixed(7295.0/65536.0,1,-nbitq), 
to_sfixed(702.0/65536.0,1,-nbitq), 
to_sfixed(156.0/65536.0,1,-nbitq), 
to_sfixed(-2092.0/65536.0,1,-nbitq), 
to_sfixed(-7081.0/65536.0,1,-nbitq), 
to_sfixed(-1600.0/65536.0,1,-nbitq), 
to_sfixed(-4688.0/65536.0,1,-nbitq), 
to_sfixed(-4281.0/65536.0,1,-nbitq), 
to_sfixed(-634.0/65536.0,1,-nbitq), 
to_sfixed(8672.0/65536.0,1,-nbitq), 
to_sfixed(-4134.0/65536.0,1,-nbitq), 
to_sfixed(5258.0/65536.0,1,-nbitq), 
to_sfixed(-4051.0/65536.0,1,-nbitq), 
to_sfixed(557.0/65536.0,1,-nbitq), 
to_sfixed(283.0/65536.0,1,-nbitq), 
to_sfixed(2088.0/65536.0,1,-nbitq), 
to_sfixed(-2473.0/65536.0,1,-nbitq), 
to_sfixed(-1182.0/65536.0,1,-nbitq), 
to_sfixed(-1358.0/65536.0,1,-nbitq), 
to_sfixed(1300.0/65536.0,1,-nbitq)  ), 
( to_sfixed(632.0/65536.0,1,-nbitq), 
to_sfixed(-829.0/65536.0,1,-nbitq), 
to_sfixed(4143.0/65536.0,1,-nbitq), 
to_sfixed(664.0/65536.0,1,-nbitq), 
to_sfixed(-8044.0/65536.0,1,-nbitq), 
to_sfixed(-5834.0/65536.0,1,-nbitq), 
to_sfixed(-2216.0/65536.0,1,-nbitq), 
to_sfixed(1326.0/65536.0,1,-nbitq), 
to_sfixed(2812.0/65536.0,1,-nbitq), 
to_sfixed(1315.0/65536.0,1,-nbitq), 
to_sfixed(970.0/65536.0,1,-nbitq), 
to_sfixed(-1894.0/65536.0,1,-nbitq), 
to_sfixed(-160.0/65536.0,1,-nbitq), 
to_sfixed(-6156.0/65536.0,1,-nbitq), 
to_sfixed(496.0/65536.0,1,-nbitq), 
to_sfixed(-187.0/65536.0,1,-nbitq), 
to_sfixed(-423.0/65536.0,1,-nbitq), 
to_sfixed(-1095.0/65536.0,1,-nbitq), 
to_sfixed(-1010.0/65536.0,1,-nbitq), 
to_sfixed(-1452.0/65536.0,1,-nbitq), 
to_sfixed(3623.0/65536.0,1,-nbitq), 
to_sfixed(1496.0/65536.0,1,-nbitq), 
to_sfixed(946.0/65536.0,1,-nbitq), 
to_sfixed(-6576.0/65536.0,1,-nbitq), 
to_sfixed(3016.0/65536.0,1,-nbitq), 
to_sfixed(-2024.0/65536.0,1,-nbitq), 
to_sfixed(-4745.0/65536.0,1,-nbitq), 
to_sfixed(-2355.0/65536.0,1,-nbitq), 
to_sfixed(2570.0/65536.0,1,-nbitq), 
to_sfixed(-1747.0/65536.0,1,-nbitq), 
to_sfixed(-6388.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(4326.0/65536.0,1,-nbitq), 
to_sfixed(698.0/65536.0,1,-nbitq), 
to_sfixed(115.0/65536.0,1,-nbitq), 
to_sfixed(1854.0/65536.0,1,-nbitq), 
to_sfixed(3116.0/65536.0,1,-nbitq), 
to_sfixed(789.0/65536.0,1,-nbitq), 
to_sfixed(2370.0/65536.0,1,-nbitq), 
to_sfixed(3303.0/65536.0,1,-nbitq), 
to_sfixed(2733.0/65536.0,1,-nbitq), 
to_sfixed(2130.0/65536.0,1,-nbitq), 
to_sfixed(-1496.0/65536.0,1,-nbitq), 
to_sfixed(-5023.0/65536.0,1,-nbitq), 
to_sfixed(2634.0/65536.0,1,-nbitq), 
to_sfixed(3240.0/65536.0,1,-nbitq), 
to_sfixed(226.0/65536.0,1,-nbitq), 
to_sfixed(-1539.0/65536.0,1,-nbitq), 
to_sfixed(2465.0/65536.0,1,-nbitq), 
to_sfixed(2488.0/65536.0,1,-nbitq), 
to_sfixed(2917.0/65536.0,1,-nbitq), 
to_sfixed(2864.0/65536.0,1,-nbitq), 
to_sfixed(-6849.0/65536.0,1,-nbitq), 
to_sfixed(3787.0/65536.0,1,-nbitq), 
to_sfixed(-4718.0/65536.0,1,-nbitq), 
to_sfixed(7308.0/65536.0,1,-nbitq), 
to_sfixed(2013.0/65536.0,1,-nbitq), 
to_sfixed(4447.0/65536.0,1,-nbitq), 
to_sfixed(89.0/65536.0,1,-nbitq), 
to_sfixed(-1622.0/65536.0,1,-nbitq), 
to_sfixed(2106.0/65536.0,1,-nbitq), 
to_sfixed(-1745.0/65536.0,1,-nbitq), 
to_sfixed(-2584.0/65536.0,1,-nbitq), 
to_sfixed(-2486.0/65536.0,1,-nbitq), 
to_sfixed(65.0/65536.0,1,-nbitq), 
to_sfixed(1788.0/65536.0,1,-nbitq), 
to_sfixed(1278.0/65536.0,1,-nbitq), 
to_sfixed(-547.0/65536.0,1,-nbitq), 
to_sfixed(6409.0/65536.0,1,-nbitq), 
to_sfixed(6842.0/65536.0,1,-nbitq), 
to_sfixed(-781.0/65536.0,1,-nbitq), 
to_sfixed(1801.0/65536.0,1,-nbitq), 
to_sfixed(-1440.0/65536.0,1,-nbitq), 
to_sfixed(-1922.0/65536.0,1,-nbitq), 
to_sfixed(-1586.0/65536.0,1,-nbitq), 
to_sfixed(2487.0/65536.0,1,-nbitq), 
to_sfixed(-2613.0/65536.0,1,-nbitq), 
to_sfixed(1842.0/65536.0,1,-nbitq), 
to_sfixed(1508.0/65536.0,1,-nbitq), 
to_sfixed(-237.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1134.0/65536.0,1,-nbitq), 
to_sfixed(-2106.0/65536.0,1,-nbitq), 
to_sfixed(-792.0/65536.0,1,-nbitq), 
to_sfixed(523.0/65536.0,1,-nbitq), 
to_sfixed(-820.0/65536.0,1,-nbitq), 
to_sfixed(-4775.0/65536.0,1,-nbitq), 
to_sfixed(-955.0/65536.0,1,-nbitq), 
to_sfixed(-1200.0/65536.0,1,-nbitq), 
to_sfixed(-2795.0/65536.0,1,-nbitq), 
to_sfixed(-2331.0/65536.0,1,-nbitq), 
to_sfixed(-2535.0/65536.0,1,-nbitq), 
to_sfixed(-21.0/65536.0,1,-nbitq), 
to_sfixed(2190.0/65536.0,1,-nbitq), 
to_sfixed(-5558.0/65536.0,1,-nbitq), 
to_sfixed(-2963.0/65536.0,1,-nbitq), 
to_sfixed(-1305.0/65536.0,1,-nbitq), 
to_sfixed(1251.0/65536.0,1,-nbitq), 
to_sfixed(-2494.0/65536.0,1,-nbitq), 
to_sfixed(-640.0/65536.0,1,-nbitq), 
to_sfixed(-1099.0/65536.0,1,-nbitq), 
to_sfixed(4264.0/65536.0,1,-nbitq), 
to_sfixed(262.0/65536.0,1,-nbitq), 
to_sfixed(-1544.0/65536.0,1,-nbitq), 
to_sfixed(-5290.0/65536.0,1,-nbitq), 
to_sfixed(3643.0/65536.0,1,-nbitq), 
to_sfixed(-5132.0/65536.0,1,-nbitq), 
to_sfixed(-7442.0/65536.0,1,-nbitq), 
to_sfixed(-3836.0/65536.0,1,-nbitq), 
to_sfixed(1749.0/65536.0,1,-nbitq), 
to_sfixed(48.0/65536.0,1,-nbitq), 
to_sfixed(-1347.0/65536.0,1,-nbitq), 
to_sfixed(825.0/65536.0,1,-nbitq), 
to_sfixed(5024.0/65536.0,1,-nbitq), 
to_sfixed(681.0/65536.0,1,-nbitq), 
to_sfixed(-1200.0/65536.0,1,-nbitq), 
to_sfixed(2859.0/65536.0,1,-nbitq), 
to_sfixed(786.0/65536.0,1,-nbitq), 
to_sfixed(972.0/65536.0,1,-nbitq), 
to_sfixed(-2360.0/65536.0,1,-nbitq), 
to_sfixed(1592.0/65536.0,1,-nbitq), 
to_sfixed(-2474.0/65536.0,1,-nbitq), 
to_sfixed(2314.0/65536.0,1,-nbitq), 
to_sfixed(2338.0/65536.0,1,-nbitq), 
to_sfixed(1729.0/65536.0,1,-nbitq), 
to_sfixed(379.0/65536.0,1,-nbitq), 
to_sfixed(5511.0/65536.0,1,-nbitq), 
to_sfixed(1995.0/65536.0,1,-nbitq), 
to_sfixed(-2989.0/65536.0,1,-nbitq), 
to_sfixed(2514.0/65536.0,1,-nbitq), 
to_sfixed(2416.0/65536.0,1,-nbitq), 
to_sfixed(-825.0/65536.0,1,-nbitq), 
to_sfixed(2989.0/65536.0,1,-nbitq), 
to_sfixed(-2037.0/65536.0,1,-nbitq), 
to_sfixed(5381.0/65536.0,1,-nbitq), 
to_sfixed(-3025.0/65536.0,1,-nbitq), 
to_sfixed(978.0/65536.0,1,-nbitq), 
to_sfixed(2829.0/65536.0,1,-nbitq), 
to_sfixed(6176.0/65536.0,1,-nbitq), 
to_sfixed(2570.0/65536.0,1,-nbitq), 
to_sfixed(-1625.0/65536.0,1,-nbitq), 
to_sfixed(-695.0/65536.0,1,-nbitq), 
to_sfixed(1182.0/65536.0,1,-nbitq), 
to_sfixed(-1214.0/65536.0,1,-nbitq), 
to_sfixed(371.0/65536.0,1,-nbitq), 
to_sfixed(-3697.0/65536.0,1,-nbitq), 
to_sfixed(-2659.0/65536.0,1,-nbitq), 
to_sfixed(1935.0/65536.0,1,-nbitq), 
to_sfixed(2796.0/65536.0,1,-nbitq), 
to_sfixed(4997.0/65536.0,1,-nbitq), 
to_sfixed(3485.0/65536.0,1,-nbitq), 
to_sfixed(-2296.0/65536.0,1,-nbitq), 
to_sfixed(-3050.0/65536.0,1,-nbitq), 
to_sfixed(3412.0/65536.0,1,-nbitq), 
to_sfixed(395.0/65536.0,1,-nbitq), 
to_sfixed(628.0/65536.0,1,-nbitq), 
to_sfixed(-503.0/65536.0,1,-nbitq), 
to_sfixed(-4985.0/65536.0,1,-nbitq), 
to_sfixed(-755.0/65536.0,1,-nbitq), 
to_sfixed(-1975.0/65536.0,1,-nbitq), 
to_sfixed(-1551.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2177.0/65536.0,1,-nbitq), 
to_sfixed(-2273.0/65536.0,1,-nbitq), 
to_sfixed(-3020.0/65536.0,1,-nbitq), 
to_sfixed(-3418.0/65536.0,1,-nbitq), 
to_sfixed(511.0/65536.0,1,-nbitq), 
to_sfixed(1469.0/65536.0,1,-nbitq), 
to_sfixed(-1703.0/65536.0,1,-nbitq), 
to_sfixed(1982.0/65536.0,1,-nbitq), 
to_sfixed(-2003.0/65536.0,1,-nbitq), 
to_sfixed(-1782.0/65536.0,1,-nbitq), 
to_sfixed(-2591.0/65536.0,1,-nbitq), 
to_sfixed(-725.0/65536.0,1,-nbitq), 
to_sfixed(2508.0/65536.0,1,-nbitq), 
to_sfixed(-3642.0/65536.0,1,-nbitq), 
to_sfixed(815.0/65536.0,1,-nbitq), 
to_sfixed(-1996.0/65536.0,1,-nbitq), 
to_sfixed(-1799.0/65536.0,1,-nbitq), 
to_sfixed(1405.0/65536.0,1,-nbitq), 
to_sfixed(-308.0/65536.0,1,-nbitq), 
to_sfixed(3396.0/65536.0,1,-nbitq), 
to_sfixed(-1895.0/65536.0,1,-nbitq), 
to_sfixed(4201.0/65536.0,1,-nbitq), 
to_sfixed(-3541.0/65536.0,1,-nbitq), 
to_sfixed(-5258.0/65536.0,1,-nbitq), 
to_sfixed(115.0/65536.0,1,-nbitq), 
to_sfixed(-5078.0/65536.0,1,-nbitq), 
to_sfixed(-1794.0/65536.0,1,-nbitq), 
to_sfixed(-2221.0/65536.0,1,-nbitq), 
to_sfixed(4226.0/65536.0,1,-nbitq), 
to_sfixed(-1186.0/65536.0,1,-nbitq), 
to_sfixed(-3072.0/65536.0,1,-nbitq), 
to_sfixed(-566.0/65536.0,1,-nbitq), 
to_sfixed(2022.0/65536.0,1,-nbitq), 
to_sfixed(929.0/65536.0,1,-nbitq), 
to_sfixed(479.0/65536.0,1,-nbitq), 
to_sfixed(-994.0/65536.0,1,-nbitq), 
to_sfixed(23.0/65536.0,1,-nbitq), 
to_sfixed(-1361.0/65536.0,1,-nbitq), 
to_sfixed(-1123.0/65536.0,1,-nbitq), 
to_sfixed(2387.0/65536.0,1,-nbitq), 
to_sfixed(802.0/65536.0,1,-nbitq), 
to_sfixed(-1491.0/65536.0,1,-nbitq), 
to_sfixed(-275.0/65536.0,1,-nbitq), 
to_sfixed(2288.0/65536.0,1,-nbitq), 
to_sfixed(2698.0/65536.0,1,-nbitq), 
to_sfixed(3519.0/65536.0,1,-nbitq), 
to_sfixed(2547.0/65536.0,1,-nbitq), 
to_sfixed(980.0/65536.0,1,-nbitq), 
to_sfixed(-2645.0/65536.0,1,-nbitq), 
to_sfixed(4474.0/65536.0,1,-nbitq), 
to_sfixed(101.0/65536.0,1,-nbitq), 
to_sfixed(-547.0/65536.0,1,-nbitq), 
to_sfixed(-3998.0/65536.0,1,-nbitq), 
to_sfixed(5774.0/65536.0,1,-nbitq), 
to_sfixed(-466.0/65536.0,1,-nbitq), 
to_sfixed(914.0/65536.0,1,-nbitq), 
to_sfixed(1526.0/65536.0,1,-nbitq), 
to_sfixed(3042.0/65536.0,1,-nbitq), 
to_sfixed(681.0/65536.0,1,-nbitq), 
to_sfixed(-3319.0/65536.0,1,-nbitq), 
to_sfixed(-289.0/65536.0,1,-nbitq), 
to_sfixed(-737.0/65536.0,1,-nbitq), 
to_sfixed(1288.0/65536.0,1,-nbitq), 
to_sfixed(-948.0/65536.0,1,-nbitq), 
to_sfixed(-955.0/65536.0,1,-nbitq), 
to_sfixed(-335.0/65536.0,1,-nbitq), 
to_sfixed(2033.0/65536.0,1,-nbitq), 
to_sfixed(3367.0/65536.0,1,-nbitq), 
to_sfixed(3553.0/65536.0,1,-nbitq), 
to_sfixed(4177.0/65536.0,1,-nbitq), 
to_sfixed(-42.0/65536.0,1,-nbitq), 
to_sfixed(1882.0/65536.0,1,-nbitq), 
to_sfixed(-287.0/65536.0,1,-nbitq), 
to_sfixed(-2593.0/65536.0,1,-nbitq), 
to_sfixed(-2658.0/65536.0,1,-nbitq), 
to_sfixed(-859.0/65536.0,1,-nbitq), 
to_sfixed(-2314.0/65536.0,1,-nbitq), 
to_sfixed(3918.0/65536.0,1,-nbitq), 
to_sfixed(-1771.0/65536.0,1,-nbitq), 
to_sfixed(2899.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3334.0/65536.0,1,-nbitq), 
to_sfixed(-2419.0/65536.0,1,-nbitq), 
to_sfixed(-2889.0/65536.0,1,-nbitq), 
to_sfixed(1850.0/65536.0,1,-nbitq), 
to_sfixed(-765.0/65536.0,1,-nbitq), 
to_sfixed(-4087.0/65536.0,1,-nbitq), 
to_sfixed(1906.0/65536.0,1,-nbitq), 
to_sfixed(3103.0/65536.0,1,-nbitq), 
to_sfixed(-1324.0/65536.0,1,-nbitq), 
to_sfixed(-299.0/65536.0,1,-nbitq), 
to_sfixed(-701.0/65536.0,1,-nbitq), 
to_sfixed(369.0/65536.0,1,-nbitq), 
to_sfixed(1459.0/65536.0,1,-nbitq), 
to_sfixed(328.0/65536.0,1,-nbitq), 
to_sfixed(-2998.0/65536.0,1,-nbitq), 
to_sfixed(787.0/65536.0,1,-nbitq), 
to_sfixed(743.0/65536.0,1,-nbitq), 
to_sfixed(1053.0/65536.0,1,-nbitq), 
to_sfixed(3155.0/65536.0,1,-nbitq), 
to_sfixed(-216.0/65536.0,1,-nbitq), 
to_sfixed(-2811.0/65536.0,1,-nbitq), 
to_sfixed(1015.0/65536.0,1,-nbitq), 
to_sfixed(-4119.0/65536.0,1,-nbitq), 
to_sfixed(-2948.0/65536.0,1,-nbitq), 
to_sfixed(2237.0/65536.0,1,-nbitq), 
to_sfixed(-2767.0/65536.0,1,-nbitq), 
to_sfixed(-587.0/65536.0,1,-nbitq), 
to_sfixed(1340.0/65536.0,1,-nbitq), 
to_sfixed(2738.0/65536.0,1,-nbitq), 
to_sfixed(-611.0/65536.0,1,-nbitq), 
to_sfixed(-1647.0/65536.0,1,-nbitq), 
to_sfixed(578.0/65536.0,1,-nbitq), 
to_sfixed(566.0/65536.0,1,-nbitq), 
to_sfixed(2672.0/65536.0,1,-nbitq), 
to_sfixed(1305.0/65536.0,1,-nbitq), 
to_sfixed(-753.0/65536.0,1,-nbitq), 
to_sfixed(-2376.0/65536.0,1,-nbitq), 
to_sfixed(-1319.0/65536.0,1,-nbitq), 
to_sfixed(463.0/65536.0,1,-nbitq), 
to_sfixed(2826.0/65536.0,1,-nbitq), 
to_sfixed(-1663.0/65536.0,1,-nbitq), 
to_sfixed(-3233.0/65536.0,1,-nbitq), 
to_sfixed(-4300.0/65536.0,1,-nbitq), 
to_sfixed(2878.0/65536.0,1,-nbitq), 
to_sfixed(3002.0/65536.0,1,-nbitq), 
to_sfixed(3821.0/65536.0,1,-nbitq), 
to_sfixed(2662.0/65536.0,1,-nbitq), 
to_sfixed(-327.0/65536.0,1,-nbitq), 
to_sfixed(893.0/65536.0,1,-nbitq), 
to_sfixed(2566.0/65536.0,1,-nbitq), 
to_sfixed(3197.0/65536.0,1,-nbitq), 
to_sfixed(1747.0/65536.0,1,-nbitq), 
to_sfixed(-2011.0/65536.0,1,-nbitq), 
to_sfixed(1264.0/65536.0,1,-nbitq), 
to_sfixed(2414.0/65536.0,1,-nbitq), 
to_sfixed(-2479.0/65536.0,1,-nbitq), 
to_sfixed(-2460.0/65536.0,1,-nbitq), 
to_sfixed(724.0/65536.0,1,-nbitq), 
to_sfixed(-2905.0/65536.0,1,-nbitq), 
to_sfixed(2143.0/65536.0,1,-nbitq), 
to_sfixed(-1998.0/65536.0,1,-nbitq), 
to_sfixed(-341.0/65536.0,1,-nbitq), 
to_sfixed(1098.0/65536.0,1,-nbitq), 
to_sfixed(-3141.0/65536.0,1,-nbitq), 
to_sfixed(1489.0/65536.0,1,-nbitq), 
to_sfixed(-2930.0/65536.0,1,-nbitq), 
to_sfixed(2015.0/65536.0,1,-nbitq), 
to_sfixed(387.0/65536.0,1,-nbitq), 
to_sfixed(1816.0/65536.0,1,-nbitq), 
to_sfixed(3259.0/65536.0,1,-nbitq), 
to_sfixed(-1108.0/65536.0,1,-nbitq), 
to_sfixed(-1572.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(1610.0/65536.0,1,-nbitq), 
to_sfixed(1228.0/65536.0,1,-nbitq), 
to_sfixed(3336.0/65536.0,1,-nbitq), 
to_sfixed(-3719.0/65536.0,1,-nbitq), 
to_sfixed(1594.0/65536.0,1,-nbitq), 
to_sfixed(777.0/65536.0,1,-nbitq), 
to_sfixed(1859.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1924.0/65536.0,1,-nbitq), 
to_sfixed(1553.0/65536.0,1,-nbitq), 
to_sfixed(359.0/65536.0,1,-nbitq), 
to_sfixed(2214.0/65536.0,1,-nbitq), 
to_sfixed(-3465.0/65536.0,1,-nbitq), 
to_sfixed(95.0/65536.0,1,-nbitq), 
to_sfixed(1558.0/65536.0,1,-nbitq), 
to_sfixed(-137.0/65536.0,1,-nbitq), 
to_sfixed(502.0/65536.0,1,-nbitq), 
to_sfixed(1859.0/65536.0,1,-nbitq), 
to_sfixed(-2626.0/65536.0,1,-nbitq), 
to_sfixed(1753.0/65536.0,1,-nbitq), 
to_sfixed(2462.0/65536.0,1,-nbitq), 
to_sfixed(1441.0/65536.0,1,-nbitq), 
to_sfixed(1863.0/65536.0,1,-nbitq), 
to_sfixed(215.0/65536.0,1,-nbitq), 
to_sfixed(-3182.0/65536.0,1,-nbitq), 
to_sfixed(-1849.0/65536.0,1,-nbitq), 
to_sfixed(-1266.0/65536.0,1,-nbitq), 
to_sfixed(2210.0/65536.0,1,-nbitq), 
to_sfixed(-962.0/65536.0,1,-nbitq), 
to_sfixed(2335.0/65536.0,1,-nbitq), 
to_sfixed(-2244.0/65536.0,1,-nbitq), 
to_sfixed(-3324.0/65536.0,1,-nbitq), 
to_sfixed(-2417.0/65536.0,1,-nbitq), 
to_sfixed(688.0/65536.0,1,-nbitq), 
to_sfixed(-4726.0/65536.0,1,-nbitq), 
to_sfixed(2930.0/65536.0,1,-nbitq), 
to_sfixed(2393.0/65536.0,1,-nbitq), 
to_sfixed(-1564.0/65536.0,1,-nbitq), 
to_sfixed(2402.0/65536.0,1,-nbitq), 
to_sfixed(503.0/65536.0,1,-nbitq), 
to_sfixed(-444.0/65536.0,1,-nbitq), 
to_sfixed(-1625.0/65536.0,1,-nbitq), 
to_sfixed(-2697.0/65536.0,1,-nbitq), 
to_sfixed(-511.0/65536.0,1,-nbitq), 
to_sfixed(-1846.0/65536.0,1,-nbitq), 
to_sfixed(1817.0/65536.0,1,-nbitq), 
to_sfixed(863.0/65536.0,1,-nbitq), 
to_sfixed(1206.0/65536.0,1,-nbitq), 
to_sfixed(-2406.0/65536.0,1,-nbitq), 
to_sfixed(-1907.0/65536.0,1,-nbitq), 
to_sfixed(-1788.0/65536.0,1,-nbitq), 
to_sfixed(750.0/65536.0,1,-nbitq), 
to_sfixed(1883.0/65536.0,1,-nbitq), 
to_sfixed(1709.0/65536.0,1,-nbitq), 
to_sfixed(-1271.0/65536.0,1,-nbitq), 
to_sfixed(-562.0/65536.0,1,-nbitq), 
to_sfixed(3147.0/65536.0,1,-nbitq), 
to_sfixed(942.0/65536.0,1,-nbitq), 
to_sfixed(301.0/65536.0,1,-nbitq), 
to_sfixed(-1424.0/65536.0,1,-nbitq), 
to_sfixed(579.0/65536.0,1,-nbitq), 
to_sfixed(-1747.0/65536.0,1,-nbitq), 
to_sfixed(105.0/65536.0,1,-nbitq), 
to_sfixed(3.0/65536.0,1,-nbitq), 
to_sfixed(233.0/65536.0,1,-nbitq), 
to_sfixed(325.0/65536.0,1,-nbitq), 
to_sfixed(2336.0/65536.0,1,-nbitq), 
to_sfixed(3710.0/65536.0,1,-nbitq), 
to_sfixed(1644.0/65536.0,1,-nbitq), 
to_sfixed(1589.0/65536.0,1,-nbitq), 
to_sfixed(-150.0/65536.0,1,-nbitq), 
to_sfixed(-2013.0/65536.0,1,-nbitq), 
to_sfixed(-1938.0/65536.0,1,-nbitq), 
to_sfixed(-872.0/65536.0,1,-nbitq), 
to_sfixed(195.0/65536.0,1,-nbitq), 
to_sfixed(-579.0/65536.0,1,-nbitq), 
to_sfixed(4497.0/65536.0,1,-nbitq), 
to_sfixed(3109.0/65536.0,1,-nbitq), 
to_sfixed(639.0/65536.0,1,-nbitq), 
to_sfixed(858.0/65536.0,1,-nbitq), 
to_sfixed(-876.0/65536.0,1,-nbitq), 
to_sfixed(-905.0/65536.0,1,-nbitq), 
to_sfixed(2470.0/65536.0,1,-nbitq), 
to_sfixed(-642.0/65536.0,1,-nbitq), 
to_sfixed(-2728.0/65536.0,1,-nbitq), 
to_sfixed(1054.0/65536.0,1,-nbitq), 
to_sfixed(549.0/65536.0,1,-nbitq), 
to_sfixed(1630.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1062.0/65536.0,1,-nbitq), 
to_sfixed(-793.0/65536.0,1,-nbitq), 
to_sfixed(4052.0/65536.0,1,-nbitq), 
to_sfixed(480.0/65536.0,1,-nbitq), 
to_sfixed(-4467.0/65536.0,1,-nbitq), 
to_sfixed(-4023.0/65536.0,1,-nbitq), 
to_sfixed(-3161.0/65536.0,1,-nbitq), 
to_sfixed(2559.0/65536.0,1,-nbitq), 
to_sfixed(-2884.0/65536.0,1,-nbitq), 
to_sfixed(-368.0/65536.0,1,-nbitq), 
to_sfixed(-557.0/65536.0,1,-nbitq), 
to_sfixed(-2932.0/65536.0,1,-nbitq), 
to_sfixed(-2839.0/65536.0,1,-nbitq), 
to_sfixed(-25.0/65536.0,1,-nbitq), 
to_sfixed(167.0/65536.0,1,-nbitq), 
to_sfixed(-1630.0/65536.0,1,-nbitq), 
to_sfixed(-2011.0/65536.0,1,-nbitq), 
to_sfixed(348.0/65536.0,1,-nbitq), 
to_sfixed(2814.0/65536.0,1,-nbitq), 
to_sfixed(734.0/65536.0,1,-nbitq), 
to_sfixed(-510.0/65536.0,1,-nbitq), 
to_sfixed(-718.0/65536.0,1,-nbitq), 
to_sfixed(195.0/65536.0,1,-nbitq), 
to_sfixed(2789.0/65536.0,1,-nbitq), 
to_sfixed(-1305.0/65536.0,1,-nbitq), 
to_sfixed(2714.0/65536.0,1,-nbitq), 
to_sfixed(-3726.0/65536.0,1,-nbitq), 
to_sfixed(-442.0/65536.0,1,-nbitq), 
to_sfixed(-1397.0/65536.0,1,-nbitq), 
to_sfixed(1731.0/65536.0,1,-nbitq), 
to_sfixed(-444.0/65536.0,1,-nbitq), 
to_sfixed(2666.0/65536.0,1,-nbitq), 
to_sfixed(-3338.0/65536.0,1,-nbitq), 
to_sfixed(-4132.0/65536.0,1,-nbitq), 
to_sfixed(2251.0/65536.0,1,-nbitq), 
to_sfixed(-91.0/65536.0,1,-nbitq), 
to_sfixed(-1017.0/65536.0,1,-nbitq), 
to_sfixed(-1264.0/65536.0,1,-nbitq), 
to_sfixed(-930.0/65536.0,1,-nbitq), 
to_sfixed(-1364.0/65536.0,1,-nbitq), 
to_sfixed(-1618.0/65536.0,1,-nbitq), 
to_sfixed(206.0/65536.0,1,-nbitq), 
to_sfixed(166.0/65536.0,1,-nbitq), 
to_sfixed(2583.0/65536.0,1,-nbitq), 
to_sfixed(1213.0/65536.0,1,-nbitq), 
to_sfixed(5717.0/65536.0,1,-nbitq), 
to_sfixed(2945.0/65536.0,1,-nbitq), 
to_sfixed(1427.0/65536.0,1,-nbitq), 
to_sfixed(2328.0/65536.0,1,-nbitq), 
to_sfixed(814.0/65536.0,1,-nbitq), 
to_sfixed(2074.0/65536.0,1,-nbitq), 
to_sfixed(-1968.0/65536.0,1,-nbitq), 
to_sfixed(46.0/65536.0,1,-nbitq), 
to_sfixed(-1632.0/65536.0,1,-nbitq), 
to_sfixed(-1059.0/65536.0,1,-nbitq), 
to_sfixed(3041.0/65536.0,1,-nbitq), 
to_sfixed(-348.0/65536.0,1,-nbitq), 
to_sfixed(-1013.0/65536.0,1,-nbitq), 
to_sfixed(1372.0/65536.0,1,-nbitq), 
to_sfixed(2375.0/65536.0,1,-nbitq), 
to_sfixed(-682.0/65536.0,1,-nbitq), 
to_sfixed(677.0/65536.0,1,-nbitq), 
to_sfixed(-2660.0/65536.0,1,-nbitq), 
to_sfixed(-982.0/65536.0,1,-nbitq), 
to_sfixed(6162.0/65536.0,1,-nbitq), 
to_sfixed(802.0/65536.0,1,-nbitq), 
to_sfixed(2962.0/65536.0,1,-nbitq), 
to_sfixed(837.0/65536.0,1,-nbitq), 
to_sfixed(2218.0/65536.0,1,-nbitq), 
to_sfixed(624.0/65536.0,1,-nbitq), 
to_sfixed(2235.0/65536.0,1,-nbitq), 
to_sfixed(-2640.0/65536.0,1,-nbitq), 
to_sfixed(2856.0/65536.0,1,-nbitq), 
to_sfixed(-2667.0/65536.0,1,-nbitq), 
to_sfixed(-2908.0/65536.0,1,-nbitq), 
to_sfixed(-840.0/65536.0,1,-nbitq), 
to_sfixed(-594.0/65536.0,1,-nbitq), 
to_sfixed(-504.0/65536.0,1,-nbitq), 
to_sfixed(2000.0/65536.0,1,-nbitq), 
to_sfixed(2118.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2659.0/65536.0,1,-nbitq), 
to_sfixed(-1044.0/65536.0,1,-nbitq), 
to_sfixed(-554.0/65536.0,1,-nbitq), 
to_sfixed(-2601.0/65536.0,1,-nbitq), 
to_sfixed(-2589.0/65536.0,1,-nbitq), 
to_sfixed(-1740.0/65536.0,1,-nbitq), 
to_sfixed(-1301.0/65536.0,1,-nbitq), 
to_sfixed(-237.0/65536.0,1,-nbitq), 
to_sfixed(-2098.0/65536.0,1,-nbitq), 
to_sfixed(433.0/65536.0,1,-nbitq), 
to_sfixed(1969.0/65536.0,1,-nbitq), 
to_sfixed(3059.0/65536.0,1,-nbitq), 
to_sfixed(-730.0/65536.0,1,-nbitq), 
to_sfixed(277.0/65536.0,1,-nbitq), 
to_sfixed(-1363.0/65536.0,1,-nbitq), 
to_sfixed(-578.0/65536.0,1,-nbitq), 
to_sfixed(-617.0/65536.0,1,-nbitq), 
to_sfixed(734.0/65536.0,1,-nbitq), 
to_sfixed(1016.0/65536.0,1,-nbitq), 
to_sfixed(1173.0/65536.0,1,-nbitq), 
to_sfixed(1581.0/65536.0,1,-nbitq), 
to_sfixed(-2599.0/65536.0,1,-nbitq), 
to_sfixed(-1475.0/65536.0,1,-nbitq), 
to_sfixed(3306.0/65536.0,1,-nbitq), 
to_sfixed(2853.0/65536.0,1,-nbitq), 
to_sfixed(249.0/65536.0,1,-nbitq), 
to_sfixed(-2983.0/65536.0,1,-nbitq), 
to_sfixed(1947.0/65536.0,1,-nbitq), 
to_sfixed(698.0/65536.0,1,-nbitq), 
to_sfixed(-1084.0/65536.0,1,-nbitq), 
to_sfixed(-769.0/65536.0,1,-nbitq), 
to_sfixed(-2023.0/65536.0,1,-nbitq), 
to_sfixed(-3930.0/65536.0,1,-nbitq), 
to_sfixed(27.0/65536.0,1,-nbitq), 
to_sfixed(-2690.0/65536.0,1,-nbitq), 
to_sfixed(967.0/65536.0,1,-nbitq), 
to_sfixed(93.0/65536.0,1,-nbitq), 
to_sfixed(-3725.0/65536.0,1,-nbitq), 
to_sfixed(757.0/65536.0,1,-nbitq), 
to_sfixed(1298.0/65536.0,1,-nbitq), 
to_sfixed(2565.0/65536.0,1,-nbitq), 
to_sfixed(-110.0/65536.0,1,-nbitq), 
to_sfixed(1176.0/65536.0,1,-nbitq), 
to_sfixed(3909.0/65536.0,1,-nbitq), 
to_sfixed(150.0/65536.0,1,-nbitq), 
to_sfixed(1655.0/65536.0,1,-nbitq), 
to_sfixed(-2337.0/65536.0,1,-nbitq), 
to_sfixed(1946.0/65536.0,1,-nbitq), 
to_sfixed(128.0/65536.0,1,-nbitq), 
to_sfixed(3071.0/65536.0,1,-nbitq), 
to_sfixed(713.0/65536.0,1,-nbitq), 
to_sfixed(802.0/65536.0,1,-nbitq), 
to_sfixed(-420.0/65536.0,1,-nbitq), 
to_sfixed(-2748.0/65536.0,1,-nbitq), 
to_sfixed(-1418.0/65536.0,1,-nbitq), 
to_sfixed(2180.0/65536.0,1,-nbitq), 
to_sfixed(-816.0/65536.0,1,-nbitq), 
to_sfixed(840.0/65536.0,1,-nbitq), 
to_sfixed(-2575.0/65536.0,1,-nbitq), 
to_sfixed(3487.0/65536.0,1,-nbitq), 
to_sfixed(-3334.0/65536.0,1,-nbitq), 
to_sfixed(-1676.0/65536.0,1,-nbitq), 
to_sfixed(-353.0/65536.0,1,-nbitq), 
to_sfixed(906.0/65536.0,1,-nbitq), 
to_sfixed(5550.0/65536.0,1,-nbitq), 
to_sfixed(2366.0/65536.0,1,-nbitq), 
to_sfixed(-1575.0/65536.0,1,-nbitq), 
to_sfixed(-3408.0/65536.0,1,-nbitq), 
to_sfixed(3542.0/65536.0,1,-nbitq), 
to_sfixed(485.0/65536.0,1,-nbitq), 
to_sfixed(-1802.0/65536.0,1,-nbitq), 
to_sfixed(686.0/65536.0,1,-nbitq), 
to_sfixed(-24.0/65536.0,1,-nbitq), 
to_sfixed(-1327.0/65536.0,1,-nbitq), 
to_sfixed(-3183.0/65536.0,1,-nbitq), 
to_sfixed(-18.0/65536.0,1,-nbitq), 
to_sfixed(-864.0/65536.0,1,-nbitq), 
to_sfixed(-357.0/65536.0,1,-nbitq), 
to_sfixed(1056.0/65536.0,1,-nbitq), 
to_sfixed(2520.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1964.0/65536.0,1,-nbitq), 
to_sfixed(-767.0/65536.0,1,-nbitq), 
to_sfixed(-1092.0/65536.0,1,-nbitq), 
to_sfixed(-38.0/65536.0,1,-nbitq), 
to_sfixed(-1723.0/65536.0,1,-nbitq), 
to_sfixed(-1681.0/65536.0,1,-nbitq), 
to_sfixed(-3615.0/65536.0,1,-nbitq), 
to_sfixed(1989.0/65536.0,1,-nbitq), 
to_sfixed(-12.0/65536.0,1,-nbitq), 
to_sfixed(-2192.0/65536.0,1,-nbitq), 
to_sfixed(-50.0/65536.0,1,-nbitq), 
to_sfixed(2941.0/65536.0,1,-nbitq), 
to_sfixed(1783.0/65536.0,1,-nbitq), 
to_sfixed(2181.0/65536.0,1,-nbitq), 
to_sfixed(-1105.0/65536.0,1,-nbitq), 
to_sfixed(1114.0/65536.0,1,-nbitq), 
to_sfixed(2361.0/65536.0,1,-nbitq), 
to_sfixed(806.0/65536.0,1,-nbitq), 
to_sfixed(2561.0/65536.0,1,-nbitq), 
to_sfixed(1647.0/65536.0,1,-nbitq), 
to_sfixed(835.0/65536.0,1,-nbitq), 
to_sfixed(1386.0/65536.0,1,-nbitq), 
to_sfixed(2389.0/65536.0,1,-nbitq), 
to_sfixed(-1735.0/65536.0,1,-nbitq), 
to_sfixed(-3072.0/65536.0,1,-nbitq), 
to_sfixed(3607.0/65536.0,1,-nbitq), 
to_sfixed(-737.0/65536.0,1,-nbitq), 
to_sfixed(-1257.0/65536.0,1,-nbitq), 
to_sfixed(-906.0/65536.0,1,-nbitq), 
to_sfixed(1030.0/65536.0,1,-nbitq), 
to_sfixed(-2270.0/65536.0,1,-nbitq), 
to_sfixed(-759.0/65536.0,1,-nbitq), 
to_sfixed(-3223.0/65536.0,1,-nbitq), 
to_sfixed(-892.0/65536.0,1,-nbitq), 
to_sfixed(809.0/65536.0,1,-nbitq), 
to_sfixed(-493.0/65536.0,1,-nbitq), 
to_sfixed(-492.0/65536.0,1,-nbitq), 
to_sfixed(-410.0/65536.0,1,-nbitq), 
to_sfixed(1760.0/65536.0,1,-nbitq), 
to_sfixed(1276.0/65536.0,1,-nbitq), 
to_sfixed(-2010.0/65536.0,1,-nbitq), 
to_sfixed(437.0/65536.0,1,-nbitq), 
to_sfixed(-431.0/65536.0,1,-nbitq), 
to_sfixed(3700.0/65536.0,1,-nbitq), 
to_sfixed(3319.0/65536.0,1,-nbitq), 
to_sfixed(3392.0/65536.0,1,-nbitq), 
to_sfixed(209.0/65536.0,1,-nbitq), 
to_sfixed(-2468.0/65536.0,1,-nbitq), 
to_sfixed(-1822.0/65536.0,1,-nbitq), 
to_sfixed(3099.0/65536.0,1,-nbitq), 
to_sfixed(2837.0/65536.0,1,-nbitq), 
to_sfixed(2023.0/65536.0,1,-nbitq), 
to_sfixed(327.0/65536.0,1,-nbitq), 
to_sfixed(3371.0/65536.0,1,-nbitq), 
to_sfixed(-1961.0/65536.0,1,-nbitq), 
to_sfixed(-1059.0/65536.0,1,-nbitq), 
to_sfixed(-2728.0/65536.0,1,-nbitq), 
to_sfixed(1495.0/65536.0,1,-nbitq), 
to_sfixed(369.0/65536.0,1,-nbitq), 
to_sfixed(-70.0/65536.0,1,-nbitq), 
to_sfixed(-593.0/65536.0,1,-nbitq), 
to_sfixed(-1034.0/65536.0,1,-nbitq), 
to_sfixed(-2709.0/65536.0,1,-nbitq), 
to_sfixed(2495.0/65536.0,1,-nbitq), 
to_sfixed(-2137.0/65536.0,1,-nbitq), 
to_sfixed(-67.0/65536.0,1,-nbitq), 
to_sfixed(1745.0/65536.0,1,-nbitq), 
to_sfixed(-609.0/65536.0,1,-nbitq), 
to_sfixed(375.0/65536.0,1,-nbitq), 
to_sfixed(3873.0/65536.0,1,-nbitq), 
to_sfixed(-575.0/65536.0,1,-nbitq), 
to_sfixed(-48.0/65536.0,1,-nbitq), 
to_sfixed(4327.0/65536.0,1,-nbitq), 
to_sfixed(-1755.0/65536.0,1,-nbitq), 
to_sfixed(2130.0/65536.0,1,-nbitq), 
to_sfixed(-2771.0/65536.0,1,-nbitq), 
to_sfixed(-3681.0/65536.0,1,-nbitq), 
to_sfixed(1856.0/65536.0,1,-nbitq), 
to_sfixed(-208.0/65536.0,1,-nbitq), 
to_sfixed(1742.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2216.0/65536.0,1,-nbitq), 
to_sfixed(-2573.0/65536.0,1,-nbitq), 
to_sfixed(-2430.0/65536.0,1,-nbitq), 
to_sfixed(2604.0/65536.0,1,-nbitq), 
to_sfixed(7378.0/65536.0,1,-nbitq), 
to_sfixed(-4605.0/65536.0,1,-nbitq), 
to_sfixed(-2599.0/65536.0,1,-nbitq), 
to_sfixed(-2747.0/65536.0,1,-nbitq), 
to_sfixed(3149.0/65536.0,1,-nbitq), 
to_sfixed(3055.0/65536.0,1,-nbitq), 
to_sfixed(41.0/65536.0,1,-nbitq), 
to_sfixed(-1321.0/65536.0,1,-nbitq), 
to_sfixed(508.0/65536.0,1,-nbitq), 
to_sfixed(3430.0/65536.0,1,-nbitq), 
to_sfixed(892.0/65536.0,1,-nbitq), 
to_sfixed(-2594.0/65536.0,1,-nbitq), 
to_sfixed(-1156.0/65536.0,1,-nbitq), 
to_sfixed(1084.0/65536.0,1,-nbitq), 
to_sfixed(-2418.0/65536.0,1,-nbitq), 
to_sfixed(-526.0/65536.0,1,-nbitq), 
to_sfixed(3656.0/65536.0,1,-nbitq), 
to_sfixed(-3026.0/65536.0,1,-nbitq), 
to_sfixed(-3607.0/65536.0,1,-nbitq), 
to_sfixed(-2091.0/65536.0,1,-nbitq), 
to_sfixed(886.0/65536.0,1,-nbitq), 
to_sfixed(-966.0/65536.0,1,-nbitq), 
to_sfixed(670.0/65536.0,1,-nbitq), 
to_sfixed(-489.0/65536.0,1,-nbitq), 
to_sfixed(4118.0/65536.0,1,-nbitq), 
to_sfixed(-5163.0/65536.0,1,-nbitq), 
to_sfixed(805.0/65536.0,1,-nbitq), 
to_sfixed(-4423.0/65536.0,1,-nbitq), 
to_sfixed(1811.0/65536.0,1,-nbitq), 
to_sfixed(1209.0/65536.0,1,-nbitq), 
to_sfixed(-657.0/65536.0,1,-nbitq), 
to_sfixed(-1995.0/65536.0,1,-nbitq), 
to_sfixed(-5560.0/65536.0,1,-nbitq), 
to_sfixed(986.0/65536.0,1,-nbitq), 
to_sfixed(-5672.0/65536.0,1,-nbitq), 
to_sfixed(3099.0/65536.0,1,-nbitq), 
to_sfixed(1904.0/65536.0,1,-nbitq), 
to_sfixed(1418.0/65536.0,1,-nbitq), 
to_sfixed(-741.0/65536.0,1,-nbitq), 
to_sfixed(769.0/65536.0,1,-nbitq), 
to_sfixed(2617.0/65536.0,1,-nbitq), 
to_sfixed(3351.0/65536.0,1,-nbitq), 
to_sfixed(-2401.0/65536.0,1,-nbitq), 
to_sfixed(-2144.0/65536.0,1,-nbitq), 
to_sfixed(-102.0/65536.0,1,-nbitq), 
to_sfixed(2250.0/65536.0,1,-nbitq), 
to_sfixed(901.0/65536.0,1,-nbitq), 
to_sfixed(702.0/65536.0,1,-nbitq), 
to_sfixed(-3520.0/65536.0,1,-nbitq), 
to_sfixed(-234.0/65536.0,1,-nbitq), 
to_sfixed(2502.0/65536.0,1,-nbitq), 
to_sfixed(145.0/65536.0,1,-nbitq), 
to_sfixed(201.0/65536.0,1,-nbitq), 
to_sfixed(161.0/65536.0,1,-nbitq), 
to_sfixed(2653.0/65536.0,1,-nbitq), 
to_sfixed(-1158.0/65536.0,1,-nbitq), 
to_sfixed(-2743.0/65536.0,1,-nbitq), 
to_sfixed(1702.0/65536.0,1,-nbitq), 
to_sfixed(1928.0/65536.0,1,-nbitq), 
to_sfixed(-763.0/65536.0,1,-nbitq), 
to_sfixed(-2453.0/65536.0,1,-nbitq), 
to_sfixed(2324.0/65536.0,1,-nbitq), 
to_sfixed(757.0/65536.0,1,-nbitq), 
to_sfixed(874.0/65536.0,1,-nbitq), 
to_sfixed(7414.0/65536.0,1,-nbitq), 
to_sfixed(4726.0/65536.0,1,-nbitq), 
to_sfixed(2222.0/65536.0,1,-nbitq), 
to_sfixed(-1157.0/65536.0,1,-nbitq), 
to_sfixed(1207.0/65536.0,1,-nbitq), 
to_sfixed(-1605.0/65536.0,1,-nbitq), 
to_sfixed(-2698.0/65536.0,1,-nbitq), 
to_sfixed(634.0/65536.0,1,-nbitq), 
to_sfixed(-7838.0/65536.0,1,-nbitq), 
to_sfixed(2914.0/65536.0,1,-nbitq), 
to_sfixed(368.0/65536.0,1,-nbitq), 
to_sfixed(1941.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1731.0/65536.0,1,-nbitq), 
to_sfixed(1504.0/65536.0,1,-nbitq), 
to_sfixed(2011.0/65536.0,1,-nbitq), 
to_sfixed(-2320.0/65536.0,1,-nbitq), 
to_sfixed(3549.0/65536.0,1,-nbitq), 
to_sfixed(-2439.0/65536.0,1,-nbitq), 
to_sfixed(1672.0/65536.0,1,-nbitq), 
to_sfixed(-5774.0/65536.0,1,-nbitq), 
to_sfixed(-3694.0/65536.0,1,-nbitq), 
to_sfixed(984.0/65536.0,1,-nbitq), 
to_sfixed(-1346.0/65536.0,1,-nbitq), 
to_sfixed(1525.0/65536.0,1,-nbitq), 
to_sfixed(2868.0/65536.0,1,-nbitq), 
to_sfixed(-2137.0/65536.0,1,-nbitq), 
to_sfixed(2822.0/65536.0,1,-nbitq), 
to_sfixed(-1373.0/65536.0,1,-nbitq), 
to_sfixed(451.0/65536.0,1,-nbitq), 
to_sfixed(-3951.0/65536.0,1,-nbitq), 
to_sfixed(-2095.0/65536.0,1,-nbitq), 
to_sfixed(2945.0/65536.0,1,-nbitq), 
to_sfixed(5028.0/65536.0,1,-nbitq), 
to_sfixed(-253.0/65536.0,1,-nbitq), 
to_sfixed(-3733.0/65536.0,1,-nbitq), 
to_sfixed(-4810.0/65536.0,1,-nbitq), 
to_sfixed(-1119.0/65536.0,1,-nbitq), 
to_sfixed(-8332.0/65536.0,1,-nbitq), 
to_sfixed(2473.0/65536.0,1,-nbitq), 
to_sfixed(-1121.0/65536.0,1,-nbitq), 
to_sfixed(5624.0/65536.0,1,-nbitq), 
to_sfixed(-3284.0/65536.0,1,-nbitq), 
to_sfixed(3054.0/65536.0,1,-nbitq), 
to_sfixed(-258.0/65536.0,1,-nbitq), 
to_sfixed(1964.0/65536.0,1,-nbitq), 
to_sfixed(247.0/65536.0,1,-nbitq), 
to_sfixed(-376.0/65536.0,1,-nbitq), 
to_sfixed(2483.0/65536.0,1,-nbitq), 
to_sfixed(-4242.0/65536.0,1,-nbitq), 
to_sfixed(3323.0/65536.0,1,-nbitq), 
to_sfixed(-2168.0/65536.0,1,-nbitq), 
to_sfixed(-565.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(1203.0/65536.0,1,-nbitq), 
to_sfixed(8139.0/65536.0,1,-nbitq), 
to_sfixed(828.0/65536.0,1,-nbitq), 
to_sfixed(653.0/65536.0,1,-nbitq), 
to_sfixed(1033.0/65536.0,1,-nbitq), 
to_sfixed(-967.0/65536.0,1,-nbitq), 
to_sfixed(-2337.0/65536.0,1,-nbitq), 
to_sfixed(2363.0/65536.0,1,-nbitq), 
to_sfixed(1441.0/65536.0,1,-nbitq), 
to_sfixed(-36.0/65536.0,1,-nbitq), 
to_sfixed(478.0/65536.0,1,-nbitq), 
to_sfixed(-3319.0/65536.0,1,-nbitq), 
to_sfixed(-578.0/65536.0,1,-nbitq), 
to_sfixed(-2158.0/65536.0,1,-nbitq), 
to_sfixed(2165.0/65536.0,1,-nbitq), 
to_sfixed(-2639.0/65536.0,1,-nbitq), 
to_sfixed(4324.0/65536.0,1,-nbitq), 
to_sfixed(-395.0/65536.0,1,-nbitq), 
to_sfixed(-4241.0/65536.0,1,-nbitq), 
to_sfixed(-4231.0/65536.0,1,-nbitq), 
to_sfixed(2147.0/65536.0,1,-nbitq), 
to_sfixed(-1481.0/65536.0,1,-nbitq), 
to_sfixed(-1170.0/65536.0,1,-nbitq), 
to_sfixed(-5899.0/65536.0,1,-nbitq), 
to_sfixed(-4395.0/65536.0,1,-nbitq), 
to_sfixed(388.0/65536.0,1,-nbitq), 
to_sfixed(4117.0/65536.0,1,-nbitq), 
to_sfixed(6697.0/65536.0,1,-nbitq), 
to_sfixed(3338.0/65536.0,1,-nbitq), 
to_sfixed(-2363.0/65536.0,1,-nbitq), 
to_sfixed(-3595.0/65536.0,1,-nbitq), 
to_sfixed(4246.0/65536.0,1,-nbitq), 
to_sfixed(-87.0/65536.0,1,-nbitq), 
to_sfixed(-2565.0/65536.0,1,-nbitq), 
to_sfixed(-289.0/65536.0,1,-nbitq), 
to_sfixed(-4774.0/65536.0,1,-nbitq), 
to_sfixed(-394.0/65536.0,1,-nbitq), 
to_sfixed(2448.0/65536.0,1,-nbitq), 
to_sfixed(-1441.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2229.0/65536.0,1,-nbitq), 
to_sfixed(-3405.0/65536.0,1,-nbitq), 
to_sfixed(-7434.0/65536.0,1,-nbitq), 
to_sfixed(719.0/65536.0,1,-nbitq), 
to_sfixed(5700.0/65536.0,1,-nbitq), 
to_sfixed(-2556.0/65536.0,1,-nbitq), 
to_sfixed(-2730.0/65536.0,1,-nbitq), 
to_sfixed(-718.0/65536.0,1,-nbitq), 
to_sfixed(-2864.0/65536.0,1,-nbitq), 
to_sfixed(383.0/65536.0,1,-nbitq), 
to_sfixed(-1846.0/65536.0,1,-nbitq), 
to_sfixed(4064.0/65536.0,1,-nbitq), 
to_sfixed(1192.0/65536.0,1,-nbitq), 
to_sfixed(349.0/65536.0,1,-nbitq), 
to_sfixed(-588.0/65536.0,1,-nbitq), 
to_sfixed(-1548.0/65536.0,1,-nbitq), 
to_sfixed(-3286.0/65536.0,1,-nbitq), 
to_sfixed(-2306.0/65536.0,1,-nbitq), 
to_sfixed(-3760.0/65536.0,1,-nbitq), 
to_sfixed(-2501.0/65536.0,1,-nbitq), 
to_sfixed(2915.0/65536.0,1,-nbitq), 
to_sfixed(3180.0/65536.0,1,-nbitq), 
to_sfixed(3483.0/65536.0,1,-nbitq), 
to_sfixed(-15769.0/65536.0,1,-nbitq), 
to_sfixed(323.0/65536.0,1,-nbitq), 
to_sfixed(-17037.0/65536.0,1,-nbitq), 
to_sfixed(-2196.0/65536.0,1,-nbitq), 
to_sfixed(3042.0/65536.0,1,-nbitq), 
to_sfixed(11028.0/65536.0,1,-nbitq), 
to_sfixed(-2061.0/65536.0,1,-nbitq), 
to_sfixed(1624.0/65536.0,1,-nbitq), 
to_sfixed(-3495.0/65536.0,1,-nbitq), 
to_sfixed(3877.0/65536.0,1,-nbitq), 
to_sfixed(2800.0/65536.0,1,-nbitq), 
to_sfixed(-610.0/65536.0,1,-nbitq), 
to_sfixed(739.0/65536.0,1,-nbitq), 
to_sfixed(-5538.0/65536.0,1,-nbitq), 
to_sfixed(1263.0/65536.0,1,-nbitq), 
to_sfixed(188.0/65536.0,1,-nbitq), 
to_sfixed(-3130.0/65536.0,1,-nbitq), 
to_sfixed(3972.0/65536.0,1,-nbitq), 
to_sfixed(495.0/65536.0,1,-nbitq), 
to_sfixed(5131.0/65536.0,1,-nbitq), 
to_sfixed(-1811.0/65536.0,1,-nbitq), 
to_sfixed(582.0/65536.0,1,-nbitq), 
to_sfixed(-2164.0/65536.0,1,-nbitq), 
to_sfixed(1230.0/65536.0,1,-nbitq), 
to_sfixed(-4760.0/65536.0,1,-nbitq), 
to_sfixed(909.0/65536.0,1,-nbitq), 
to_sfixed(944.0/65536.0,1,-nbitq), 
to_sfixed(2354.0/65536.0,1,-nbitq), 
to_sfixed(-2099.0/65536.0,1,-nbitq), 
to_sfixed(-5074.0/65536.0,1,-nbitq), 
to_sfixed(1207.0/65536.0,1,-nbitq), 
to_sfixed(-4354.0/65536.0,1,-nbitq), 
to_sfixed(-1408.0/65536.0,1,-nbitq), 
to_sfixed(-692.0/65536.0,1,-nbitq), 
to_sfixed(3671.0/65536.0,1,-nbitq), 
to_sfixed(1196.0/65536.0,1,-nbitq), 
to_sfixed(-11148.0/65536.0,1,-nbitq), 
to_sfixed(-4338.0/65536.0,1,-nbitq), 
to_sfixed(-1909.0/65536.0,1,-nbitq), 
to_sfixed(1721.0/65536.0,1,-nbitq), 
to_sfixed(-1377.0/65536.0,1,-nbitq), 
to_sfixed(-8033.0/65536.0,1,-nbitq), 
to_sfixed(-1959.0/65536.0,1,-nbitq), 
to_sfixed(-913.0/65536.0,1,-nbitq), 
to_sfixed(3250.0/65536.0,1,-nbitq), 
to_sfixed(9343.0/65536.0,1,-nbitq), 
to_sfixed(951.0/65536.0,1,-nbitq), 
to_sfixed(1215.0/65536.0,1,-nbitq), 
to_sfixed(-2037.0/65536.0,1,-nbitq), 
to_sfixed(-2046.0/65536.0,1,-nbitq), 
to_sfixed(-2154.0/65536.0,1,-nbitq), 
to_sfixed(2368.0/65536.0,1,-nbitq), 
to_sfixed(591.0/65536.0,1,-nbitq), 
to_sfixed(-650.0/65536.0,1,-nbitq), 
to_sfixed(80.0/65536.0,1,-nbitq), 
to_sfixed(997.0/65536.0,1,-nbitq), 
to_sfixed(-2591.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2996.0/65536.0,1,-nbitq), 
to_sfixed(-845.0/65536.0,1,-nbitq), 
to_sfixed(-6465.0/65536.0,1,-nbitq), 
to_sfixed(-67.0/65536.0,1,-nbitq), 
to_sfixed(-4339.0/65536.0,1,-nbitq), 
to_sfixed(4214.0/65536.0,1,-nbitq), 
to_sfixed(-3488.0/65536.0,1,-nbitq), 
to_sfixed(3469.0/65536.0,1,-nbitq), 
to_sfixed(-1044.0/65536.0,1,-nbitq), 
to_sfixed(-643.0/65536.0,1,-nbitq), 
to_sfixed(-1999.0/65536.0,1,-nbitq), 
to_sfixed(-3436.0/65536.0,1,-nbitq), 
to_sfixed(1784.0/65536.0,1,-nbitq), 
to_sfixed(5725.0/65536.0,1,-nbitq), 
to_sfixed(702.0/65536.0,1,-nbitq), 
to_sfixed(-843.0/65536.0,1,-nbitq), 
to_sfixed(1198.0/65536.0,1,-nbitq), 
to_sfixed(4429.0/65536.0,1,-nbitq), 
to_sfixed(1251.0/65536.0,1,-nbitq), 
to_sfixed(-2099.0/65536.0,1,-nbitq), 
to_sfixed(3163.0/65536.0,1,-nbitq), 
to_sfixed(-410.0/65536.0,1,-nbitq), 
to_sfixed(4265.0/65536.0,1,-nbitq), 
to_sfixed(-12142.0/65536.0,1,-nbitq), 
to_sfixed(4711.0/65536.0,1,-nbitq), 
to_sfixed(-16220.0/65536.0,1,-nbitq), 
to_sfixed(-1874.0/65536.0,1,-nbitq), 
to_sfixed(1088.0/65536.0,1,-nbitq), 
to_sfixed(1633.0/65536.0,1,-nbitq), 
to_sfixed(2093.0/65536.0,1,-nbitq), 
to_sfixed(3174.0/65536.0,1,-nbitq), 
to_sfixed(-3054.0/65536.0,1,-nbitq), 
to_sfixed(4713.0/65536.0,1,-nbitq), 
to_sfixed(-3048.0/65536.0,1,-nbitq), 
to_sfixed(2443.0/65536.0,1,-nbitq), 
to_sfixed(1131.0/65536.0,1,-nbitq), 
to_sfixed(-5048.0/65536.0,1,-nbitq), 
to_sfixed(-170.0/65536.0,1,-nbitq), 
to_sfixed(4263.0/65536.0,1,-nbitq), 
to_sfixed(-7349.0/65536.0,1,-nbitq), 
to_sfixed(7220.0/65536.0,1,-nbitq), 
to_sfixed(-1089.0/65536.0,1,-nbitq), 
to_sfixed(4946.0/65536.0,1,-nbitq), 
to_sfixed(2416.0/65536.0,1,-nbitq), 
to_sfixed(700.0/65536.0,1,-nbitq), 
to_sfixed(930.0/65536.0,1,-nbitq), 
to_sfixed(2241.0/65536.0,1,-nbitq), 
to_sfixed(-10588.0/65536.0,1,-nbitq), 
to_sfixed(1651.0/65536.0,1,-nbitq), 
to_sfixed(2746.0/65536.0,1,-nbitq), 
to_sfixed(1400.0/65536.0,1,-nbitq), 
to_sfixed(1778.0/65536.0,1,-nbitq), 
to_sfixed(-3700.0/65536.0,1,-nbitq), 
to_sfixed(6116.0/65536.0,1,-nbitq), 
to_sfixed(-4298.0/65536.0,1,-nbitq), 
to_sfixed(-4297.0/65536.0,1,-nbitq), 
to_sfixed(1708.0/65536.0,1,-nbitq), 
to_sfixed(86.0/65536.0,1,-nbitq), 
to_sfixed(-1220.0/65536.0,1,-nbitq), 
to_sfixed(-11578.0/65536.0,1,-nbitq), 
to_sfixed(-1237.0/65536.0,1,-nbitq), 
to_sfixed(-3026.0/65536.0,1,-nbitq), 
to_sfixed(2586.0/65536.0,1,-nbitq), 
to_sfixed(421.0/65536.0,1,-nbitq), 
to_sfixed(-5930.0/65536.0,1,-nbitq), 
to_sfixed(5103.0/65536.0,1,-nbitq), 
to_sfixed(2419.0/65536.0,1,-nbitq), 
to_sfixed(401.0/65536.0,1,-nbitq), 
to_sfixed(4427.0/65536.0,1,-nbitq), 
to_sfixed(-3057.0/65536.0,1,-nbitq), 
to_sfixed(-2786.0/65536.0,1,-nbitq), 
to_sfixed(-1260.0/65536.0,1,-nbitq), 
to_sfixed(-2547.0/65536.0,1,-nbitq), 
to_sfixed(-788.0/65536.0,1,-nbitq), 
to_sfixed(-1652.0/65536.0,1,-nbitq), 
to_sfixed(-1697.0/65536.0,1,-nbitq), 
to_sfixed(1306.0/65536.0,1,-nbitq), 
to_sfixed(-1374.0/65536.0,1,-nbitq), 
to_sfixed(-1289.0/65536.0,1,-nbitq), 
to_sfixed(-6481.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3552.0/65536.0,1,-nbitq), 
to_sfixed(-747.0/65536.0,1,-nbitq), 
to_sfixed(-1803.0/65536.0,1,-nbitq), 
to_sfixed(-2856.0/65536.0,1,-nbitq), 
to_sfixed(-265.0/65536.0,1,-nbitq), 
to_sfixed(4927.0/65536.0,1,-nbitq), 
to_sfixed(-6978.0/65536.0,1,-nbitq), 
to_sfixed(6602.0/65536.0,1,-nbitq), 
to_sfixed(-3655.0/65536.0,1,-nbitq), 
to_sfixed(2793.0/65536.0,1,-nbitq), 
to_sfixed(-5389.0/65536.0,1,-nbitq), 
to_sfixed(-6764.0/65536.0,1,-nbitq), 
to_sfixed(1760.0/65536.0,1,-nbitq), 
to_sfixed(4668.0/65536.0,1,-nbitq), 
to_sfixed(436.0/65536.0,1,-nbitq), 
to_sfixed(1471.0/65536.0,1,-nbitq), 
to_sfixed(-712.0/65536.0,1,-nbitq), 
to_sfixed(7888.0/65536.0,1,-nbitq), 
to_sfixed(1476.0/65536.0,1,-nbitq), 
to_sfixed(1780.0/65536.0,1,-nbitq), 
to_sfixed(3089.0/65536.0,1,-nbitq), 
to_sfixed(-7426.0/65536.0,1,-nbitq), 
to_sfixed(-2655.0/65536.0,1,-nbitq), 
to_sfixed(-11648.0/65536.0,1,-nbitq), 
to_sfixed(558.0/65536.0,1,-nbitq), 
to_sfixed(-14954.0/65536.0,1,-nbitq), 
to_sfixed(2731.0/65536.0,1,-nbitq), 
to_sfixed(45.0/65536.0,1,-nbitq), 
to_sfixed(2761.0/65536.0,1,-nbitq), 
to_sfixed(5113.0/65536.0,1,-nbitq), 
to_sfixed(2653.0/65536.0,1,-nbitq), 
to_sfixed(44.0/65536.0,1,-nbitq), 
to_sfixed(2405.0/65536.0,1,-nbitq), 
to_sfixed(1538.0/65536.0,1,-nbitq), 
to_sfixed(1763.0/65536.0,1,-nbitq), 
to_sfixed(618.0/65536.0,1,-nbitq), 
to_sfixed(-6867.0/65536.0,1,-nbitq), 
to_sfixed(330.0/65536.0,1,-nbitq), 
to_sfixed(3076.0/65536.0,1,-nbitq), 
to_sfixed(-1819.0/65536.0,1,-nbitq), 
to_sfixed(5242.0/65536.0,1,-nbitq), 
to_sfixed(-3053.0/65536.0,1,-nbitq), 
to_sfixed(4065.0/65536.0,1,-nbitq), 
to_sfixed(4316.0/65536.0,1,-nbitq), 
to_sfixed(1205.0/65536.0,1,-nbitq), 
to_sfixed(-3083.0/65536.0,1,-nbitq), 
to_sfixed(2381.0/65536.0,1,-nbitq), 
to_sfixed(-11423.0/65536.0,1,-nbitq), 
to_sfixed(1810.0/65536.0,1,-nbitq), 
to_sfixed(3015.0/65536.0,1,-nbitq), 
to_sfixed(1034.0/65536.0,1,-nbitq), 
to_sfixed(-2898.0/65536.0,1,-nbitq), 
to_sfixed(-5784.0/65536.0,1,-nbitq), 
to_sfixed(1643.0/65536.0,1,-nbitq), 
to_sfixed(-2874.0/65536.0,1,-nbitq), 
to_sfixed(-2442.0/65536.0,1,-nbitq), 
to_sfixed(2512.0/65536.0,1,-nbitq), 
to_sfixed(-1181.0/65536.0,1,-nbitq), 
to_sfixed(-2659.0/65536.0,1,-nbitq), 
to_sfixed(-8572.0/65536.0,1,-nbitq), 
to_sfixed(9854.0/65536.0,1,-nbitq), 
to_sfixed(-2757.0/65536.0,1,-nbitq), 
to_sfixed(2449.0/65536.0,1,-nbitq), 
to_sfixed(-2600.0/65536.0,1,-nbitq), 
to_sfixed(-7147.0/65536.0,1,-nbitq), 
to_sfixed(5008.0/65536.0,1,-nbitq), 
to_sfixed(-869.0/65536.0,1,-nbitq), 
to_sfixed(3648.0/65536.0,1,-nbitq), 
to_sfixed(8511.0/65536.0,1,-nbitq), 
to_sfixed(-3214.0/65536.0,1,-nbitq), 
to_sfixed(-875.0/65536.0,1,-nbitq), 
to_sfixed(2427.0/65536.0,1,-nbitq), 
to_sfixed(-1559.0/65536.0,1,-nbitq), 
to_sfixed(589.0/65536.0,1,-nbitq), 
to_sfixed(2708.0/65536.0,1,-nbitq), 
to_sfixed(-935.0/65536.0,1,-nbitq), 
to_sfixed(4862.0/65536.0,1,-nbitq), 
to_sfixed(-3532.0/65536.0,1,-nbitq), 
to_sfixed(2606.0/65536.0,1,-nbitq), 
to_sfixed(-3821.0/65536.0,1,-nbitq)  ), 
( to_sfixed(602.0/65536.0,1,-nbitq), 
to_sfixed(-4297.0/65536.0,1,-nbitq), 
to_sfixed(3055.0/65536.0,1,-nbitq), 
to_sfixed(-3771.0/65536.0,1,-nbitq), 
to_sfixed(1209.0/65536.0,1,-nbitq), 
to_sfixed(2398.0/65536.0,1,-nbitq), 
to_sfixed(-12417.0/65536.0,1,-nbitq), 
to_sfixed(4487.0/65536.0,1,-nbitq), 
to_sfixed(-2833.0/65536.0,1,-nbitq), 
to_sfixed(-682.0/65536.0,1,-nbitq), 
to_sfixed(-1744.0/65536.0,1,-nbitq), 
to_sfixed(-3838.0/65536.0,1,-nbitq), 
to_sfixed(2443.0/65536.0,1,-nbitq), 
to_sfixed(-3307.0/65536.0,1,-nbitq), 
to_sfixed(3968.0/65536.0,1,-nbitq), 
to_sfixed(3176.0/65536.0,1,-nbitq), 
to_sfixed(-2094.0/65536.0,1,-nbitq), 
to_sfixed(9956.0/65536.0,1,-nbitq), 
to_sfixed(8376.0/65536.0,1,-nbitq), 
to_sfixed(-2461.0/65536.0,1,-nbitq), 
to_sfixed(4982.0/65536.0,1,-nbitq), 
to_sfixed(-3268.0/65536.0,1,-nbitq), 
to_sfixed(1997.0/65536.0,1,-nbitq), 
to_sfixed(-4586.0/65536.0,1,-nbitq), 
to_sfixed(-813.0/65536.0,1,-nbitq), 
to_sfixed(-8179.0/65536.0,1,-nbitq), 
to_sfixed(-3819.0/65536.0,1,-nbitq), 
to_sfixed(-689.0/65536.0,1,-nbitq), 
to_sfixed(-2902.0/65536.0,1,-nbitq), 
to_sfixed(6440.0/65536.0,1,-nbitq), 
to_sfixed(-381.0/65536.0,1,-nbitq), 
to_sfixed(552.0/65536.0,1,-nbitq), 
to_sfixed(8172.0/65536.0,1,-nbitq), 
to_sfixed(6552.0/65536.0,1,-nbitq), 
to_sfixed(-391.0/65536.0,1,-nbitq), 
to_sfixed(2152.0/65536.0,1,-nbitq), 
to_sfixed(-8957.0/65536.0,1,-nbitq), 
to_sfixed(604.0/65536.0,1,-nbitq), 
to_sfixed(-399.0/65536.0,1,-nbitq), 
to_sfixed(5118.0/65536.0,1,-nbitq), 
to_sfixed(120.0/65536.0,1,-nbitq), 
to_sfixed(1033.0/65536.0,1,-nbitq), 
to_sfixed(4421.0/65536.0,1,-nbitq), 
to_sfixed(-1908.0/65536.0,1,-nbitq), 
to_sfixed(-2030.0/65536.0,1,-nbitq), 
to_sfixed(-4800.0/65536.0,1,-nbitq), 
to_sfixed(-929.0/65536.0,1,-nbitq), 
to_sfixed(-11701.0/65536.0,1,-nbitq), 
to_sfixed(-1635.0/65536.0,1,-nbitq), 
to_sfixed(4285.0/65536.0,1,-nbitq), 
to_sfixed(-753.0/65536.0,1,-nbitq), 
to_sfixed(-6472.0/65536.0,1,-nbitq), 
to_sfixed(-4946.0/65536.0,1,-nbitq), 
to_sfixed(-11224.0/65536.0,1,-nbitq), 
to_sfixed(-3762.0/65536.0,1,-nbitq), 
to_sfixed(-6142.0/65536.0,1,-nbitq), 
to_sfixed(-461.0/65536.0,1,-nbitq), 
to_sfixed(2571.0/65536.0,1,-nbitq), 
to_sfixed(830.0/65536.0,1,-nbitq), 
to_sfixed(4251.0/65536.0,1,-nbitq), 
to_sfixed(16269.0/65536.0,1,-nbitq), 
to_sfixed(-1930.0/65536.0,1,-nbitq), 
to_sfixed(672.0/65536.0,1,-nbitq), 
to_sfixed(-615.0/65536.0,1,-nbitq), 
to_sfixed(-5159.0/65536.0,1,-nbitq), 
to_sfixed(1411.0/65536.0,1,-nbitq), 
to_sfixed(3863.0/65536.0,1,-nbitq), 
to_sfixed(-2837.0/65536.0,1,-nbitq), 
to_sfixed(2310.0/65536.0,1,-nbitq), 
to_sfixed(-3100.0/65536.0,1,-nbitq), 
to_sfixed(-2097.0/65536.0,1,-nbitq), 
to_sfixed(1932.0/65536.0,1,-nbitq), 
to_sfixed(-1268.0/65536.0,1,-nbitq), 
to_sfixed(2378.0/65536.0,1,-nbitq), 
to_sfixed(-260.0/65536.0,1,-nbitq), 
to_sfixed(2822.0/65536.0,1,-nbitq), 
to_sfixed(11419.0/65536.0,1,-nbitq), 
to_sfixed(-6635.0/65536.0,1,-nbitq), 
to_sfixed(-1901.0/65536.0,1,-nbitq), 
to_sfixed(-4917.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4837.0/65536.0,1,-nbitq), 
to_sfixed(2683.0/65536.0,1,-nbitq), 
to_sfixed(-3387.0/65536.0,1,-nbitq), 
to_sfixed(-2079.0/65536.0,1,-nbitq), 
to_sfixed(-8011.0/65536.0,1,-nbitq), 
to_sfixed(879.0/65536.0,1,-nbitq), 
to_sfixed(-10336.0/65536.0,1,-nbitq), 
to_sfixed(6625.0/65536.0,1,-nbitq), 
to_sfixed(1352.0/65536.0,1,-nbitq), 
to_sfixed(-1198.0/65536.0,1,-nbitq), 
to_sfixed(-407.0/65536.0,1,-nbitq), 
to_sfixed(-3796.0/65536.0,1,-nbitq), 
to_sfixed(4578.0/65536.0,1,-nbitq), 
to_sfixed(-4517.0/65536.0,1,-nbitq), 
to_sfixed(2296.0/65536.0,1,-nbitq), 
to_sfixed(-1863.0/65536.0,1,-nbitq), 
to_sfixed(694.0/65536.0,1,-nbitq), 
to_sfixed(11679.0/65536.0,1,-nbitq), 
to_sfixed(7345.0/65536.0,1,-nbitq), 
to_sfixed(814.0/65536.0,1,-nbitq), 
to_sfixed(1882.0/65536.0,1,-nbitq), 
to_sfixed(4457.0/65536.0,1,-nbitq), 
to_sfixed(-1809.0/65536.0,1,-nbitq), 
to_sfixed(-6175.0/65536.0,1,-nbitq), 
to_sfixed(-1648.0/65536.0,1,-nbitq), 
to_sfixed(-9721.0/65536.0,1,-nbitq), 
to_sfixed(-5430.0/65536.0,1,-nbitq), 
to_sfixed(4776.0/65536.0,1,-nbitq), 
to_sfixed(-6489.0/65536.0,1,-nbitq), 
to_sfixed(6016.0/65536.0,1,-nbitq), 
to_sfixed(-4782.0/65536.0,1,-nbitq), 
to_sfixed(-3605.0/65536.0,1,-nbitq), 
to_sfixed(2861.0/65536.0,1,-nbitq), 
to_sfixed(6948.0/65536.0,1,-nbitq), 
to_sfixed(243.0/65536.0,1,-nbitq), 
to_sfixed(2529.0/65536.0,1,-nbitq), 
to_sfixed(-14199.0/65536.0,1,-nbitq), 
to_sfixed(3860.0/65536.0,1,-nbitq), 
to_sfixed(1677.0/65536.0,1,-nbitq), 
to_sfixed(2107.0/65536.0,1,-nbitq), 
to_sfixed(549.0/65536.0,1,-nbitq), 
to_sfixed(-3091.0/65536.0,1,-nbitq), 
to_sfixed(842.0/65536.0,1,-nbitq), 
to_sfixed(-3829.0/65536.0,1,-nbitq), 
to_sfixed(-353.0/65536.0,1,-nbitq), 
to_sfixed(-6431.0/65536.0,1,-nbitq), 
to_sfixed(-2343.0/65536.0,1,-nbitq), 
to_sfixed(-4821.0/65536.0,1,-nbitq), 
to_sfixed(-1596.0/65536.0,1,-nbitq), 
to_sfixed(-1541.0/65536.0,1,-nbitq), 
to_sfixed(1216.0/65536.0,1,-nbitq), 
to_sfixed(-34.0/65536.0,1,-nbitq), 
to_sfixed(-6513.0/65536.0,1,-nbitq), 
to_sfixed(-14901.0/65536.0,1,-nbitq), 
to_sfixed(-1814.0/65536.0,1,-nbitq), 
to_sfixed(-2298.0/65536.0,1,-nbitq), 
to_sfixed(3117.0/65536.0,1,-nbitq), 
to_sfixed(4300.0/65536.0,1,-nbitq), 
to_sfixed(2618.0/65536.0,1,-nbitq), 
to_sfixed(5434.0/65536.0,1,-nbitq), 
to_sfixed(13332.0/65536.0,1,-nbitq), 
to_sfixed(1108.0/65536.0,1,-nbitq), 
to_sfixed(2134.0/65536.0,1,-nbitq), 
to_sfixed(400.0/65536.0,1,-nbitq), 
to_sfixed(-5508.0/65536.0,1,-nbitq), 
to_sfixed(1212.0/65536.0,1,-nbitq), 
to_sfixed(1923.0/65536.0,1,-nbitq), 
to_sfixed(3141.0/65536.0,1,-nbitq), 
to_sfixed(4166.0/65536.0,1,-nbitq), 
to_sfixed(3763.0/65536.0,1,-nbitq), 
to_sfixed(-824.0/65536.0,1,-nbitq), 
to_sfixed(1213.0/65536.0,1,-nbitq), 
to_sfixed(-3759.0/65536.0,1,-nbitq), 
to_sfixed(-1106.0/65536.0,1,-nbitq), 
to_sfixed(-1469.0/65536.0,1,-nbitq), 
to_sfixed(4960.0/65536.0,1,-nbitq), 
to_sfixed(6193.0/65536.0,1,-nbitq), 
to_sfixed(-2364.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(-7434.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3836.0/65536.0,1,-nbitq), 
to_sfixed(5985.0/65536.0,1,-nbitq), 
to_sfixed(-8442.0/65536.0,1,-nbitq), 
to_sfixed(-2353.0/65536.0,1,-nbitq), 
to_sfixed(-4705.0/65536.0,1,-nbitq), 
to_sfixed(1405.0/65536.0,1,-nbitq), 
to_sfixed(-6118.0/65536.0,1,-nbitq), 
to_sfixed(-5737.0/65536.0,1,-nbitq), 
to_sfixed(1980.0/65536.0,1,-nbitq), 
to_sfixed(-962.0/65536.0,1,-nbitq), 
to_sfixed(-5513.0/65536.0,1,-nbitq), 
to_sfixed(-4059.0/65536.0,1,-nbitq), 
to_sfixed(-758.0/65536.0,1,-nbitq), 
to_sfixed(-5303.0/65536.0,1,-nbitq), 
to_sfixed(1433.0/65536.0,1,-nbitq), 
to_sfixed(-2204.0/65536.0,1,-nbitq), 
to_sfixed(-1213.0/65536.0,1,-nbitq), 
to_sfixed(174.0/65536.0,1,-nbitq), 
to_sfixed(4904.0/65536.0,1,-nbitq), 
to_sfixed(-2399.0/65536.0,1,-nbitq), 
to_sfixed(3310.0/65536.0,1,-nbitq), 
to_sfixed(8893.0/65536.0,1,-nbitq), 
to_sfixed(-3776.0/65536.0,1,-nbitq), 
to_sfixed(-3125.0/65536.0,1,-nbitq), 
to_sfixed(-3075.0/65536.0,1,-nbitq), 
to_sfixed(-4429.0/65536.0,1,-nbitq), 
to_sfixed(1009.0/65536.0,1,-nbitq), 
to_sfixed(2765.0/65536.0,1,-nbitq), 
to_sfixed(-4883.0/65536.0,1,-nbitq), 
to_sfixed(4393.0/65536.0,1,-nbitq), 
to_sfixed(-2634.0/65536.0,1,-nbitq), 
to_sfixed(-4547.0/65536.0,1,-nbitq), 
to_sfixed(3091.0/65536.0,1,-nbitq), 
to_sfixed(-9067.0/65536.0,1,-nbitq), 
to_sfixed(-1753.0/65536.0,1,-nbitq), 
to_sfixed(1324.0/65536.0,1,-nbitq), 
to_sfixed(-18211.0/65536.0,1,-nbitq), 
to_sfixed(1276.0/65536.0,1,-nbitq), 
to_sfixed(1535.0/65536.0,1,-nbitq), 
to_sfixed(191.0/65536.0,1,-nbitq), 
to_sfixed(-2412.0/65536.0,1,-nbitq), 
to_sfixed(1925.0/65536.0,1,-nbitq), 
to_sfixed(-12928.0/65536.0,1,-nbitq), 
to_sfixed(-3886.0/65536.0,1,-nbitq), 
to_sfixed(-2054.0/65536.0,1,-nbitq), 
to_sfixed(-755.0/65536.0,1,-nbitq), 
to_sfixed(-68.0/65536.0,1,-nbitq), 
to_sfixed(168.0/65536.0,1,-nbitq), 
to_sfixed(2367.0/65536.0,1,-nbitq), 
to_sfixed(1553.0/65536.0,1,-nbitq), 
to_sfixed(-1595.0/65536.0,1,-nbitq), 
to_sfixed(-2723.0/65536.0,1,-nbitq), 
to_sfixed(-3031.0/65536.0,1,-nbitq), 
to_sfixed(-17.0/65536.0,1,-nbitq), 
to_sfixed(73.0/65536.0,1,-nbitq), 
to_sfixed(-3865.0/65536.0,1,-nbitq), 
to_sfixed(2750.0/65536.0,1,-nbitq), 
to_sfixed(1224.0/65536.0,1,-nbitq), 
to_sfixed(-2973.0/65536.0,1,-nbitq), 
to_sfixed(5608.0/65536.0,1,-nbitq), 
to_sfixed(1905.0/65536.0,1,-nbitq), 
to_sfixed(-1292.0/65536.0,1,-nbitq), 
to_sfixed(471.0/65536.0,1,-nbitq), 
to_sfixed(891.0/65536.0,1,-nbitq), 
to_sfixed(-4732.0/65536.0,1,-nbitq), 
to_sfixed(23563.0/65536.0,1,-nbitq), 
to_sfixed(1463.0/65536.0,1,-nbitq), 
to_sfixed(1062.0/65536.0,1,-nbitq), 
to_sfixed(138.0/65536.0,1,-nbitq), 
to_sfixed(-2825.0/65536.0,1,-nbitq), 
to_sfixed(-3529.0/65536.0,1,-nbitq), 
to_sfixed(1015.0/65536.0,1,-nbitq), 
to_sfixed(-8694.0/65536.0,1,-nbitq), 
to_sfixed(86.0/65536.0,1,-nbitq), 
to_sfixed(-2786.0/65536.0,1,-nbitq), 
to_sfixed(2931.0/65536.0,1,-nbitq), 
to_sfixed(3591.0/65536.0,1,-nbitq), 
to_sfixed(2803.0/65536.0,1,-nbitq), 
to_sfixed(-2431.0/65536.0,1,-nbitq), 
to_sfixed(-11619.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-7097.0/65536.0,1,-nbitq), 
to_sfixed(7858.0/65536.0,1,-nbitq), 
to_sfixed(-11306.0/65536.0,1,-nbitq), 
to_sfixed(-984.0/65536.0,1,-nbitq), 
to_sfixed(-1308.0/65536.0,1,-nbitq), 
to_sfixed(1967.0/65536.0,1,-nbitq), 
to_sfixed(-125.0/65536.0,1,-nbitq), 
to_sfixed(-9920.0/65536.0,1,-nbitq), 
to_sfixed(-19.0/65536.0,1,-nbitq), 
to_sfixed(-930.0/65536.0,1,-nbitq), 
to_sfixed(-5291.0/65536.0,1,-nbitq), 
to_sfixed(-9107.0/65536.0,1,-nbitq), 
to_sfixed(3221.0/65536.0,1,-nbitq), 
to_sfixed(1879.0/65536.0,1,-nbitq), 
to_sfixed(1349.0/65536.0,1,-nbitq), 
to_sfixed(2232.0/65536.0,1,-nbitq), 
to_sfixed(2251.0/65536.0,1,-nbitq), 
to_sfixed(-16640.0/65536.0,1,-nbitq), 
to_sfixed(1113.0/65536.0,1,-nbitq), 
to_sfixed(2205.0/65536.0,1,-nbitq), 
to_sfixed(-376.0/65536.0,1,-nbitq), 
to_sfixed(3020.0/65536.0,1,-nbitq), 
to_sfixed(-5031.0/65536.0,1,-nbitq), 
to_sfixed(-402.0/65536.0,1,-nbitq), 
to_sfixed(-4182.0/65536.0,1,-nbitq), 
to_sfixed(-43.0/65536.0,1,-nbitq), 
to_sfixed(-3030.0/65536.0,1,-nbitq), 
to_sfixed(3082.0/65536.0,1,-nbitq), 
to_sfixed(-9529.0/65536.0,1,-nbitq), 
to_sfixed(6434.0/65536.0,1,-nbitq), 
to_sfixed(-8784.0/65536.0,1,-nbitq), 
to_sfixed(-3186.0/65536.0,1,-nbitq), 
to_sfixed(-1006.0/65536.0,1,-nbitq), 
to_sfixed(-4723.0/65536.0,1,-nbitq), 
to_sfixed(744.0/65536.0,1,-nbitq), 
to_sfixed(-223.0/65536.0,1,-nbitq), 
to_sfixed(-7867.0/65536.0,1,-nbitq), 
to_sfixed(5034.0/65536.0,1,-nbitq), 
to_sfixed(8361.0/65536.0,1,-nbitq), 
to_sfixed(3683.0/65536.0,1,-nbitq), 
to_sfixed(1139.0/65536.0,1,-nbitq), 
to_sfixed(1079.0/65536.0,1,-nbitq), 
to_sfixed(-11171.0/65536.0,1,-nbitq), 
to_sfixed(1292.0/65536.0,1,-nbitq), 
to_sfixed(-895.0/65536.0,1,-nbitq), 
to_sfixed(-281.0/65536.0,1,-nbitq), 
to_sfixed(-5413.0/65536.0,1,-nbitq), 
to_sfixed(-1995.0/65536.0,1,-nbitq), 
to_sfixed(3294.0/65536.0,1,-nbitq), 
to_sfixed(976.0/65536.0,1,-nbitq), 
to_sfixed(-1509.0/65536.0,1,-nbitq), 
to_sfixed(-614.0/65536.0,1,-nbitq), 
to_sfixed(-3111.0/65536.0,1,-nbitq), 
to_sfixed(5839.0/65536.0,1,-nbitq), 
to_sfixed(3056.0/65536.0,1,-nbitq), 
to_sfixed(-4963.0/65536.0,1,-nbitq), 
to_sfixed(1696.0/65536.0,1,-nbitq), 
to_sfixed(5551.0/65536.0,1,-nbitq), 
to_sfixed(-289.0/65536.0,1,-nbitq), 
to_sfixed(4333.0/65536.0,1,-nbitq), 
to_sfixed(-4550.0/65536.0,1,-nbitq), 
to_sfixed(1682.0/65536.0,1,-nbitq), 
to_sfixed(-2417.0/65536.0,1,-nbitq), 
to_sfixed(-843.0/65536.0,1,-nbitq), 
to_sfixed(-5559.0/65536.0,1,-nbitq), 
to_sfixed(16055.0/65536.0,1,-nbitq), 
to_sfixed(596.0/65536.0,1,-nbitq), 
to_sfixed(-2768.0/65536.0,1,-nbitq), 
to_sfixed(-5118.0/65536.0,1,-nbitq), 
to_sfixed(-6638.0/65536.0,1,-nbitq), 
to_sfixed(-4720.0/65536.0,1,-nbitq), 
to_sfixed(-2975.0/65536.0,1,-nbitq), 
to_sfixed(-7161.0/65536.0,1,-nbitq), 
to_sfixed(-2875.0/65536.0,1,-nbitq), 
to_sfixed(1739.0/65536.0,1,-nbitq), 
to_sfixed(-6071.0/65536.0,1,-nbitq), 
to_sfixed(2377.0/65536.0,1,-nbitq), 
to_sfixed(5540.0/65536.0,1,-nbitq), 
to_sfixed(236.0/65536.0,1,-nbitq), 
to_sfixed(-6754.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4205.0/65536.0,1,-nbitq), 
to_sfixed(10599.0/65536.0,1,-nbitq), 
to_sfixed(-5945.0/65536.0,1,-nbitq), 
to_sfixed(-2216.0/65536.0,1,-nbitq), 
to_sfixed(-11423.0/65536.0,1,-nbitq), 
to_sfixed(5175.0/65536.0,1,-nbitq), 
to_sfixed(-4606.0/65536.0,1,-nbitq), 
to_sfixed(-8100.0/65536.0,1,-nbitq), 
to_sfixed(-2742.0/65536.0,1,-nbitq), 
to_sfixed(-1156.0/65536.0,1,-nbitq), 
to_sfixed(-1343.0/65536.0,1,-nbitq), 
to_sfixed(-5786.0/65536.0,1,-nbitq), 
to_sfixed(2778.0/65536.0,1,-nbitq), 
to_sfixed(4683.0/65536.0,1,-nbitq), 
to_sfixed(3413.0/65536.0,1,-nbitq), 
to_sfixed(-2905.0/65536.0,1,-nbitq), 
to_sfixed(2321.0/65536.0,1,-nbitq), 
to_sfixed(-16948.0/65536.0,1,-nbitq), 
to_sfixed(4197.0/65536.0,1,-nbitq), 
to_sfixed(1980.0/65536.0,1,-nbitq), 
to_sfixed(-5531.0/65536.0,1,-nbitq), 
to_sfixed(11085.0/65536.0,1,-nbitq), 
to_sfixed(2624.0/65536.0,1,-nbitq), 
to_sfixed(-4335.0/65536.0,1,-nbitq), 
to_sfixed(-3635.0/65536.0,1,-nbitq), 
to_sfixed(-4131.0/65536.0,1,-nbitq), 
to_sfixed(5927.0/65536.0,1,-nbitq), 
to_sfixed(-584.0/65536.0,1,-nbitq), 
to_sfixed(-12626.0/65536.0,1,-nbitq), 
to_sfixed(2385.0/65536.0,1,-nbitq), 
to_sfixed(-31.0/65536.0,1,-nbitq), 
to_sfixed(4088.0/65536.0,1,-nbitq), 
to_sfixed(-5210.0/65536.0,1,-nbitq), 
to_sfixed(7093.0/65536.0,1,-nbitq), 
to_sfixed(-1107.0/65536.0,1,-nbitq), 
to_sfixed(-955.0/65536.0,1,-nbitq), 
to_sfixed(169.0/65536.0,1,-nbitq), 
to_sfixed(6567.0/65536.0,1,-nbitq), 
to_sfixed(15717.0/65536.0,1,-nbitq), 
to_sfixed(891.0/65536.0,1,-nbitq), 
to_sfixed(5791.0/65536.0,1,-nbitq), 
to_sfixed(1614.0/65536.0,1,-nbitq), 
to_sfixed(-8923.0/65536.0,1,-nbitq), 
to_sfixed(-1043.0/65536.0,1,-nbitq), 
to_sfixed(2955.0/65536.0,1,-nbitq), 
to_sfixed(439.0/65536.0,1,-nbitq), 
to_sfixed(-4242.0/65536.0,1,-nbitq), 
to_sfixed(-179.0/65536.0,1,-nbitq), 
to_sfixed(672.0/65536.0,1,-nbitq), 
to_sfixed(-1313.0/65536.0,1,-nbitq), 
to_sfixed(2803.0/65536.0,1,-nbitq), 
to_sfixed(382.0/65536.0,1,-nbitq), 
to_sfixed(-1849.0/65536.0,1,-nbitq), 
to_sfixed(-2155.0/65536.0,1,-nbitq), 
to_sfixed(7420.0/65536.0,1,-nbitq), 
to_sfixed(-7030.0/65536.0,1,-nbitq), 
to_sfixed(-676.0/65536.0,1,-nbitq), 
to_sfixed(1238.0/65536.0,1,-nbitq), 
to_sfixed(2048.0/65536.0,1,-nbitq), 
to_sfixed(3874.0/65536.0,1,-nbitq), 
to_sfixed(-9276.0/65536.0,1,-nbitq), 
to_sfixed(-2766.0/65536.0,1,-nbitq), 
to_sfixed(-1568.0/65536.0,1,-nbitq), 
to_sfixed(-1534.0/65536.0,1,-nbitq), 
to_sfixed(-2204.0/65536.0,1,-nbitq), 
to_sfixed(1187.0/65536.0,1,-nbitq), 
to_sfixed(-9512.0/65536.0,1,-nbitq), 
to_sfixed(8267.0/65536.0,1,-nbitq), 
to_sfixed(-4252.0/65536.0,1,-nbitq), 
to_sfixed(-8096.0/65536.0,1,-nbitq), 
to_sfixed(-5876.0/65536.0,1,-nbitq), 
to_sfixed(-1589.0/65536.0,1,-nbitq), 
to_sfixed(-7062.0/65536.0,1,-nbitq), 
to_sfixed(-599.0/65536.0,1,-nbitq), 
to_sfixed(-593.0/65536.0,1,-nbitq), 
to_sfixed(-11413.0/65536.0,1,-nbitq), 
to_sfixed(4409.0/65536.0,1,-nbitq), 
to_sfixed(-2966.0/65536.0,1,-nbitq), 
to_sfixed(141.0/65536.0,1,-nbitq), 
to_sfixed(4894.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4588.0/65536.0,1,-nbitq), 
to_sfixed(4882.0/65536.0,1,-nbitq), 
to_sfixed(-2507.0/65536.0,1,-nbitq), 
to_sfixed(-1190.0/65536.0,1,-nbitq), 
to_sfixed(7479.0/65536.0,1,-nbitq), 
to_sfixed(3909.0/65536.0,1,-nbitq), 
to_sfixed(259.0/65536.0,1,-nbitq), 
to_sfixed(-12080.0/65536.0,1,-nbitq), 
to_sfixed(-116.0/65536.0,1,-nbitq), 
to_sfixed(-868.0/65536.0,1,-nbitq), 
to_sfixed(-2713.0/65536.0,1,-nbitq), 
to_sfixed(-5347.0/65536.0,1,-nbitq), 
to_sfixed(-419.0/65536.0,1,-nbitq), 
to_sfixed(-4156.0/65536.0,1,-nbitq), 
to_sfixed(-608.0/65536.0,1,-nbitq), 
to_sfixed(-2705.0/65536.0,1,-nbitq), 
to_sfixed(1955.0/65536.0,1,-nbitq), 
to_sfixed(-8562.0/65536.0,1,-nbitq), 
to_sfixed(-852.0/65536.0,1,-nbitq), 
to_sfixed(-2504.0/65536.0,1,-nbitq), 
to_sfixed(-1165.0/65536.0,1,-nbitq), 
to_sfixed(5842.0/65536.0,1,-nbitq), 
to_sfixed(3.0/65536.0,1,-nbitq), 
to_sfixed(-887.0/65536.0,1,-nbitq), 
to_sfixed(662.0/65536.0,1,-nbitq), 
to_sfixed(-2418.0/65536.0,1,-nbitq), 
to_sfixed(1701.0/65536.0,1,-nbitq), 
to_sfixed(758.0/65536.0,1,-nbitq), 
to_sfixed(-13238.0/65536.0,1,-nbitq), 
to_sfixed(485.0/65536.0,1,-nbitq), 
to_sfixed(7444.0/65536.0,1,-nbitq), 
to_sfixed(6091.0/65536.0,1,-nbitq), 
to_sfixed(-10737.0/65536.0,1,-nbitq), 
to_sfixed(6628.0/65536.0,1,-nbitq), 
to_sfixed(-2781.0/65536.0,1,-nbitq), 
to_sfixed(-2307.0/65536.0,1,-nbitq), 
to_sfixed(-4863.0/65536.0,1,-nbitq), 
to_sfixed(5557.0/65536.0,1,-nbitq), 
to_sfixed(17918.0/65536.0,1,-nbitq), 
to_sfixed(-2555.0/65536.0,1,-nbitq), 
to_sfixed(4636.0/65536.0,1,-nbitq), 
to_sfixed(2103.0/65536.0,1,-nbitq), 
to_sfixed(-2738.0/65536.0,1,-nbitq), 
to_sfixed(-3015.0/65536.0,1,-nbitq), 
to_sfixed(2251.0/65536.0,1,-nbitq), 
to_sfixed(869.0/65536.0,1,-nbitq), 
to_sfixed(-1176.0/65536.0,1,-nbitq), 
to_sfixed(1273.0/65536.0,1,-nbitq), 
to_sfixed(-2133.0/65536.0,1,-nbitq), 
to_sfixed(-370.0/65536.0,1,-nbitq), 
to_sfixed(-1409.0/65536.0,1,-nbitq), 
to_sfixed(4993.0/65536.0,1,-nbitq), 
to_sfixed(693.0/65536.0,1,-nbitq), 
to_sfixed(-6073.0/65536.0,1,-nbitq), 
to_sfixed(4420.0/65536.0,1,-nbitq), 
to_sfixed(-1261.0/65536.0,1,-nbitq), 
to_sfixed(897.0/65536.0,1,-nbitq), 
to_sfixed(641.0/65536.0,1,-nbitq), 
to_sfixed(1293.0/65536.0,1,-nbitq), 
to_sfixed(5990.0/65536.0,1,-nbitq), 
to_sfixed(-5424.0/65536.0,1,-nbitq), 
to_sfixed(-150.0/65536.0,1,-nbitq), 
to_sfixed(2934.0/65536.0,1,-nbitq), 
to_sfixed(-3010.0/65536.0,1,-nbitq), 
to_sfixed(-8903.0/65536.0,1,-nbitq), 
to_sfixed(-6448.0/65536.0,1,-nbitq), 
to_sfixed(-8748.0/65536.0,1,-nbitq), 
to_sfixed(588.0/65536.0,1,-nbitq), 
to_sfixed(-3672.0/65536.0,1,-nbitq), 
to_sfixed(4861.0/65536.0,1,-nbitq), 
to_sfixed(195.0/65536.0,1,-nbitq), 
to_sfixed(5264.0/65536.0,1,-nbitq), 
to_sfixed(-8392.0/65536.0,1,-nbitq), 
to_sfixed(897.0/65536.0,1,-nbitq), 
to_sfixed(151.0/65536.0,1,-nbitq), 
to_sfixed(-14658.0/65536.0,1,-nbitq), 
to_sfixed(9245.0/65536.0,1,-nbitq), 
to_sfixed(-2518.0/65536.0,1,-nbitq), 
to_sfixed(-1439.0/65536.0,1,-nbitq), 
to_sfixed(6421.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3660.0/65536.0,1,-nbitq), 
to_sfixed(1064.0/65536.0,1,-nbitq), 
to_sfixed(5935.0/65536.0,1,-nbitq), 
to_sfixed(-197.0/65536.0,1,-nbitq), 
to_sfixed(4610.0/65536.0,1,-nbitq), 
to_sfixed(3504.0/65536.0,1,-nbitq), 
to_sfixed(3253.0/65536.0,1,-nbitq), 
to_sfixed(-11385.0/65536.0,1,-nbitq), 
to_sfixed(-971.0/65536.0,1,-nbitq), 
to_sfixed(3144.0/65536.0,1,-nbitq), 
to_sfixed(1228.0/65536.0,1,-nbitq), 
to_sfixed(5472.0/65536.0,1,-nbitq), 
to_sfixed(404.0/65536.0,1,-nbitq), 
to_sfixed(-10269.0/65536.0,1,-nbitq), 
to_sfixed(824.0/65536.0,1,-nbitq), 
to_sfixed(1448.0/65536.0,1,-nbitq), 
to_sfixed(-2446.0/65536.0,1,-nbitq), 
to_sfixed(2645.0/65536.0,1,-nbitq), 
to_sfixed(-3797.0/65536.0,1,-nbitq), 
to_sfixed(1067.0/65536.0,1,-nbitq), 
to_sfixed(1815.0/65536.0,1,-nbitq), 
to_sfixed(7225.0/65536.0,1,-nbitq), 
to_sfixed(9648.0/65536.0,1,-nbitq), 
to_sfixed(-646.0/65536.0,1,-nbitq), 
to_sfixed(1738.0/65536.0,1,-nbitq), 
to_sfixed(-6346.0/65536.0,1,-nbitq), 
to_sfixed(2930.0/65536.0,1,-nbitq), 
to_sfixed(-1390.0/65536.0,1,-nbitq), 
to_sfixed(-6226.0/65536.0,1,-nbitq), 
to_sfixed(915.0/65536.0,1,-nbitq), 
to_sfixed(14645.0/65536.0,1,-nbitq), 
to_sfixed(11543.0/65536.0,1,-nbitq), 
to_sfixed(-3153.0/65536.0,1,-nbitq), 
to_sfixed(12159.0/65536.0,1,-nbitq), 
to_sfixed(-869.0/65536.0,1,-nbitq), 
to_sfixed(1005.0/65536.0,1,-nbitq), 
to_sfixed(-3020.0/65536.0,1,-nbitq), 
to_sfixed(5127.0/65536.0,1,-nbitq), 
to_sfixed(11059.0/65536.0,1,-nbitq), 
to_sfixed(3388.0/65536.0,1,-nbitq), 
to_sfixed(-5401.0/65536.0,1,-nbitq), 
to_sfixed(-1049.0/65536.0,1,-nbitq), 
to_sfixed(2408.0/65536.0,1,-nbitq), 
to_sfixed(-7710.0/65536.0,1,-nbitq), 
to_sfixed(-169.0/65536.0,1,-nbitq), 
to_sfixed(-1091.0/65536.0,1,-nbitq), 
to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(-1458.0/65536.0,1,-nbitq), 
to_sfixed(-1106.0/65536.0,1,-nbitq), 
to_sfixed(605.0/65536.0,1,-nbitq), 
to_sfixed(1114.0/65536.0,1,-nbitq), 
to_sfixed(-2780.0/65536.0,1,-nbitq), 
to_sfixed(-2086.0/65536.0,1,-nbitq), 
to_sfixed(7042.0/65536.0,1,-nbitq), 
to_sfixed(3558.0/65536.0,1,-nbitq), 
to_sfixed(-1555.0/65536.0,1,-nbitq), 
to_sfixed(-1254.0/65536.0,1,-nbitq), 
to_sfixed(-6752.0/65536.0,1,-nbitq), 
to_sfixed(1158.0/65536.0,1,-nbitq), 
to_sfixed(1950.0/65536.0,1,-nbitq), 
to_sfixed(-672.0/65536.0,1,-nbitq), 
to_sfixed(2247.0/65536.0,1,-nbitq), 
to_sfixed(255.0/65536.0,1,-nbitq), 
to_sfixed(1911.0/65536.0,1,-nbitq), 
to_sfixed(-10736.0/65536.0,1,-nbitq), 
to_sfixed(-8456.0/65536.0,1,-nbitq), 
to_sfixed(-2455.0/65536.0,1,-nbitq), 
to_sfixed(-4656.0/65536.0,1,-nbitq), 
to_sfixed(-545.0/65536.0,1,-nbitq), 
to_sfixed(3272.0/65536.0,1,-nbitq), 
to_sfixed(-2891.0/65536.0,1,-nbitq), 
to_sfixed(1747.0/65536.0,1,-nbitq), 
to_sfixed(-4956.0/65536.0,1,-nbitq), 
to_sfixed(-660.0/65536.0,1,-nbitq), 
to_sfixed(-2630.0/65536.0,1,-nbitq), 
to_sfixed(4472.0/65536.0,1,-nbitq), 
to_sfixed(3439.0/65536.0,1,-nbitq), 
to_sfixed(6604.0/65536.0,1,-nbitq), 
to_sfixed(-1897.0/65536.0,1,-nbitq), 
to_sfixed(-385.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3654.0/65536.0,1,-nbitq), 
to_sfixed(-2425.0/65536.0,1,-nbitq), 
to_sfixed(2755.0/65536.0,1,-nbitq), 
to_sfixed(-3156.0/65536.0,1,-nbitq), 
to_sfixed(3719.0/65536.0,1,-nbitq), 
to_sfixed(4512.0/65536.0,1,-nbitq), 
to_sfixed(2399.0/65536.0,1,-nbitq), 
to_sfixed(-10764.0/65536.0,1,-nbitq), 
to_sfixed(-7233.0/65536.0,1,-nbitq), 
to_sfixed(3137.0/65536.0,1,-nbitq), 
to_sfixed(-1.0/65536.0,1,-nbitq), 
to_sfixed(-2222.0/65536.0,1,-nbitq), 
to_sfixed(-1265.0/65536.0,1,-nbitq), 
to_sfixed(-5116.0/65536.0,1,-nbitq), 
to_sfixed(2196.0/65536.0,1,-nbitq), 
to_sfixed(-1300.0/65536.0,1,-nbitq), 
to_sfixed(2020.0/65536.0,1,-nbitq), 
to_sfixed(8159.0/65536.0,1,-nbitq), 
to_sfixed(-362.0/65536.0,1,-nbitq), 
to_sfixed(-1539.0/65536.0,1,-nbitq), 
to_sfixed(-1018.0/65536.0,1,-nbitq), 
to_sfixed(6635.0/65536.0,1,-nbitq), 
to_sfixed(1253.0/65536.0,1,-nbitq), 
to_sfixed(2719.0/65536.0,1,-nbitq), 
to_sfixed(2587.0/65536.0,1,-nbitq), 
to_sfixed(-518.0/65536.0,1,-nbitq), 
to_sfixed(3567.0/65536.0,1,-nbitq), 
to_sfixed(-3270.0/65536.0,1,-nbitq), 
to_sfixed(-3420.0/65536.0,1,-nbitq), 
to_sfixed(3228.0/65536.0,1,-nbitq), 
to_sfixed(8559.0/65536.0,1,-nbitq), 
to_sfixed(15880.0/65536.0,1,-nbitq), 
to_sfixed(-4777.0/65536.0,1,-nbitq), 
to_sfixed(7642.0/65536.0,1,-nbitq), 
to_sfixed(-3252.0/65536.0,1,-nbitq), 
to_sfixed(-1195.0/65536.0,1,-nbitq), 
to_sfixed(1677.0/65536.0,1,-nbitq), 
to_sfixed(4880.0/65536.0,1,-nbitq), 
to_sfixed(-1620.0/65536.0,1,-nbitq), 
to_sfixed(3879.0/65536.0,1,-nbitq), 
to_sfixed(3325.0/65536.0,1,-nbitq), 
to_sfixed(-12.0/65536.0,1,-nbitq), 
to_sfixed(2017.0/65536.0,1,-nbitq), 
to_sfixed(-12035.0/65536.0,1,-nbitq), 
to_sfixed(-1724.0/65536.0,1,-nbitq), 
to_sfixed(-1664.0/65536.0,1,-nbitq), 
to_sfixed(-494.0/65536.0,1,-nbitq), 
to_sfixed(-8483.0/65536.0,1,-nbitq), 
to_sfixed(1431.0/65536.0,1,-nbitq), 
to_sfixed(1785.0/65536.0,1,-nbitq), 
to_sfixed(-2719.0/65536.0,1,-nbitq), 
to_sfixed(-2497.0/65536.0,1,-nbitq), 
to_sfixed(2206.0/65536.0,1,-nbitq), 
to_sfixed(2036.0/65536.0,1,-nbitq), 
to_sfixed(5487.0/65536.0,1,-nbitq), 
to_sfixed(6132.0/65536.0,1,-nbitq), 
to_sfixed(-1414.0/65536.0,1,-nbitq), 
to_sfixed(-5394.0/65536.0,1,-nbitq), 
to_sfixed(867.0/65536.0,1,-nbitq), 
to_sfixed(6878.0/65536.0,1,-nbitq), 
to_sfixed(-1003.0/65536.0,1,-nbitq), 
to_sfixed(-207.0/65536.0,1,-nbitq), 
to_sfixed(243.0/65536.0,1,-nbitq), 
to_sfixed(-523.0/65536.0,1,-nbitq), 
to_sfixed(-12888.0/65536.0,1,-nbitq), 
to_sfixed(-3724.0/65536.0,1,-nbitq), 
to_sfixed(2077.0/65536.0,1,-nbitq), 
to_sfixed(-4226.0/65536.0,1,-nbitq), 
to_sfixed(-6480.0/65536.0,1,-nbitq), 
to_sfixed(-4085.0/65536.0,1,-nbitq), 
to_sfixed(-70.0/65536.0,1,-nbitq), 
to_sfixed(-2025.0/65536.0,1,-nbitq), 
to_sfixed(1568.0/65536.0,1,-nbitq), 
to_sfixed(1419.0/65536.0,1,-nbitq), 
to_sfixed(-1292.0/65536.0,1,-nbitq), 
to_sfixed(8594.0/65536.0,1,-nbitq), 
to_sfixed(11063.0/65536.0,1,-nbitq), 
to_sfixed(-2305.0/65536.0,1,-nbitq), 
to_sfixed(-1863.0/65536.0,1,-nbitq), 
to_sfixed(-862.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3436.0/65536.0,1,-nbitq), 
to_sfixed(1747.0/65536.0,1,-nbitq), 
to_sfixed(-2756.0/65536.0,1,-nbitq), 
to_sfixed(2368.0/65536.0,1,-nbitq), 
to_sfixed(-3002.0/65536.0,1,-nbitq), 
to_sfixed(-7098.0/65536.0,1,-nbitq), 
to_sfixed(10082.0/65536.0,1,-nbitq), 
to_sfixed(-6248.0/65536.0,1,-nbitq), 
to_sfixed(-5626.0/65536.0,1,-nbitq), 
to_sfixed(535.0/65536.0,1,-nbitq), 
to_sfixed(-1395.0/65536.0,1,-nbitq), 
to_sfixed(-8619.0/65536.0,1,-nbitq), 
to_sfixed(-2051.0/65536.0,1,-nbitq), 
to_sfixed(-1514.0/65536.0,1,-nbitq), 
to_sfixed(2250.0/65536.0,1,-nbitq), 
to_sfixed(-1882.0/65536.0,1,-nbitq), 
to_sfixed(390.0/65536.0,1,-nbitq), 
to_sfixed(14138.0/65536.0,1,-nbitq), 
to_sfixed(-1479.0/65536.0,1,-nbitq), 
to_sfixed(1222.0/65536.0,1,-nbitq), 
to_sfixed(-1792.0/65536.0,1,-nbitq), 
to_sfixed(10152.0/65536.0,1,-nbitq), 
to_sfixed(1555.0/65536.0,1,-nbitq), 
to_sfixed(-4000.0/65536.0,1,-nbitq), 
to_sfixed(4690.0/65536.0,1,-nbitq), 
to_sfixed(-3822.0/65536.0,1,-nbitq), 
to_sfixed(1446.0/65536.0,1,-nbitq), 
to_sfixed(745.0/65536.0,1,-nbitq), 
to_sfixed(-10726.0/65536.0,1,-nbitq), 
to_sfixed(1572.0/65536.0,1,-nbitq), 
to_sfixed(-5234.0/65536.0,1,-nbitq), 
to_sfixed(11398.0/65536.0,1,-nbitq), 
to_sfixed(1005.0/65536.0,1,-nbitq), 
to_sfixed(-5231.0/65536.0,1,-nbitq), 
to_sfixed(-2788.0/65536.0,1,-nbitq), 
to_sfixed(3019.0/65536.0,1,-nbitq), 
to_sfixed(-2662.0/65536.0,1,-nbitq), 
to_sfixed(3187.0/65536.0,1,-nbitq), 
to_sfixed(-7251.0/65536.0,1,-nbitq), 
to_sfixed(2605.0/65536.0,1,-nbitq), 
to_sfixed(5023.0/65536.0,1,-nbitq), 
to_sfixed(1318.0/65536.0,1,-nbitq), 
to_sfixed(-4101.0/65536.0,1,-nbitq), 
to_sfixed(-15735.0/65536.0,1,-nbitq), 
to_sfixed(672.0/65536.0,1,-nbitq), 
to_sfixed(-7872.0/65536.0,1,-nbitq), 
to_sfixed(126.0/65536.0,1,-nbitq), 
to_sfixed(-7770.0/65536.0,1,-nbitq), 
to_sfixed(3315.0/65536.0,1,-nbitq), 
to_sfixed(3958.0/65536.0,1,-nbitq), 
to_sfixed(2997.0/65536.0,1,-nbitq), 
to_sfixed(136.0/65536.0,1,-nbitq), 
to_sfixed(-4818.0/65536.0,1,-nbitq), 
to_sfixed(-1159.0/65536.0,1,-nbitq), 
to_sfixed(3036.0/65536.0,1,-nbitq), 
to_sfixed(145.0/65536.0,1,-nbitq), 
to_sfixed(1592.0/65536.0,1,-nbitq), 
to_sfixed(-7231.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(495.0/65536.0,1,-nbitq), 
to_sfixed(-2369.0/65536.0,1,-nbitq), 
to_sfixed(-2263.0/65536.0,1,-nbitq), 
to_sfixed(2852.0/65536.0,1,-nbitq), 
to_sfixed(-994.0/65536.0,1,-nbitq), 
to_sfixed(-17896.0/65536.0,1,-nbitq), 
to_sfixed(-9971.0/65536.0,1,-nbitq), 
to_sfixed(3800.0/65536.0,1,-nbitq), 
to_sfixed(-2687.0/65536.0,1,-nbitq), 
to_sfixed(-7010.0/65536.0,1,-nbitq), 
to_sfixed(-449.0/65536.0,1,-nbitq), 
to_sfixed(2417.0/65536.0,1,-nbitq), 
to_sfixed(2751.0/65536.0,1,-nbitq), 
to_sfixed(553.0/65536.0,1,-nbitq), 
to_sfixed(-1799.0/65536.0,1,-nbitq), 
to_sfixed(-2046.0/65536.0,1,-nbitq), 
to_sfixed(3458.0/65536.0,1,-nbitq), 
to_sfixed(9971.0/65536.0,1,-nbitq), 
to_sfixed(-5380.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(-969.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1345.0/65536.0,1,-nbitq), 
to_sfixed(534.0/65536.0,1,-nbitq), 
to_sfixed(3690.0/65536.0,1,-nbitq), 
to_sfixed(2319.0/65536.0,1,-nbitq), 
to_sfixed(-11667.0/65536.0,1,-nbitq), 
to_sfixed(-1652.0/65536.0,1,-nbitq), 
to_sfixed(4870.0/65536.0,1,-nbitq), 
to_sfixed(361.0/65536.0,1,-nbitq), 
to_sfixed(-3822.0/65536.0,1,-nbitq), 
to_sfixed(1138.0/65536.0,1,-nbitq), 
to_sfixed(-2491.0/65536.0,1,-nbitq), 
to_sfixed(-3989.0/65536.0,1,-nbitq), 
to_sfixed(2189.0/65536.0,1,-nbitq), 
to_sfixed(-1865.0/65536.0,1,-nbitq), 
to_sfixed(-1533.0/65536.0,1,-nbitq), 
to_sfixed(704.0/65536.0,1,-nbitq), 
to_sfixed(-1087.0/65536.0,1,-nbitq), 
to_sfixed(2094.0/65536.0,1,-nbitq), 
to_sfixed(-3784.0/65536.0,1,-nbitq), 
to_sfixed(2902.0/65536.0,1,-nbitq), 
to_sfixed(3580.0/65536.0,1,-nbitq), 
to_sfixed(10119.0/65536.0,1,-nbitq), 
to_sfixed(4471.0/65536.0,1,-nbitq), 
to_sfixed(1207.0/65536.0,1,-nbitq), 
to_sfixed(5352.0/65536.0,1,-nbitq), 
to_sfixed(-10447.0/65536.0,1,-nbitq), 
to_sfixed(8665.0/65536.0,1,-nbitq), 
to_sfixed(824.0/65536.0,1,-nbitq), 
to_sfixed(-4701.0/65536.0,1,-nbitq), 
to_sfixed(1888.0/65536.0,1,-nbitq), 
to_sfixed(-10618.0/65536.0,1,-nbitq), 
to_sfixed(7930.0/65536.0,1,-nbitq), 
to_sfixed(2764.0/65536.0,1,-nbitq), 
to_sfixed(-5734.0/65536.0,1,-nbitq), 
to_sfixed(1677.0/65536.0,1,-nbitq), 
to_sfixed(2971.0/65536.0,1,-nbitq), 
to_sfixed(-5163.0/65536.0,1,-nbitq), 
to_sfixed(-4079.0/65536.0,1,-nbitq), 
to_sfixed(-7094.0/65536.0,1,-nbitq), 
to_sfixed(2701.0/65536.0,1,-nbitq), 
to_sfixed(2109.0/65536.0,1,-nbitq), 
to_sfixed(2275.0/65536.0,1,-nbitq), 
to_sfixed(2471.0/65536.0,1,-nbitq), 
to_sfixed(-15629.0/65536.0,1,-nbitq), 
to_sfixed(-1720.0/65536.0,1,-nbitq), 
to_sfixed(-3407.0/65536.0,1,-nbitq), 
to_sfixed(-2091.0/65536.0,1,-nbitq), 
to_sfixed(-1659.0/65536.0,1,-nbitq), 
to_sfixed(-1956.0/65536.0,1,-nbitq), 
to_sfixed(5081.0/65536.0,1,-nbitq), 
to_sfixed(2777.0/65536.0,1,-nbitq), 
to_sfixed(222.0/65536.0,1,-nbitq), 
to_sfixed(-4077.0/65536.0,1,-nbitq), 
to_sfixed(-61.0/65536.0,1,-nbitq), 
to_sfixed(2128.0/65536.0,1,-nbitq), 
to_sfixed(-540.0/65536.0,1,-nbitq), 
to_sfixed(-844.0/65536.0,1,-nbitq), 
to_sfixed(-7732.0/65536.0,1,-nbitq), 
to_sfixed(1989.0/65536.0,1,-nbitq), 
to_sfixed(441.0/65536.0,1,-nbitq), 
to_sfixed(240.0/65536.0,1,-nbitq), 
to_sfixed(1696.0/65536.0,1,-nbitq), 
to_sfixed(-275.0/65536.0,1,-nbitq), 
to_sfixed(-161.0/65536.0,1,-nbitq), 
to_sfixed(-12465.0/65536.0,1,-nbitq), 
to_sfixed(-10157.0/65536.0,1,-nbitq), 
to_sfixed(-3977.0/65536.0,1,-nbitq), 
to_sfixed(-1455.0/65536.0,1,-nbitq), 
to_sfixed(-5239.0/65536.0,1,-nbitq), 
to_sfixed(647.0/65536.0,1,-nbitq), 
to_sfixed(2980.0/65536.0,1,-nbitq), 
to_sfixed(-2534.0/65536.0,1,-nbitq), 
to_sfixed(-3805.0/65536.0,1,-nbitq), 
to_sfixed(-676.0/65536.0,1,-nbitq), 
to_sfixed(-1416.0/65536.0,1,-nbitq), 
to_sfixed(1994.0/65536.0,1,-nbitq), 
to_sfixed(7015.0/65536.0,1,-nbitq), 
to_sfixed(-4029.0/65536.0,1,-nbitq), 
to_sfixed(-1545.0/65536.0,1,-nbitq), 
to_sfixed(-4201.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2195.0/65536.0,1,-nbitq), 
to_sfixed(-2882.0/65536.0,1,-nbitq), 
to_sfixed(-1476.0/65536.0,1,-nbitq), 
to_sfixed(962.0/65536.0,1,-nbitq), 
to_sfixed(-9476.0/65536.0,1,-nbitq), 
to_sfixed(-6648.0/65536.0,1,-nbitq), 
to_sfixed(1859.0/65536.0,1,-nbitq), 
to_sfixed(1828.0/65536.0,1,-nbitq), 
to_sfixed(-1285.0/65536.0,1,-nbitq), 
to_sfixed(-640.0/65536.0,1,-nbitq), 
to_sfixed(-561.0/65536.0,1,-nbitq), 
to_sfixed(-5998.0/65536.0,1,-nbitq), 
to_sfixed(2486.0/65536.0,1,-nbitq), 
to_sfixed(-7446.0/65536.0,1,-nbitq), 
to_sfixed(-3317.0/65536.0,1,-nbitq), 
to_sfixed(-2484.0/65536.0,1,-nbitq), 
to_sfixed(-2550.0/65536.0,1,-nbitq), 
to_sfixed(2107.0/65536.0,1,-nbitq), 
to_sfixed(-8891.0/65536.0,1,-nbitq), 
to_sfixed(-221.0/65536.0,1,-nbitq), 
to_sfixed(4974.0/65536.0,1,-nbitq), 
to_sfixed(11153.0/65536.0,1,-nbitq), 
to_sfixed(3582.0/65536.0,1,-nbitq), 
to_sfixed(-422.0/65536.0,1,-nbitq), 
to_sfixed(3928.0/65536.0,1,-nbitq), 
to_sfixed(-11963.0/65536.0,1,-nbitq), 
to_sfixed(-3524.0/65536.0,1,-nbitq), 
to_sfixed(-1201.0/65536.0,1,-nbitq), 
to_sfixed(-10830.0/65536.0,1,-nbitq), 
to_sfixed(77.0/65536.0,1,-nbitq), 
to_sfixed(-7801.0/65536.0,1,-nbitq), 
to_sfixed(7479.0/65536.0,1,-nbitq), 
to_sfixed(1230.0/65536.0,1,-nbitq), 
to_sfixed(-5840.0/65536.0,1,-nbitq), 
to_sfixed(1688.0/65536.0,1,-nbitq), 
to_sfixed(2011.0/65536.0,1,-nbitq), 
to_sfixed(-7614.0/65536.0,1,-nbitq), 
to_sfixed(-6816.0/65536.0,1,-nbitq), 
to_sfixed(-3210.0/65536.0,1,-nbitq), 
to_sfixed(2025.0/65536.0,1,-nbitq), 
to_sfixed(5531.0/65536.0,1,-nbitq), 
to_sfixed(-2040.0/65536.0,1,-nbitq), 
to_sfixed(4000.0/65536.0,1,-nbitq), 
to_sfixed(-12695.0/65536.0,1,-nbitq), 
to_sfixed(2592.0/65536.0,1,-nbitq), 
to_sfixed(4612.0/65536.0,1,-nbitq), 
to_sfixed(-3889.0/65536.0,1,-nbitq), 
to_sfixed(-5590.0/65536.0,1,-nbitq), 
to_sfixed(-2975.0/65536.0,1,-nbitq), 
to_sfixed(3842.0/65536.0,1,-nbitq), 
to_sfixed(-1208.0/65536.0,1,-nbitq), 
to_sfixed(-2557.0/65536.0,1,-nbitq), 
to_sfixed(-5394.0/65536.0,1,-nbitq), 
to_sfixed(1248.0/65536.0,1,-nbitq), 
to_sfixed(2994.0/65536.0,1,-nbitq), 
to_sfixed(-4902.0/65536.0,1,-nbitq), 
to_sfixed(1316.0/65536.0,1,-nbitq), 
to_sfixed(-4651.0/65536.0,1,-nbitq), 
to_sfixed(-1584.0/65536.0,1,-nbitq), 
to_sfixed(-4086.0/65536.0,1,-nbitq), 
to_sfixed(-2914.0/65536.0,1,-nbitq), 
to_sfixed(-2490.0/65536.0,1,-nbitq), 
to_sfixed(51.0/65536.0,1,-nbitq), 
to_sfixed(-1021.0/65536.0,1,-nbitq), 
to_sfixed(-8045.0/65536.0,1,-nbitq), 
to_sfixed(-10991.0/65536.0,1,-nbitq), 
to_sfixed(-4005.0/65536.0,1,-nbitq), 
to_sfixed(-3618.0/65536.0,1,-nbitq), 
to_sfixed(-1634.0/65536.0,1,-nbitq), 
to_sfixed(4826.0/65536.0,1,-nbitq), 
to_sfixed(-1055.0/65536.0,1,-nbitq), 
to_sfixed(2156.0/65536.0,1,-nbitq), 
to_sfixed(-2755.0/65536.0,1,-nbitq), 
to_sfixed(2789.0/65536.0,1,-nbitq), 
to_sfixed(1943.0/65536.0,1,-nbitq), 
to_sfixed(-5245.0/65536.0,1,-nbitq), 
to_sfixed(278.0/65536.0,1,-nbitq), 
to_sfixed(1810.0/65536.0,1,-nbitq), 
to_sfixed(661.0/65536.0,1,-nbitq), 
to_sfixed(236.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1331.0/65536.0,1,-nbitq), 
to_sfixed(-4040.0/65536.0,1,-nbitq), 
to_sfixed(7077.0/65536.0,1,-nbitq), 
to_sfixed(185.0/65536.0,1,-nbitq), 
to_sfixed(-4756.0/65536.0,1,-nbitq), 
to_sfixed(-3669.0/65536.0,1,-nbitq), 
to_sfixed(795.0/65536.0,1,-nbitq), 
to_sfixed(-3991.0/65536.0,1,-nbitq), 
to_sfixed(-2288.0/65536.0,1,-nbitq), 
to_sfixed(-740.0/65536.0,1,-nbitq), 
to_sfixed(-870.0/65536.0,1,-nbitq), 
to_sfixed(652.0/65536.0,1,-nbitq), 
to_sfixed(-66.0/65536.0,1,-nbitq), 
to_sfixed(-6674.0/65536.0,1,-nbitq), 
to_sfixed(2817.0/65536.0,1,-nbitq), 
to_sfixed(2050.0/65536.0,1,-nbitq), 
to_sfixed(-2425.0/65536.0,1,-nbitq), 
to_sfixed(573.0/65536.0,1,-nbitq), 
to_sfixed(-3413.0/65536.0,1,-nbitq), 
to_sfixed(-933.0/65536.0,1,-nbitq), 
to_sfixed(1915.0/65536.0,1,-nbitq), 
to_sfixed(5631.0/65536.0,1,-nbitq), 
to_sfixed(-406.0/65536.0,1,-nbitq), 
to_sfixed(-145.0/65536.0,1,-nbitq), 
to_sfixed(4506.0/65536.0,1,-nbitq), 
to_sfixed(-5908.0/65536.0,1,-nbitq), 
to_sfixed(-7920.0/65536.0,1,-nbitq), 
to_sfixed(-2173.0/65536.0,1,-nbitq), 
to_sfixed(-6785.0/65536.0,1,-nbitq), 
to_sfixed(13.0/65536.0,1,-nbitq), 
to_sfixed(-1964.0/65536.0,1,-nbitq), 
to_sfixed(7401.0/65536.0,1,-nbitq), 
to_sfixed(1300.0/65536.0,1,-nbitq), 
to_sfixed(3621.0/65536.0,1,-nbitq), 
to_sfixed(-1602.0/65536.0,1,-nbitq), 
to_sfixed(-1124.0/65536.0,1,-nbitq), 
to_sfixed(152.0/65536.0,1,-nbitq), 
to_sfixed(-3730.0/65536.0,1,-nbitq), 
to_sfixed(3760.0/65536.0,1,-nbitq), 
to_sfixed(4761.0/65536.0,1,-nbitq), 
to_sfixed(3091.0/65536.0,1,-nbitq), 
to_sfixed(9.0/65536.0,1,-nbitq), 
to_sfixed(928.0/65536.0,1,-nbitq), 
to_sfixed(-9556.0/65536.0,1,-nbitq), 
to_sfixed(-1388.0/65536.0,1,-nbitq), 
to_sfixed(304.0/65536.0,1,-nbitq), 
to_sfixed(-2983.0/65536.0,1,-nbitq), 
to_sfixed(-5112.0/65536.0,1,-nbitq), 
to_sfixed(-724.0/65536.0,1,-nbitq), 
to_sfixed(529.0/65536.0,1,-nbitq), 
to_sfixed(-1566.0/65536.0,1,-nbitq), 
to_sfixed(-30.0/65536.0,1,-nbitq), 
to_sfixed(-2965.0/65536.0,1,-nbitq), 
to_sfixed(2939.0/65536.0,1,-nbitq), 
to_sfixed(1654.0/65536.0,1,-nbitq), 
to_sfixed(-918.0/65536.0,1,-nbitq), 
to_sfixed(-487.0/65536.0,1,-nbitq), 
to_sfixed(-695.0/65536.0,1,-nbitq), 
to_sfixed(782.0/65536.0,1,-nbitq), 
to_sfixed(-441.0/65536.0,1,-nbitq), 
to_sfixed(-835.0/65536.0,1,-nbitq), 
to_sfixed(-337.0/65536.0,1,-nbitq), 
to_sfixed(-571.0/65536.0,1,-nbitq), 
to_sfixed(-1308.0/65536.0,1,-nbitq), 
to_sfixed(-6807.0/65536.0,1,-nbitq), 
to_sfixed(-6407.0/65536.0,1,-nbitq), 
to_sfixed(-793.0/65536.0,1,-nbitq), 
to_sfixed(-9440.0/65536.0,1,-nbitq), 
to_sfixed(-1012.0/65536.0,1,-nbitq), 
to_sfixed(2500.0/65536.0,1,-nbitq), 
to_sfixed(-2117.0/65536.0,1,-nbitq), 
to_sfixed(2746.0/65536.0,1,-nbitq), 
to_sfixed(-546.0/65536.0,1,-nbitq), 
to_sfixed(-2415.0/65536.0,1,-nbitq), 
to_sfixed(342.0/65536.0,1,-nbitq), 
to_sfixed(-1835.0/65536.0,1,-nbitq), 
to_sfixed(-6371.0/65536.0,1,-nbitq), 
to_sfixed(131.0/65536.0,1,-nbitq), 
to_sfixed(-3280.0/65536.0,1,-nbitq), 
to_sfixed(-1160.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3926.0/65536.0,1,-nbitq), 
to_sfixed(-1443.0/65536.0,1,-nbitq), 
to_sfixed(2088.0/65536.0,1,-nbitq), 
to_sfixed(-3019.0/65536.0,1,-nbitq), 
to_sfixed(-3691.0/65536.0,1,-nbitq), 
to_sfixed(-4483.0/65536.0,1,-nbitq), 
to_sfixed(2454.0/65536.0,1,-nbitq), 
to_sfixed(-2387.0/65536.0,1,-nbitq), 
to_sfixed(4340.0/65536.0,1,-nbitq), 
to_sfixed(1150.0/65536.0,1,-nbitq), 
to_sfixed(-2505.0/65536.0,1,-nbitq), 
to_sfixed(4043.0/65536.0,1,-nbitq), 
to_sfixed(-614.0/65536.0,1,-nbitq), 
to_sfixed(-4548.0/65536.0,1,-nbitq), 
to_sfixed(497.0/65536.0,1,-nbitq), 
to_sfixed(-2425.0/65536.0,1,-nbitq), 
to_sfixed(-123.0/65536.0,1,-nbitq), 
to_sfixed(528.0/65536.0,1,-nbitq), 
to_sfixed(-3079.0/65536.0,1,-nbitq), 
to_sfixed(3200.0/65536.0,1,-nbitq), 
to_sfixed(1611.0/65536.0,1,-nbitq), 
to_sfixed(-621.0/65536.0,1,-nbitq), 
to_sfixed(152.0/65536.0,1,-nbitq), 
to_sfixed(-6771.0/65536.0,1,-nbitq), 
to_sfixed(4522.0/65536.0,1,-nbitq), 
to_sfixed(-3569.0/65536.0,1,-nbitq), 
to_sfixed(-6649.0/65536.0,1,-nbitq), 
to_sfixed(846.0/65536.0,1,-nbitq), 
to_sfixed(-3672.0/65536.0,1,-nbitq), 
to_sfixed(1983.0/65536.0,1,-nbitq), 
to_sfixed(-2106.0/65536.0,1,-nbitq), 
to_sfixed(3709.0/65536.0,1,-nbitq), 
to_sfixed(2181.0/65536.0,1,-nbitq), 
to_sfixed(6955.0/65536.0,1,-nbitq), 
to_sfixed(-1110.0/65536.0,1,-nbitq), 
to_sfixed(-748.0/65536.0,1,-nbitq), 
to_sfixed(730.0/65536.0,1,-nbitq), 
to_sfixed(-2288.0/65536.0,1,-nbitq), 
to_sfixed(4447.0/65536.0,1,-nbitq), 
to_sfixed(-372.0/65536.0,1,-nbitq), 
to_sfixed(1218.0/65536.0,1,-nbitq), 
to_sfixed(-1692.0/65536.0,1,-nbitq), 
to_sfixed(3079.0/65536.0,1,-nbitq), 
to_sfixed(-6890.0/65536.0,1,-nbitq), 
to_sfixed(-1161.0/65536.0,1,-nbitq), 
to_sfixed(-2312.0/65536.0,1,-nbitq), 
to_sfixed(-2045.0/65536.0,1,-nbitq), 
to_sfixed(-1620.0/65536.0,1,-nbitq), 
to_sfixed(1976.0/65536.0,1,-nbitq), 
to_sfixed(2899.0/65536.0,1,-nbitq), 
to_sfixed(556.0/65536.0,1,-nbitq), 
to_sfixed(2219.0/65536.0,1,-nbitq), 
to_sfixed(-3169.0/65536.0,1,-nbitq), 
to_sfixed(3924.0/65536.0,1,-nbitq), 
to_sfixed(329.0/65536.0,1,-nbitq), 
to_sfixed(609.0/65536.0,1,-nbitq), 
to_sfixed(1830.0/65536.0,1,-nbitq), 
to_sfixed(4386.0/65536.0,1,-nbitq), 
to_sfixed(-2118.0/65536.0,1,-nbitq), 
to_sfixed(-6360.0/65536.0,1,-nbitq), 
to_sfixed(3185.0/65536.0,1,-nbitq), 
to_sfixed(-643.0/65536.0,1,-nbitq), 
to_sfixed(781.0/65536.0,1,-nbitq), 
to_sfixed(-1747.0/65536.0,1,-nbitq), 
to_sfixed(-5450.0/65536.0,1,-nbitq), 
to_sfixed(-2535.0/65536.0,1,-nbitq), 
to_sfixed(373.0/65536.0,1,-nbitq), 
to_sfixed(-2375.0/65536.0,1,-nbitq), 
to_sfixed(260.0/65536.0,1,-nbitq), 
to_sfixed(5592.0/65536.0,1,-nbitq), 
to_sfixed(-248.0/65536.0,1,-nbitq), 
to_sfixed(1145.0/65536.0,1,-nbitq), 
to_sfixed(-1248.0/65536.0,1,-nbitq), 
to_sfixed(966.0/65536.0,1,-nbitq), 
to_sfixed(2529.0/65536.0,1,-nbitq), 
to_sfixed(323.0/65536.0,1,-nbitq), 
to_sfixed(-3542.0/65536.0,1,-nbitq), 
to_sfixed(2785.0/65536.0,1,-nbitq), 
to_sfixed(-2392.0/65536.0,1,-nbitq), 
to_sfixed(-5608.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-741.0/65536.0,1,-nbitq), 
to_sfixed(-2136.0/65536.0,1,-nbitq), 
to_sfixed(5352.0/65536.0,1,-nbitq), 
to_sfixed(2216.0/65536.0,1,-nbitq), 
to_sfixed(-5507.0/65536.0,1,-nbitq), 
to_sfixed(-7817.0/65536.0,1,-nbitq), 
to_sfixed(-1278.0/65536.0,1,-nbitq), 
to_sfixed(-233.0/65536.0,1,-nbitq), 
to_sfixed(3880.0/65536.0,1,-nbitq), 
to_sfixed(830.0/65536.0,1,-nbitq), 
to_sfixed(-2656.0/65536.0,1,-nbitq), 
to_sfixed(-5696.0/65536.0,1,-nbitq), 
to_sfixed(-189.0/65536.0,1,-nbitq), 
to_sfixed(-8145.0/65536.0,1,-nbitq), 
to_sfixed(4188.0/65536.0,1,-nbitq), 
to_sfixed(611.0/65536.0,1,-nbitq), 
to_sfixed(-1091.0/65536.0,1,-nbitq), 
to_sfixed(77.0/65536.0,1,-nbitq), 
to_sfixed(-1204.0/65536.0,1,-nbitq), 
to_sfixed(-2054.0/65536.0,1,-nbitq), 
to_sfixed(1357.0/65536.0,1,-nbitq), 
to_sfixed(3805.0/65536.0,1,-nbitq), 
to_sfixed(4872.0/65536.0,1,-nbitq), 
to_sfixed(-9732.0/65536.0,1,-nbitq), 
to_sfixed(52.0/65536.0,1,-nbitq), 
to_sfixed(1112.0/65536.0,1,-nbitq), 
to_sfixed(-6365.0/65536.0,1,-nbitq), 
to_sfixed(1094.0/65536.0,1,-nbitq), 
to_sfixed(-705.0/65536.0,1,-nbitq), 
to_sfixed(2003.0/65536.0,1,-nbitq), 
to_sfixed(-5176.0/65536.0,1,-nbitq), 
to_sfixed(1487.0/65536.0,1,-nbitq), 
to_sfixed(1586.0/65536.0,1,-nbitq), 
to_sfixed(2136.0/65536.0,1,-nbitq), 
to_sfixed(1743.0/65536.0,1,-nbitq), 
to_sfixed(-1035.0/65536.0,1,-nbitq), 
to_sfixed(2361.0/65536.0,1,-nbitq), 
to_sfixed(-135.0/65536.0,1,-nbitq), 
to_sfixed(-2568.0/65536.0,1,-nbitq), 
to_sfixed(3838.0/65536.0,1,-nbitq), 
to_sfixed(740.0/65536.0,1,-nbitq), 
to_sfixed(-622.0/65536.0,1,-nbitq), 
to_sfixed(4473.0/65536.0,1,-nbitq), 
to_sfixed(-1567.0/65536.0,1,-nbitq), 
to_sfixed(317.0/65536.0,1,-nbitq), 
to_sfixed(2184.0/65536.0,1,-nbitq), 
to_sfixed(1374.0/65536.0,1,-nbitq), 
to_sfixed(-2661.0/65536.0,1,-nbitq), 
to_sfixed(139.0/65536.0,1,-nbitq), 
to_sfixed(4133.0/65536.0,1,-nbitq), 
to_sfixed(-1559.0/65536.0,1,-nbitq), 
to_sfixed(3712.0/65536.0,1,-nbitq), 
to_sfixed(-906.0/65536.0,1,-nbitq), 
to_sfixed(7970.0/65536.0,1,-nbitq), 
to_sfixed(-3517.0/65536.0,1,-nbitq), 
to_sfixed(6505.0/65536.0,1,-nbitq), 
to_sfixed(1403.0/65536.0,1,-nbitq), 
to_sfixed(2785.0/65536.0,1,-nbitq), 
to_sfixed(-3018.0/65536.0,1,-nbitq), 
to_sfixed(-4891.0/65536.0,1,-nbitq), 
to_sfixed(4634.0/65536.0,1,-nbitq), 
to_sfixed(-1845.0/65536.0,1,-nbitq), 
to_sfixed(2645.0/65536.0,1,-nbitq), 
to_sfixed(-2536.0/65536.0,1,-nbitq), 
to_sfixed(-53.0/65536.0,1,-nbitq), 
to_sfixed(2760.0/65536.0,1,-nbitq), 
to_sfixed(538.0/65536.0,1,-nbitq), 
to_sfixed(2757.0/65536.0,1,-nbitq), 
to_sfixed(6205.0/65536.0,1,-nbitq), 
to_sfixed(4549.0/65536.0,1,-nbitq), 
to_sfixed(-1225.0/65536.0,1,-nbitq), 
to_sfixed(3390.0/65536.0,1,-nbitq), 
to_sfixed(2229.0/65536.0,1,-nbitq), 
to_sfixed(-665.0/65536.0,1,-nbitq), 
to_sfixed(-2814.0/65536.0,1,-nbitq), 
to_sfixed(2940.0/65536.0,1,-nbitq), 
to_sfixed(-939.0/65536.0,1,-nbitq), 
to_sfixed(2815.0/65536.0,1,-nbitq), 
to_sfixed(-1008.0/65536.0,1,-nbitq), 
to_sfixed(-979.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2908.0/65536.0,1,-nbitq), 
to_sfixed(1608.0/65536.0,1,-nbitq), 
to_sfixed(3302.0/65536.0,1,-nbitq), 
to_sfixed(-1501.0/65536.0,1,-nbitq), 
to_sfixed(-79.0/65536.0,1,-nbitq), 
to_sfixed(-2925.0/65536.0,1,-nbitq), 
to_sfixed(-979.0/65536.0,1,-nbitq), 
to_sfixed(-1026.0/65536.0,1,-nbitq), 
to_sfixed(1168.0/65536.0,1,-nbitq), 
to_sfixed(2281.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(-4332.0/65536.0,1,-nbitq), 
to_sfixed(3837.0/65536.0,1,-nbitq), 
to_sfixed(-8394.0/65536.0,1,-nbitq), 
to_sfixed(2488.0/65536.0,1,-nbitq), 
to_sfixed(-875.0/65536.0,1,-nbitq), 
to_sfixed(2283.0/65536.0,1,-nbitq), 
to_sfixed(-5759.0/65536.0,1,-nbitq), 
to_sfixed(-1640.0/65536.0,1,-nbitq), 
to_sfixed(-2294.0/65536.0,1,-nbitq), 
to_sfixed(612.0/65536.0,1,-nbitq), 
to_sfixed(3955.0/65536.0,1,-nbitq), 
to_sfixed(-2280.0/65536.0,1,-nbitq), 
to_sfixed(-8499.0/65536.0,1,-nbitq), 
to_sfixed(1335.0/65536.0,1,-nbitq), 
to_sfixed(1350.0/65536.0,1,-nbitq), 
to_sfixed(-8250.0/65536.0,1,-nbitq), 
to_sfixed(-3456.0/65536.0,1,-nbitq), 
to_sfixed(529.0/65536.0,1,-nbitq), 
to_sfixed(2902.0/65536.0,1,-nbitq), 
to_sfixed(-5207.0/65536.0,1,-nbitq), 
to_sfixed(-657.0/65536.0,1,-nbitq), 
to_sfixed(5093.0/65536.0,1,-nbitq), 
to_sfixed(3460.0/65536.0,1,-nbitq), 
to_sfixed(236.0/65536.0,1,-nbitq), 
to_sfixed(-1267.0/65536.0,1,-nbitq), 
to_sfixed(1268.0/65536.0,1,-nbitq), 
to_sfixed(116.0/65536.0,1,-nbitq), 
to_sfixed(-254.0/65536.0,1,-nbitq), 
to_sfixed(-1712.0/65536.0,1,-nbitq), 
to_sfixed(4228.0/65536.0,1,-nbitq), 
to_sfixed(2166.0/65536.0,1,-nbitq), 
to_sfixed(4323.0/65536.0,1,-nbitq), 
to_sfixed(-1578.0/65536.0,1,-nbitq), 
to_sfixed(1741.0/65536.0,1,-nbitq), 
to_sfixed(1339.0/65536.0,1,-nbitq), 
to_sfixed(-2284.0/65536.0,1,-nbitq), 
to_sfixed(2369.0/65536.0,1,-nbitq), 
to_sfixed(1989.0/65536.0,1,-nbitq), 
to_sfixed(-928.0/65536.0,1,-nbitq), 
to_sfixed(1816.0/65536.0,1,-nbitq), 
to_sfixed(369.0/65536.0,1,-nbitq), 
to_sfixed(-4718.0/65536.0,1,-nbitq), 
to_sfixed(8436.0/65536.0,1,-nbitq), 
to_sfixed(-5825.0/65536.0,1,-nbitq), 
to_sfixed(7270.0/65536.0,1,-nbitq), 
to_sfixed(-2822.0/65536.0,1,-nbitq), 
to_sfixed(5299.0/65536.0,1,-nbitq), 
to_sfixed(2905.0/65536.0,1,-nbitq), 
to_sfixed(-3300.0/65536.0,1,-nbitq), 
to_sfixed(2878.0/65536.0,1,-nbitq), 
to_sfixed(1473.0/65536.0,1,-nbitq), 
to_sfixed(-1912.0/65536.0,1,-nbitq), 
to_sfixed(2154.0/65536.0,1,-nbitq), 
to_sfixed(986.0/65536.0,1,-nbitq), 
to_sfixed(2941.0/65536.0,1,-nbitq), 
to_sfixed(-718.0/65536.0,1,-nbitq), 
to_sfixed(2822.0/65536.0,1,-nbitq), 
to_sfixed(7700.0/65536.0,1,-nbitq), 
to_sfixed(3282.0/65536.0,1,-nbitq), 
to_sfixed(668.0/65536.0,1,-nbitq), 
to_sfixed(-3604.0/65536.0,1,-nbitq), 
to_sfixed(4837.0/65536.0,1,-nbitq), 
to_sfixed(111.0/65536.0,1,-nbitq), 
to_sfixed(1906.0/65536.0,1,-nbitq), 
to_sfixed(4680.0/65536.0,1,-nbitq), 
to_sfixed(-2516.0/65536.0,1,-nbitq), 
to_sfixed(2935.0/65536.0,1,-nbitq), 
to_sfixed(2319.0/65536.0,1,-nbitq), 
to_sfixed(-1545.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1962.0/65536.0,1,-nbitq), 
to_sfixed(2605.0/65536.0,1,-nbitq), 
to_sfixed(2733.0/65536.0,1,-nbitq), 
to_sfixed(-3478.0/65536.0,1,-nbitq), 
to_sfixed(-2049.0/65536.0,1,-nbitq), 
to_sfixed(-785.0/65536.0,1,-nbitq), 
to_sfixed(-2728.0/65536.0,1,-nbitq), 
to_sfixed(3907.0/65536.0,1,-nbitq), 
to_sfixed(386.0/65536.0,1,-nbitq), 
to_sfixed(-2381.0/65536.0,1,-nbitq), 
to_sfixed(808.0/65536.0,1,-nbitq), 
to_sfixed(-1163.0/65536.0,1,-nbitq), 
to_sfixed(2860.0/65536.0,1,-nbitq), 
to_sfixed(-7783.0/65536.0,1,-nbitq), 
to_sfixed(-190.0/65536.0,1,-nbitq), 
to_sfixed(-255.0/65536.0,1,-nbitq), 
to_sfixed(-656.0/65536.0,1,-nbitq), 
to_sfixed(-3432.0/65536.0,1,-nbitq), 
to_sfixed(-3415.0/65536.0,1,-nbitq), 
to_sfixed(706.0/65536.0,1,-nbitq), 
to_sfixed(4170.0/65536.0,1,-nbitq), 
to_sfixed(5111.0/65536.0,1,-nbitq), 
to_sfixed(-5914.0/65536.0,1,-nbitq), 
to_sfixed(-7790.0/65536.0,1,-nbitq), 
to_sfixed(2126.0/65536.0,1,-nbitq), 
to_sfixed(-2966.0/65536.0,1,-nbitq), 
to_sfixed(-3018.0/65536.0,1,-nbitq), 
to_sfixed(937.0/65536.0,1,-nbitq), 
to_sfixed(1027.0/65536.0,1,-nbitq), 
to_sfixed(2269.0/65536.0,1,-nbitq), 
to_sfixed(-3760.0/65536.0,1,-nbitq), 
to_sfixed(1930.0/65536.0,1,-nbitq), 
to_sfixed(2654.0/65536.0,1,-nbitq), 
to_sfixed(5137.0/65536.0,1,-nbitq), 
to_sfixed(-1513.0/65536.0,1,-nbitq), 
to_sfixed(2480.0/65536.0,1,-nbitq), 
to_sfixed(2443.0/65536.0,1,-nbitq), 
to_sfixed(-2704.0/65536.0,1,-nbitq), 
to_sfixed(-1470.0/65536.0,1,-nbitq), 
to_sfixed(-1231.0/65536.0,1,-nbitq), 
to_sfixed(878.0/65536.0,1,-nbitq), 
to_sfixed(17.0/65536.0,1,-nbitq), 
to_sfixed(1022.0/65536.0,1,-nbitq), 
to_sfixed(1641.0/65536.0,1,-nbitq), 
to_sfixed(1810.0/65536.0,1,-nbitq), 
to_sfixed(3759.0/65536.0,1,-nbitq), 
to_sfixed(-663.0/65536.0,1,-nbitq), 
to_sfixed(-538.0/65536.0,1,-nbitq), 
to_sfixed(2937.0/65536.0,1,-nbitq), 
to_sfixed(-983.0/65536.0,1,-nbitq), 
to_sfixed(709.0/65536.0,1,-nbitq), 
to_sfixed(-1283.0/65536.0,1,-nbitq), 
to_sfixed(2047.0/65536.0,1,-nbitq), 
to_sfixed(5732.0/65536.0,1,-nbitq), 
to_sfixed(-2435.0/65536.0,1,-nbitq), 
to_sfixed(4614.0/65536.0,1,-nbitq), 
to_sfixed(1445.0/65536.0,1,-nbitq), 
to_sfixed(2476.0/65536.0,1,-nbitq), 
to_sfixed(-2441.0/65536.0,1,-nbitq), 
to_sfixed(-4112.0/65536.0,1,-nbitq), 
to_sfixed(-160.0/65536.0,1,-nbitq), 
to_sfixed(-436.0/65536.0,1,-nbitq), 
to_sfixed(-1746.0/65536.0,1,-nbitq), 
to_sfixed(-2933.0/65536.0,1,-nbitq), 
to_sfixed(736.0/65536.0,1,-nbitq), 
to_sfixed(-1290.0/65536.0,1,-nbitq), 
to_sfixed(1285.0/65536.0,1,-nbitq), 
to_sfixed(1498.0/65536.0,1,-nbitq), 
to_sfixed(7999.0/65536.0,1,-nbitq), 
to_sfixed(684.0/65536.0,1,-nbitq), 
to_sfixed(471.0/65536.0,1,-nbitq), 
to_sfixed(886.0/65536.0,1,-nbitq), 
to_sfixed(2307.0/65536.0,1,-nbitq), 
to_sfixed(2572.0/65536.0,1,-nbitq), 
to_sfixed(-191.0/65536.0,1,-nbitq), 
to_sfixed(4872.0/65536.0,1,-nbitq), 
to_sfixed(-5102.0/65536.0,1,-nbitq), 
to_sfixed(-472.0/65536.0,1,-nbitq), 
to_sfixed(-985.0/65536.0,1,-nbitq), 
to_sfixed(2189.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1509.0/65536.0,1,-nbitq), 
to_sfixed(2816.0/65536.0,1,-nbitq), 
to_sfixed(-3324.0/65536.0,1,-nbitq), 
to_sfixed(-1230.0/65536.0,1,-nbitq), 
to_sfixed(-2702.0/65536.0,1,-nbitq), 
to_sfixed(328.0/65536.0,1,-nbitq), 
to_sfixed(1149.0/65536.0,1,-nbitq), 
to_sfixed(-301.0/65536.0,1,-nbitq), 
to_sfixed(925.0/65536.0,1,-nbitq), 
to_sfixed(-1678.0/65536.0,1,-nbitq), 
to_sfixed(1339.0/65536.0,1,-nbitq), 
to_sfixed(-530.0/65536.0,1,-nbitq), 
to_sfixed(-491.0/65536.0,1,-nbitq), 
to_sfixed(-6420.0/65536.0,1,-nbitq), 
to_sfixed(-503.0/65536.0,1,-nbitq), 
to_sfixed(-993.0/65536.0,1,-nbitq), 
to_sfixed(772.0/65536.0,1,-nbitq), 
to_sfixed(1859.0/65536.0,1,-nbitq), 
to_sfixed(331.0/65536.0,1,-nbitq), 
to_sfixed(-980.0/65536.0,1,-nbitq), 
to_sfixed(1856.0/65536.0,1,-nbitq), 
to_sfixed(1056.0/65536.0,1,-nbitq), 
to_sfixed(-3548.0/65536.0,1,-nbitq), 
to_sfixed(-1978.0/65536.0,1,-nbitq), 
to_sfixed(-1915.0/65536.0,1,-nbitq), 
to_sfixed(-748.0/65536.0,1,-nbitq), 
to_sfixed(-3381.0/65536.0,1,-nbitq), 
to_sfixed(-478.0/65536.0,1,-nbitq), 
to_sfixed(358.0/65536.0,1,-nbitq), 
to_sfixed(-2849.0/65536.0,1,-nbitq), 
to_sfixed(-2502.0/65536.0,1,-nbitq), 
to_sfixed(630.0/65536.0,1,-nbitq), 
to_sfixed(-1515.0/65536.0,1,-nbitq), 
to_sfixed(4064.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(-453.0/65536.0,1,-nbitq), 
to_sfixed(-521.0/65536.0,1,-nbitq), 
to_sfixed(1223.0/65536.0,1,-nbitq), 
to_sfixed(-3223.0/65536.0,1,-nbitq), 
to_sfixed(-217.0/65536.0,1,-nbitq), 
to_sfixed(2579.0/65536.0,1,-nbitq), 
to_sfixed(-2576.0/65536.0,1,-nbitq), 
to_sfixed(-3819.0/65536.0,1,-nbitq), 
to_sfixed(1010.0/65536.0,1,-nbitq), 
to_sfixed(-839.0/65536.0,1,-nbitq), 
to_sfixed(5334.0/65536.0,1,-nbitq), 
to_sfixed(-2356.0/65536.0,1,-nbitq), 
to_sfixed(277.0/65536.0,1,-nbitq), 
to_sfixed(1059.0/65536.0,1,-nbitq), 
to_sfixed(1628.0/65536.0,1,-nbitq), 
to_sfixed(163.0/65536.0,1,-nbitq), 
to_sfixed(-3406.0/65536.0,1,-nbitq), 
to_sfixed(-1790.0/65536.0,1,-nbitq), 
to_sfixed(4186.0/65536.0,1,-nbitq), 
to_sfixed(3122.0/65536.0,1,-nbitq), 
to_sfixed(-40.0/65536.0,1,-nbitq), 
to_sfixed(1002.0/65536.0,1,-nbitq), 
to_sfixed(2180.0/65536.0,1,-nbitq), 
to_sfixed(2731.0/65536.0,1,-nbitq), 
to_sfixed(-279.0/65536.0,1,-nbitq), 
to_sfixed(-178.0/65536.0,1,-nbitq), 
to_sfixed(-2366.0/65536.0,1,-nbitq), 
to_sfixed(-2380.0/65536.0,1,-nbitq), 
to_sfixed(-132.0/65536.0,1,-nbitq), 
to_sfixed(1046.0/65536.0,1,-nbitq), 
to_sfixed(1720.0/65536.0,1,-nbitq), 
to_sfixed(2701.0/65536.0,1,-nbitq), 
to_sfixed(-1964.0/65536.0,1,-nbitq), 
to_sfixed(3713.0/65536.0,1,-nbitq), 
to_sfixed(-359.0/65536.0,1,-nbitq), 
to_sfixed(-2298.0/65536.0,1,-nbitq), 
to_sfixed(-3309.0/65536.0,1,-nbitq), 
to_sfixed(-1114.0/65536.0,1,-nbitq), 
to_sfixed(-2014.0/65536.0,1,-nbitq), 
to_sfixed(-847.0/65536.0,1,-nbitq), 
to_sfixed(-77.0/65536.0,1,-nbitq), 
to_sfixed(-5513.0/65536.0,1,-nbitq), 
to_sfixed(3023.0/65536.0,1,-nbitq), 
to_sfixed(-2349.0/65536.0,1,-nbitq), 
to_sfixed(2641.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1641.0/65536.0,1,-nbitq), 
to_sfixed(-431.0/65536.0,1,-nbitq), 
to_sfixed(-196.0/65536.0,1,-nbitq), 
to_sfixed(-719.0/65536.0,1,-nbitq), 
to_sfixed(85.0/65536.0,1,-nbitq), 
to_sfixed(-1366.0/65536.0,1,-nbitq), 
to_sfixed(-2659.0/65536.0,1,-nbitq), 
to_sfixed(-1030.0/65536.0,1,-nbitq), 
to_sfixed(-2712.0/65536.0,1,-nbitq), 
to_sfixed(-748.0/65536.0,1,-nbitq), 
to_sfixed(-1732.0/65536.0,1,-nbitq), 
to_sfixed(-177.0/65536.0,1,-nbitq), 
to_sfixed(-2192.0/65536.0,1,-nbitq), 
to_sfixed(-258.0/65536.0,1,-nbitq), 
to_sfixed(-1155.0/65536.0,1,-nbitq), 
to_sfixed(1066.0/65536.0,1,-nbitq), 
to_sfixed(-597.0/65536.0,1,-nbitq), 
to_sfixed(2760.0/65536.0,1,-nbitq), 
to_sfixed(-434.0/65536.0,1,-nbitq), 
to_sfixed(-1409.0/65536.0,1,-nbitq), 
to_sfixed(-3310.0/65536.0,1,-nbitq), 
to_sfixed(4002.0/65536.0,1,-nbitq), 
to_sfixed(1894.0/65536.0,1,-nbitq), 
to_sfixed(2200.0/65536.0,1,-nbitq), 
to_sfixed(-273.0/65536.0,1,-nbitq), 
to_sfixed(-1802.0/65536.0,1,-nbitq), 
to_sfixed(-1754.0/65536.0,1,-nbitq), 
to_sfixed(1599.0/65536.0,1,-nbitq), 
to_sfixed(2205.0/65536.0,1,-nbitq), 
to_sfixed(1058.0/65536.0,1,-nbitq), 
to_sfixed(2476.0/65536.0,1,-nbitq), 
to_sfixed(-2209.0/65536.0,1,-nbitq), 
to_sfixed(-4238.0/65536.0,1,-nbitq), 
to_sfixed(-3056.0/65536.0,1,-nbitq), 
to_sfixed(-1536.0/65536.0,1,-nbitq), 
to_sfixed(1075.0/65536.0,1,-nbitq), 
to_sfixed(-2968.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(-3519.0/65536.0,1,-nbitq), 
to_sfixed(591.0/65536.0,1,-nbitq), 
to_sfixed(-1076.0/65536.0,1,-nbitq), 
to_sfixed(2043.0/65536.0,1,-nbitq), 
to_sfixed(-4943.0/65536.0,1,-nbitq), 
to_sfixed(441.0/65536.0,1,-nbitq), 
to_sfixed(-1664.0/65536.0,1,-nbitq), 
to_sfixed(22.0/65536.0,1,-nbitq), 
to_sfixed(2416.0/65536.0,1,-nbitq), 
to_sfixed(-84.0/65536.0,1,-nbitq), 
to_sfixed(863.0/65536.0,1,-nbitq), 
to_sfixed(-767.0/65536.0,1,-nbitq), 
to_sfixed(927.0/65536.0,1,-nbitq), 
to_sfixed(-606.0/65536.0,1,-nbitq), 
to_sfixed(688.0/65536.0,1,-nbitq), 
to_sfixed(-2465.0/65536.0,1,-nbitq), 
to_sfixed(-1586.0/65536.0,1,-nbitq), 
to_sfixed(-617.0/65536.0,1,-nbitq), 
to_sfixed(2051.0/65536.0,1,-nbitq), 
to_sfixed(1612.0/65536.0,1,-nbitq), 
to_sfixed(162.0/65536.0,1,-nbitq), 
to_sfixed(216.0/65536.0,1,-nbitq), 
to_sfixed(-206.0/65536.0,1,-nbitq), 
to_sfixed(-2858.0/65536.0,1,-nbitq), 
to_sfixed(1502.0/65536.0,1,-nbitq), 
to_sfixed(-866.0/65536.0,1,-nbitq), 
to_sfixed(602.0/65536.0,1,-nbitq), 
to_sfixed(3221.0/65536.0,1,-nbitq), 
to_sfixed(2212.0/65536.0,1,-nbitq), 
to_sfixed(2434.0/65536.0,1,-nbitq), 
to_sfixed(3073.0/65536.0,1,-nbitq), 
to_sfixed(-30.0/65536.0,1,-nbitq), 
to_sfixed(-309.0/65536.0,1,-nbitq), 
to_sfixed(100.0/65536.0,1,-nbitq), 
to_sfixed(-206.0/65536.0,1,-nbitq), 
to_sfixed(-665.0/65536.0,1,-nbitq), 
to_sfixed(-2308.0/65536.0,1,-nbitq), 
to_sfixed(1379.0/65536.0,1,-nbitq), 
to_sfixed(-1627.0/65536.0,1,-nbitq), 
to_sfixed(-533.0/65536.0,1,-nbitq), 
to_sfixed(-990.0/65536.0,1,-nbitq), 
to_sfixed(-476.0/65536.0,1,-nbitq)  ), 
( to_sfixed(259.0/65536.0,1,-nbitq), 
to_sfixed(-1886.0/65536.0,1,-nbitq), 
to_sfixed(1996.0/65536.0,1,-nbitq), 
to_sfixed(-1546.0/65536.0,1,-nbitq), 
to_sfixed(216.0/65536.0,1,-nbitq), 
to_sfixed(125.0/65536.0,1,-nbitq), 
to_sfixed(-2738.0/65536.0,1,-nbitq), 
to_sfixed(-220.0/65536.0,1,-nbitq), 
to_sfixed(-2683.0/65536.0,1,-nbitq), 
to_sfixed(-2255.0/65536.0,1,-nbitq), 
to_sfixed(-935.0/65536.0,1,-nbitq), 
to_sfixed(-3076.0/65536.0,1,-nbitq), 
to_sfixed(1165.0/65536.0,1,-nbitq), 
to_sfixed(-3870.0/65536.0,1,-nbitq), 
to_sfixed(-1481.0/65536.0,1,-nbitq), 
to_sfixed(2323.0/65536.0,1,-nbitq), 
to_sfixed(1898.0/65536.0,1,-nbitq), 
to_sfixed(-166.0/65536.0,1,-nbitq), 
to_sfixed(1238.0/65536.0,1,-nbitq), 
to_sfixed(691.0/65536.0,1,-nbitq), 
to_sfixed(-3093.0/65536.0,1,-nbitq), 
to_sfixed(2759.0/65536.0,1,-nbitq), 
to_sfixed(-1442.0/65536.0,1,-nbitq), 
to_sfixed(4283.0/65536.0,1,-nbitq), 
to_sfixed(1033.0/65536.0,1,-nbitq), 
to_sfixed(1745.0/65536.0,1,-nbitq), 
to_sfixed(-755.0/65536.0,1,-nbitq), 
to_sfixed(1836.0/65536.0,1,-nbitq), 
to_sfixed(-2198.0/65536.0,1,-nbitq), 
to_sfixed(-3037.0/65536.0,1,-nbitq), 
to_sfixed(-985.0/65536.0,1,-nbitq), 
to_sfixed(-2592.0/65536.0,1,-nbitq), 
to_sfixed(-3387.0/65536.0,1,-nbitq), 
to_sfixed(-43.0/65536.0,1,-nbitq), 
to_sfixed(637.0/65536.0,1,-nbitq), 
to_sfixed(150.0/65536.0,1,-nbitq), 
to_sfixed(-1137.0/65536.0,1,-nbitq), 
to_sfixed(-1498.0/65536.0,1,-nbitq), 
to_sfixed(-2017.0/65536.0,1,-nbitq), 
to_sfixed(2592.0/65536.0,1,-nbitq), 
to_sfixed(-1403.0/65536.0,1,-nbitq), 
to_sfixed(812.0/65536.0,1,-nbitq), 
to_sfixed(-4899.0/65536.0,1,-nbitq), 
to_sfixed(-761.0/65536.0,1,-nbitq), 
to_sfixed(-2079.0/65536.0,1,-nbitq), 
to_sfixed(892.0/65536.0,1,-nbitq), 
to_sfixed(-1743.0/65536.0,1,-nbitq), 
to_sfixed(96.0/65536.0,1,-nbitq), 
to_sfixed(-1386.0/65536.0,1,-nbitq), 
to_sfixed(1826.0/65536.0,1,-nbitq), 
to_sfixed(1441.0/65536.0,1,-nbitq), 
to_sfixed(2494.0/65536.0,1,-nbitq), 
to_sfixed(1525.0/65536.0,1,-nbitq), 
to_sfixed(2901.0/65536.0,1,-nbitq), 
to_sfixed(-615.0/65536.0,1,-nbitq), 
to_sfixed(-1620.0/65536.0,1,-nbitq), 
to_sfixed(2664.0/65536.0,1,-nbitq), 
to_sfixed(2884.0/65536.0,1,-nbitq), 
to_sfixed(-901.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(-3446.0/65536.0,1,-nbitq), 
to_sfixed(-3086.0/65536.0,1,-nbitq), 
to_sfixed(2029.0/65536.0,1,-nbitq), 
to_sfixed(1575.0/65536.0,1,-nbitq), 
to_sfixed(3068.0/65536.0,1,-nbitq), 
to_sfixed(188.0/65536.0,1,-nbitq), 
to_sfixed(338.0/65536.0,1,-nbitq), 
to_sfixed(-130.0/65536.0,1,-nbitq), 
to_sfixed(1719.0/65536.0,1,-nbitq), 
to_sfixed(3070.0/65536.0,1,-nbitq), 
to_sfixed(956.0/65536.0,1,-nbitq), 
to_sfixed(2922.0/65536.0,1,-nbitq), 
to_sfixed(3940.0/65536.0,1,-nbitq), 
to_sfixed(2657.0/65536.0,1,-nbitq), 
to_sfixed(-1565.0/65536.0,1,-nbitq), 
to_sfixed(3871.0/65536.0,1,-nbitq), 
to_sfixed(-2949.0/65536.0,1,-nbitq), 
to_sfixed(4767.0/65536.0,1,-nbitq), 
to_sfixed(-2532.0/65536.0,1,-nbitq), 
to_sfixed(4629.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(384.0/65536.0,1,-nbitq), 
to_sfixed(146.0/65536.0,1,-nbitq), 
to_sfixed(1171.0/65536.0,1,-nbitq), 
to_sfixed(-832.0/65536.0,1,-nbitq), 
to_sfixed(411.0/65536.0,1,-nbitq), 
to_sfixed(-2488.0/65536.0,1,-nbitq), 
to_sfixed(-108.0/65536.0,1,-nbitq), 
to_sfixed(-1675.0/65536.0,1,-nbitq), 
to_sfixed(-95.0/65536.0,1,-nbitq), 
to_sfixed(879.0/65536.0,1,-nbitq), 
to_sfixed(-917.0/65536.0,1,-nbitq), 
to_sfixed(-2944.0/65536.0,1,-nbitq), 
to_sfixed(1800.0/65536.0,1,-nbitq), 
to_sfixed(1202.0/65536.0,1,-nbitq), 
to_sfixed(-1557.0/65536.0,1,-nbitq), 
to_sfixed(-1888.0/65536.0,1,-nbitq), 
to_sfixed(2069.0/65536.0,1,-nbitq), 
to_sfixed(-64.0/65536.0,1,-nbitq), 
to_sfixed(-162.0/65536.0,1,-nbitq), 
to_sfixed(2658.0/65536.0,1,-nbitq), 
to_sfixed(489.0/65536.0,1,-nbitq), 
to_sfixed(-1452.0/65536.0,1,-nbitq), 
to_sfixed(2497.0/65536.0,1,-nbitq), 
to_sfixed(395.0/65536.0,1,-nbitq), 
to_sfixed(1713.0/65536.0,1,-nbitq), 
to_sfixed(1477.0/65536.0,1,-nbitq), 
to_sfixed(-2809.0/65536.0,1,-nbitq), 
to_sfixed(-1892.0/65536.0,1,-nbitq), 
to_sfixed(-4775.0/65536.0,1,-nbitq), 
to_sfixed(-2739.0/65536.0,1,-nbitq), 
to_sfixed(1304.0/65536.0,1,-nbitq), 
to_sfixed(-101.0/65536.0,1,-nbitq), 
to_sfixed(-2810.0/65536.0,1,-nbitq), 
to_sfixed(2272.0/65536.0,1,-nbitq), 
to_sfixed(-1716.0/65536.0,1,-nbitq), 
to_sfixed(-2493.0/65536.0,1,-nbitq), 
to_sfixed(-278.0/65536.0,1,-nbitq), 
to_sfixed(-2511.0/65536.0,1,-nbitq), 
to_sfixed(-3717.0/65536.0,1,-nbitq), 
to_sfixed(-683.0/65536.0,1,-nbitq), 
to_sfixed(-4254.0/65536.0,1,-nbitq), 
to_sfixed(-2254.0/65536.0,1,-nbitq), 
to_sfixed(-3443.0/65536.0,1,-nbitq), 
to_sfixed(4335.0/65536.0,1,-nbitq), 
to_sfixed(2505.0/65536.0,1,-nbitq), 
to_sfixed(3496.0/65536.0,1,-nbitq), 
to_sfixed(656.0/65536.0,1,-nbitq), 
to_sfixed(-617.0/65536.0,1,-nbitq), 
to_sfixed(-955.0/65536.0,1,-nbitq), 
to_sfixed(-1181.0/65536.0,1,-nbitq), 
to_sfixed(2272.0/65536.0,1,-nbitq), 
to_sfixed(1555.0/65536.0,1,-nbitq), 
to_sfixed(1865.0/65536.0,1,-nbitq), 
to_sfixed(-2177.0/65536.0,1,-nbitq), 
to_sfixed(2990.0/65536.0,1,-nbitq), 
to_sfixed(286.0/65536.0,1,-nbitq), 
to_sfixed(-2120.0/65536.0,1,-nbitq), 
to_sfixed(2985.0/65536.0,1,-nbitq), 
to_sfixed(-1960.0/65536.0,1,-nbitq), 
to_sfixed(1645.0/65536.0,1,-nbitq), 
to_sfixed(-2958.0/65536.0,1,-nbitq), 
to_sfixed(1996.0/65536.0,1,-nbitq), 
to_sfixed(-1886.0/65536.0,1,-nbitq), 
to_sfixed(954.0/65536.0,1,-nbitq), 
to_sfixed(1544.0/65536.0,1,-nbitq), 
to_sfixed(2420.0/65536.0,1,-nbitq), 
to_sfixed(2070.0/65536.0,1,-nbitq), 
to_sfixed(1057.0/65536.0,1,-nbitq), 
to_sfixed(2938.0/65536.0,1,-nbitq), 
to_sfixed(-107.0/65536.0,1,-nbitq), 
to_sfixed(3029.0/65536.0,1,-nbitq), 
to_sfixed(419.0/65536.0,1,-nbitq), 
to_sfixed(3638.0/65536.0,1,-nbitq), 
to_sfixed(2418.0/65536.0,1,-nbitq), 
to_sfixed(1646.0/65536.0,1,-nbitq), 
to_sfixed(1252.0/65536.0,1,-nbitq), 
to_sfixed(1758.0/65536.0,1,-nbitq), 
to_sfixed(3162.0/65536.0,1,-nbitq), 
to_sfixed(469.0/65536.0,1,-nbitq), 
to_sfixed(326.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-330.0/65536.0,1,-nbitq), 
to_sfixed(-485.0/65536.0,1,-nbitq), 
to_sfixed(4173.0/65536.0,1,-nbitq), 
to_sfixed(-452.0/65536.0,1,-nbitq), 
to_sfixed(-2694.0/65536.0,1,-nbitq), 
to_sfixed(-5319.0/65536.0,1,-nbitq), 
to_sfixed(228.0/65536.0,1,-nbitq), 
to_sfixed(-1563.0/65536.0,1,-nbitq), 
to_sfixed(1025.0/65536.0,1,-nbitq), 
to_sfixed(1468.0/65536.0,1,-nbitq), 
to_sfixed(70.0/65536.0,1,-nbitq), 
to_sfixed(115.0/65536.0,1,-nbitq), 
to_sfixed(1638.0/65536.0,1,-nbitq), 
to_sfixed(-892.0/65536.0,1,-nbitq), 
to_sfixed(-3668.0/65536.0,1,-nbitq), 
to_sfixed(1589.0/65536.0,1,-nbitq), 
to_sfixed(1182.0/65536.0,1,-nbitq), 
to_sfixed(-1384.0/65536.0,1,-nbitq), 
to_sfixed(3281.0/65536.0,1,-nbitq), 
to_sfixed(-2118.0/65536.0,1,-nbitq), 
to_sfixed(1389.0/65536.0,1,-nbitq), 
to_sfixed(2263.0/65536.0,1,-nbitq), 
to_sfixed(695.0/65536.0,1,-nbitq), 
to_sfixed(4148.0/65536.0,1,-nbitq), 
to_sfixed(-2604.0/65536.0,1,-nbitq), 
to_sfixed(-572.0/65536.0,1,-nbitq), 
to_sfixed(-4208.0/65536.0,1,-nbitq), 
to_sfixed(1622.0/65536.0,1,-nbitq), 
to_sfixed(-3049.0/65536.0,1,-nbitq), 
to_sfixed(852.0/65536.0,1,-nbitq), 
to_sfixed(199.0/65536.0,1,-nbitq), 
to_sfixed(-1230.0/65536.0,1,-nbitq), 
to_sfixed(207.0/65536.0,1,-nbitq), 
to_sfixed(1249.0/65536.0,1,-nbitq), 
to_sfixed(179.0/65536.0,1,-nbitq), 
to_sfixed(-2518.0/65536.0,1,-nbitq), 
to_sfixed(-2683.0/65536.0,1,-nbitq), 
to_sfixed(399.0/65536.0,1,-nbitq), 
to_sfixed(-866.0/65536.0,1,-nbitq), 
to_sfixed(3216.0/65536.0,1,-nbitq), 
to_sfixed(660.0/65536.0,1,-nbitq), 
to_sfixed(-884.0/65536.0,1,-nbitq), 
to_sfixed(-3713.0/65536.0,1,-nbitq), 
to_sfixed(1017.0/65536.0,1,-nbitq), 
to_sfixed(2668.0/65536.0,1,-nbitq), 
to_sfixed(2745.0/65536.0,1,-nbitq), 
to_sfixed(916.0/65536.0,1,-nbitq), 
to_sfixed(3553.0/65536.0,1,-nbitq), 
to_sfixed(-965.0/65536.0,1,-nbitq), 
to_sfixed(457.0/65536.0,1,-nbitq), 
to_sfixed(-889.0/65536.0,1,-nbitq), 
to_sfixed(3088.0/65536.0,1,-nbitq), 
to_sfixed(2219.0/65536.0,1,-nbitq), 
to_sfixed(2154.0/65536.0,1,-nbitq), 
to_sfixed(-898.0/65536.0,1,-nbitq), 
to_sfixed(1941.0/65536.0,1,-nbitq), 
to_sfixed(-654.0/65536.0,1,-nbitq), 
to_sfixed(928.0/65536.0,1,-nbitq), 
to_sfixed(-1340.0/65536.0,1,-nbitq), 
to_sfixed(4380.0/65536.0,1,-nbitq), 
to_sfixed(-2724.0/65536.0,1,-nbitq), 
to_sfixed(830.0/65536.0,1,-nbitq), 
to_sfixed(2183.0/65536.0,1,-nbitq), 
to_sfixed(-3185.0/65536.0,1,-nbitq), 
to_sfixed(2572.0/65536.0,1,-nbitq), 
to_sfixed(-1036.0/65536.0,1,-nbitq), 
to_sfixed(-2294.0/65536.0,1,-nbitq), 
to_sfixed(1098.0/65536.0,1,-nbitq), 
to_sfixed(375.0/65536.0,1,-nbitq), 
to_sfixed(5263.0/65536.0,1,-nbitq), 
to_sfixed(1387.0/65536.0,1,-nbitq), 
to_sfixed(1505.0/65536.0,1,-nbitq), 
to_sfixed(-790.0/65536.0,1,-nbitq), 
to_sfixed(-2664.0/65536.0,1,-nbitq), 
to_sfixed(2454.0/65536.0,1,-nbitq), 
to_sfixed(2178.0/65536.0,1,-nbitq), 
to_sfixed(-2413.0/65536.0,1,-nbitq), 
to_sfixed(-210.0/65536.0,1,-nbitq), 
to_sfixed(-2552.0/65536.0,1,-nbitq), 
to_sfixed(783.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1821.0/65536.0,1,-nbitq), 
to_sfixed(-3176.0/65536.0,1,-nbitq), 
to_sfixed(551.0/65536.0,1,-nbitq), 
to_sfixed(2200.0/65536.0,1,-nbitq), 
to_sfixed(5449.0/65536.0,1,-nbitq), 
to_sfixed(-1657.0/65536.0,1,-nbitq), 
to_sfixed(-3780.0/65536.0,1,-nbitq), 
to_sfixed(-906.0/65536.0,1,-nbitq), 
to_sfixed(-71.0/65536.0,1,-nbitq), 
to_sfixed(-348.0/65536.0,1,-nbitq), 
to_sfixed(2086.0/65536.0,1,-nbitq), 
to_sfixed(-4148.0/65536.0,1,-nbitq), 
to_sfixed(491.0/65536.0,1,-nbitq), 
to_sfixed(775.0/65536.0,1,-nbitq), 
to_sfixed(419.0/65536.0,1,-nbitq), 
to_sfixed(2660.0/65536.0,1,-nbitq), 
to_sfixed(-2971.0/65536.0,1,-nbitq), 
to_sfixed(3623.0/65536.0,1,-nbitq), 
to_sfixed(-3895.0/65536.0,1,-nbitq), 
to_sfixed(1678.0/65536.0,1,-nbitq), 
to_sfixed(1480.0/65536.0,1,-nbitq), 
to_sfixed(-2280.0/65536.0,1,-nbitq), 
to_sfixed(1605.0/65536.0,1,-nbitq), 
to_sfixed(-749.0/65536.0,1,-nbitq), 
to_sfixed(2402.0/65536.0,1,-nbitq), 
to_sfixed(-134.0/65536.0,1,-nbitq), 
to_sfixed(585.0/65536.0,1,-nbitq), 
to_sfixed(1595.0/65536.0,1,-nbitq), 
to_sfixed(-1713.0/65536.0,1,-nbitq), 
to_sfixed(-3999.0/65536.0,1,-nbitq), 
to_sfixed(-2138.0/65536.0,1,-nbitq), 
to_sfixed(1881.0/65536.0,1,-nbitq), 
to_sfixed(-824.0/65536.0,1,-nbitq), 
to_sfixed(3749.0/65536.0,1,-nbitq), 
to_sfixed(-1666.0/65536.0,1,-nbitq), 
to_sfixed(572.0/65536.0,1,-nbitq), 
to_sfixed(-1382.0/65536.0,1,-nbitq), 
to_sfixed(-308.0/65536.0,1,-nbitq), 
to_sfixed(-1014.0/65536.0,1,-nbitq), 
to_sfixed(-2326.0/65536.0,1,-nbitq), 
to_sfixed(-4590.0/65536.0,1,-nbitq), 
to_sfixed(-1245.0/65536.0,1,-nbitq), 
to_sfixed(-2866.0/65536.0,1,-nbitq), 
to_sfixed(-270.0/65536.0,1,-nbitq), 
to_sfixed(3279.0/65536.0,1,-nbitq), 
to_sfixed(3804.0/65536.0,1,-nbitq), 
to_sfixed(770.0/65536.0,1,-nbitq), 
to_sfixed(2055.0/65536.0,1,-nbitq), 
to_sfixed(-155.0/65536.0,1,-nbitq), 
to_sfixed(1192.0/65536.0,1,-nbitq), 
to_sfixed(2029.0/65536.0,1,-nbitq), 
to_sfixed(241.0/65536.0,1,-nbitq), 
to_sfixed(-2200.0/65536.0,1,-nbitq), 
to_sfixed(3506.0/65536.0,1,-nbitq), 
to_sfixed(-2381.0/65536.0,1,-nbitq), 
to_sfixed(1011.0/65536.0,1,-nbitq), 
to_sfixed(1532.0/65536.0,1,-nbitq), 
to_sfixed(-1282.0/65536.0,1,-nbitq), 
to_sfixed(1639.0/65536.0,1,-nbitq), 
to_sfixed(4262.0/65536.0,1,-nbitq), 
to_sfixed(-1735.0/65536.0,1,-nbitq), 
to_sfixed(-479.0/65536.0,1,-nbitq), 
to_sfixed(1936.0/65536.0,1,-nbitq), 
to_sfixed(-1729.0/65536.0,1,-nbitq), 
to_sfixed(708.0/65536.0,1,-nbitq), 
to_sfixed(3669.0/65536.0,1,-nbitq), 
to_sfixed(-148.0/65536.0,1,-nbitq), 
to_sfixed(4339.0/65536.0,1,-nbitq), 
to_sfixed(1642.0/65536.0,1,-nbitq), 
to_sfixed(2220.0/65536.0,1,-nbitq), 
to_sfixed(2234.0/65536.0,1,-nbitq), 
to_sfixed(-232.0/65536.0,1,-nbitq), 
to_sfixed(939.0/65536.0,1,-nbitq), 
to_sfixed(1797.0/65536.0,1,-nbitq), 
to_sfixed(-792.0/65536.0,1,-nbitq), 
to_sfixed(3168.0/65536.0,1,-nbitq), 
to_sfixed(-2801.0/65536.0,1,-nbitq), 
to_sfixed(-52.0/65536.0,1,-nbitq), 
to_sfixed(2011.0/65536.0,1,-nbitq), 
to_sfixed(3659.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1157.0/65536.0,1,-nbitq), 
to_sfixed(2141.0/65536.0,1,-nbitq), 
to_sfixed(-4238.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(6385.0/65536.0,1,-nbitq), 
to_sfixed(-2443.0/65536.0,1,-nbitq), 
to_sfixed(1059.0/65536.0,1,-nbitq), 
to_sfixed(-2368.0/65536.0,1,-nbitq), 
to_sfixed(-4471.0/65536.0,1,-nbitq), 
to_sfixed(1881.0/65536.0,1,-nbitq), 
to_sfixed(-83.0/65536.0,1,-nbitq), 
to_sfixed(134.0/65536.0,1,-nbitq), 
to_sfixed(-300.0/65536.0,1,-nbitq), 
to_sfixed(2435.0/65536.0,1,-nbitq), 
to_sfixed(-1191.0/65536.0,1,-nbitq), 
to_sfixed(1569.0/65536.0,1,-nbitq), 
to_sfixed(-1421.0/65536.0,1,-nbitq), 
to_sfixed(2196.0/65536.0,1,-nbitq), 
to_sfixed(502.0/65536.0,1,-nbitq), 
to_sfixed(2003.0/65536.0,1,-nbitq), 
to_sfixed(-304.0/65536.0,1,-nbitq), 
to_sfixed(944.0/65536.0,1,-nbitq), 
to_sfixed(-1123.0/65536.0,1,-nbitq), 
to_sfixed(-103.0/65536.0,1,-nbitq), 
to_sfixed(2847.0/65536.0,1,-nbitq), 
to_sfixed(1701.0/65536.0,1,-nbitq), 
to_sfixed(-4327.0/65536.0,1,-nbitq), 
to_sfixed(-1011.0/65536.0,1,-nbitq), 
to_sfixed(2336.0/65536.0,1,-nbitq), 
to_sfixed(-1234.0/65536.0,1,-nbitq), 
to_sfixed(-962.0/65536.0,1,-nbitq), 
to_sfixed(-5268.0/65536.0,1,-nbitq), 
to_sfixed(1484.0/65536.0,1,-nbitq), 
to_sfixed(-1712.0/65536.0,1,-nbitq), 
to_sfixed(1162.0/65536.0,1,-nbitq), 
to_sfixed(1588.0/65536.0,1,-nbitq), 
to_sfixed(-6707.0/65536.0,1,-nbitq), 
to_sfixed(3494.0/65536.0,1,-nbitq), 
to_sfixed(-3059.0/65536.0,1,-nbitq), 
to_sfixed(-853.0/65536.0,1,-nbitq), 
to_sfixed(-2434.0/65536.0,1,-nbitq), 
to_sfixed(909.0/65536.0,1,-nbitq), 
to_sfixed(1117.0/65536.0,1,-nbitq), 
to_sfixed(2538.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(4678.0/65536.0,1,-nbitq), 
to_sfixed(-2511.0/65536.0,1,-nbitq), 
to_sfixed(-2087.0/65536.0,1,-nbitq), 
to_sfixed(1294.0/65536.0,1,-nbitq), 
to_sfixed(-2301.0/65536.0,1,-nbitq), 
to_sfixed(-2259.0/65536.0,1,-nbitq), 
to_sfixed(1055.0/65536.0,1,-nbitq), 
to_sfixed(669.0/65536.0,1,-nbitq), 
to_sfixed(-2618.0/65536.0,1,-nbitq), 
to_sfixed(272.0/65536.0,1,-nbitq), 
to_sfixed(269.0/65536.0,1,-nbitq), 
to_sfixed(236.0/65536.0,1,-nbitq), 
to_sfixed(4144.0/65536.0,1,-nbitq), 
to_sfixed(-862.0/65536.0,1,-nbitq), 
to_sfixed(-780.0/65536.0,1,-nbitq), 
to_sfixed(-4446.0/65536.0,1,-nbitq), 
to_sfixed(-2607.0/65536.0,1,-nbitq), 
to_sfixed(1151.0/65536.0,1,-nbitq), 
to_sfixed(-3260.0/65536.0,1,-nbitq), 
to_sfixed(-2874.0/65536.0,1,-nbitq), 
to_sfixed(-2075.0/65536.0,1,-nbitq), 
to_sfixed(-1465.0/65536.0,1,-nbitq), 
to_sfixed(1058.0/65536.0,1,-nbitq), 
to_sfixed(5253.0/65536.0,1,-nbitq), 
to_sfixed(3144.0/65536.0,1,-nbitq), 
to_sfixed(1211.0/65536.0,1,-nbitq), 
to_sfixed(-904.0/65536.0,1,-nbitq), 
to_sfixed(1384.0/65536.0,1,-nbitq), 
to_sfixed(-1161.0/65536.0,1,-nbitq), 
to_sfixed(2511.0/65536.0,1,-nbitq), 
to_sfixed(2944.0/65536.0,1,-nbitq), 
to_sfixed(-6007.0/65536.0,1,-nbitq), 
to_sfixed(1579.0/65536.0,1,-nbitq), 
to_sfixed(-3033.0/65536.0,1,-nbitq), 
to_sfixed(-1478.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2263.0/65536.0,1,-nbitq), 
to_sfixed(-1155.0/65536.0,1,-nbitq), 
to_sfixed(-6354.0/65536.0,1,-nbitq), 
to_sfixed(1473.0/65536.0,1,-nbitq), 
to_sfixed(7688.0/65536.0,1,-nbitq), 
to_sfixed(-687.0/65536.0,1,-nbitq), 
to_sfixed(-2806.0/65536.0,1,-nbitq), 
to_sfixed(-5295.0/65536.0,1,-nbitq), 
to_sfixed(-2216.0/65536.0,1,-nbitq), 
to_sfixed(2965.0/65536.0,1,-nbitq), 
to_sfixed(3558.0/65536.0,1,-nbitq), 
to_sfixed(4252.0/65536.0,1,-nbitq), 
to_sfixed(-57.0/65536.0,1,-nbitq), 
to_sfixed(4192.0/65536.0,1,-nbitq), 
to_sfixed(-433.0/65536.0,1,-nbitq), 
to_sfixed(-454.0/65536.0,1,-nbitq), 
to_sfixed(131.0/65536.0,1,-nbitq), 
to_sfixed(-1884.0/65536.0,1,-nbitq), 
to_sfixed(433.0/65536.0,1,-nbitq), 
to_sfixed(-2127.0/65536.0,1,-nbitq), 
to_sfixed(1359.0/65536.0,1,-nbitq), 
to_sfixed(2272.0/65536.0,1,-nbitq), 
to_sfixed(-819.0/65536.0,1,-nbitq), 
to_sfixed(-8396.0/65536.0,1,-nbitq), 
to_sfixed(-522.0/65536.0,1,-nbitq), 
to_sfixed(-10302.0/65536.0,1,-nbitq), 
to_sfixed(-3274.0/65536.0,1,-nbitq), 
to_sfixed(816.0/65536.0,1,-nbitq), 
to_sfixed(7084.0/65536.0,1,-nbitq), 
to_sfixed(-2890.0/65536.0,1,-nbitq), 
to_sfixed(-1551.0/65536.0,1,-nbitq), 
to_sfixed(-1218.0/65536.0,1,-nbitq), 
to_sfixed(-1606.0/65536.0,1,-nbitq), 
to_sfixed(-5043.0/65536.0,1,-nbitq), 
to_sfixed(3319.0/65536.0,1,-nbitq), 
to_sfixed(795.0/65536.0,1,-nbitq), 
to_sfixed(-8351.0/65536.0,1,-nbitq), 
to_sfixed(2286.0/65536.0,1,-nbitq), 
to_sfixed(-1436.0/65536.0,1,-nbitq), 
to_sfixed(-3852.0/65536.0,1,-nbitq), 
to_sfixed(962.0/65536.0,1,-nbitq), 
to_sfixed(-1012.0/65536.0,1,-nbitq), 
to_sfixed(1704.0/65536.0,1,-nbitq), 
to_sfixed(4304.0/65536.0,1,-nbitq), 
to_sfixed(2057.0/65536.0,1,-nbitq), 
to_sfixed(1905.0/65536.0,1,-nbitq), 
to_sfixed(-1979.0/65536.0,1,-nbitq), 
to_sfixed(-4485.0/65536.0,1,-nbitq), 
to_sfixed(2619.0/65536.0,1,-nbitq), 
to_sfixed(1481.0/65536.0,1,-nbitq), 
to_sfixed(-1242.0/65536.0,1,-nbitq), 
to_sfixed(-1666.0/65536.0,1,-nbitq), 
to_sfixed(-2825.0/65536.0,1,-nbitq), 
to_sfixed(-231.0/65536.0,1,-nbitq), 
to_sfixed(-2793.0/65536.0,1,-nbitq), 
to_sfixed(3704.0/65536.0,1,-nbitq), 
to_sfixed(-2691.0/65536.0,1,-nbitq), 
to_sfixed(751.0/65536.0,1,-nbitq), 
to_sfixed(554.0/65536.0,1,-nbitq), 
to_sfixed(-9493.0/65536.0,1,-nbitq), 
to_sfixed(-3565.0/65536.0,1,-nbitq), 
to_sfixed(936.0/65536.0,1,-nbitq), 
to_sfixed(-372.0/65536.0,1,-nbitq), 
to_sfixed(-1971.0/65536.0,1,-nbitq), 
to_sfixed(-5087.0/65536.0,1,-nbitq), 
to_sfixed(1618.0/65536.0,1,-nbitq), 
to_sfixed(1275.0/65536.0,1,-nbitq), 
to_sfixed(311.0/65536.0,1,-nbitq), 
to_sfixed(3791.0/65536.0,1,-nbitq), 
to_sfixed(6001.0/65536.0,1,-nbitq), 
to_sfixed(2277.0/65536.0,1,-nbitq), 
to_sfixed(-882.0/65536.0,1,-nbitq), 
to_sfixed(-656.0/65536.0,1,-nbitq), 
to_sfixed(-2896.0/65536.0,1,-nbitq), 
to_sfixed(-2490.0/65536.0,1,-nbitq), 
to_sfixed(-1029.0/65536.0,1,-nbitq), 
to_sfixed(-5949.0/65536.0,1,-nbitq), 
to_sfixed(-2241.0/65536.0,1,-nbitq), 
to_sfixed(1129.0/65536.0,1,-nbitq), 
to_sfixed(-3991.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2652.0/65536.0,1,-nbitq), 
to_sfixed(-1568.0/65536.0,1,-nbitq), 
to_sfixed(-7502.0/65536.0,1,-nbitq), 
to_sfixed(-4927.0/65536.0,1,-nbitq), 
to_sfixed(-2296.0/65536.0,1,-nbitq), 
to_sfixed(-3648.0/65536.0,1,-nbitq), 
to_sfixed(-5984.0/65536.0,1,-nbitq), 
to_sfixed(-180.0/65536.0,1,-nbitq), 
to_sfixed(2956.0/65536.0,1,-nbitq), 
to_sfixed(-2323.0/65536.0,1,-nbitq), 
to_sfixed(-2417.0/65536.0,1,-nbitq), 
to_sfixed(5573.0/65536.0,1,-nbitq), 
to_sfixed(791.0/65536.0,1,-nbitq), 
to_sfixed(1139.0/65536.0,1,-nbitq), 
to_sfixed(-92.0/65536.0,1,-nbitq), 
to_sfixed(-38.0/65536.0,1,-nbitq), 
to_sfixed(505.0/65536.0,1,-nbitq), 
to_sfixed(1608.0/65536.0,1,-nbitq), 
to_sfixed(-3375.0/65536.0,1,-nbitq), 
to_sfixed(2968.0/65536.0,1,-nbitq), 
to_sfixed(4308.0/65536.0,1,-nbitq), 
to_sfixed(8748.0/65536.0,1,-nbitq), 
to_sfixed(2609.0/65536.0,1,-nbitq), 
to_sfixed(-10554.0/65536.0,1,-nbitq), 
to_sfixed(3135.0/65536.0,1,-nbitq), 
to_sfixed(-18318.0/65536.0,1,-nbitq), 
to_sfixed(-1228.0/65536.0,1,-nbitq), 
to_sfixed(487.0/65536.0,1,-nbitq), 
to_sfixed(3642.0/65536.0,1,-nbitq), 
to_sfixed(-5758.0/65536.0,1,-nbitq), 
to_sfixed(1354.0/65536.0,1,-nbitq), 
to_sfixed(-1564.0/65536.0,1,-nbitq), 
to_sfixed(1312.0/65536.0,1,-nbitq), 
to_sfixed(-1406.0/65536.0,1,-nbitq), 
to_sfixed(722.0/65536.0,1,-nbitq), 
to_sfixed(-838.0/65536.0,1,-nbitq), 
to_sfixed(-6189.0/65536.0,1,-nbitq), 
to_sfixed(4322.0/65536.0,1,-nbitq), 
to_sfixed(-10.0/65536.0,1,-nbitq), 
to_sfixed(-8474.0/65536.0,1,-nbitq), 
to_sfixed(-1268.0/65536.0,1,-nbitq), 
to_sfixed(-2344.0/65536.0,1,-nbitq), 
to_sfixed(7818.0/65536.0,1,-nbitq), 
to_sfixed(5357.0/65536.0,1,-nbitq), 
to_sfixed(2948.0/65536.0,1,-nbitq), 
to_sfixed(5118.0/65536.0,1,-nbitq), 
to_sfixed(2610.0/65536.0,1,-nbitq), 
to_sfixed(-502.0/65536.0,1,-nbitq), 
to_sfixed(2581.0/65536.0,1,-nbitq), 
to_sfixed(2591.0/65536.0,1,-nbitq), 
to_sfixed(-40.0/65536.0,1,-nbitq), 
to_sfixed(-2191.0/65536.0,1,-nbitq), 
to_sfixed(-69.0/65536.0,1,-nbitq), 
to_sfixed(1245.0/65536.0,1,-nbitq), 
to_sfixed(-7101.0/65536.0,1,-nbitq), 
to_sfixed(515.0/65536.0,1,-nbitq), 
to_sfixed(3716.0/65536.0,1,-nbitq), 
to_sfixed(2646.0/65536.0,1,-nbitq), 
to_sfixed(330.0/65536.0,1,-nbitq), 
to_sfixed(-11462.0/65536.0,1,-nbitq), 
to_sfixed(-8866.0/65536.0,1,-nbitq), 
to_sfixed(-2120.0/65536.0,1,-nbitq), 
to_sfixed(2613.0/65536.0,1,-nbitq), 
to_sfixed(1248.0/65536.0,1,-nbitq), 
to_sfixed(-7462.0/65536.0,1,-nbitq), 
to_sfixed(2616.0/65536.0,1,-nbitq), 
to_sfixed(3382.0/65536.0,1,-nbitq), 
to_sfixed(3435.0/65536.0,1,-nbitq), 
to_sfixed(4731.0/65536.0,1,-nbitq), 
to_sfixed(387.0/65536.0,1,-nbitq), 
to_sfixed(-333.0/65536.0,1,-nbitq), 
to_sfixed(566.0/65536.0,1,-nbitq), 
to_sfixed(946.0/65536.0,1,-nbitq), 
to_sfixed(-3320.0/65536.0,1,-nbitq), 
to_sfixed(-1349.0/65536.0,1,-nbitq), 
to_sfixed(-4670.0/65536.0,1,-nbitq), 
to_sfixed(82.0/65536.0,1,-nbitq), 
to_sfixed(-4574.0/65536.0,1,-nbitq), 
to_sfixed(67.0/65536.0,1,-nbitq), 
to_sfixed(-1441.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1432.0/65536.0,1,-nbitq), 
to_sfixed(-4689.0/65536.0,1,-nbitq), 
to_sfixed(-10589.0/65536.0,1,-nbitq), 
to_sfixed(-5658.0/65536.0,1,-nbitq), 
to_sfixed(-4829.0/65536.0,1,-nbitq), 
to_sfixed(7702.0/65536.0,1,-nbitq), 
to_sfixed(-5694.0/65536.0,1,-nbitq), 
to_sfixed(-57.0/65536.0,1,-nbitq), 
to_sfixed(-1526.0/65536.0,1,-nbitq), 
to_sfixed(-119.0/65536.0,1,-nbitq), 
to_sfixed(-1402.0/65536.0,1,-nbitq), 
to_sfixed(-3121.0/65536.0,1,-nbitq), 
to_sfixed(810.0/65536.0,1,-nbitq), 
to_sfixed(4924.0/65536.0,1,-nbitq), 
to_sfixed(-654.0/65536.0,1,-nbitq), 
to_sfixed(2656.0/65536.0,1,-nbitq), 
to_sfixed(-1021.0/65536.0,1,-nbitq), 
to_sfixed(6035.0/65536.0,1,-nbitq), 
to_sfixed(-1941.0/65536.0,1,-nbitq), 
to_sfixed(3316.0/65536.0,1,-nbitq), 
to_sfixed(1379.0/65536.0,1,-nbitq), 
to_sfixed(-3722.0/65536.0,1,-nbitq), 
to_sfixed(121.0/65536.0,1,-nbitq), 
to_sfixed(-15215.0/65536.0,1,-nbitq), 
to_sfixed(135.0/65536.0,1,-nbitq), 
to_sfixed(-21993.0/65536.0,1,-nbitq), 
to_sfixed(-1227.0/65536.0,1,-nbitq), 
to_sfixed(-1053.0/65536.0,1,-nbitq), 
to_sfixed(3728.0/65536.0,1,-nbitq), 
to_sfixed(-2554.0/65536.0,1,-nbitq), 
to_sfixed(5163.0/65536.0,1,-nbitq), 
to_sfixed(959.0/65536.0,1,-nbitq), 
to_sfixed(2764.0/65536.0,1,-nbitq), 
to_sfixed(-884.0/65536.0,1,-nbitq), 
to_sfixed(2465.0/65536.0,1,-nbitq), 
to_sfixed(1225.0/65536.0,1,-nbitq), 
to_sfixed(-9756.0/65536.0,1,-nbitq), 
to_sfixed(5438.0/65536.0,1,-nbitq), 
to_sfixed(2477.0/65536.0,1,-nbitq), 
to_sfixed(-9676.0/65536.0,1,-nbitq), 
to_sfixed(3220.0/65536.0,1,-nbitq), 
to_sfixed(2527.0/65536.0,1,-nbitq), 
to_sfixed(5621.0/65536.0,1,-nbitq), 
to_sfixed(5421.0/65536.0,1,-nbitq), 
to_sfixed(178.0/65536.0,1,-nbitq), 
to_sfixed(-1876.0/65536.0,1,-nbitq), 
to_sfixed(1425.0/65536.0,1,-nbitq), 
to_sfixed(-4062.0/65536.0,1,-nbitq), 
to_sfixed(1392.0/65536.0,1,-nbitq), 
to_sfixed(286.0/65536.0,1,-nbitq), 
to_sfixed(773.0/65536.0,1,-nbitq), 
to_sfixed(553.0/65536.0,1,-nbitq), 
to_sfixed(-4753.0/65536.0,1,-nbitq), 
to_sfixed(5700.0/65536.0,1,-nbitq), 
to_sfixed(-4139.0/65536.0,1,-nbitq), 
to_sfixed(-746.0/65536.0,1,-nbitq), 
to_sfixed(3819.0/65536.0,1,-nbitq), 
to_sfixed(1708.0/65536.0,1,-nbitq), 
to_sfixed(2740.0/65536.0,1,-nbitq), 
to_sfixed(-11468.0/65536.0,1,-nbitq), 
to_sfixed(-2242.0/65536.0,1,-nbitq), 
to_sfixed(-3045.0/65536.0,1,-nbitq), 
to_sfixed(2344.0/65536.0,1,-nbitq), 
to_sfixed(-1562.0/65536.0,1,-nbitq), 
to_sfixed(-9565.0/65536.0,1,-nbitq), 
to_sfixed(4939.0/65536.0,1,-nbitq), 
to_sfixed(-672.0/65536.0,1,-nbitq), 
to_sfixed(1335.0/65536.0,1,-nbitq), 
to_sfixed(7031.0/65536.0,1,-nbitq), 
to_sfixed(-2643.0/65536.0,1,-nbitq), 
to_sfixed(1923.0/65536.0,1,-nbitq), 
to_sfixed(-75.0/65536.0,1,-nbitq), 
to_sfixed(-713.0/65536.0,1,-nbitq), 
to_sfixed(-167.0/65536.0,1,-nbitq), 
to_sfixed(1536.0/65536.0,1,-nbitq), 
to_sfixed(-1530.0/65536.0,1,-nbitq), 
to_sfixed(-4448.0/65536.0,1,-nbitq), 
to_sfixed(-2172.0/65536.0,1,-nbitq), 
to_sfixed(-473.0/65536.0,1,-nbitq), 
to_sfixed(-3992.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3079.0/65536.0,1,-nbitq), 
to_sfixed(-1791.0/65536.0,1,-nbitq), 
to_sfixed(-5964.0/65536.0,1,-nbitq), 
to_sfixed(-3239.0/65536.0,1,-nbitq), 
to_sfixed(233.0/65536.0,1,-nbitq), 
to_sfixed(2238.0/65536.0,1,-nbitq), 
to_sfixed(-5732.0/65536.0,1,-nbitq), 
to_sfixed(6475.0/65536.0,1,-nbitq), 
to_sfixed(-4760.0/65536.0,1,-nbitq), 
to_sfixed(491.0/65536.0,1,-nbitq), 
to_sfixed(-4382.0/65536.0,1,-nbitq), 
to_sfixed(-5587.0/65536.0,1,-nbitq), 
to_sfixed(-1421.0/65536.0,1,-nbitq), 
to_sfixed(70.0/65536.0,1,-nbitq), 
to_sfixed(1132.0/65536.0,1,-nbitq), 
to_sfixed(413.0/65536.0,1,-nbitq), 
to_sfixed(1325.0/65536.0,1,-nbitq), 
to_sfixed(4366.0/65536.0,1,-nbitq), 
to_sfixed(1335.0/65536.0,1,-nbitq), 
to_sfixed(1681.0/65536.0,1,-nbitq), 
to_sfixed(3980.0/65536.0,1,-nbitq), 
to_sfixed(-5932.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(-9258.0/65536.0,1,-nbitq), 
to_sfixed(-1980.0/65536.0,1,-nbitq), 
to_sfixed(-13590.0/65536.0,1,-nbitq), 
to_sfixed(-468.0/65536.0,1,-nbitq), 
to_sfixed(2880.0/65536.0,1,-nbitq), 
to_sfixed(2618.0/65536.0,1,-nbitq), 
to_sfixed(2991.0/65536.0,1,-nbitq), 
to_sfixed(2018.0/65536.0,1,-nbitq), 
to_sfixed(-1007.0/65536.0,1,-nbitq), 
to_sfixed(5301.0/65536.0,1,-nbitq), 
to_sfixed(1463.0/65536.0,1,-nbitq), 
to_sfixed(-3036.0/65536.0,1,-nbitq), 
to_sfixed(-1105.0/65536.0,1,-nbitq), 
to_sfixed(-3846.0/65536.0,1,-nbitq), 
to_sfixed(3913.0/65536.0,1,-nbitq), 
to_sfixed(1859.0/65536.0,1,-nbitq), 
to_sfixed(-4907.0/65536.0,1,-nbitq), 
to_sfixed(4325.0/65536.0,1,-nbitq), 
to_sfixed(1073.0/65536.0,1,-nbitq), 
to_sfixed(7806.0/65536.0,1,-nbitq), 
to_sfixed(4098.0/65536.0,1,-nbitq), 
to_sfixed(163.0/65536.0,1,-nbitq), 
to_sfixed(-752.0/65536.0,1,-nbitq), 
to_sfixed(122.0/65536.0,1,-nbitq), 
to_sfixed(-1691.0/65536.0,1,-nbitq), 
to_sfixed(2346.0/65536.0,1,-nbitq), 
to_sfixed(9.0/65536.0,1,-nbitq), 
to_sfixed(-2592.0/65536.0,1,-nbitq), 
to_sfixed(-4232.0/65536.0,1,-nbitq), 
to_sfixed(-1736.0/65536.0,1,-nbitq), 
to_sfixed(7232.0/65536.0,1,-nbitq), 
to_sfixed(-7378.0/65536.0,1,-nbitq), 
to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(-1197.0/65536.0,1,-nbitq), 
to_sfixed(-2204.0/65536.0,1,-nbitq), 
to_sfixed(175.0/65536.0,1,-nbitq), 
to_sfixed(-4477.0/65536.0,1,-nbitq), 
to_sfixed(7890.0/65536.0,1,-nbitq), 
to_sfixed(2310.0/65536.0,1,-nbitq), 
to_sfixed(42.0/65536.0,1,-nbitq), 
to_sfixed(-2840.0/65536.0,1,-nbitq), 
to_sfixed(-1223.0/65536.0,1,-nbitq), 
to_sfixed(8577.0/65536.0,1,-nbitq), 
to_sfixed(3184.0/65536.0,1,-nbitq), 
to_sfixed(-931.0/65536.0,1,-nbitq), 
to_sfixed(8244.0/65536.0,1,-nbitq), 
to_sfixed(-4117.0/65536.0,1,-nbitq), 
to_sfixed(-359.0/65536.0,1,-nbitq), 
to_sfixed(1711.0/65536.0,1,-nbitq), 
to_sfixed(-329.0/65536.0,1,-nbitq), 
to_sfixed(-829.0/65536.0,1,-nbitq), 
to_sfixed(-1944.0/65536.0,1,-nbitq), 
to_sfixed(-478.0/65536.0,1,-nbitq), 
to_sfixed(1764.0/65536.0,1,-nbitq), 
to_sfixed(1114.0/65536.0,1,-nbitq), 
to_sfixed(1694.0/65536.0,1,-nbitq), 
to_sfixed(-2877.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1047.0/65536.0,1,-nbitq), 
to_sfixed(-2932.0/65536.0,1,-nbitq), 
to_sfixed(-3272.0/65536.0,1,-nbitq), 
to_sfixed(-1745.0/65536.0,1,-nbitq), 
to_sfixed(1093.0/65536.0,1,-nbitq), 
to_sfixed(3983.0/65536.0,1,-nbitq), 
to_sfixed(-11862.0/65536.0,1,-nbitq), 
to_sfixed(12509.0/65536.0,1,-nbitq), 
to_sfixed(3741.0/65536.0,1,-nbitq), 
to_sfixed(-2753.0/65536.0,1,-nbitq), 
to_sfixed(-3014.0/65536.0,1,-nbitq), 
to_sfixed(-11101.0/65536.0,1,-nbitq), 
to_sfixed(-1078.0/65536.0,1,-nbitq), 
to_sfixed(2595.0/65536.0,1,-nbitq), 
to_sfixed(2495.0/65536.0,1,-nbitq), 
to_sfixed(3000.0/65536.0,1,-nbitq), 
to_sfixed(696.0/65536.0,1,-nbitq), 
to_sfixed(9360.0/65536.0,1,-nbitq), 
to_sfixed(-223.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(-907.0/65536.0,1,-nbitq), 
to_sfixed(-4454.0/65536.0,1,-nbitq), 
to_sfixed(-869.0/65536.0,1,-nbitq), 
to_sfixed(-152.0/65536.0,1,-nbitq), 
to_sfixed(-2050.0/65536.0,1,-nbitq), 
to_sfixed(-16454.0/65536.0,1,-nbitq), 
to_sfixed(-3638.0/65536.0,1,-nbitq), 
to_sfixed(1815.0/65536.0,1,-nbitq), 
to_sfixed(94.0/65536.0,1,-nbitq), 
to_sfixed(5090.0/65536.0,1,-nbitq), 
to_sfixed(3355.0/65536.0,1,-nbitq), 
to_sfixed(3642.0/65536.0,1,-nbitq), 
to_sfixed(3177.0/65536.0,1,-nbitq), 
to_sfixed(1748.0/65536.0,1,-nbitq), 
to_sfixed(-2952.0/65536.0,1,-nbitq), 
to_sfixed(-370.0/65536.0,1,-nbitq), 
to_sfixed(-14797.0/65536.0,1,-nbitq), 
to_sfixed(2278.0/65536.0,1,-nbitq), 
to_sfixed(-2960.0/65536.0,1,-nbitq), 
to_sfixed(2484.0/65536.0,1,-nbitq), 
to_sfixed(976.0/65536.0,1,-nbitq), 
to_sfixed(-571.0/65536.0,1,-nbitq), 
to_sfixed(5664.0/65536.0,1,-nbitq), 
to_sfixed(3049.0/65536.0,1,-nbitq), 
to_sfixed(-564.0/65536.0,1,-nbitq), 
to_sfixed(-8357.0/65536.0,1,-nbitq), 
to_sfixed(3674.0/65536.0,1,-nbitq), 
to_sfixed(-1299.0/65536.0,1,-nbitq), 
to_sfixed(3988.0/65536.0,1,-nbitq), 
to_sfixed(1410.0/65536.0,1,-nbitq), 
to_sfixed(-2205.0/65536.0,1,-nbitq), 
to_sfixed(2073.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(-298.0/65536.0,1,-nbitq), 
to_sfixed(-4900.0/65536.0,1,-nbitq), 
to_sfixed(-5223.0/65536.0,1,-nbitq), 
to_sfixed(1055.0/65536.0,1,-nbitq), 
to_sfixed(-4544.0/65536.0,1,-nbitq), 
to_sfixed(-1845.0/65536.0,1,-nbitq), 
to_sfixed(3015.0/65536.0,1,-nbitq), 
to_sfixed(20071.0/65536.0,1,-nbitq), 
to_sfixed(-824.0/65536.0,1,-nbitq), 
to_sfixed(542.0/65536.0,1,-nbitq), 
to_sfixed(-911.0/65536.0,1,-nbitq), 
to_sfixed(585.0/65536.0,1,-nbitq), 
to_sfixed(-1060.0/65536.0,1,-nbitq), 
to_sfixed(-358.0/65536.0,1,-nbitq), 
to_sfixed(-2996.0/65536.0,1,-nbitq), 
to_sfixed(5394.0/65536.0,1,-nbitq), 
to_sfixed(-9521.0/65536.0,1,-nbitq), 
to_sfixed(-1991.0/65536.0,1,-nbitq), 
to_sfixed(4282.0/65536.0,1,-nbitq), 
to_sfixed(-2085.0/65536.0,1,-nbitq), 
to_sfixed(473.0/65536.0,1,-nbitq), 
to_sfixed(-2383.0/65536.0,1,-nbitq), 
to_sfixed(-3362.0/65536.0,1,-nbitq), 
to_sfixed(7678.0/65536.0,1,-nbitq), 
to_sfixed(-4783.0/65536.0,1,-nbitq), 
to_sfixed(2650.0/65536.0,1,-nbitq), 
to_sfixed(-2687.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-288.0/65536.0,1,-nbitq), 
to_sfixed(2887.0/65536.0,1,-nbitq), 
to_sfixed(-7949.0/65536.0,1,-nbitq), 
to_sfixed(-1868.0/65536.0,1,-nbitq), 
to_sfixed(-5801.0/65536.0,1,-nbitq), 
to_sfixed(4148.0/65536.0,1,-nbitq), 
to_sfixed(-7755.0/65536.0,1,-nbitq), 
to_sfixed(7905.0/65536.0,1,-nbitq), 
to_sfixed(668.0/65536.0,1,-nbitq), 
to_sfixed(-448.0/65536.0,1,-nbitq), 
to_sfixed(-67.0/65536.0,1,-nbitq), 
to_sfixed(3283.0/65536.0,1,-nbitq), 
to_sfixed(1607.0/65536.0,1,-nbitq), 
to_sfixed(-4736.0/65536.0,1,-nbitq), 
to_sfixed(1087.0/65536.0,1,-nbitq), 
to_sfixed(1761.0/65536.0,1,-nbitq), 
to_sfixed(417.0/65536.0,1,-nbitq), 
to_sfixed(7931.0/65536.0,1,-nbitq), 
to_sfixed(5646.0/65536.0,1,-nbitq), 
to_sfixed(-2561.0/65536.0,1,-nbitq), 
to_sfixed(68.0/65536.0,1,-nbitq), 
to_sfixed(-2351.0/65536.0,1,-nbitq), 
to_sfixed(910.0/65536.0,1,-nbitq), 
to_sfixed(-8566.0/65536.0,1,-nbitq), 
to_sfixed(1219.0/65536.0,1,-nbitq), 
to_sfixed(-12571.0/65536.0,1,-nbitq), 
to_sfixed(-10865.0/65536.0,1,-nbitq), 
to_sfixed(1422.0/65536.0,1,-nbitq), 
to_sfixed(-6736.0/65536.0,1,-nbitq), 
to_sfixed(3484.0/65536.0,1,-nbitq), 
to_sfixed(-1770.0/65536.0,1,-nbitq), 
to_sfixed(-5182.0/65536.0,1,-nbitq), 
to_sfixed(2901.0/65536.0,1,-nbitq), 
to_sfixed(-9584.0/65536.0,1,-nbitq), 
to_sfixed(-2965.0/65536.0,1,-nbitq), 
to_sfixed(2758.0/65536.0,1,-nbitq), 
to_sfixed(-6356.0/65536.0,1,-nbitq), 
to_sfixed(-506.0/65536.0,1,-nbitq), 
to_sfixed(-3212.0/65536.0,1,-nbitq), 
to_sfixed(2868.0/65536.0,1,-nbitq), 
to_sfixed(-4552.0/65536.0,1,-nbitq), 
to_sfixed(-1705.0/65536.0,1,-nbitq), 
to_sfixed(3007.0/65536.0,1,-nbitq), 
to_sfixed(436.0/65536.0,1,-nbitq), 
to_sfixed(375.0/65536.0,1,-nbitq), 
to_sfixed(-800.0/65536.0,1,-nbitq), 
to_sfixed(-1560.0/65536.0,1,-nbitq), 
to_sfixed(-1720.0/65536.0,1,-nbitq), 
to_sfixed(-540.0/65536.0,1,-nbitq), 
to_sfixed(1434.0/65536.0,1,-nbitq), 
to_sfixed(-2159.0/65536.0,1,-nbitq), 
to_sfixed(-1074.0/65536.0,1,-nbitq), 
to_sfixed(-2402.0/65536.0,1,-nbitq), 
to_sfixed(-17973.0/65536.0,1,-nbitq), 
to_sfixed(-4719.0/65536.0,1,-nbitq), 
to_sfixed(-6496.0/65536.0,1,-nbitq), 
to_sfixed(-261.0/65536.0,1,-nbitq), 
to_sfixed(2703.0/65536.0,1,-nbitq), 
to_sfixed(1676.0/65536.0,1,-nbitq), 
to_sfixed(3873.0/65536.0,1,-nbitq), 
to_sfixed(17813.0/65536.0,1,-nbitq), 
to_sfixed(-1633.0/65536.0,1,-nbitq), 
to_sfixed(2345.0/65536.0,1,-nbitq), 
to_sfixed(481.0/65536.0,1,-nbitq), 
to_sfixed(-2274.0/65536.0,1,-nbitq), 
to_sfixed(940.0/65536.0,1,-nbitq), 
to_sfixed(-1931.0/65536.0,1,-nbitq), 
to_sfixed(-2244.0/65536.0,1,-nbitq), 
to_sfixed(6078.0/65536.0,1,-nbitq), 
to_sfixed(1404.0/65536.0,1,-nbitq), 
to_sfixed(-1015.0/65536.0,1,-nbitq), 
to_sfixed(1747.0/65536.0,1,-nbitq), 
to_sfixed(-5062.0/65536.0,1,-nbitq), 
to_sfixed(-1293.0/65536.0,1,-nbitq), 
to_sfixed(-2652.0/65536.0,1,-nbitq), 
to_sfixed(-2508.0/65536.0,1,-nbitq), 
to_sfixed(86.0/65536.0,1,-nbitq), 
to_sfixed(-5794.0/65536.0,1,-nbitq), 
to_sfixed(2336.0/65536.0,1,-nbitq), 
to_sfixed(-9732.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2400.0/65536.0,1,-nbitq), 
to_sfixed(1059.0/65536.0,1,-nbitq), 
to_sfixed(-1079.0/65536.0,1,-nbitq), 
to_sfixed(-2774.0/65536.0,1,-nbitq), 
to_sfixed(-4486.0/65536.0,1,-nbitq), 
to_sfixed(1696.0/65536.0,1,-nbitq), 
to_sfixed(-1710.0/65536.0,1,-nbitq), 
to_sfixed(2869.0/65536.0,1,-nbitq), 
to_sfixed(2191.0/65536.0,1,-nbitq), 
to_sfixed(1373.0/65536.0,1,-nbitq), 
to_sfixed(-727.0/65536.0,1,-nbitq), 
to_sfixed(-1867.0/65536.0,1,-nbitq), 
to_sfixed(3518.0/65536.0,1,-nbitq), 
to_sfixed(-10070.0/65536.0,1,-nbitq), 
to_sfixed(3096.0/65536.0,1,-nbitq), 
to_sfixed(2568.0/65536.0,1,-nbitq), 
to_sfixed(2515.0/65536.0,1,-nbitq), 
to_sfixed(992.0/65536.0,1,-nbitq), 
to_sfixed(2409.0/65536.0,1,-nbitq), 
to_sfixed(1833.0/65536.0,1,-nbitq), 
to_sfixed(751.0/65536.0,1,-nbitq), 
to_sfixed(5614.0/65536.0,1,-nbitq), 
to_sfixed(191.0/65536.0,1,-nbitq), 
to_sfixed(-10247.0/65536.0,1,-nbitq), 
to_sfixed(-3055.0/65536.0,1,-nbitq), 
to_sfixed(-9046.0/65536.0,1,-nbitq), 
to_sfixed(-8890.0/65536.0,1,-nbitq), 
to_sfixed(1330.0/65536.0,1,-nbitq), 
to_sfixed(-8840.0/65536.0,1,-nbitq), 
to_sfixed(3663.0/65536.0,1,-nbitq), 
to_sfixed(-2128.0/65536.0,1,-nbitq), 
to_sfixed(-6980.0/65536.0,1,-nbitq), 
to_sfixed(237.0/65536.0,1,-nbitq), 
to_sfixed(-6458.0/65536.0,1,-nbitq), 
to_sfixed(-1960.0/65536.0,1,-nbitq), 
to_sfixed(1888.0/65536.0,1,-nbitq), 
to_sfixed(-7206.0/65536.0,1,-nbitq), 
to_sfixed(4834.0/65536.0,1,-nbitq), 
to_sfixed(-5314.0/65536.0,1,-nbitq), 
to_sfixed(1707.0/65536.0,1,-nbitq), 
to_sfixed(-3109.0/65536.0,1,-nbitq), 
to_sfixed(350.0/65536.0,1,-nbitq), 
to_sfixed(-4963.0/65536.0,1,-nbitq), 
to_sfixed(-1104.0/65536.0,1,-nbitq), 
to_sfixed(411.0/65536.0,1,-nbitq), 
to_sfixed(224.0/65536.0,1,-nbitq), 
to_sfixed(-4097.0/65536.0,1,-nbitq), 
to_sfixed(3799.0/65536.0,1,-nbitq), 
to_sfixed(-2343.0/65536.0,1,-nbitq), 
to_sfixed(-215.0/65536.0,1,-nbitq), 
to_sfixed(-1675.0/65536.0,1,-nbitq), 
to_sfixed(-1332.0/65536.0,1,-nbitq), 
to_sfixed(3155.0/65536.0,1,-nbitq), 
to_sfixed(-9658.0/65536.0,1,-nbitq), 
to_sfixed(-3539.0/65536.0,1,-nbitq), 
to_sfixed(2326.0/65536.0,1,-nbitq), 
to_sfixed(137.0/65536.0,1,-nbitq), 
to_sfixed(3630.0/65536.0,1,-nbitq), 
to_sfixed(1632.0/65536.0,1,-nbitq), 
to_sfixed(2594.0/65536.0,1,-nbitq), 
to_sfixed(5217.0/65536.0,1,-nbitq), 
to_sfixed(-489.0/65536.0,1,-nbitq), 
to_sfixed(1315.0/65536.0,1,-nbitq), 
to_sfixed(-2770.0/65536.0,1,-nbitq), 
to_sfixed(757.0/65536.0,1,-nbitq), 
to_sfixed(21343.0/65536.0,1,-nbitq), 
to_sfixed(2624.0/65536.0,1,-nbitq), 
to_sfixed(5796.0/65536.0,1,-nbitq), 
to_sfixed(1860.0/65536.0,1,-nbitq), 
to_sfixed(2734.0/65536.0,1,-nbitq), 
to_sfixed(-2254.0/65536.0,1,-nbitq), 
to_sfixed(-1551.0/65536.0,1,-nbitq), 
to_sfixed(-4426.0/65536.0,1,-nbitq), 
to_sfixed(-156.0/65536.0,1,-nbitq), 
to_sfixed(2232.0/65536.0,1,-nbitq), 
to_sfixed(-3789.0/65536.0,1,-nbitq), 
to_sfixed(-2423.0/65536.0,1,-nbitq), 
to_sfixed(4871.0/65536.0,1,-nbitq), 
to_sfixed(1809.0/65536.0,1,-nbitq), 
to_sfixed(-8163.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-5292.0/65536.0,1,-nbitq), 
to_sfixed(4100.0/65536.0,1,-nbitq), 
to_sfixed(-9812.0/65536.0,1,-nbitq), 
to_sfixed(1823.0/65536.0,1,-nbitq), 
to_sfixed(-5887.0/65536.0,1,-nbitq), 
to_sfixed(5031.0/65536.0,1,-nbitq), 
to_sfixed(-2222.0/65536.0,1,-nbitq), 
to_sfixed(-4872.0/65536.0,1,-nbitq), 
to_sfixed(-4215.0/65536.0,1,-nbitq), 
to_sfixed(1309.0/65536.0,1,-nbitq), 
to_sfixed(-2014.0/65536.0,1,-nbitq), 
to_sfixed(-5866.0/65536.0,1,-nbitq), 
to_sfixed(3443.0/65536.0,1,-nbitq), 
to_sfixed(-5433.0/65536.0,1,-nbitq), 
to_sfixed(244.0/65536.0,1,-nbitq), 
to_sfixed(2006.0/65536.0,1,-nbitq), 
to_sfixed(552.0/65536.0,1,-nbitq), 
to_sfixed(-13503.0/65536.0,1,-nbitq), 
to_sfixed(5898.0/65536.0,1,-nbitq), 
to_sfixed(470.0/65536.0,1,-nbitq), 
to_sfixed(862.0/65536.0,1,-nbitq), 
to_sfixed(5987.0/65536.0,1,-nbitq), 
to_sfixed(-12496.0/65536.0,1,-nbitq), 
to_sfixed(-1498.0/65536.0,1,-nbitq), 
to_sfixed(-8875.0/65536.0,1,-nbitq), 
to_sfixed(-4101.0/65536.0,1,-nbitq), 
to_sfixed(-9773.0/65536.0,1,-nbitq), 
to_sfixed(-508.0/65536.0,1,-nbitq), 
to_sfixed(-12408.0/65536.0,1,-nbitq), 
to_sfixed(5933.0/65536.0,1,-nbitq), 
to_sfixed(-5719.0/65536.0,1,-nbitq), 
to_sfixed(-5197.0/65536.0,1,-nbitq), 
to_sfixed(-2041.0/65536.0,1,-nbitq), 
to_sfixed(10172.0/65536.0,1,-nbitq), 
to_sfixed(911.0/65536.0,1,-nbitq), 
to_sfixed(-111.0/65536.0,1,-nbitq), 
to_sfixed(1739.0/65536.0,1,-nbitq), 
to_sfixed(1769.0/65536.0,1,-nbitq), 
to_sfixed(110.0/65536.0,1,-nbitq), 
to_sfixed(2829.0/65536.0,1,-nbitq), 
to_sfixed(6409.0/65536.0,1,-nbitq), 
to_sfixed(224.0/65536.0,1,-nbitq), 
to_sfixed(-10797.0/65536.0,1,-nbitq), 
to_sfixed(2930.0/65536.0,1,-nbitq), 
to_sfixed(145.0/65536.0,1,-nbitq), 
to_sfixed(-3938.0/65536.0,1,-nbitq), 
to_sfixed(-2883.0/65536.0,1,-nbitq), 
to_sfixed(4783.0/65536.0,1,-nbitq), 
to_sfixed(3882.0/65536.0,1,-nbitq), 
to_sfixed(-229.0/65536.0,1,-nbitq), 
to_sfixed(-1880.0/65536.0,1,-nbitq), 
to_sfixed(-3713.0/65536.0,1,-nbitq), 
to_sfixed(-3011.0/65536.0,1,-nbitq), 
to_sfixed(-5088.0/65536.0,1,-nbitq), 
to_sfixed(7.0/65536.0,1,-nbitq), 
to_sfixed(-1114.0/65536.0,1,-nbitq), 
to_sfixed(551.0/65536.0,1,-nbitq), 
to_sfixed(1330.0/65536.0,1,-nbitq), 
to_sfixed(-1997.0/65536.0,1,-nbitq), 
to_sfixed(3342.0/65536.0,1,-nbitq), 
to_sfixed(-7774.0/65536.0,1,-nbitq), 
to_sfixed(-2249.0/65536.0,1,-nbitq), 
to_sfixed(-891.0/65536.0,1,-nbitq), 
to_sfixed(-182.0/65536.0,1,-nbitq), 
to_sfixed(1786.0/65536.0,1,-nbitq), 
to_sfixed(9190.0/65536.0,1,-nbitq), 
to_sfixed(2122.0/65536.0,1,-nbitq), 
to_sfixed(10608.0/65536.0,1,-nbitq), 
to_sfixed(1407.0/65536.0,1,-nbitq), 
to_sfixed(2330.0/65536.0,1,-nbitq), 
to_sfixed(-4201.0/65536.0,1,-nbitq), 
to_sfixed(2440.0/65536.0,1,-nbitq), 
to_sfixed(-8652.0/65536.0,1,-nbitq), 
to_sfixed(-2425.0/65536.0,1,-nbitq), 
to_sfixed(2560.0/65536.0,1,-nbitq), 
to_sfixed(-8741.0/65536.0,1,-nbitq), 
to_sfixed(6780.0/65536.0,1,-nbitq), 
to_sfixed(9404.0/65536.0,1,-nbitq), 
to_sfixed(2777.0/65536.0,1,-nbitq), 
to_sfixed(-2847.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-8697.0/65536.0,1,-nbitq), 
to_sfixed(2430.0/65536.0,1,-nbitq), 
to_sfixed(-10289.0/65536.0,1,-nbitq), 
to_sfixed(2210.0/65536.0,1,-nbitq), 
to_sfixed(-10539.0/65536.0,1,-nbitq), 
to_sfixed(6494.0/65536.0,1,-nbitq), 
to_sfixed(-2090.0/65536.0,1,-nbitq), 
to_sfixed(-8303.0/65536.0,1,-nbitq), 
to_sfixed(2501.0/65536.0,1,-nbitq), 
to_sfixed(1931.0/65536.0,1,-nbitq), 
to_sfixed(2946.0/65536.0,1,-nbitq), 
to_sfixed(-7830.0/65536.0,1,-nbitq), 
to_sfixed(362.0/65536.0,1,-nbitq), 
to_sfixed(47.0/65536.0,1,-nbitq), 
to_sfixed(-1156.0/65536.0,1,-nbitq), 
to_sfixed(-2785.0/65536.0,1,-nbitq), 
to_sfixed(2755.0/65536.0,1,-nbitq), 
to_sfixed(-9379.0/65536.0,1,-nbitq), 
to_sfixed(-671.0/65536.0,1,-nbitq), 
to_sfixed(-2576.0/65536.0,1,-nbitq), 
to_sfixed(-5757.0/65536.0,1,-nbitq), 
to_sfixed(11032.0/65536.0,1,-nbitq), 
to_sfixed(-5218.0/65536.0,1,-nbitq), 
to_sfixed(-987.0/65536.0,1,-nbitq), 
to_sfixed(-11454.0/65536.0,1,-nbitq), 
to_sfixed(-6578.0/65536.0,1,-nbitq), 
to_sfixed(-6470.0/65536.0,1,-nbitq), 
to_sfixed(3108.0/65536.0,1,-nbitq), 
to_sfixed(-13600.0/65536.0,1,-nbitq), 
to_sfixed(9621.0/65536.0,1,-nbitq), 
to_sfixed(505.0/65536.0,1,-nbitq), 
to_sfixed(-1889.0/65536.0,1,-nbitq), 
to_sfixed(-4763.0/65536.0,1,-nbitq), 
to_sfixed(11741.0/65536.0,1,-nbitq), 
to_sfixed(-2270.0/65536.0,1,-nbitq), 
to_sfixed(3514.0/65536.0,1,-nbitq), 
to_sfixed(-4321.0/65536.0,1,-nbitq), 
to_sfixed(8612.0/65536.0,1,-nbitq), 
to_sfixed(9623.0/65536.0,1,-nbitq), 
to_sfixed(1092.0/65536.0,1,-nbitq), 
to_sfixed(9449.0/65536.0,1,-nbitq), 
to_sfixed(197.0/65536.0,1,-nbitq), 
to_sfixed(-2950.0/65536.0,1,-nbitq), 
to_sfixed(-364.0/65536.0,1,-nbitq), 
to_sfixed(1660.0/65536.0,1,-nbitq), 
to_sfixed(1200.0/65536.0,1,-nbitq), 
to_sfixed(-6402.0/65536.0,1,-nbitq), 
to_sfixed(7079.0/65536.0,1,-nbitq), 
to_sfixed(3589.0/65536.0,1,-nbitq), 
to_sfixed(-3695.0/65536.0,1,-nbitq), 
to_sfixed(2756.0/65536.0,1,-nbitq), 
to_sfixed(5109.0/65536.0,1,-nbitq), 
to_sfixed(-3269.0/65536.0,1,-nbitq), 
to_sfixed(-3697.0/65536.0,1,-nbitq), 
to_sfixed(1282.0/65536.0,1,-nbitq), 
to_sfixed(-1123.0/65536.0,1,-nbitq), 
to_sfixed(1380.0/65536.0,1,-nbitq), 
to_sfixed(5812.0/65536.0,1,-nbitq), 
to_sfixed(-738.0/65536.0,1,-nbitq), 
to_sfixed(4446.0/65536.0,1,-nbitq), 
to_sfixed(-11785.0/65536.0,1,-nbitq), 
to_sfixed(-2185.0/65536.0,1,-nbitq), 
to_sfixed(740.0/65536.0,1,-nbitq), 
to_sfixed(2078.0/65536.0,1,-nbitq), 
to_sfixed(622.0/65536.0,1,-nbitq), 
to_sfixed(-9321.0/65536.0,1,-nbitq), 
to_sfixed(-648.0/65536.0,1,-nbitq), 
to_sfixed(4243.0/65536.0,1,-nbitq), 
to_sfixed(4334.0/65536.0,1,-nbitq), 
to_sfixed(1526.0/65536.0,1,-nbitq), 
to_sfixed(-5603.0/65536.0,1,-nbitq), 
to_sfixed(-8582.0/65536.0,1,-nbitq), 
to_sfixed(-6285.0/65536.0,1,-nbitq), 
to_sfixed(1510.0/65536.0,1,-nbitq), 
to_sfixed(-832.0/65536.0,1,-nbitq), 
to_sfixed(-8862.0/65536.0,1,-nbitq), 
to_sfixed(6486.0/65536.0,1,-nbitq), 
to_sfixed(4886.0/65536.0,1,-nbitq), 
to_sfixed(-1965.0/65536.0,1,-nbitq), 
to_sfixed(-173.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-5013.0/65536.0,1,-nbitq), 
to_sfixed(796.0/65536.0,1,-nbitq), 
to_sfixed(-7826.0/65536.0,1,-nbitq), 
to_sfixed(-1599.0/65536.0,1,-nbitq), 
to_sfixed(2384.0/65536.0,1,-nbitq), 
to_sfixed(6484.0/65536.0,1,-nbitq), 
to_sfixed(722.0/65536.0,1,-nbitq), 
to_sfixed(-5153.0/65536.0,1,-nbitq), 
to_sfixed(4031.0/65536.0,1,-nbitq), 
to_sfixed(1542.0/65536.0,1,-nbitq), 
to_sfixed(619.0/65536.0,1,-nbitq), 
to_sfixed(-7550.0/65536.0,1,-nbitq), 
to_sfixed(4094.0/65536.0,1,-nbitq), 
to_sfixed(-7645.0/65536.0,1,-nbitq), 
to_sfixed(1789.0/65536.0,1,-nbitq), 
to_sfixed(1391.0/65536.0,1,-nbitq), 
to_sfixed(2139.0/65536.0,1,-nbitq), 
to_sfixed(879.0/65536.0,1,-nbitq), 
to_sfixed(1013.0/65536.0,1,-nbitq), 
to_sfixed(-2773.0/65536.0,1,-nbitq), 
to_sfixed(-3863.0/65536.0,1,-nbitq), 
to_sfixed(6189.0/65536.0,1,-nbitq), 
to_sfixed(1380.0/65536.0,1,-nbitq), 
to_sfixed(-3483.0/65536.0,1,-nbitq), 
to_sfixed(-13810.0/65536.0,1,-nbitq), 
to_sfixed(-7079.0/65536.0,1,-nbitq), 
to_sfixed(-83.0/65536.0,1,-nbitq), 
to_sfixed(35.0/65536.0,1,-nbitq), 
to_sfixed(-6369.0/65536.0,1,-nbitq), 
to_sfixed(3052.0/65536.0,1,-nbitq), 
to_sfixed(1678.0/65536.0,1,-nbitq), 
to_sfixed(560.0/65536.0,1,-nbitq), 
to_sfixed(-1660.0/65536.0,1,-nbitq), 
to_sfixed(12599.0/65536.0,1,-nbitq), 
to_sfixed(-3481.0/65536.0,1,-nbitq), 
to_sfixed(668.0/65536.0,1,-nbitq), 
to_sfixed(-9972.0/65536.0,1,-nbitq), 
to_sfixed(6587.0/65536.0,1,-nbitq), 
to_sfixed(19721.0/65536.0,1,-nbitq), 
to_sfixed(1741.0/65536.0,1,-nbitq), 
to_sfixed(8842.0/65536.0,1,-nbitq), 
to_sfixed(-919.0/65536.0,1,-nbitq), 
to_sfixed(-3777.0/65536.0,1,-nbitq), 
to_sfixed(1069.0/65536.0,1,-nbitq), 
to_sfixed(-2564.0/65536.0,1,-nbitq), 
to_sfixed(138.0/65536.0,1,-nbitq), 
to_sfixed(-3773.0/65536.0,1,-nbitq), 
to_sfixed(-289.0/65536.0,1,-nbitq), 
to_sfixed(3616.0/65536.0,1,-nbitq), 
to_sfixed(1527.0/65536.0,1,-nbitq), 
to_sfixed(2579.0/65536.0,1,-nbitq), 
to_sfixed(10081.0/65536.0,1,-nbitq), 
to_sfixed(-1422.0/65536.0,1,-nbitq), 
to_sfixed(-3894.0/65536.0,1,-nbitq), 
to_sfixed(-878.0/65536.0,1,-nbitq), 
to_sfixed(-2625.0/65536.0,1,-nbitq), 
to_sfixed(259.0/65536.0,1,-nbitq), 
to_sfixed(302.0/65536.0,1,-nbitq), 
to_sfixed(966.0/65536.0,1,-nbitq), 
to_sfixed(-855.0/65536.0,1,-nbitq), 
to_sfixed(-4530.0/65536.0,1,-nbitq), 
to_sfixed(2523.0/65536.0,1,-nbitq), 
to_sfixed(2128.0/65536.0,1,-nbitq), 
to_sfixed(2032.0/65536.0,1,-nbitq), 
to_sfixed(-6206.0/65536.0,1,-nbitq), 
to_sfixed(-9027.0/65536.0,1,-nbitq), 
to_sfixed(-2093.0/65536.0,1,-nbitq), 
to_sfixed(211.0/65536.0,1,-nbitq), 
to_sfixed(4510.0/65536.0,1,-nbitq), 
to_sfixed(3791.0/65536.0,1,-nbitq), 
to_sfixed(-3443.0/65536.0,1,-nbitq), 
to_sfixed(-9615.0/65536.0,1,-nbitq), 
to_sfixed(-13172.0/65536.0,1,-nbitq), 
to_sfixed(2537.0/65536.0,1,-nbitq), 
to_sfixed(1509.0/65536.0,1,-nbitq), 
to_sfixed(-7293.0/65536.0,1,-nbitq), 
to_sfixed(8216.0/65536.0,1,-nbitq), 
to_sfixed(1429.0/65536.0,1,-nbitq), 
to_sfixed(-104.0/65536.0,1,-nbitq), 
to_sfixed(3171.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-7847.0/65536.0,1,-nbitq), 
to_sfixed(2692.0/65536.0,1,-nbitq), 
to_sfixed(2129.0/65536.0,1,-nbitq), 
to_sfixed(-3887.0/65536.0,1,-nbitq), 
to_sfixed(4543.0/65536.0,1,-nbitq), 
to_sfixed(6611.0/65536.0,1,-nbitq), 
to_sfixed(1765.0/65536.0,1,-nbitq), 
to_sfixed(3468.0/65536.0,1,-nbitq), 
to_sfixed(2166.0/65536.0,1,-nbitq), 
to_sfixed(889.0/65536.0,1,-nbitq), 
to_sfixed(-796.0/65536.0,1,-nbitq), 
to_sfixed(739.0/65536.0,1,-nbitq), 
to_sfixed(3811.0/65536.0,1,-nbitq), 
to_sfixed(-7451.0/65536.0,1,-nbitq), 
to_sfixed(1171.0/65536.0,1,-nbitq), 
to_sfixed(-2099.0/65536.0,1,-nbitq), 
to_sfixed(-1510.0/65536.0,1,-nbitq), 
to_sfixed(171.0/65536.0,1,-nbitq), 
to_sfixed(-2480.0/65536.0,1,-nbitq), 
to_sfixed(2471.0/65536.0,1,-nbitq), 
to_sfixed(4188.0/65536.0,1,-nbitq), 
to_sfixed(5633.0/65536.0,1,-nbitq), 
to_sfixed(1816.0/65536.0,1,-nbitq), 
to_sfixed(-368.0/65536.0,1,-nbitq), 
to_sfixed(-11813.0/65536.0,1,-nbitq), 
to_sfixed(-7647.0/65536.0,1,-nbitq), 
to_sfixed(-2099.0/65536.0,1,-nbitq), 
to_sfixed(3712.0/65536.0,1,-nbitq), 
to_sfixed(1490.0/65536.0,1,-nbitq), 
to_sfixed(-719.0/65536.0,1,-nbitq), 
to_sfixed(6170.0/65536.0,1,-nbitq), 
to_sfixed(7039.0/65536.0,1,-nbitq), 
to_sfixed(-3510.0/65536.0,1,-nbitq), 
to_sfixed(8500.0/65536.0,1,-nbitq), 
to_sfixed(-2549.0/65536.0,1,-nbitq), 
to_sfixed(-1120.0/65536.0,1,-nbitq), 
to_sfixed(-8474.0/65536.0,1,-nbitq), 
to_sfixed(6973.0/65536.0,1,-nbitq), 
to_sfixed(16268.0/65536.0,1,-nbitq), 
to_sfixed(1336.0/65536.0,1,-nbitq), 
to_sfixed(5235.0/65536.0,1,-nbitq), 
to_sfixed(659.0/65536.0,1,-nbitq), 
to_sfixed(476.0/65536.0,1,-nbitq), 
to_sfixed(-5403.0/65536.0,1,-nbitq), 
to_sfixed(-2712.0/65536.0,1,-nbitq), 
to_sfixed(-4038.0/65536.0,1,-nbitq), 
to_sfixed(-2097.0/65536.0,1,-nbitq), 
to_sfixed(-5861.0/65536.0,1,-nbitq), 
to_sfixed(-3005.0/65536.0,1,-nbitq), 
to_sfixed(-2149.0/65536.0,1,-nbitq), 
to_sfixed(-2688.0/65536.0,1,-nbitq), 
to_sfixed(91.0/65536.0,1,-nbitq), 
to_sfixed(-1658.0/65536.0,1,-nbitq), 
to_sfixed(2930.0/65536.0,1,-nbitq), 
to_sfixed(5382.0/65536.0,1,-nbitq), 
to_sfixed(-6459.0/65536.0,1,-nbitq), 
to_sfixed(-302.0/65536.0,1,-nbitq), 
to_sfixed(-4045.0/65536.0,1,-nbitq), 
to_sfixed(-3419.0/65536.0,1,-nbitq), 
to_sfixed(1440.0/65536.0,1,-nbitq), 
to_sfixed(2455.0/65536.0,1,-nbitq), 
to_sfixed(-2716.0/65536.0,1,-nbitq), 
to_sfixed(-973.0/65536.0,1,-nbitq), 
to_sfixed(1971.0/65536.0,1,-nbitq), 
to_sfixed(-7509.0/65536.0,1,-nbitq), 
to_sfixed(-5627.0/65536.0,1,-nbitq), 
to_sfixed(-3695.0/65536.0,1,-nbitq), 
to_sfixed(578.0/65536.0,1,-nbitq), 
to_sfixed(441.0/65536.0,1,-nbitq), 
to_sfixed(-7567.0/65536.0,1,-nbitq), 
to_sfixed(820.0/65536.0,1,-nbitq), 
to_sfixed(-1827.0/65536.0,1,-nbitq), 
to_sfixed(-7827.0/65536.0,1,-nbitq), 
to_sfixed(-2382.0/65536.0,1,-nbitq), 
to_sfixed(-2427.0/65536.0,1,-nbitq), 
to_sfixed(1380.0/65536.0,1,-nbitq), 
to_sfixed(4729.0/65536.0,1,-nbitq), 
to_sfixed(1382.0/65536.0,1,-nbitq), 
to_sfixed(1877.0/65536.0,1,-nbitq), 
to_sfixed(-2554.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4303.0/65536.0,1,-nbitq), 
to_sfixed(1390.0/65536.0,1,-nbitq), 
to_sfixed(3182.0/65536.0,1,-nbitq), 
to_sfixed(-3854.0/65536.0,1,-nbitq), 
to_sfixed(-6691.0/65536.0,1,-nbitq), 
to_sfixed(-2349.0/65536.0,1,-nbitq), 
to_sfixed(5718.0/65536.0,1,-nbitq), 
to_sfixed(-680.0/65536.0,1,-nbitq), 
to_sfixed(-6947.0/65536.0,1,-nbitq), 
to_sfixed(-597.0/65536.0,1,-nbitq), 
to_sfixed(-404.0/65536.0,1,-nbitq), 
to_sfixed(-8485.0/65536.0,1,-nbitq), 
to_sfixed(2323.0/65536.0,1,-nbitq), 
to_sfixed(-1663.0/65536.0,1,-nbitq), 
to_sfixed(1655.0/65536.0,1,-nbitq), 
to_sfixed(368.0/65536.0,1,-nbitq), 
to_sfixed(-1099.0/65536.0,1,-nbitq), 
to_sfixed(-622.0/65536.0,1,-nbitq), 
to_sfixed(-4613.0/65536.0,1,-nbitq), 
to_sfixed(13.0/65536.0,1,-nbitq), 
to_sfixed(-487.0/65536.0,1,-nbitq), 
to_sfixed(10195.0/65536.0,1,-nbitq), 
to_sfixed(3721.0/65536.0,1,-nbitq), 
to_sfixed(-1624.0/65536.0,1,-nbitq), 
to_sfixed(-10323.0/65536.0,1,-nbitq), 
to_sfixed(-1758.0/65536.0,1,-nbitq), 
to_sfixed(2928.0/65536.0,1,-nbitq), 
to_sfixed(1513.0/65536.0,1,-nbitq), 
to_sfixed(4939.0/65536.0,1,-nbitq), 
to_sfixed(1801.0/65536.0,1,-nbitq), 
to_sfixed(7126.0/65536.0,1,-nbitq), 
to_sfixed(15057.0/65536.0,1,-nbitq), 
to_sfixed(-1204.0/65536.0,1,-nbitq), 
to_sfixed(-2301.0/65536.0,1,-nbitq), 
to_sfixed(-2157.0/65536.0,1,-nbitq), 
to_sfixed(2909.0/65536.0,1,-nbitq), 
to_sfixed(-10662.0/65536.0,1,-nbitq), 
to_sfixed(9018.0/65536.0,1,-nbitq), 
to_sfixed(-1851.0/65536.0,1,-nbitq), 
to_sfixed(4354.0/65536.0,1,-nbitq), 
to_sfixed(5219.0/65536.0,1,-nbitq), 
to_sfixed(-49.0/65536.0,1,-nbitq), 
to_sfixed(5098.0/65536.0,1,-nbitq), 
to_sfixed(-11049.0/65536.0,1,-nbitq), 
to_sfixed(-1083.0/65536.0,1,-nbitq), 
to_sfixed(328.0/65536.0,1,-nbitq), 
to_sfixed(1425.0/65536.0,1,-nbitq), 
to_sfixed(-5810.0/65536.0,1,-nbitq), 
to_sfixed(380.0/65536.0,1,-nbitq), 
to_sfixed(2335.0/65536.0,1,-nbitq), 
to_sfixed(-1968.0/65536.0,1,-nbitq), 
to_sfixed(-4798.0/65536.0,1,-nbitq), 
to_sfixed(-4131.0/65536.0,1,-nbitq), 
to_sfixed(3483.0/65536.0,1,-nbitq), 
to_sfixed(2466.0/65536.0,1,-nbitq), 
to_sfixed(-261.0/65536.0,1,-nbitq), 
to_sfixed(1502.0/65536.0,1,-nbitq), 
to_sfixed(-2233.0/65536.0,1,-nbitq), 
to_sfixed(590.0/65536.0,1,-nbitq), 
to_sfixed(4718.0/65536.0,1,-nbitq), 
to_sfixed(365.0/65536.0,1,-nbitq), 
to_sfixed(-2639.0/65536.0,1,-nbitq), 
to_sfixed(-2437.0/65536.0,1,-nbitq), 
to_sfixed(2483.0/65536.0,1,-nbitq), 
to_sfixed(-7921.0/65536.0,1,-nbitq), 
to_sfixed(-8858.0/65536.0,1,-nbitq), 
to_sfixed(-339.0/65536.0,1,-nbitq), 
to_sfixed(-4541.0/65536.0,1,-nbitq), 
to_sfixed(-1218.0/65536.0,1,-nbitq), 
to_sfixed(-10098.0/65536.0,1,-nbitq), 
to_sfixed(2262.0/65536.0,1,-nbitq), 
to_sfixed(-5175.0/65536.0,1,-nbitq), 
to_sfixed(3568.0/65536.0,1,-nbitq), 
to_sfixed(-2429.0/65536.0,1,-nbitq), 
to_sfixed(1779.0/65536.0,1,-nbitq), 
to_sfixed(5896.0/65536.0,1,-nbitq), 
to_sfixed(3708.0/65536.0,1,-nbitq), 
to_sfixed(-3002.0/65536.0,1,-nbitq), 
to_sfixed(-488.0/65536.0,1,-nbitq), 
to_sfixed(-2793.0/65536.0,1,-nbitq)  ), 
( to_sfixed(221.0/65536.0,1,-nbitq), 
to_sfixed(-487.0/65536.0,1,-nbitq), 
to_sfixed(2911.0/65536.0,1,-nbitq), 
to_sfixed(-818.0/65536.0,1,-nbitq), 
to_sfixed(-6920.0/65536.0,1,-nbitq), 
to_sfixed(-1014.0/65536.0,1,-nbitq), 
to_sfixed(3805.0/65536.0,1,-nbitq), 
to_sfixed(-2225.0/65536.0,1,-nbitq), 
to_sfixed(-4971.0/65536.0,1,-nbitq), 
to_sfixed(-1165.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(-5972.0/65536.0,1,-nbitq), 
to_sfixed(3233.0/65536.0,1,-nbitq), 
to_sfixed(-476.0/65536.0,1,-nbitq), 
to_sfixed(3436.0/65536.0,1,-nbitq), 
to_sfixed(-1686.0/65536.0,1,-nbitq), 
to_sfixed(1835.0/65536.0,1,-nbitq), 
to_sfixed(-5322.0/65536.0,1,-nbitq), 
to_sfixed(-5572.0/65536.0,1,-nbitq), 
to_sfixed(1035.0/65536.0,1,-nbitq), 
to_sfixed(-2382.0/65536.0,1,-nbitq), 
to_sfixed(5054.0/65536.0,1,-nbitq), 
to_sfixed(7335.0/65536.0,1,-nbitq), 
to_sfixed(-6512.0/65536.0,1,-nbitq), 
to_sfixed(-10341.0/65536.0,1,-nbitq), 
to_sfixed(-5043.0/65536.0,1,-nbitq), 
to_sfixed(4075.0/65536.0,1,-nbitq), 
to_sfixed(2176.0/65536.0,1,-nbitq), 
to_sfixed(5620.0/65536.0,1,-nbitq), 
to_sfixed(5518.0/65536.0,1,-nbitq), 
to_sfixed(1674.0/65536.0,1,-nbitq), 
to_sfixed(17234.0/65536.0,1,-nbitq), 
to_sfixed(795.0/65536.0,1,-nbitq), 
to_sfixed(-6648.0/65536.0,1,-nbitq), 
to_sfixed(-2844.0/65536.0,1,-nbitq), 
to_sfixed(-2271.0/65536.0,1,-nbitq), 
to_sfixed(-6839.0/65536.0,1,-nbitq), 
to_sfixed(1674.0/65536.0,1,-nbitq), 
to_sfixed(-5882.0/65536.0,1,-nbitq), 
to_sfixed(-989.0/65536.0,1,-nbitq), 
to_sfixed(3644.0/65536.0,1,-nbitq), 
to_sfixed(-1302.0/65536.0,1,-nbitq), 
to_sfixed(5461.0/65536.0,1,-nbitq), 
to_sfixed(-7979.0/65536.0,1,-nbitq), 
to_sfixed(2458.0/65536.0,1,-nbitq), 
to_sfixed(-5781.0/65536.0,1,-nbitq), 
to_sfixed(499.0/65536.0,1,-nbitq), 
to_sfixed(-9148.0/65536.0,1,-nbitq), 
to_sfixed(2434.0/65536.0,1,-nbitq), 
to_sfixed(486.0/65536.0,1,-nbitq), 
to_sfixed(2776.0/65536.0,1,-nbitq), 
to_sfixed(-3408.0/65536.0,1,-nbitq), 
to_sfixed(2579.0/65536.0,1,-nbitq), 
to_sfixed(-7555.0/65536.0,1,-nbitq), 
to_sfixed(4184.0/65536.0,1,-nbitq), 
to_sfixed(135.0/65536.0,1,-nbitq), 
to_sfixed(227.0/65536.0,1,-nbitq), 
to_sfixed(-6328.0/65536.0,1,-nbitq), 
to_sfixed(-453.0/65536.0,1,-nbitq), 
to_sfixed(-1457.0/65536.0,1,-nbitq), 
to_sfixed(1335.0/65536.0,1,-nbitq), 
to_sfixed(2132.0/65536.0,1,-nbitq), 
to_sfixed(-1753.0/65536.0,1,-nbitq), 
to_sfixed(-688.0/65536.0,1,-nbitq), 
to_sfixed(-11992.0/65536.0,1,-nbitq), 
to_sfixed(-12116.0/65536.0,1,-nbitq), 
to_sfixed(2993.0/65536.0,1,-nbitq), 
to_sfixed(317.0/65536.0,1,-nbitq), 
to_sfixed(-5337.0/65536.0,1,-nbitq), 
to_sfixed(-8588.0/65536.0,1,-nbitq), 
to_sfixed(2427.0/65536.0,1,-nbitq), 
to_sfixed(-2777.0/65536.0,1,-nbitq), 
to_sfixed(4648.0/65536.0,1,-nbitq), 
to_sfixed(2248.0/65536.0,1,-nbitq), 
to_sfixed(-1716.0/65536.0,1,-nbitq), 
to_sfixed(2648.0/65536.0,1,-nbitq), 
to_sfixed(5764.0/65536.0,1,-nbitq), 
to_sfixed(-3383.0/65536.0,1,-nbitq), 
to_sfixed(-1550.0/65536.0,1,-nbitq), 
to_sfixed(945.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1775.0/65536.0,1,-nbitq), 
to_sfixed(-1343.0/65536.0,1,-nbitq), 
to_sfixed(6127.0/65536.0,1,-nbitq), 
to_sfixed(4399.0/65536.0,1,-nbitq), 
to_sfixed(-11458.0/65536.0,1,-nbitq), 
to_sfixed(-1758.0/65536.0,1,-nbitq), 
to_sfixed(8205.0/65536.0,1,-nbitq), 
to_sfixed(2500.0/65536.0,1,-nbitq), 
to_sfixed(-915.0/65536.0,1,-nbitq), 
to_sfixed(-2226.0/65536.0,1,-nbitq), 
to_sfixed(2426.0/65536.0,1,-nbitq), 
to_sfixed(-1938.0/65536.0,1,-nbitq), 
to_sfixed(224.0/65536.0,1,-nbitq), 
to_sfixed(1936.0/65536.0,1,-nbitq), 
to_sfixed(-2965.0/65536.0,1,-nbitq), 
to_sfixed(-2161.0/65536.0,1,-nbitq), 
to_sfixed(-1181.0/65536.0,1,-nbitq), 
to_sfixed(-5975.0/65536.0,1,-nbitq), 
to_sfixed(-4325.0/65536.0,1,-nbitq), 
to_sfixed(2080.0/65536.0,1,-nbitq), 
to_sfixed(-3025.0/65536.0,1,-nbitq), 
to_sfixed(7735.0/65536.0,1,-nbitq), 
to_sfixed(6485.0/65536.0,1,-nbitq), 
to_sfixed(-572.0/65536.0,1,-nbitq), 
to_sfixed(-10513.0/65536.0,1,-nbitq), 
to_sfixed(-11398.0/65536.0,1,-nbitq), 
to_sfixed(695.0/65536.0,1,-nbitq), 
to_sfixed(3237.0/65536.0,1,-nbitq), 
to_sfixed(2512.0/65536.0,1,-nbitq), 
to_sfixed(513.0/65536.0,1,-nbitq), 
to_sfixed(-9824.0/65536.0,1,-nbitq), 
to_sfixed(6012.0/65536.0,1,-nbitq), 
to_sfixed(253.0/65536.0,1,-nbitq), 
to_sfixed(-10611.0/65536.0,1,-nbitq), 
to_sfixed(-3338.0/65536.0,1,-nbitq), 
to_sfixed(-2540.0/65536.0,1,-nbitq), 
to_sfixed(-3047.0/65536.0,1,-nbitq), 
to_sfixed(1541.0/65536.0,1,-nbitq), 
to_sfixed(-2448.0/65536.0,1,-nbitq), 
to_sfixed(3834.0/65536.0,1,-nbitq), 
to_sfixed(103.0/65536.0,1,-nbitq), 
to_sfixed(-1656.0/65536.0,1,-nbitq), 
to_sfixed(663.0/65536.0,1,-nbitq), 
to_sfixed(-5023.0/65536.0,1,-nbitq), 
to_sfixed(2795.0/65536.0,1,-nbitq), 
to_sfixed(-423.0/65536.0,1,-nbitq), 
to_sfixed(-3955.0/65536.0,1,-nbitq), 
to_sfixed(-2980.0/65536.0,1,-nbitq), 
to_sfixed(-1367.0/65536.0,1,-nbitq), 
to_sfixed(2920.0/65536.0,1,-nbitq), 
to_sfixed(1209.0/65536.0,1,-nbitq), 
to_sfixed(5441.0/65536.0,1,-nbitq), 
to_sfixed(224.0/65536.0,1,-nbitq), 
to_sfixed(-6176.0/65536.0,1,-nbitq), 
to_sfixed(598.0/65536.0,1,-nbitq), 
to_sfixed(-1389.0/65536.0,1,-nbitq), 
to_sfixed(933.0/65536.0,1,-nbitq), 
to_sfixed(-8948.0/65536.0,1,-nbitq), 
to_sfixed(-3382.0/65536.0,1,-nbitq), 
to_sfixed(-8394.0/65536.0,1,-nbitq), 
to_sfixed(3224.0/65536.0,1,-nbitq), 
to_sfixed(-2650.0/65536.0,1,-nbitq), 
to_sfixed(2898.0/65536.0,1,-nbitq), 
to_sfixed(-2747.0/65536.0,1,-nbitq), 
to_sfixed(-7733.0/65536.0,1,-nbitq), 
to_sfixed(-9147.0/65536.0,1,-nbitq), 
to_sfixed(-1565.0/65536.0,1,-nbitq), 
to_sfixed(-1585.0/65536.0,1,-nbitq), 
to_sfixed(833.0/65536.0,1,-nbitq), 
to_sfixed(2470.0/65536.0,1,-nbitq), 
to_sfixed(6789.0/65536.0,1,-nbitq), 
to_sfixed(-5640.0/65536.0,1,-nbitq), 
to_sfixed(503.0/65536.0,1,-nbitq), 
to_sfixed(-2677.0/65536.0,1,-nbitq), 
to_sfixed(-121.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(4945.0/65536.0,1,-nbitq), 
to_sfixed(-3988.0/65536.0,1,-nbitq), 
to_sfixed(702.0/65536.0,1,-nbitq), 
to_sfixed(-923.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1136.0/65536.0,1,-nbitq), 
to_sfixed(-3448.0/65536.0,1,-nbitq), 
to_sfixed(10196.0/65536.0,1,-nbitq), 
to_sfixed(1788.0/65536.0,1,-nbitq), 
to_sfixed(-11564.0/65536.0,1,-nbitq), 
to_sfixed(-5292.0/65536.0,1,-nbitq), 
to_sfixed(6137.0/65536.0,1,-nbitq), 
to_sfixed(3293.0/65536.0,1,-nbitq), 
to_sfixed(-2795.0/65536.0,1,-nbitq), 
to_sfixed(-1952.0/65536.0,1,-nbitq), 
to_sfixed(-4789.0/65536.0,1,-nbitq), 
to_sfixed(-952.0/65536.0,1,-nbitq), 
to_sfixed(-1306.0/65536.0,1,-nbitq), 
to_sfixed(-3171.0/65536.0,1,-nbitq), 
to_sfixed(25.0/65536.0,1,-nbitq), 
to_sfixed(1949.0/65536.0,1,-nbitq), 
to_sfixed(-1265.0/65536.0,1,-nbitq), 
to_sfixed(-7394.0/65536.0,1,-nbitq), 
to_sfixed(-8079.0/65536.0,1,-nbitq), 
to_sfixed(1779.0/65536.0,1,-nbitq), 
to_sfixed(2264.0/65536.0,1,-nbitq), 
to_sfixed(7759.0/65536.0,1,-nbitq), 
to_sfixed(6972.0/65536.0,1,-nbitq), 
to_sfixed(-3124.0/65536.0,1,-nbitq), 
to_sfixed(-2620.0/65536.0,1,-nbitq), 
to_sfixed(-14064.0/65536.0,1,-nbitq), 
to_sfixed(-6860.0/65536.0,1,-nbitq), 
to_sfixed(493.0/65536.0,1,-nbitq), 
to_sfixed(-626.0/65536.0,1,-nbitq), 
to_sfixed(4098.0/65536.0,1,-nbitq), 
to_sfixed(-1050.0/65536.0,1,-nbitq), 
to_sfixed(7915.0/65536.0,1,-nbitq), 
to_sfixed(-2225.0/65536.0,1,-nbitq), 
to_sfixed(-7925.0/65536.0,1,-nbitq), 
to_sfixed(2162.0/65536.0,1,-nbitq), 
to_sfixed(-1182.0/65536.0,1,-nbitq), 
to_sfixed(-576.0/65536.0,1,-nbitq), 
to_sfixed(-5792.0/65536.0,1,-nbitq), 
to_sfixed(-980.0/65536.0,1,-nbitq), 
to_sfixed(2562.0/65536.0,1,-nbitq), 
to_sfixed(4906.0/65536.0,1,-nbitq), 
to_sfixed(1699.0/65536.0,1,-nbitq), 
to_sfixed(1258.0/65536.0,1,-nbitq), 
to_sfixed(-6402.0/65536.0,1,-nbitq), 
to_sfixed(12.0/65536.0,1,-nbitq), 
to_sfixed(2157.0/65536.0,1,-nbitq), 
to_sfixed(-4852.0/65536.0,1,-nbitq), 
to_sfixed(1159.0/65536.0,1,-nbitq), 
to_sfixed(-2758.0/65536.0,1,-nbitq), 
to_sfixed(-23.0/65536.0,1,-nbitq), 
to_sfixed(2267.0/65536.0,1,-nbitq), 
to_sfixed(5967.0/65536.0,1,-nbitq), 
to_sfixed(638.0/65536.0,1,-nbitq), 
to_sfixed(-2608.0/65536.0,1,-nbitq), 
to_sfixed(600.0/65536.0,1,-nbitq), 
to_sfixed(2683.0/65536.0,1,-nbitq), 
to_sfixed(1614.0/65536.0,1,-nbitq), 
to_sfixed(-6466.0/65536.0,1,-nbitq), 
to_sfixed(-806.0/65536.0,1,-nbitq), 
to_sfixed(-9460.0/65536.0,1,-nbitq), 
to_sfixed(3513.0/65536.0,1,-nbitq), 
to_sfixed(-1371.0/65536.0,1,-nbitq), 
to_sfixed(1187.0/65536.0,1,-nbitq), 
to_sfixed(-470.0/65536.0,1,-nbitq), 
to_sfixed(-322.0/65536.0,1,-nbitq), 
to_sfixed(-6939.0/65536.0,1,-nbitq), 
to_sfixed(-432.0/65536.0,1,-nbitq), 
to_sfixed(-7788.0/65536.0,1,-nbitq), 
to_sfixed(2647.0/65536.0,1,-nbitq), 
to_sfixed(3603.0/65536.0,1,-nbitq), 
to_sfixed(3059.0/65536.0,1,-nbitq), 
to_sfixed(4878.0/65536.0,1,-nbitq), 
to_sfixed(1186.0/65536.0,1,-nbitq), 
to_sfixed(-2736.0/65536.0,1,-nbitq), 
to_sfixed(-533.0/65536.0,1,-nbitq), 
to_sfixed(-6242.0/65536.0,1,-nbitq), 
to_sfixed(-5313.0/65536.0,1,-nbitq), 
to_sfixed(4796.0/65536.0,1,-nbitq), 
to_sfixed(-1466.0/65536.0,1,-nbitq), 
to_sfixed(-2384.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2476.0/65536.0,1,-nbitq), 
to_sfixed(-2428.0/65536.0,1,-nbitq), 
to_sfixed(8502.0/65536.0,1,-nbitq), 
to_sfixed(1607.0/65536.0,1,-nbitq), 
to_sfixed(1448.0/65536.0,1,-nbitq), 
to_sfixed(-2499.0/65536.0,1,-nbitq), 
to_sfixed(4338.0/65536.0,1,-nbitq), 
to_sfixed(716.0/65536.0,1,-nbitq), 
to_sfixed(-3206.0/65536.0,1,-nbitq), 
to_sfixed(-2485.0/65536.0,1,-nbitq), 
to_sfixed(-1914.0/65536.0,1,-nbitq), 
to_sfixed(1787.0/65536.0,1,-nbitq), 
to_sfixed(1256.0/65536.0,1,-nbitq), 
to_sfixed(-4705.0/65536.0,1,-nbitq), 
to_sfixed(2807.0/65536.0,1,-nbitq), 
to_sfixed(1300.0/65536.0,1,-nbitq), 
to_sfixed(263.0/65536.0,1,-nbitq), 
to_sfixed(-8059.0/65536.0,1,-nbitq), 
to_sfixed(-9809.0/65536.0,1,-nbitq), 
to_sfixed(-2051.0/65536.0,1,-nbitq), 
to_sfixed(1701.0/65536.0,1,-nbitq), 
to_sfixed(8934.0/65536.0,1,-nbitq), 
to_sfixed(-1263.0/65536.0,1,-nbitq), 
to_sfixed(-10783.0/65536.0,1,-nbitq), 
to_sfixed(-3385.0/65536.0,1,-nbitq), 
to_sfixed(-10780.0/65536.0,1,-nbitq), 
to_sfixed(-4149.0/65536.0,1,-nbitq), 
to_sfixed(-2295.0/65536.0,1,-nbitq), 
to_sfixed(6188.0/65536.0,1,-nbitq), 
to_sfixed(2074.0/65536.0,1,-nbitq), 
to_sfixed(-1620.0/65536.0,1,-nbitq), 
to_sfixed(5565.0/65536.0,1,-nbitq), 
to_sfixed(951.0/65536.0,1,-nbitq), 
to_sfixed(188.0/65536.0,1,-nbitq), 
to_sfixed(2924.0/65536.0,1,-nbitq), 
to_sfixed(-3235.0/65536.0,1,-nbitq), 
to_sfixed(2153.0/65536.0,1,-nbitq), 
to_sfixed(-4976.0/65536.0,1,-nbitq), 
to_sfixed(-412.0/65536.0,1,-nbitq), 
to_sfixed(2358.0/65536.0,1,-nbitq), 
to_sfixed(3812.0/65536.0,1,-nbitq), 
to_sfixed(556.0/65536.0,1,-nbitq), 
to_sfixed(-552.0/65536.0,1,-nbitq), 
to_sfixed(-8318.0/65536.0,1,-nbitq), 
to_sfixed(1660.0/65536.0,1,-nbitq), 
to_sfixed(-1675.0/65536.0,1,-nbitq), 
to_sfixed(775.0/65536.0,1,-nbitq), 
to_sfixed(2338.0/65536.0,1,-nbitq), 
to_sfixed(476.0/65536.0,1,-nbitq), 
to_sfixed(397.0/65536.0,1,-nbitq), 
to_sfixed(202.0/65536.0,1,-nbitq), 
to_sfixed(3993.0/65536.0,1,-nbitq), 
to_sfixed(-8561.0/65536.0,1,-nbitq), 
to_sfixed(1420.0/65536.0,1,-nbitq), 
to_sfixed(-1529.0/65536.0,1,-nbitq), 
to_sfixed(-2293.0/65536.0,1,-nbitq), 
to_sfixed(1161.0/65536.0,1,-nbitq), 
to_sfixed(2277.0/65536.0,1,-nbitq), 
to_sfixed(-653.0/65536.0,1,-nbitq), 
to_sfixed(-3715.0/65536.0,1,-nbitq), 
to_sfixed(4387.0/65536.0,1,-nbitq), 
to_sfixed(2256.0/65536.0,1,-nbitq), 
to_sfixed(936.0/65536.0,1,-nbitq), 
to_sfixed(866.0/65536.0,1,-nbitq), 
to_sfixed(-6589.0/65536.0,1,-nbitq), 
to_sfixed(-6278.0/65536.0,1,-nbitq), 
to_sfixed(-1663.0/65536.0,1,-nbitq), 
to_sfixed(-7852.0/65536.0,1,-nbitq), 
to_sfixed(2251.0/65536.0,1,-nbitq), 
to_sfixed(11600.0/65536.0,1,-nbitq), 
to_sfixed(-691.0/65536.0,1,-nbitq), 
to_sfixed(5549.0/65536.0,1,-nbitq), 
to_sfixed(1857.0/65536.0,1,-nbitq), 
to_sfixed(-1532.0/65536.0,1,-nbitq), 
to_sfixed(2328.0/65536.0,1,-nbitq), 
to_sfixed(148.0/65536.0,1,-nbitq), 
to_sfixed(-11760.0/65536.0,1,-nbitq), 
to_sfixed(1968.0/65536.0,1,-nbitq), 
to_sfixed(-3039.0/65536.0,1,-nbitq), 
to_sfixed(-4609.0/65536.0,1,-nbitq)  ), 
( to_sfixed(416.0/65536.0,1,-nbitq), 
to_sfixed(-1476.0/65536.0,1,-nbitq), 
to_sfixed(9351.0/65536.0,1,-nbitq), 
to_sfixed(-846.0/65536.0,1,-nbitq), 
to_sfixed(-2175.0/65536.0,1,-nbitq), 
to_sfixed(-6569.0/65536.0,1,-nbitq), 
to_sfixed(1712.0/65536.0,1,-nbitq), 
to_sfixed(-1083.0/65536.0,1,-nbitq), 
to_sfixed(-988.0/65536.0,1,-nbitq), 
to_sfixed(1031.0/65536.0,1,-nbitq), 
to_sfixed(-4436.0/65536.0,1,-nbitq), 
to_sfixed(-1486.0/65536.0,1,-nbitq), 
to_sfixed(-2182.0/65536.0,1,-nbitq), 
to_sfixed(-9524.0/65536.0,1,-nbitq), 
to_sfixed(457.0/65536.0,1,-nbitq), 
to_sfixed(630.0/65536.0,1,-nbitq), 
to_sfixed(1770.0/65536.0,1,-nbitq), 
to_sfixed(-2677.0/65536.0,1,-nbitq), 
to_sfixed(-3393.0/65536.0,1,-nbitq), 
to_sfixed(-896.0/65536.0,1,-nbitq), 
to_sfixed(3456.0/65536.0,1,-nbitq), 
to_sfixed(2077.0/65536.0,1,-nbitq), 
to_sfixed(5740.0/65536.0,1,-nbitq), 
to_sfixed(-5876.0/65536.0,1,-nbitq), 
to_sfixed(-3591.0/65536.0,1,-nbitq), 
to_sfixed(-9718.0/65536.0,1,-nbitq), 
to_sfixed(-4981.0/65536.0,1,-nbitq), 
to_sfixed(-626.0/65536.0,1,-nbitq), 
to_sfixed(4393.0/65536.0,1,-nbitq), 
to_sfixed(2946.0/65536.0,1,-nbitq), 
to_sfixed(-5130.0/65536.0,1,-nbitq), 
to_sfixed(1250.0/65536.0,1,-nbitq), 
to_sfixed(-1873.0/65536.0,1,-nbitq), 
to_sfixed(164.0/65536.0,1,-nbitq), 
to_sfixed(414.0/65536.0,1,-nbitq), 
to_sfixed(-435.0/65536.0,1,-nbitq), 
to_sfixed(1214.0/65536.0,1,-nbitq), 
to_sfixed(-3233.0/65536.0,1,-nbitq), 
to_sfixed(3507.0/65536.0,1,-nbitq), 
to_sfixed(3515.0/65536.0,1,-nbitq), 
to_sfixed(1848.0/65536.0,1,-nbitq), 
to_sfixed(-1745.0/65536.0,1,-nbitq), 
to_sfixed(860.0/65536.0,1,-nbitq), 
to_sfixed(-4666.0/65536.0,1,-nbitq), 
to_sfixed(1495.0/65536.0,1,-nbitq), 
to_sfixed(-5419.0/65536.0,1,-nbitq), 
to_sfixed(789.0/65536.0,1,-nbitq), 
to_sfixed(1035.0/65536.0,1,-nbitq), 
to_sfixed(-834.0/65536.0,1,-nbitq), 
to_sfixed(63.0/65536.0,1,-nbitq), 
to_sfixed(569.0/65536.0,1,-nbitq), 
to_sfixed(2322.0/65536.0,1,-nbitq), 
to_sfixed(-11938.0/65536.0,1,-nbitq), 
to_sfixed(5417.0/65536.0,1,-nbitq), 
to_sfixed(-1279.0/65536.0,1,-nbitq), 
to_sfixed(-1865.0/65536.0,1,-nbitq), 
to_sfixed(296.0/65536.0,1,-nbitq), 
to_sfixed(5396.0/65536.0,1,-nbitq), 
to_sfixed(-2762.0/65536.0,1,-nbitq), 
to_sfixed(-8405.0/65536.0,1,-nbitq), 
to_sfixed(1058.0/65536.0,1,-nbitq), 
to_sfixed(784.0/65536.0,1,-nbitq), 
to_sfixed(1747.0/65536.0,1,-nbitq), 
to_sfixed(-2341.0/65536.0,1,-nbitq), 
to_sfixed(349.0/65536.0,1,-nbitq), 
to_sfixed(-3318.0/65536.0,1,-nbitq), 
to_sfixed(51.0/65536.0,1,-nbitq), 
to_sfixed(921.0/65536.0,1,-nbitq), 
to_sfixed(3490.0/65536.0,1,-nbitq), 
to_sfixed(8217.0/65536.0,1,-nbitq), 
to_sfixed(-2472.0/65536.0,1,-nbitq), 
to_sfixed(6871.0/65536.0,1,-nbitq), 
to_sfixed(901.0/65536.0,1,-nbitq), 
to_sfixed(-668.0/65536.0,1,-nbitq), 
to_sfixed(1571.0/65536.0,1,-nbitq), 
to_sfixed(2783.0/65536.0,1,-nbitq), 
to_sfixed(-8598.0/65536.0,1,-nbitq), 
to_sfixed(3521.0/65536.0,1,-nbitq), 
to_sfixed(285.0/65536.0,1,-nbitq), 
to_sfixed(-2443.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2242.0/65536.0,1,-nbitq), 
to_sfixed(-1438.0/65536.0,1,-nbitq), 
to_sfixed(7304.0/65536.0,1,-nbitq), 
to_sfixed(4935.0/65536.0,1,-nbitq), 
to_sfixed(-3456.0/65536.0,1,-nbitq), 
to_sfixed(-1464.0/65536.0,1,-nbitq), 
to_sfixed(221.0/65536.0,1,-nbitq), 
to_sfixed(1328.0/65536.0,1,-nbitq), 
to_sfixed(-2129.0/65536.0,1,-nbitq), 
to_sfixed(-2711.0/65536.0,1,-nbitq), 
to_sfixed(1254.0/65536.0,1,-nbitq), 
to_sfixed(-4203.0/65536.0,1,-nbitq), 
to_sfixed(2854.0/65536.0,1,-nbitq), 
to_sfixed(-5425.0/65536.0,1,-nbitq), 
to_sfixed(555.0/65536.0,1,-nbitq), 
to_sfixed(1470.0/65536.0,1,-nbitq), 
to_sfixed(-2815.0/65536.0,1,-nbitq), 
to_sfixed(-2489.0/65536.0,1,-nbitq), 
to_sfixed(-1108.0/65536.0,1,-nbitq), 
to_sfixed(-1059.0/65536.0,1,-nbitq), 
to_sfixed(122.0/65536.0,1,-nbitq), 
to_sfixed(2061.0/65536.0,1,-nbitq), 
to_sfixed(4056.0/65536.0,1,-nbitq), 
to_sfixed(-2896.0/65536.0,1,-nbitq), 
to_sfixed(-3688.0/65536.0,1,-nbitq), 
to_sfixed(-4969.0/65536.0,1,-nbitq), 
to_sfixed(-660.0/65536.0,1,-nbitq), 
to_sfixed(522.0/65536.0,1,-nbitq), 
to_sfixed(2337.0/65536.0,1,-nbitq), 
to_sfixed(1878.0/65536.0,1,-nbitq), 
to_sfixed(-9204.0/65536.0,1,-nbitq), 
to_sfixed(-1123.0/65536.0,1,-nbitq), 
to_sfixed(2337.0/65536.0,1,-nbitq), 
to_sfixed(-1989.0/65536.0,1,-nbitq), 
to_sfixed(1823.0/65536.0,1,-nbitq), 
to_sfixed(1558.0/65536.0,1,-nbitq), 
to_sfixed(-2948.0/65536.0,1,-nbitq), 
to_sfixed(-3249.0/65536.0,1,-nbitq), 
to_sfixed(2452.0/65536.0,1,-nbitq), 
to_sfixed(-344.0/65536.0,1,-nbitq), 
to_sfixed(-471.0/65536.0,1,-nbitq), 
to_sfixed(-3192.0/65536.0,1,-nbitq), 
to_sfixed(-813.0/65536.0,1,-nbitq), 
to_sfixed(-5192.0/65536.0,1,-nbitq), 
to_sfixed(-714.0/65536.0,1,-nbitq), 
to_sfixed(2741.0/65536.0,1,-nbitq), 
to_sfixed(354.0/65536.0,1,-nbitq), 
to_sfixed(2248.0/65536.0,1,-nbitq), 
to_sfixed(-210.0/65536.0,1,-nbitq), 
to_sfixed(4095.0/65536.0,1,-nbitq), 
to_sfixed(-1183.0/65536.0,1,-nbitq), 
to_sfixed(3124.0/65536.0,1,-nbitq), 
to_sfixed(-5625.0/65536.0,1,-nbitq), 
to_sfixed(6415.0/65536.0,1,-nbitq), 
to_sfixed(-2327.0/65536.0,1,-nbitq), 
to_sfixed(-3573.0/65536.0,1,-nbitq), 
to_sfixed(-2571.0/65536.0,1,-nbitq), 
to_sfixed(5061.0/65536.0,1,-nbitq), 
to_sfixed(880.0/65536.0,1,-nbitq), 
to_sfixed(-4465.0/65536.0,1,-nbitq), 
to_sfixed(6002.0/65536.0,1,-nbitq), 
to_sfixed(-655.0/65536.0,1,-nbitq), 
to_sfixed(183.0/65536.0,1,-nbitq), 
to_sfixed(664.0/65536.0,1,-nbitq), 
to_sfixed(2539.0/65536.0,1,-nbitq), 
to_sfixed(631.0/65536.0,1,-nbitq), 
to_sfixed(1957.0/65536.0,1,-nbitq), 
to_sfixed(783.0/65536.0,1,-nbitq), 
to_sfixed(3056.0/65536.0,1,-nbitq), 
to_sfixed(8721.0/65536.0,1,-nbitq), 
to_sfixed(-1368.0/65536.0,1,-nbitq), 
to_sfixed(4090.0/65536.0,1,-nbitq), 
to_sfixed(4236.0/65536.0,1,-nbitq), 
to_sfixed(1717.0/65536.0,1,-nbitq), 
to_sfixed(-2050.0/65536.0,1,-nbitq), 
to_sfixed(-1238.0/65536.0,1,-nbitq), 
to_sfixed(-7337.0/65536.0,1,-nbitq), 
to_sfixed(4999.0/65536.0,1,-nbitq), 
to_sfixed(1338.0/65536.0,1,-nbitq), 
to_sfixed(-3616.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-153.0/65536.0,1,-nbitq), 
to_sfixed(1617.0/65536.0,1,-nbitq), 
to_sfixed(4997.0/65536.0,1,-nbitq), 
to_sfixed(1161.0/65536.0,1,-nbitq), 
to_sfixed(-2163.0/65536.0,1,-nbitq), 
to_sfixed(-68.0/65536.0,1,-nbitq), 
to_sfixed(2301.0/65536.0,1,-nbitq), 
to_sfixed(4819.0/65536.0,1,-nbitq), 
to_sfixed(-3773.0/65536.0,1,-nbitq), 
to_sfixed(-326.0/65536.0,1,-nbitq), 
to_sfixed(4121.0/65536.0,1,-nbitq), 
to_sfixed(-4739.0/65536.0,1,-nbitq), 
to_sfixed(884.0/65536.0,1,-nbitq), 
to_sfixed(-5461.0/65536.0,1,-nbitq), 
to_sfixed(2219.0/65536.0,1,-nbitq), 
to_sfixed(-310.0/65536.0,1,-nbitq), 
to_sfixed(2118.0/65536.0,1,-nbitq), 
to_sfixed(-7146.0/65536.0,1,-nbitq), 
to_sfixed(-6006.0/65536.0,1,-nbitq), 
to_sfixed(-468.0/65536.0,1,-nbitq), 
to_sfixed(2173.0/65536.0,1,-nbitq), 
to_sfixed(3275.0/65536.0,1,-nbitq), 
to_sfixed(3811.0/65536.0,1,-nbitq), 
to_sfixed(-8042.0/65536.0,1,-nbitq), 
to_sfixed(-4501.0/65536.0,1,-nbitq), 
to_sfixed(-4166.0/65536.0,1,-nbitq), 
to_sfixed(-6513.0/65536.0,1,-nbitq), 
to_sfixed(-1037.0/65536.0,1,-nbitq), 
to_sfixed(5296.0/65536.0,1,-nbitq), 
to_sfixed(887.0/65536.0,1,-nbitq), 
to_sfixed(-2813.0/65536.0,1,-nbitq), 
to_sfixed(-4655.0/65536.0,1,-nbitq), 
to_sfixed(3083.0/65536.0,1,-nbitq), 
to_sfixed(-744.0/65536.0,1,-nbitq), 
to_sfixed(-1455.0/65536.0,1,-nbitq), 
to_sfixed(889.0/65536.0,1,-nbitq), 
to_sfixed(-64.0/65536.0,1,-nbitq), 
to_sfixed(-5097.0/65536.0,1,-nbitq), 
to_sfixed(-1518.0/65536.0,1,-nbitq), 
to_sfixed(1018.0/65536.0,1,-nbitq), 
to_sfixed(476.0/65536.0,1,-nbitq), 
to_sfixed(389.0/65536.0,1,-nbitq), 
to_sfixed(5194.0/65536.0,1,-nbitq), 
to_sfixed(-9485.0/65536.0,1,-nbitq), 
to_sfixed(-822.0/65536.0,1,-nbitq), 
to_sfixed(3724.0/65536.0,1,-nbitq), 
to_sfixed(-504.0/65536.0,1,-nbitq), 
to_sfixed(5004.0/65536.0,1,-nbitq), 
to_sfixed(1305.0/65536.0,1,-nbitq), 
to_sfixed(3073.0/65536.0,1,-nbitq), 
to_sfixed(1086.0/65536.0,1,-nbitq), 
to_sfixed(-670.0/65536.0,1,-nbitq), 
to_sfixed(-3580.0/65536.0,1,-nbitq), 
to_sfixed(8961.0/65536.0,1,-nbitq), 
to_sfixed(-7412.0/65536.0,1,-nbitq), 
to_sfixed(-2017.0/65536.0,1,-nbitq), 
to_sfixed(2346.0/65536.0,1,-nbitq), 
to_sfixed(2997.0/65536.0,1,-nbitq), 
to_sfixed(-204.0/65536.0,1,-nbitq), 
to_sfixed(-3950.0/65536.0,1,-nbitq), 
to_sfixed(3244.0/65536.0,1,-nbitq), 
to_sfixed(-1592.0/65536.0,1,-nbitq), 
to_sfixed(1350.0/65536.0,1,-nbitq), 
to_sfixed(-2935.0/65536.0,1,-nbitq), 
to_sfixed(5704.0/65536.0,1,-nbitq), 
to_sfixed(1538.0/65536.0,1,-nbitq), 
to_sfixed(2911.0/65536.0,1,-nbitq), 
to_sfixed(1817.0/65536.0,1,-nbitq), 
to_sfixed(3693.0/65536.0,1,-nbitq), 
to_sfixed(6525.0/65536.0,1,-nbitq), 
to_sfixed(-1837.0/65536.0,1,-nbitq), 
to_sfixed(2154.0/65536.0,1,-nbitq), 
to_sfixed(2966.0/65536.0,1,-nbitq), 
to_sfixed(1740.0/65536.0,1,-nbitq), 
to_sfixed(1900.0/65536.0,1,-nbitq), 
to_sfixed(1869.0/65536.0,1,-nbitq), 
to_sfixed(-4636.0/65536.0,1,-nbitq), 
to_sfixed(1080.0/65536.0,1,-nbitq), 
to_sfixed(-1190.0/65536.0,1,-nbitq), 
to_sfixed(-193.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1661.0/65536.0,1,-nbitq), 
to_sfixed(-3052.0/65536.0,1,-nbitq), 
to_sfixed(96.0/65536.0,1,-nbitq), 
to_sfixed(453.0/65536.0,1,-nbitq), 
to_sfixed(214.0/65536.0,1,-nbitq), 
to_sfixed(-41.0/65536.0,1,-nbitq), 
to_sfixed(1797.0/65536.0,1,-nbitq), 
to_sfixed(-474.0/65536.0,1,-nbitq), 
to_sfixed(674.0/65536.0,1,-nbitq), 
to_sfixed(-1032.0/65536.0,1,-nbitq), 
to_sfixed(991.0/65536.0,1,-nbitq), 
to_sfixed(-4139.0/65536.0,1,-nbitq), 
to_sfixed(2412.0/65536.0,1,-nbitq), 
to_sfixed(-4861.0/65536.0,1,-nbitq), 
to_sfixed(-4415.0/65536.0,1,-nbitq), 
to_sfixed(2177.0/65536.0,1,-nbitq), 
to_sfixed(1865.0/65536.0,1,-nbitq), 
to_sfixed(-11147.0/65536.0,1,-nbitq), 
to_sfixed(-1361.0/65536.0,1,-nbitq), 
to_sfixed(1253.0/65536.0,1,-nbitq), 
to_sfixed(1544.0/65536.0,1,-nbitq), 
to_sfixed(3523.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(-7868.0/65536.0,1,-nbitq), 
to_sfixed(-4064.0/65536.0,1,-nbitq), 
to_sfixed(-3153.0/65536.0,1,-nbitq), 
to_sfixed(-2110.0/65536.0,1,-nbitq), 
to_sfixed(-1333.0/65536.0,1,-nbitq), 
to_sfixed(2415.0/65536.0,1,-nbitq), 
to_sfixed(2956.0/65536.0,1,-nbitq), 
to_sfixed(936.0/65536.0,1,-nbitq), 
to_sfixed(-2834.0/65536.0,1,-nbitq), 
to_sfixed(5357.0/65536.0,1,-nbitq), 
to_sfixed(-259.0/65536.0,1,-nbitq), 
to_sfixed(-2244.0/65536.0,1,-nbitq), 
to_sfixed(-1628.0/65536.0,1,-nbitq), 
to_sfixed(-2552.0/65536.0,1,-nbitq), 
to_sfixed(-1332.0/65536.0,1,-nbitq), 
to_sfixed(-2684.0/65536.0,1,-nbitq), 
to_sfixed(-1757.0/65536.0,1,-nbitq), 
to_sfixed(3292.0/65536.0,1,-nbitq), 
to_sfixed(-33.0/65536.0,1,-nbitq), 
to_sfixed(3490.0/65536.0,1,-nbitq), 
to_sfixed(-1330.0/65536.0,1,-nbitq), 
to_sfixed(3135.0/65536.0,1,-nbitq), 
to_sfixed(2808.0/65536.0,1,-nbitq), 
to_sfixed(2181.0/65536.0,1,-nbitq), 
to_sfixed(2601.0/65536.0,1,-nbitq), 
to_sfixed(-1077.0/65536.0,1,-nbitq), 
to_sfixed(-927.0/65536.0,1,-nbitq), 
to_sfixed(1451.0/65536.0,1,-nbitq), 
to_sfixed(2434.0/65536.0,1,-nbitq), 
to_sfixed(-3028.0/65536.0,1,-nbitq), 
to_sfixed(5534.0/65536.0,1,-nbitq), 
to_sfixed(-1874.0/65536.0,1,-nbitq), 
to_sfixed(-200.0/65536.0,1,-nbitq), 
to_sfixed(657.0/65536.0,1,-nbitq), 
to_sfixed(-74.0/65536.0,1,-nbitq), 
to_sfixed(2781.0/65536.0,1,-nbitq), 
to_sfixed(-1320.0/65536.0,1,-nbitq), 
to_sfixed(3566.0/65536.0,1,-nbitq), 
to_sfixed(270.0/65536.0,1,-nbitq), 
to_sfixed(749.0/65536.0,1,-nbitq), 
to_sfixed(-2534.0/65536.0,1,-nbitq), 
to_sfixed(-266.0/65536.0,1,-nbitq), 
to_sfixed(-1929.0/65536.0,1,-nbitq), 
to_sfixed(1174.0/65536.0,1,-nbitq), 
to_sfixed(1653.0/65536.0,1,-nbitq), 
to_sfixed(9217.0/65536.0,1,-nbitq), 
to_sfixed(5365.0/65536.0,1,-nbitq), 
to_sfixed(2624.0/65536.0,1,-nbitq), 
to_sfixed(-2996.0/65536.0,1,-nbitq), 
to_sfixed(4480.0/65536.0,1,-nbitq), 
to_sfixed(2064.0/65536.0,1,-nbitq), 
to_sfixed(817.0/65536.0,1,-nbitq), 
to_sfixed(3374.0/65536.0,1,-nbitq), 
to_sfixed(-8480.0/65536.0,1,-nbitq), 
to_sfixed(-882.0/65536.0,1,-nbitq), 
to_sfixed(2719.0/65536.0,1,-nbitq), 
to_sfixed(1465.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1452.0/65536.0,1,-nbitq), 
to_sfixed(2724.0/65536.0,1,-nbitq), 
to_sfixed(1077.0/65536.0,1,-nbitq), 
to_sfixed(1301.0/65536.0,1,-nbitq), 
to_sfixed(-5245.0/65536.0,1,-nbitq), 
to_sfixed(-2298.0/65536.0,1,-nbitq), 
to_sfixed(-359.0/65536.0,1,-nbitq), 
to_sfixed(-1333.0/65536.0,1,-nbitq), 
to_sfixed(-2140.0/65536.0,1,-nbitq), 
to_sfixed(1477.0/65536.0,1,-nbitq), 
to_sfixed(-1006.0/65536.0,1,-nbitq), 
to_sfixed(165.0/65536.0,1,-nbitq), 
to_sfixed(458.0/65536.0,1,-nbitq), 
to_sfixed(-994.0/65536.0,1,-nbitq), 
to_sfixed(-1851.0/65536.0,1,-nbitq), 
to_sfixed(-2831.0/65536.0,1,-nbitq), 
to_sfixed(2157.0/65536.0,1,-nbitq), 
to_sfixed(2057.0/65536.0,1,-nbitq), 
to_sfixed(-1088.0/65536.0,1,-nbitq), 
to_sfixed(-1656.0/65536.0,1,-nbitq), 
to_sfixed(-1178.0/65536.0,1,-nbitq), 
to_sfixed(3633.0/65536.0,1,-nbitq), 
to_sfixed(-1719.0/65536.0,1,-nbitq), 
to_sfixed(-1790.0/65536.0,1,-nbitq), 
to_sfixed(-2942.0/65536.0,1,-nbitq), 
to_sfixed(-1007.0/65536.0,1,-nbitq), 
to_sfixed(-2483.0/65536.0,1,-nbitq), 
to_sfixed(-2125.0/65536.0,1,-nbitq), 
to_sfixed(4215.0/65536.0,1,-nbitq), 
to_sfixed(-2747.0/65536.0,1,-nbitq), 
to_sfixed(-3809.0/65536.0,1,-nbitq), 
to_sfixed(-1193.0/65536.0,1,-nbitq), 
to_sfixed(232.0/65536.0,1,-nbitq), 
to_sfixed(885.0/65536.0,1,-nbitq), 
to_sfixed(-2296.0/65536.0,1,-nbitq), 
to_sfixed(2426.0/65536.0,1,-nbitq), 
to_sfixed(-3631.0/65536.0,1,-nbitq), 
to_sfixed(-687.0/65536.0,1,-nbitq), 
to_sfixed(-3863.0/65536.0,1,-nbitq), 
to_sfixed(217.0/65536.0,1,-nbitq), 
to_sfixed(2871.0/65536.0,1,-nbitq), 
to_sfixed(-454.0/65536.0,1,-nbitq), 
to_sfixed(1444.0/65536.0,1,-nbitq), 
to_sfixed(-155.0/65536.0,1,-nbitq), 
to_sfixed(640.0/65536.0,1,-nbitq), 
to_sfixed(2822.0/65536.0,1,-nbitq), 
to_sfixed(-1162.0/65536.0,1,-nbitq), 
to_sfixed(2878.0/65536.0,1,-nbitq), 
to_sfixed(1321.0/65536.0,1,-nbitq), 
to_sfixed(-313.0/65536.0,1,-nbitq), 
to_sfixed(3319.0/65536.0,1,-nbitq), 
to_sfixed(-1219.0/65536.0,1,-nbitq), 
to_sfixed(-2506.0/65536.0,1,-nbitq), 
to_sfixed(5836.0/65536.0,1,-nbitq), 
to_sfixed(29.0/65536.0,1,-nbitq), 
to_sfixed(322.0/65536.0,1,-nbitq), 
to_sfixed(-1580.0/65536.0,1,-nbitq), 
to_sfixed(820.0/65536.0,1,-nbitq), 
to_sfixed(-1001.0/65536.0,1,-nbitq), 
to_sfixed(1688.0/65536.0,1,-nbitq), 
to_sfixed(2640.0/65536.0,1,-nbitq), 
to_sfixed(-1451.0/65536.0,1,-nbitq), 
to_sfixed(3042.0/65536.0,1,-nbitq), 
to_sfixed(231.0/65536.0,1,-nbitq), 
to_sfixed(-1466.0/65536.0,1,-nbitq), 
to_sfixed(-592.0/65536.0,1,-nbitq), 
to_sfixed(173.0/65536.0,1,-nbitq), 
to_sfixed(1359.0/65536.0,1,-nbitq), 
to_sfixed(4720.0/65536.0,1,-nbitq), 
to_sfixed(2907.0/65536.0,1,-nbitq), 
to_sfixed(752.0/65536.0,1,-nbitq), 
to_sfixed(-1156.0/65536.0,1,-nbitq), 
to_sfixed(767.0/65536.0,1,-nbitq), 
to_sfixed(-2451.0/65536.0,1,-nbitq), 
to_sfixed(-295.0/65536.0,1,-nbitq), 
to_sfixed(4940.0/65536.0,1,-nbitq), 
to_sfixed(-2273.0/65536.0,1,-nbitq), 
to_sfixed(-623.0/65536.0,1,-nbitq), 
to_sfixed(2568.0/65536.0,1,-nbitq), 
to_sfixed(3523.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2624.0/65536.0,1,-nbitq), 
to_sfixed(2918.0/65536.0,1,-nbitq), 
to_sfixed(-936.0/65536.0,1,-nbitq), 
to_sfixed(395.0/65536.0,1,-nbitq), 
to_sfixed(-2733.0/65536.0,1,-nbitq), 
to_sfixed(-1568.0/65536.0,1,-nbitq), 
to_sfixed(-1934.0/65536.0,1,-nbitq), 
to_sfixed(-1999.0/65536.0,1,-nbitq), 
to_sfixed(-2886.0/65536.0,1,-nbitq), 
to_sfixed(1080.0/65536.0,1,-nbitq), 
to_sfixed(259.0/65536.0,1,-nbitq), 
to_sfixed(868.0/65536.0,1,-nbitq), 
to_sfixed(-1572.0/65536.0,1,-nbitq), 
to_sfixed(-4817.0/65536.0,1,-nbitq), 
to_sfixed(683.0/65536.0,1,-nbitq), 
to_sfixed(-1662.0/65536.0,1,-nbitq), 
to_sfixed(2455.0/65536.0,1,-nbitq), 
to_sfixed(-345.0/65536.0,1,-nbitq), 
to_sfixed(-500.0/65536.0,1,-nbitq), 
to_sfixed(585.0/65536.0,1,-nbitq), 
to_sfixed(-2607.0/65536.0,1,-nbitq), 
to_sfixed(-1049.0/65536.0,1,-nbitq), 
to_sfixed(1885.0/65536.0,1,-nbitq), 
to_sfixed(1931.0/65536.0,1,-nbitq), 
to_sfixed(2852.0/65536.0,1,-nbitq), 
to_sfixed(2479.0/65536.0,1,-nbitq), 
to_sfixed(-1755.0/65536.0,1,-nbitq), 
to_sfixed(-2580.0/65536.0,1,-nbitq), 
to_sfixed(1583.0/65536.0,1,-nbitq), 
to_sfixed(31.0/65536.0,1,-nbitq), 
to_sfixed(-452.0/65536.0,1,-nbitq), 
to_sfixed(-2391.0/65536.0,1,-nbitq), 
to_sfixed(-3312.0/65536.0,1,-nbitq), 
to_sfixed(-1402.0/65536.0,1,-nbitq), 
to_sfixed(-36.0/65536.0,1,-nbitq), 
to_sfixed(1178.0/65536.0,1,-nbitq), 
to_sfixed(-19.0/65536.0,1,-nbitq), 
to_sfixed(-3393.0/65536.0,1,-nbitq), 
to_sfixed(1404.0/65536.0,1,-nbitq), 
to_sfixed(-1826.0/65536.0,1,-nbitq), 
to_sfixed(-1002.0/65536.0,1,-nbitq), 
to_sfixed(83.0/65536.0,1,-nbitq), 
to_sfixed(-939.0/65536.0,1,-nbitq), 
to_sfixed(3049.0/65536.0,1,-nbitq), 
to_sfixed(2011.0/65536.0,1,-nbitq), 
to_sfixed(1988.0/65536.0,1,-nbitq), 
to_sfixed(-1879.0/65536.0,1,-nbitq), 
to_sfixed(2399.0/65536.0,1,-nbitq), 
to_sfixed(1508.0/65536.0,1,-nbitq), 
to_sfixed(2338.0/65536.0,1,-nbitq), 
to_sfixed(268.0/65536.0,1,-nbitq), 
to_sfixed(600.0/65536.0,1,-nbitq), 
to_sfixed(-957.0/65536.0,1,-nbitq), 
to_sfixed(2937.0/65536.0,1,-nbitq), 
to_sfixed(578.0/65536.0,1,-nbitq), 
to_sfixed(-286.0/65536.0,1,-nbitq), 
to_sfixed(-1094.0/65536.0,1,-nbitq), 
to_sfixed(639.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(-587.0/65536.0,1,-nbitq), 
to_sfixed(97.0/65536.0,1,-nbitq), 
to_sfixed(-1952.0/65536.0,1,-nbitq), 
to_sfixed(-1169.0/65536.0,1,-nbitq), 
to_sfixed(807.0/65536.0,1,-nbitq), 
to_sfixed(-757.0/65536.0,1,-nbitq), 
to_sfixed(332.0/65536.0,1,-nbitq), 
to_sfixed(-638.0/65536.0,1,-nbitq), 
to_sfixed(-3016.0/65536.0,1,-nbitq), 
to_sfixed(4064.0/65536.0,1,-nbitq), 
to_sfixed(-985.0/65536.0,1,-nbitq), 
to_sfixed(-329.0/65536.0,1,-nbitq), 
to_sfixed(-2282.0/65536.0,1,-nbitq), 
to_sfixed(-1174.0/65536.0,1,-nbitq), 
to_sfixed(-1393.0/65536.0,1,-nbitq), 
to_sfixed(-1289.0/65536.0,1,-nbitq), 
to_sfixed(-113.0/65536.0,1,-nbitq), 
to_sfixed(-527.0/65536.0,1,-nbitq), 
to_sfixed(1942.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(4914.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-110.0/65536.0,1,-nbitq), 
to_sfixed(-1188.0/65536.0,1,-nbitq), 
to_sfixed(1769.0/65536.0,1,-nbitq), 
to_sfixed(-1967.0/65536.0,1,-nbitq), 
to_sfixed(-2126.0/65536.0,1,-nbitq), 
to_sfixed(535.0/65536.0,1,-nbitq), 
to_sfixed(1686.0/65536.0,1,-nbitq), 
to_sfixed(-2316.0/65536.0,1,-nbitq), 
to_sfixed(2100.0/65536.0,1,-nbitq), 
to_sfixed(-2752.0/65536.0,1,-nbitq), 
to_sfixed(-3520.0/65536.0,1,-nbitq), 
to_sfixed(479.0/65536.0,1,-nbitq), 
to_sfixed(-916.0/65536.0,1,-nbitq), 
to_sfixed(-2850.0/65536.0,1,-nbitq), 
to_sfixed(2638.0/65536.0,1,-nbitq), 
to_sfixed(2381.0/65536.0,1,-nbitq), 
to_sfixed(1544.0/65536.0,1,-nbitq), 
to_sfixed(750.0/65536.0,1,-nbitq), 
to_sfixed(4181.0/65536.0,1,-nbitq), 
to_sfixed(-581.0/65536.0,1,-nbitq), 
to_sfixed(-874.0/65536.0,1,-nbitq), 
to_sfixed(-1327.0/65536.0,1,-nbitq), 
to_sfixed(385.0/65536.0,1,-nbitq), 
to_sfixed(507.0/65536.0,1,-nbitq), 
to_sfixed(1183.0/65536.0,1,-nbitq), 
to_sfixed(-1508.0/65536.0,1,-nbitq), 
to_sfixed(-3409.0/65536.0,1,-nbitq), 
to_sfixed(-1660.0/65536.0,1,-nbitq), 
to_sfixed(-2382.0/65536.0,1,-nbitq), 
to_sfixed(-2802.0/65536.0,1,-nbitq), 
to_sfixed(-1489.0/65536.0,1,-nbitq), 
to_sfixed(-2083.0/65536.0,1,-nbitq), 
to_sfixed(-5367.0/65536.0,1,-nbitq), 
to_sfixed(-5409.0/65536.0,1,-nbitq), 
to_sfixed(-2955.0/65536.0,1,-nbitq), 
to_sfixed(371.0/65536.0,1,-nbitq), 
to_sfixed(-2291.0/65536.0,1,-nbitq), 
to_sfixed(-1357.0/65536.0,1,-nbitq), 
to_sfixed(-3437.0/65536.0,1,-nbitq), 
to_sfixed(2048.0/65536.0,1,-nbitq), 
to_sfixed(-3826.0/65536.0,1,-nbitq), 
to_sfixed(-204.0/65536.0,1,-nbitq), 
to_sfixed(458.0/65536.0,1,-nbitq), 
to_sfixed(2677.0/65536.0,1,-nbitq), 
to_sfixed(2030.0/65536.0,1,-nbitq), 
to_sfixed(2381.0/65536.0,1,-nbitq), 
to_sfixed(2907.0/65536.0,1,-nbitq), 
to_sfixed(-575.0/65536.0,1,-nbitq), 
to_sfixed(2778.0/65536.0,1,-nbitq), 
to_sfixed(3105.0/65536.0,1,-nbitq), 
to_sfixed(-57.0/65536.0,1,-nbitq), 
to_sfixed(293.0/65536.0,1,-nbitq), 
to_sfixed(-1002.0/65536.0,1,-nbitq), 
to_sfixed(-2234.0/65536.0,1,-nbitq), 
to_sfixed(2791.0/65536.0,1,-nbitq), 
to_sfixed(168.0/65536.0,1,-nbitq), 
to_sfixed(-1992.0/65536.0,1,-nbitq), 
to_sfixed(308.0/65536.0,1,-nbitq), 
to_sfixed(2336.0/65536.0,1,-nbitq), 
to_sfixed(1809.0/65536.0,1,-nbitq), 
to_sfixed(-436.0/65536.0,1,-nbitq), 
to_sfixed(-428.0/65536.0,1,-nbitq), 
to_sfixed(-2158.0/65536.0,1,-nbitq), 
to_sfixed(-1316.0/65536.0,1,-nbitq), 
to_sfixed(-622.0/65536.0,1,-nbitq), 
to_sfixed(-1889.0/65536.0,1,-nbitq), 
to_sfixed(-1313.0/65536.0,1,-nbitq), 
to_sfixed(1270.0/65536.0,1,-nbitq), 
to_sfixed(2031.0/65536.0,1,-nbitq), 
to_sfixed(-2336.0/65536.0,1,-nbitq), 
to_sfixed(-1851.0/65536.0,1,-nbitq), 
to_sfixed(3025.0/65536.0,1,-nbitq), 
to_sfixed(3622.0/65536.0,1,-nbitq), 
to_sfixed(-1347.0/65536.0,1,-nbitq), 
to_sfixed(-399.0/65536.0,1,-nbitq), 
to_sfixed(2456.0/65536.0,1,-nbitq), 
to_sfixed(-1096.0/65536.0,1,-nbitq), 
to_sfixed(2743.0/65536.0,1,-nbitq), 
to_sfixed(2527.0/65536.0,1,-nbitq), 
to_sfixed(2107.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1518.0/65536.0,1,-nbitq), 
to_sfixed(1110.0/65536.0,1,-nbitq), 
to_sfixed(-578.0/65536.0,1,-nbitq), 
to_sfixed(727.0/65536.0,1,-nbitq), 
to_sfixed(-3832.0/65536.0,1,-nbitq), 
to_sfixed(-1304.0/65536.0,1,-nbitq), 
to_sfixed(-321.0/65536.0,1,-nbitq), 
to_sfixed(-625.0/65536.0,1,-nbitq), 
to_sfixed(1978.0/65536.0,1,-nbitq), 
to_sfixed(1319.0/65536.0,1,-nbitq), 
to_sfixed(-1346.0/65536.0,1,-nbitq), 
to_sfixed(3480.0/65536.0,1,-nbitq), 
to_sfixed(1722.0/65536.0,1,-nbitq), 
to_sfixed(1157.0/65536.0,1,-nbitq), 
to_sfixed(-1102.0/65536.0,1,-nbitq), 
to_sfixed(-1857.0/65536.0,1,-nbitq), 
to_sfixed(391.0/65536.0,1,-nbitq), 
to_sfixed(3425.0/65536.0,1,-nbitq), 
to_sfixed(778.0/65536.0,1,-nbitq), 
to_sfixed(-409.0/65536.0,1,-nbitq), 
to_sfixed(-2351.0/65536.0,1,-nbitq), 
to_sfixed(1528.0/65536.0,1,-nbitq), 
to_sfixed(1457.0/65536.0,1,-nbitq), 
to_sfixed(642.0/65536.0,1,-nbitq), 
to_sfixed(1936.0/65536.0,1,-nbitq), 
to_sfixed(-2226.0/65536.0,1,-nbitq), 
to_sfixed(-4457.0/65536.0,1,-nbitq), 
to_sfixed(3009.0/65536.0,1,-nbitq), 
to_sfixed(-792.0/65536.0,1,-nbitq), 
to_sfixed(1117.0/65536.0,1,-nbitq), 
to_sfixed(-2239.0/65536.0,1,-nbitq), 
to_sfixed(-1665.0/65536.0,1,-nbitq), 
to_sfixed(-5755.0/65536.0,1,-nbitq), 
to_sfixed(-1051.0/65536.0,1,-nbitq), 
to_sfixed(2557.0/65536.0,1,-nbitq), 
to_sfixed(-605.0/65536.0,1,-nbitq), 
to_sfixed(-883.0/65536.0,1,-nbitq), 
to_sfixed(-880.0/65536.0,1,-nbitq), 
to_sfixed(-4065.0/65536.0,1,-nbitq), 
to_sfixed(2054.0/65536.0,1,-nbitq), 
to_sfixed(-2257.0/65536.0,1,-nbitq), 
to_sfixed(-2428.0/65536.0,1,-nbitq), 
to_sfixed(-3072.0/65536.0,1,-nbitq), 
to_sfixed(-242.0/65536.0,1,-nbitq), 
to_sfixed(-848.0/65536.0,1,-nbitq), 
to_sfixed(-503.0/65536.0,1,-nbitq), 
to_sfixed(-1445.0/65536.0,1,-nbitq), 
to_sfixed(94.0/65536.0,1,-nbitq), 
to_sfixed(-1545.0/65536.0,1,-nbitq), 
to_sfixed(940.0/65536.0,1,-nbitq), 
to_sfixed(104.0/65536.0,1,-nbitq), 
to_sfixed(322.0/65536.0,1,-nbitq), 
to_sfixed(590.0/65536.0,1,-nbitq), 
to_sfixed(-1808.0/65536.0,1,-nbitq), 
to_sfixed(-543.0/65536.0,1,-nbitq), 
to_sfixed(-1912.0/65536.0,1,-nbitq), 
to_sfixed(514.0/65536.0,1,-nbitq), 
to_sfixed(-409.0/65536.0,1,-nbitq), 
to_sfixed(903.0/65536.0,1,-nbitq), 
to_sfixed(4575.0/65536.0,1,-nbitq), 
to_sfixed(428.0/65536.0,1,-nbitq), 
to_sfixed(867.0/65536.0,1,-nbitq), 
to_sfixed(-1149.0/65536.0,1,-nbitq), 
to_sfixed(-274.0/65536.0,1,-nbitq), 
to_sfixed(637.0/65536.0,1,-nbitq), 
to_sfixed(750.0/65536.0,1,-nbitq), 
to_sfixed(-1779.0/65536.0,1,-nbitq), 
to_sfixed(-1843.0/65536.0,1,-nbitq), 
to_sfixed(3238.0/65536.0,1,-nbitq), 
to_sfixed(736.0/65536.0,1,-nbitq), 
to_sfixed(-1497.0/65536.0,1,-nbitq), 
to_sfixed(-471.0/65536.0,1,-nbitq), 
to_sfixed(665.0/65536.0,1,-nbitq), 
to_sfixed(1743.0/65536.0,1,-nbitq), 
to_sfixed(1072.0/65536.0,1,-nbitq), 
to_sfixed(1396.0/65536.0,1,-nbitq), 
to_sfixed(-684.0/65536.0,1,-nbitq), 
to_sfixed(-294.0/65536.0,1,-nbitq), 
to_sfixed(-1243.0/65536.0,1,-nbitq), 
to_sfixed(3871.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1868.0/65536.0,1,-nbitq), 
to_sfixed(2446.0/65536.0,1,-nbitq), 
to_sfixed(-1021.0/65536.0,1,-nbitq), 
to_sfixed(1310.0/65536.0,1,-nbitq), 
to_sfixed(-2035.0/65536.0,1,-nbitq), 
to_sfixed(-3444.0/65536.0,1,-nbitq), 
to_sfixed(-908.0/65536.0,1,-nbitq), 
to_sfixed(303.0/65536.0,1,-nbitq), 
to_sfixed(241.0/65536.0,1,-nbitq), 
to_sfixed(2763.0/65536.0,1,-nbitq), 
to_sfixed(-1096.0/65536.0,1,-nbitq), 
to_sfixed(239.0/65536.0,1,-nbitq), 
to_sfixed(714.0/65536.0,1,-nbitq), 
to_sfixed(18.0/65536.0,1,-nbitq), 
to_sfixed(91.0/65536.0,1,-nbitq), 
to_sfixed(1390.0/65536.0,1,-nbitq), 
to_sfixed(-1385.0/65536.0,1,-nbitq), 
to_sfixed(220.0/65536.0,1,-nbitq), 
to_sfixed(2134.0/65536.0,1,-nbitq), 
to_sfixed(432.0/65536.0,1,-nbitq), 
to_sfixed(995.0/65536.0,1,-nbitq), 
to_sfixed(-649.0/65536.0,1,-nbitq), 
to_sfixed(-2062.0/65536.0,1,-nbitq), 
to_sfixed(1120.0/65536.0,1,-nbitq), 
to_sfixed(43.0/65536.0,1,-nbitq), 
to_sfixed(-536.0/65536.0,1,-nbitq), 
to_sfixed(-779.0/65536.0,1,-nbitq), 
to_sfixed(145.0/65536.0,1,-nbitq), 
to_sfixed(-2608.0/65536.0,1,-nbitq), 
to_sfixed(-3622.0/65536.0,1,-nbitq), 
to_sfixed(-1154.0/65536.0,1,-nbitq), 
to_sfixed(3159.0/65536.0,1,-nbitq), 
to_sfixed(-1439.0/65536.0,1,-nbitq), 
to_sfixed(-533.0/65536.0,1,-nbitq), 
to_sfixed(-1379.0/65536.0,1,-nbitq), 
to_sfixed(-133.0/65536.0,1,-nbitq), 
to_sfixed(-3591.0/65536.0,1,-nbitq), 
to_sfixed(951.0/65536.0,1,-nbitq), 
to_sfixed(-3361.0/65536.0,1,-nbitq), 
to_sfixed(1205.0/65536.0,1,-nbitq), 
to_sfixed(-914.0/65536.0,1,-nbitq), 
to_sfixed(-2358.0/65536.0,1,-nbitq), 
to_sfixed(311.0/65536.0,1,-nbitq), 
to_sfixed(96.0/65536.0,1,-nbitq), 
to_sfixed(-1224.0/65536.0,1,-nbitq), 
to_sfixed(4610.0/65536.0,1,-nbitq), 
to_sfixed(-899.0/65536.0,1,-nbitq), 
to_sfixed(605.0/65536.0,1,-nbitq), 
to_sfixed(155.0/65536.0,1,-nbitq), 
to_sfixed(3371.0/65536.0,1,-nbitq), 
to_sfixed(644.0/65536.0,1,-nbitq), 
to_sfixed(2835.0/65536.0,1,-nbitq), 
to_sfixed(-1546.0/65536.0,1,-nbitq), 
to_sfixed(1572.0/65536.0,1,-nbitq), 
to_sfixed(-391.0/65536.0,1,-nbitq), 
to_sfixed(2770.0/65536.0,1,-nbitq), 
to_sfixed(-2440.0/65536.0,1,-nbitq), 
to_sfixed(958.0/65536.0,1,-nbitq), 
to_sfixed(-2936.0/65536.0,1,-nbitq), 
to_sfixed(399.0/65536.0,1,-nbitq), 
to_sfixed(794.0/65536.0,1,-nbitq), 
to_sfixed(608.0/65536.0,1,-nbitq), 
to_sfixed(2162.0/65536.0,1,-nbitq), 
to_sfixed(807.0/65536.0,1,-nbitq), 
to_sfixed(-1960.0/65536.0,1,-nbitq), 
to_sfixed(2964.0/65536.0,1,-nbitq), 
to_sfixed(-274.0/65536.0,1,-nbitq), 
to_sfixed(2044.0/65536.0,1,-nbitq), 
to_sfixed(2722.0/65536.0,1,-nbitq), 
to_sfixed(2711.0/65536.0,1,-nbitq), 
to_sfixed(1241.0/65536.0,1,-nbitq), 
to_sfixed(-1664.0/65536.0,1,-nbitq), 
to_sfixed(2593.0/65536.0,1,-nbitq), 
to_sfixed(1094.0/65536.0,1,-nbitq), 
to_sfixed(1403.0/65536.0,1,-nbitq), 
to_sfixed(675.0/65536.0,1,-nbitq), 
to_sfixed(-3193.0/65536.0,1,-nbitq), 
to_sfixed(3063.0/65536.0,1,-nbitq), 
to_sfixed(-820.0/65536.0,1,-nbitq), 
to_sfixed(4141.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1348.0/65536.0,1,-nbitq), 
to_sfixed(2306.0/65536.0,1,-nbitq), 
to_sfixed(2601.0/65536.0,1,-nbitq), 
to_sfixed(-2362.0/65536.0,1,-nbitq), 
to_sfixed(4401.0/65536.0,1,-nbitq), 
to_sfixed(-668.0/65536.0,1,-nbitq), 
to_sfixed(-555.0/65536.0,1,-nbitq), 
to_sfixed(-3418.0/65536.0,1,-nbitq), 
to_sfixed(-4112.0/65536.0,1,-nbitq), 
to_sfixed(2208.0/65536.0,1,-nbitq), 
to_sfixed(213.0/65536.0,1,-nbitq), 
to_sfixed(-4669.0/65536.0,1,-nbitq), 
to_sfixed(-1489.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(-1567.0/65536.0,1,-nbitq), 
to_sfixed(2129.0/65536.0,1,-nbitq), 
to_sfixed(2125.0/65536.0,1,-nbitq), 
to_sfixed(-295.0/65536.0,1,-nbitq), 
to_sfixed(-1381.0/65536.0,1,-nbitq), 
to_sfixed(2232.0/65536.0,1,-nbitq), 
to_sfixed(280.0/65536.0,1,-nbitq), 
to_sfixed(2076.0/65536.0,1,-nbitq), 
to_sfixed(640.0/65536.0,1,-nbitq), 
to_sfixed(2202.0/65536.0,1,-nbitq), 
to_sfixed(-147.0/65536.0,1,-nbitq), 
to_sfixed(2738.0/65536.0,1,-nbitq), 
to_sfixed(-2347.0/65536.0,1,-nbitq), 
to_sfixed(-2125.0/65536.0,1,-nbitq), 
to_sfixed(2254.0/65536.0,1,-nbitq), 
to_sfixed(-3115.0/65536.0,1,-nbitq), 
to_sfixed(-1150.0/65536.0,1,-nbitq), 
to_sfixed(2401.0/65536.0,1,-nbitq), 
to_sfixed(394.0/65536.0,1,-nbitq), 
to_sfixed(-1519.0/65536.0,1,-nbitq), 
to_sfixed(-1485.0/65536.0,1,-nbitq), 
to_sfixed(1134.0/65536.0,1,-nbitq), 
to_sfixed(-1028.0/65536.0,1,-nbitq), 
to_sfixed(-1319.0/65536.0,1,-nbitq), 
to_sfixed(-4286.0/65536.0,1,-nbitq), 
to_sfixed(880.0/65536.0,1,-nbitq), 
to_sfixed(-3102.0/65536.0,1,-nbitq), 
to_sfixed(-1971.0/65536.0,1,-nbitq), 
to_sfixed(-164.0/65536.0,1,-nbitq), 
to_sfixed(1232.0/65536.0,1,-nbitq), 
to_sfixed(976.0/65536.0,1,-nbitq), 
to_sfixed(2851.0/65536.0,1,-nbitq), 
to_sfixed(485.0/65536.0,1,-nbitq), 
to_sfixed(905.0/65536.0,1,-nbitq), 
to_sfixed(361.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(-246.0/65536.0,1,-nbitq), 
to_sfixed(2449.0/65536.0,1,-nbitq), 
to_sfixed(1932.0/65536.0,1,-nbitq), 
to_sfixed(-1250.0/65536.0,1,-nbitq), 
to_sfixed(2944.0/65536.0,1,-nbitq), 
to_sfixed(-2207.0/65536.0,1,-nbitq), 
to_sfixed(-1516.0/65536.0,1,-nbitq), 
to_sfixed(3735.0/65536.0,1,-nbitq), 
to_sfixed(1790.0/65536.0,1,-nbitq), 
to_sfixed(-58.0/65536.0,1,-nbitq), 
to_sfixed(340.0/65536.0,1,-nbitq), 
to_sfixed(2294.0/65536.0,1,-nbitq), 
to_sfixed(1683.0/65536.0,1,-nbitq), 
to_sfixed(-763.0/65536.0,1,-nbitq), 
to_sfixed(-1019.0/65536.0,1,-nbitq), 
to_sfixed(3633.0/65536.0,1,-nbitq), 
to_sfixed(2530.0/65536.0,1,-nbitq), 
to_sfixed(987.0/65536.0,1,-nbitq), 
to_sfixed(1639.0/65536.0,1,-nbitq), 
to_sfixed(4024.0/65536.0,1,-nbitq), 
to_sfixed(1686.0/65536.0,1,-nbitq), 
to_sfixed(-603.0/65536.0,1,-nbitq), 
to_sfixed(1520.0/65536.0,1,-nbitq), 
to_sfixed(524.0/65536.0,1,-nbitq), 
to_sfixed(-1176.0/65536.0,1,-nbitq), 
to_sfixed(1511.0/65536.0,1,-nbitq), 
to_sfixed(-5316.0/65536.0,1,-nbitq), 
to_sfixed(1913.0/65536.0,1,-nbitq), 
to_sfixed(-1042.0/65536.0,1,-nbitq), 
to_sfixed(1861.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2693.0/65536.0,1,-nbitq), 
to_sfixed(-2551.0/65536.0,1,-nbitq), 
to_sfixed(-544.0/65536.0,1,-nbitq), 
to_sfixed(1494.0/65536.0,1,-nbitq), 
to_sfixed(8237.0/65536.0,1,-nbitq), 
to_sfixed(-318.0/65536.0,1,-nbitq), 
to_sfixed(-2071.0/65536.0,1,-nbitq), 
to_sfixed(-738.0/65536.0,1,-nbitq), 
to_sfixed(-3306.0/65536.0,1,-nbitq), 
to_sfixed(-377.0/65536.0,1,-nbitq), 
to_sfixed(301.0/65536.0,1,-nbitq), 
to_sfixed(-146.0/65536.0,1,-nbitq), 
to_sfixed(2435.0/65536.0,1,-nbitq), 
to_sfixed(1611.0/65536.0,1,-nbitq), 
to_sfixed(-751.0/65536.0,1,-nbitq), 
to_sfixed(530.0/65536.0,1,-nbitq), 
to_sfixed(1527.0/65536.0,1,-nbitq), 
to_sfixed(-1344.0/65536.0,1,-nbitq), 
to_sfixed(-2942.0/65536.0,1,-nbitq), 
to_sfixed(1962.0/65536.0,1,-nbitq), 
to_sfixed(4560.0/65536.0,1,-nbitq), 
to_sfixed(-972.0/65536.0,1,-nbitq), 
to_sfixed(442.0/65536.0,1,-nbitq), 
to_sfixed(-2712.0/65536.0,1,-nbitq), 
to_sfixed(-291.0/65536.0,1,-nbitq), 
to_sfixed(2420.0/65536.0,1,-nbitq), 
to_sfixed(1325.0/65536.0,1,-nbitq), 
to_sfixed(1887.0/65536.0,1,-nbitq), 
to_sfixed(6650.0/65536.0,1,-nbitq), 
to_sfixed(-3321.0/65536.0,1,-nbitq), 
to_sfixed(-1103.0/65536.0,1,-nbitq), 
to_sfixed(-385.0/65536.0,1,-nbitq), 
to_sfixed(1013.0/65536.0,1,-nbitq), 
to_sfixed(-5669.0/65536.0,1,-nbitq), 
to_sfixed(2355.0/65536.0,1,-nbitq), 
to_sfixed(-3084.0/65536.0,1,-nbitq), 
to_sfixed(-8329.0/65536.0,1,-nbitq), 
to_sfixed(1299.0/65536.0,1,-nbitq), 
to_sfixed(-4923.0/65536.0,1,-nbitq), 
to_sfixed(-2840.0/65536.0,1,-nbitq), 
to_sfixed(-294.0/65536.0,1,-nbitq), 
to_sfixed(-988.0/65536.0,1,-nbitq), 
to_sfixed(1671.0/65536.0,1,-nbitq), 
to_sfixed(4361.0/65536.0,1,-nbitq), 
to_sfixed(-1185.0/65536.0,1,-nbitq), 
to_sfixed(-665.0/65536.0,1,-nbitq), 
to_sfixed(2747.0/65536.0,1,-nbitq), 
to_sfixed(-277.0/65536.0,1,-nbitq), 
to_sfixed(-1872.0/65536.0,1,-nbitq), 
to_sfixed(-730.0/65536.0,1,-nbitq), 
to_sfixed(-946.0/65536.0,1,-nbitq), 
to_sfixed(1480.0/65536.0,1,-nbitq), 
to_sfixed(1558.0/65536.0,1,-nbitq), 
to_sfixed(-2645.0/65536.0,1,-nbitq), 
to_sfixed(-3815.0/65536.0,1,-nbitq), 
to_sfixed(1689.0/65536.0,1,-nbitq), 
to_sfixed(-2198.0/65536.0,1,-nbitq), 
to_sfixed(5631.0/65536.0,1,-nbitq), 
to_sfixed(-661.0/65536.0,1,-nbitq), 
to_sfixed(-3319.0/65536.0,1,-nbitq), 
to_sfixed(-6073.0/65536.0,1,-nbitq), 
to_sfixed(2020.0/65536.0,1,-nbitq), 
to_sfixed(2432.0/65536.0,1,-nbitq), 
to_sfixed(-2866.0/65536.0,1,-nbitq), 
to_sfixed(-1593.0/65536.0,1,-nbitq), 
to_sfixed(3413.0/65536.0,1,-nbitq), 
to_sfixed(-1833.0/65536.0,1,-nbitq), 
to_sfixed(24.0/65536.0,1,-nbitq), 
to_sfixed(2092.0/65536.0,1,-nbitq), 
to_sfixed(-775.0/65536.0,1,-nbitq), 
to_sfixed(2247.0/65536.0,1,-nbitq), 
to_sfixed(-2613.0/65536.0,1,-nbitq), 
to_sfixed(-1102.0/65536.0,1,-nbitq), 
to_sfixed(2455.0/65536.0,1,-nbitq), 
to_sfixed(-327.0/65536.0,1,-nbitq), 
to_sfixed(4241.0/65536.0,1,-nbitq), 
to_sfixed(-7760.0/65536.0,1,-nbitq), 
to_sfixed(-2867.0/65536.0,1,-nbitq), 
to_sfixed(137.0/65536.0,1,-nbitq), 
to_sfixed(-925.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3376.0/65536.0,1,-nbitq), 
to_sfixed(-360.0/65536.0,1,-nbitq), 
to_sfixed(-6400.0/65536.0,1,-nbitq), 
to_sfixed(-167.0/65536.0,1,-nbitq), 
to_sfixed(510.0/65536.0,1,-nbitq), 
to_sfixed(539.0/65536.0,1,-nbitq), 
to_sfixed(-1407.0/65536.0,1,-nbitq), 
to_sfixed(-691.0/65536.0,1,-nbitq), 
to_sfixed(-4611.0/65536.0,1,-nbitq), 
to_sfixed(-19.0/65536.0,1,-nbitq), 
to_sfixed(6419.0/65536.0,1,-nbitq), 
to_sfixed(-3982.0/65536.0,1,-nbitq), 
to_sfixed(1088.0/65536.0,1,-nbitq), 
to_sfixed(2814.0/65536.0,1,-nbitq), 
to_sfixed(-536.0/65536.0,1,-nbitq), 
to_sfixed(-957.0/65536.0,1,-nbitq), 
to_sfixed(2562.0/65536.0,1,-nbitq), 
to_sfixed(-607.0/65536.0,1,-nbitq), 
to_sfixed(825.0/65536.0,1,-nbitq), 
to_sfixed(-1898.0/65536.0,1,-nbitq), 
to_sfixed(3586.0/65536.0,1,-nbitq), 
to_sfixed(4580.0/65536.0,1,-nbitq), 
to_sfixed(985.0/65536.0,1,-nbitq), 
to_sfixed(-4019.0/65536.0,1,-nbitq), 
to_sfixed(92.0/65536.0,1,-nbitq), 
to_sfixed(-4816.0/65536.0,1,-nbitq), 
to_sfixed(-542.0/65536.0,1,-nbitq), 
to_sfixed(3738.0/65536.0,1,-nbitq), 
to_sfixed(488.0/65536.0,1,-nbitq), 
to_sfixed(-5526.0/65536.0,1,-nbitq), 
to_sfixed(-469.0/65536.0,1,-nbitq), 
to_sfixed(-2348.0/65536.0,1,-nbitq), 
to_sfixed(1567.0/65536.0,1,-nbitq), 
to_sfixed(-9457.0/65536.0,1,-nbitq), 
to_sfixed(1594.0/65536.0,1,-nbitq), 
to_sfixed(-2898.0/65536.0,1,-nbitq), 
to_sfixed(-12269.0/65536.0,1,-nbitq), 
to_sfixed(4222.0/65536.0,1,-nbitq), 
to_sfixed(-8361.0/65536.0,1,-nbitq), 
to_sfixed(128.0/65536.0,1,-nbitq), 
to_sfixed(7071.0/65536.0,1,-nbitq), 
to_sfixed(1215.0/65536.0,1,-nbitq), 
to_sfixed(674.0/65536.0,1,-nbitq), 
to_sfixed(5111.0/65536.0,1,-nbitq), 
to_sfixed(-611.0/65536.0,1,-nbitq), 
to_sfixed(6004.0/65536.0,1,-nbitq), 
to_sfixed(-1766.0/65536.0,1,-nbitq), 
to_sfixed(-372.0/65536.0,1,-nbitq), 
to_sfixed(-1740.0/65536.0,1,-nbitq), 
to_sfixed(2053.0/65536.0,1,-nbitq), 
to_sfixed(-1618.0/65536.0,1,-nbitq), 
to_sfixed(606.0/65536.0,1,-nbitq), 
to_sfixed(-1530.0/65536.0,1,-nbitq), 
to_sfixed(1094.0/65536.0,1,-nbitq), 
to_sfixed(-1585.0/65536.0,1,-nbitq), 
to_sfixed(4454.0/65536.0,1,-nbitq), 
to_sfixed(151.0/65536.0,1,-nbitq), 
to_sfixed(-236.0/65536.0,1,-nbitq), 
to_sfixed(-584.0/65536.0,1,-nbitq), 
to_sfixed(-9404.0/65536.0,1,-nbitq), 
to_sfixed(-4396.0/65536.0,1,-nbitq), 
to_sfixed(-1008.0/65536.0,1,-nbitq), 
to_sfixed(-2122.0/65536.0,1,-nbitq), 
to_sfixed(-1894.0/65536.0,1,-nbitq), 
to_sfixed(1750.0/65536.0,1,-nbitq), 
to_sfixed(5435.0/65536.0,1,-nbitq), 
to_sfixed(1825.0/65536.0,1,-nbitq), 
to_sfixed(2051.0/65536.0,1,-nbitq), 
to_sfixed(8192.0/65536.0,1,-nbitq), 
to_sfixed(3425.0/65536.0,1,-nbitq), 
to_sfixed(-125.0/65536.0,1,-nbitq), 
to_sfixed(2129.0/65536.0,1,-nbitq), 
to_sfixed(2629.0/65536.0,1,-nbitq), 
to_sfixed(281.0/65536.0,1,-nbitq), 
to_sfixed(2134.0/65536.0,1,-nbitq), 
to_sfixed(-3057.0/65536.0,1,-nbitq), 
to_sfixed(-6129.0/65536.0,1,-nbitq), 
to_sfixed(-2656.0/65536.0,1,-nbitq), 
to_sfixed(-744.0/65536.0,1,-nbitq), 
to_sfixed(-2540.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3657.0/65536.0,1,-nbitq), 
to_sfixed(-3484.0/65536.0,1,-nbitq), 
to_sfixed(-4400.0/65536.0,1,-nbitq), 
to_sfixed(-5087.0/65536.0,1,-nbitq), 
to_sfixed(-3188.0/65536.0,1,-nbitq), 
to_sfixed(-1841.0/65536.0,1,-nbitq), 
to_sfixed(-7426.0/65536.0,1,-nbitq), 
to_sfixed(-5508.0/65536.0,1,-nbitq), 
to_sfixed(-3037.0/65536.0,1,-nbitq), 
to_sfixed(2499.0/65536.0,1,-nbitq), 
to_sfixed(4427.0/65536.0,1,-nbitq), 
to_sfixed(3809.0/65536.0,1,-nbitq), 
to_sfixed(972.0/65536.0,1,-nbitq), 
to_sfixed(-255.0/65536.0,1,-nbitq), 
to_sfixed(-3968.0/65536.0,1,-nbitq), 
to_sfixed(1705.0/65536.0,1,-nbitq), 
to_sfixed(980.0/65536.0,1,-nbitq), 
to_sfixed(-1512.0/65536.0,1,-nbitq), 
to_sfixed(123.0/65536.0,1,-nbitq), 
to_sfixed(1612.0/65536.0,1,-nbitq), 
to_sfixed(-526.0/65536.0,1,-nbitq), 
to_sfixed(4439.0/65536.0,1,-nbitq), 
to_sfixed(4752.0/65536.0,1,-nbitq), 
to_sfixed(-12483.0/65536.0,1,-nbitq), 
to_sfixed(2065.0/65536.0,1,-nbitq), 
to_sfixed(-13631.0/65536.0,1,-nbitq), 
to_sfixed(-6601.0/65536.0,1,-nbitq), 
to_sfixed(134.0/65536.0,1,-nbitq), 
to_sfixed(113.0/65536.0,1,-nbitq), 
to_sfixed(-4981.0/65536.0,1,-nbitq), 
to_sfixed(4614.0/65536.0,1,-nbitq), 
to_sfixed(1828.0/65536.0,1,-nbitq), 
to_sfixed(2071.0/65536.0,1,-nbitq), 
to_sfixed(-7103.0/65536.0,1,-nbitq), 
to_sfixed(466.0/65536.0,1,-nbitq), 
to_sfixed(2728.0/65536.0,1,-nbitq), 
to_sfixed(-12470.0/65536.0,1,-nbitq), 
to_sfixed(5658.0/65536.0,1,-nbitq), 
to_sfixed(-5296.0/65536.0,1,-nbitq), 
to_sfixed(-9845.0/65536.0,1,-nbitq), 
to_sfixed(5028.0/65536.0,1,-nbitq), 
to_sfixed(1067.0/65536.0,1,-nbitq), 
to_sfixed(4297.0/65536.0,1,-nbitq), 
to_sfixed(7955.0/65536.0,1,-nbitq), 
to_sfixed(-1397.0/65536.0,1,-nbitq), 
to_sfixed(2776.0/65536.0,1,-nbitq), 
to_sfixed(687.0/65536.0,1,-nbitq), 
to_sfixed(1481.0/65536.0,1,-nbitq), 
to_sfixed(1619.0/65536.0,1,-nbitq), 
to_sfixed(1458.0/65536.0,1,-nbitq), 
to_sfixed(1423.0/65536.0,1,-nbitq), 
to_sfixed(-548.0/65536.0,1,-nbitq), 
to_sfixed(-59.0/65536.0,1,-nbitq), 
to_sfixed(-2097.0/65536.0,1,-nbitq), 
to_sfixed(-3217.0/65536.0,1,-nbitq), 
to_sfixed(4739.0/65536.0,1,-nbitq), 
to_sfixed(902.0/65536.0,1,-nbitq), 
to_sfixed(3041.0/65536.0,1,-nbitq), 
to_sfixed(1756.0/65536.0,1,-nbitq), 
to_sfixed(-15008.0/65536.0,1,-nbitq), 
to_sfixed(-7840.0/65536.0,1,-nbitq), 
to_sfixed(1710.0/65536.0,1,-nbitq), 
to_sfixed(1811.0/65536.0,1,-nbitq), 
to_sfixed(-3493.0/65536.0,1,-nbitq), 
to_sfixed(-6456.0/65536.0,1,-nbitq), 
to_sfixed(3719.0/65536.0,1,-nbitq), 
to_sfixed(-597.0/65536.0,1,-nbitq), 
to_sfixed(5083.0/65536.0,1,-nbitq), 
to_sfixed(4771.0/65536.0,1,-nbitq), 
to_sfixed(538.0/65536.0,1,-nbitq), 
to_sfixed(612.0/65536.0,1,-nbitq), 
to_sfixed(2968.0/65536.0,1,-nbitq), 
to_sfixed(-461.0/65536.0,1,-nbitq), 
to_sfixed(-2169.0/65536.0,1,-nbitq), 
to_sfixed(190.0/65536.0,1,-nbitq), 
to_sfixed(351.0/65536.0,1,-nbitq), 
to_sfixed(-3174.0/65536.0,1,-nbitq), 
to_sfixed(2506.0/65536.0,1,-nbitq), 
to_sfixed(-119.0/65536.0,1,-nbitq), 
to_sfixed(-2634.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3952.0/65536.0,1,-nbitq), 
to_sfixed(-1329.0/65536.0,1,-nbitq), 
to_sfixed(-4065.0/65536.0,1,-nbitq), 
to_sfixed(-2481.0/65536.0,1,-nbitq), 
to_sfixed(-10084.0/65536.0,1,-nbitq), 
to_sfixed(970.0/65536.0,1,-nbitq), 
to_sfixed(-8911.0/65536.0,1,-nbitq), 
to_sfixed(-2818.0/65536.0,1,-nbitq), 
to_sfixed(-4237.0/65536.0,1,-nbitq), 
to_sfixed(2840.0/65536.0,1,-nbitq), 
to_sfixed(-2570.0/65536.0,1,-nbitq), 
to_sfixed(138.0/65536.0,1,-nbitq), 
to_sfixed(-574.0/65536.0,1,-nbitq), 
to_sfixed(-2553.0/65536.0,1,-nbitq), 
to_sfixed(-1250.0/65536.0,1,-nbitq), 
to_sfixed(-1518.0/65536.0,1,-nbitq), 
to_sfixed(-1206.0/65536.0,1,-nbitq), 
to_sfixed(4600.0/65536.0,1,-nbitq), 
to_sfixed(-6472.0/65536.0,1,-nbitq), 
to_sfixed(-1697.0/65536.0,1,-nbitq), 
to_sfixed(-2431.0/65536.0,1,-nbitq), 
to_sfixed(-5847.0/65536.0,1,-nbitq), 
to_sfixed(-940.0/65536.0,1,-nbitq), 
to_sfixed(-11602.0/65536.0,1,-nbitq), 
to_sfixed(4226.0/65536.0,1,-nbitq), 
to_sfixed(-17208.0/65536.0,1,-nbitq), 
to_sfixed(-2098.0/65536.0,1,-nbitq), 
to_sfixed(1059.0/65536.0,1,-nbitq), 
to_sfixed(-1904.0/65536.0,1,-nbitq), 
to_sfixed(-4178.0/65536.0,1,-nbitq), 
to_sfixed(3888.0/65536.0,1,-nbitq), 
to_sfixed(2893.0/65536.0,1,-nbitq), 
to_sfixed(1120.0/65536.0,1,-nbitq), 
to_sfixed(-4276.0/65536.0,1,-nbitq), 
to_sfixed(-2197.0/65536.0,1,-nbitq), 
to_sfixed(-343.0/65536.0,1,-nbitq), 
to_sfixed(-14317.0/65536.0,1,-nbitq), 
to_sfixed(5339.0/65536.0,1,-nbitq), 
to_sfixed(-2815.0/65536.0,1,-nbitq), 
to_sfixed(-11028.0/65536.0,1,-nbitq), 
to_sfixed(4306.0/65536.0,1,-nbitq), 
to_sfixed(-2766.0/65536.0,1,-nbitq), 
to_sfixed(6880.0/65536.0,1,-nbitq), 
to_sfixed(4429.0/65536.0,1,-nbitq), 
to_sfixed(-2137.0/65536.0,1,-nbitq), 
to_sfixed(2653.0/65536.0,1,-nbitq), 
to_sfixed(2837.0/65536.0,1,-nbitq), 
to_sfixed(865.0/65536.0,1,-nbitq), 
to_sfixed(1062.0/65536.0,1,-nbitq), 
to_sfixed(3249.0/65536.0,1,-nbitq), 
to_sfixed(1958.0/65536.0,1,-nbitq), 
to_sfixed(2107.0/65536.0,1,-nbitq), 
to_sfixed(1760.0/65536.0,1,-nbitq), 
to_sfixed(-1974.0/65536.0,1,-nbitq), 
to_sfixed(-9565.0/65536.0,1,-nbitq), 
to_sfixed(819.0/65536.0,1,-nbitq), 
to_sfixed(1330.0/65536.0,1,-nbitq), 
to_sfixed(-392.0/65536.0,1,-nbitq), 
to_sfixed(-1843.0/65536.0,1,-nbitq), 
to_sfixed(-9041.0/65536.0,1,-nbitq), 
to_sfixed(-4506.0/65536.0,1,-nbitq), 
to_sfixed(675.0/65536.0,1,-nbitq), 
to_sfixed(-2328.0/65536.0,1,-nbitq), 
to_sfixed(-2144.0/65536.0,1,-nbitq), 
to_sfixed(-4377.0/65536.0,1,-nbitq), 
to_sfixed(10382.0/65536.0,1,-nbitq), 
to_sfixed(1243.0/65536.0,1,-nbitq), 
to_sfixed(4519.0/65536.0,1,-nbitq), 
to_sfixed(3951.0/65536.0,1,-nbitq), 
to_sfixed(-1604.0/65536.0,1,-nbitq), 
to_sfixed(376.0/65536.0,1,-nbitq), 
to_sfixed(238.0/65536.0,1,-nbitq), 
to_sfixed(-355.0/65536.0,1,-nbitq), 
to_sfixed(-690.0/65536.0,1,-nbitq), 
to_sfixed(2052.0/65536.0,1,-nbitq), 
to_sfixed(-2428.0/65536.0,1,-nbitq), 
to_sfixed(-3142.0/65536.0,1,-nbitq), 
to_sfixed(1614.0/65536.0,1,-nbitq), 
to_sfixed(2556.0/65536.0,1,-nbitq), 
to_sfixed(1409.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2456.0/65536.0,1,-nbitq), 
to_sfixed(-3056.0/65536.0,1,-nbitq), 
to_sfixed(-4936.0/65536.0,1,-nbitq), 
to_sfixed(-3832.0/65536.0,1,-nbitq), 
to_sfixed(5492.0/65536.0,1,-nbitq), 
to_sfixed(3264.0/65536.0,1,-nbitq), 
to_sfixed(-8496.0/65536.0,1,-nbitq), 
to_sfixed(3645.0/65536.0,1,-nbitq), 
to_sfixed(1591.0/65536.0,1,-nbitq), 
to_sfixed(-749.0/65536.0,1,-nbitq), 
to_sfixed(-104.0/65536.0,1,-nbitq), 
to_sfixed(-8506.0/65536.0,1,-nbitq), 
to_sfixed(2081.0/65536.0,1,-nbitq), 
to_sfixed(3801.0/65536.0,1,-nbitq), 
to_sfixed(-2073.0/65536.0,1,-nbitq), 
to_sfixed(2725.0/65536.0,1,-nbitq), 
to_sfixed(-710.0/65536.0,1,-nbitq), 
to_sfixed(1843.0/65536.0,1,-nbitq), 
to_sfixed(-2238.0/65536.0,1,-nbitq), 
to_sfixed(734.0/65536.0,1,-nbitq), 
to_sfixed(939.0/65536.0,1,-nbitq), 
to_sfixed(-16819.0/65536.0,1,-nbitq), 
to_sfixed(-2276.0/65536.0,1,-nbitq), 
to_sfixed(6633.0/65536.0,1,-nbitq), 
to_sfixed(-1672.0/65536.0,1,-nbitq), 
to_sfixed(-13608.0/65536.0,1,-nbitq), 
to_sfixed(-189.0/65536.0,1,-nbitq), 
to_sfixed(4301.0/65536.0,1,-nbitq), 
to_sfixed(-3667.0/65536.0,1,-nbitq), 
to_sfixed(973.0/65536.0,1,-nbitq), 
to_sfixed(3709.0/65536.0,1,-nbitq), 
to_sfixed(2739.0/65536.0,1,-nbitq), 
to_sfixed(2301.0/65536.0,1,-nbitq), 
to_sfixed(1654.0/65536.0,1,-nbitq), 
to_sfixed(-457.0/65536.0,1,-nbitq), 
to_sfixed(2326.0/65536.0,1,-nbitq), 
to_sfixed(-11733.0/65536.0,1,-nbitq), 
to_sfixed(3185.0/65536.0,1,-nbitq), 
to_sfixed(1877.0/65536.0,1,-nbitq), 
to_sfixed(-3942.0/65536.0,1,-nbitq), 
to_sfixed(6480.0/65536.0,1,-nbitq), 
to_sfixed(-1451.0/65536.0,1,-nbitq), 
to_sfixed(1515.0/65536.0,1,-nbitq), 
to_sfixed(11178.0/65536.0,1,-nbitq), 
to_sfixed(-403.0/65536.0,1,-nbitq), 
to_sfixed(-6574.0/65536.0,1,-nbitq), 
to_sfixed(1425.0/65536.0,1,-nbitq), 
to_sfixed(4049.0/65536.0,1,-nbitq), 
to_sfixed(871.0/65536.0,1,-nbitq), 
to_sfixed(855.0/65536.0,1,-nbitq), 
to_sfixed(2828.0/65536.0,1,-nbitq), 
to_sfixed(3494.0/65536.0,1,-nbitq), 
to_sfixed(-1781.0/65536.0,1,-nbitq), 
to_sfixed(4176.0/65536.0,1,-nbitq), 
to_sfixed(-10373.0/65536.0,1,-nbitq), 
to_sfixed(-652.0/65536.0,1,-nbitq), 
to_sfixed(-753.0/65536.0,1,-nbitq), 
to_sfixed(-9379.0/65536.0,1,-nbitq), 
to_sfixed(-496.0/65536.0,1,-nbitq), 
to_sfixed(813.0/65536.0,1,-nbitq), 
to_sfixed(9743.0/65536.0,1,-nbitq), 
to_sfixed(-2319.0/65536.0,1,-nbitq), 
to_sfixed(-243.0/65536.0,1,-nbitq), 
to_sfixed(2456.0/65536.0,1,-nbitq), 
to_sfixed(4885.0/65536.0,1,-nbitq), 
to_sfixed(9209.0/65536.0,1,-nbitq), 
to_sfixed(-3126.0/65536.0,1,-nbitq), 
to_sfixed(6967.0/65536.0,1,-nbitq), 
to_sfixed(736.0/65536.0,1,-nbitq), 
to_sfixed(-6893.0/65536.0,1,-nbitq), 
to_sfixed(642.0/65536.0,1,-nbitq), 
to_sfixed(-984.0/65536.0,1,-nbitq), 
to_sfixed(-980.0/65536.0,1,-nbitq), 
to_sfixed(2409.0/65536.0,1,-nbitq), 
to_sfixed(-2356.0/65536.0,1,-nbitq), 
to_sfixed(-2059.0/65536.0,1,-nbitq), 
to_sfixed(-2385.0/65536.0,1,-nbitq), 
to_sfixed(-4363.0/65536.0,1,-nbitq), 
to_sfixed(2128.0/65536.0,1,-nbitq), 
to_sfixed(-1817.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5657.0/65536.0,1,-nbitq), 
to_sfixed(-789.0/65536.0,1,-nbitq), 
to_sfixed(-5890.0/65536.0,1,-nbitq), 
to_sfixed(-6279.0/65536.0,1,-nbitq), 
to_sfixed(449.0/65536.0,1,-nbitq), 
to_sfixed(4740.0/65536.0,1,-nbitq), 
to_sfixed(-8047.0/65536.0,1,-nbitq), 
to_sfixed(11632.0/65536.0,1,-nbitq), 
to_sfixed(3550.0/65536.0,1,-nbitq), 
to_sfixed(1564.0/65536.0,1,-nbitq), 
to_sfixed(-3049.0/65536.0,1,-nbitq), 
to_sfixed(-10071.0/65536.0,1,-nbitq), 
to_sfixed(899.0/65536.0,1,-nbitq), 
to_sfixed(3627.0/65536.0,1,-nbitq), 
to_sfixed(1817.0/65536.0,1,-nbitq), 
to_sfixed(1866.0/65536.0,1,-nbitq), 
to_sfixed(-2264.0/65536.0,1,-nbitq), 
to_sfixed(10048.0/65536.0,1,-nbitq), 
to_sfixed(-4145.0/65536.0,1,-nbitq), 
to_sfixed(-89.0/65536.0,1,-nbitq), 
to_sfixed(834.0/65536.0,1,-nbitq), 
to_sfixed(-12440.0/65536.0,1,-nbitq), 
to_sfixed(-1060.0/65536.0,1,-nbitq), 
to_sfixed(8580.0/65536.0,1,-nbitq), 
to_sfixed(1225.0/65536.0,1,-nbitq), 
to_sfixed(-12090.0/65536.0,1,-nbitq), 
to_sfixed(-12774.0/65536.0,1,-nbitq), 
to_sfixed(5188.0/65536.0,1,-nbitq), 
to_sfixed(-4432.0/65536.0,1,-nbitq), 
to_sfixed(-1428.0/65536.0,1,-nbitq), 
to_sfixed(5331.0/65536.0,1,-nbitq), 
to_sfixed(171.0/65536.0,1,-nbitq), 
to_sfixed(2770.0/65536.0,1,-nbitq), 
to_sfixed(-11961.0/65536.0,1,-nbitq), 
to_sfixed(912.0/65536.0,1,-nbitq), 
to_sfixed(-2277.0/65536.0,1,-nbitq), 
to_sfixed(-10315.0/65536.0,1,-nbitq), 
to_sfixed(4431.0/65536.0,1,-nbitq), 
to_sfixed(2580.0/65536.0,1,-nbitq), 
to_sfixed(-599.0/65536.0,1,-nbitq), 
to_sfixed(5984.0/65536.0,1,-nbitq), 
to_sfixed(1472.0/65536.0,1,-nbitq), 
to_sfixed(3957.0/65536.0,1,-nbitq), 
to_sfixed(8341.0/65536.0,1,-nbitq), 
to_sfixed(1504.0/65536.0,1,-nbitq), 
to_sfixed(-7728.0/65536.0,1,-nbitq), 
to_sfixed(5726.0/65536.0,1,-nbitq), 
to_sfixed(6310.0/65536.0,1,-nbitq), 
to_sfixed(-318.0/65536.0,1,-nbitq), 
to_sfixed(1039.0/65536.0,1,-nbitq), 
to_sfixed(1144.0/65536.0,1,-nbitq), 
to_sfixed(234.0/65536.0,1,-nbitq), 
to_sfixed(254.0/65536.0,1,-nbitq), 
to_sfixed(3421.0/65536.0,1,-nbitq), 
to_sfixed(-9717.0/65536.0,1,-nbitq), 
to_sfixed(-7044.0/65536.0,1,-nbitq), 
to_sfixed(433.0/65536.0,1,-nbitq), 
to_sfixed(-6052.0/65536.0,1,-nbitq), 
to_sfixed(1149.0/65536.0,1,-nbitq), 
to_sfixed(3539.0/65536.0,1,-nbitq), 
to_sfixed(17259.0/65536.0,1,-nbitq), 
to_sfixed(728.0/65536.0,1,-nbitq), 
to_sfixed(-2493.0/65536.0,1,-nbitq), 
to_sfixed(1135.0/65536.0,1,-nbitq), 
to_sfixed(8187.0/65536.0,1,-nbitq), 
to_sfixed(6082.0/65536.0,1,-nbitq), 
to_sfixed(-2425.0/65536.0,1,-nbitq), 
to_sfixed(9857.0/65536.0,1,-nbitq), 
to_sfixed(4357.0/65536.0,1,-nbitq), 
to_sfixed(-3738.0/65536.0,1,-nbitq), 
to_sfixed(32.0/65536.0,1,-nbitq), 
to_sfixed(4364.0/65536.0,1,-nbitq), 
to_sfixed(-2581.0/65536.0,1,-nbitq), 
to_sfixed(486.0/65536.0,1,-nbitq), 
to_sfixed(-1892.0/65536.0,1,-nbitq), 
to_sfixed(666.0/65536.0,1,-nbitq), 
to_sfixed(2806.0/65536.0,1,-nbitq), 
to_sfixed(-8164.0/65536.0,1,-nbitq), 
to_sfixed(1895.0/65536.0,1,-nbitq), 
to_sfixed(-2233.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1451.0/65536.0,1,-nbitq), 
to_sfixed(-5762.0/65536.0,1,-nbitq), 
to_sfixed(-6991.0/65536.0,1,-nbitq), 
to_sfixed(-5030.0/65536.0,1,-nbitq), 
to_sfixed(-3452.0/65536.0,1,-nbitq), 
to_sfixed(-1583.0/65536.0,1,-nbitq), 
to_sfixed(-4200.0/65536.0,1,-nbitq), 
to_sfixed(8307.0/65536.0,1,-nbitq), 
to_sfixed(-178.0/65536.0,1,-nbitq), 
to_sfixed(1534.0/65536.0,1,-nbitq), 
to_sfixed(-1154.0/65536.0,1,-nbitq), 
to_sfixed(-6470.0/65536.0,1,-nbitq), 
to_sfixed(2740.0/65536.0,1,-nbitq), 
to_sfixed(-4179.0/65536.0,1,-nbitq), 
to_sfixed(-2971.0/65536.0,1,-nbitq), 
to_sfixed(528.0/65536.0,1,-nbitq), 
to_sfixed(-1670.0/65536.0,1,-nbitq), 
to_sfixed(17070.0/65536.0,1,-nbitq), 
to_sfixed(-3677.0/65536.0,1,-nbitq), 
to_sfixed(-1590.0/65536.0,1,-nbitq), 
to_sfixed(-1648.0/65536.0,1,-nbitq), 
to_sfixed(-1402.0/65536.0,1,-nbitq), 
to_sfixed(5735.0/65536.0,1,-nbitq), 
to_sfixed(2091.0/65536.0,1,-nbitq), 
to_sfixed(1157.0/65536.0,1,-nbitq), 
to_sfixed(-8178.0/65536.0,1,-nbitq), 
to_sfixed(-16997.0/65536.0,1,-nbitq), 
to_sfixed(1129.0/65536.0,1,-nbitq), 
to_sfixed(-5036.0/65536.0,1,-nbitq), 
to_sfixed(857.0/65536.0,1,-nbitq), 
to_sfixed(3898.0/65536.0,1,-nbitq), 
to_sfixed(-213.0/65536.0,1,-nbitq), 
to_sfixed(4878.0/65536.0,1,-nbitq), 
to_sfixed(-8152.0/65536.0,1,-nbitq), 
to_sfixed(1690.0/65536.0,1,-nbitq), 
to_sfixed(-494.0/65536.0,1,-nbitq), 
to_sfixed(-1759.0/65536.0,1,-nbitq), 
to_sfixed(2251.0/65536.0,1,-nbitq), 
to_sfixed(214.0/65536.0,1,-nbitq), 
to_sfixed(4093.0/65536.0,1,-nbitq), 
to_sfixed(-2136.0/65536.0,1,-nbitq), 
to_sfixed(-2588.0/65536.0,1,-nbitq), 
to_sfixed(4032.0/65536.0,1,-nbitq), 
to_sfixed(3036.0/65536.0,1,-nbitq), 
to_sfixed(131.0/65536.0,1,-nbitq), 
to_sfixed(-6995.0/65536.0,1,-nbitq), 
to_sfixed(933.0/65536.0,1,-nbitq), 
to_sfixed(11859.0/65536.0,1,-nbitq), 
to_sfixed(2637.0/65536.0,1,-nbitq), 
to_sfixed(-1252.0/65536.0,1,-nbitq), 
to_sfixed(2499.0/65536.0,1,-nbitq), 
to_sfixed(1466.0/65536.0,1,-nbitq), 
to_sfixed(-371.0/65536.0,1,-nbitq), 
to_sfixed(-7502.0/65536.0,1,-nbitq), 
to_sfixed(-4659.0/65536.0,1,-nbitq), 
to_sfixed(-7767.0/65536.0,1,-nbitq), 
to_sfixed(1755.0/65536.0,1,-nbitq), 
to_sfixed(458.0/65536.0,1,-nbitq), 
to_sfixed(2375.0/65536.0,1,-nbitq), 
to_sfixed(4275.0/65536.0,1,-nbitq), 
to_sfixed(18110.0/65536.0,1,-nbitq), 
to_sfixed(1942.0/65536.0,1,-nbitq), 
to_sfixed(-1927.0/65536.0,1,-nbitq), 
to_sfixed(-458.0/65536.0,1,-nbitq), 
to_sfixed(10383.0/65536.0,1,-nbitq), 
to_sfixed(5525.0/65536.0,1,-nbitq), 
to_sfixed(-1898.0/65536.0,1,-nbitq), 
to_sfixed(2896.0/65536.0,1,-nbitq), 
to_sfixed(2458.0/65536.0,1,-nbitq), 
to_sfixed(3153.0/65536.0,1,-nbitq), 
to_sfixed(546.0/65536.0,1,-nbitq), 
to_sfixed(-3146.0/65536.0,1,-nbitq), 
to_sfixed(-4366.0/65536.0,1,-nbitq), 
to_sfixed(1616.0/65536.0,1,-nbitq), 
to_sfixed(-2266.0/65536.0,1,-nbitq), 
to_sfixed(-5079.0/65536.0,1,-nbitq), 
to_sfixed(-2255.0/65536.0,1,-nbitq), 
to_sfixed(-10951.0/65536.0,1,-nbitq), 
to_sfixed(633.0/65536.0,1,-nbitq), 
to_sfixed(-2585.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-387.0/65536.0,1,-nbitq), 
to_sfixed(-7468.0/65536.0,1,-nbitq), 
to_sfixed(-2660.0/65536.0,1,-nbitq), 
to_sfixed(-3508.0/65536.0,1,-nbitq), 
to_sfixed(-12506.0/65536.0,1,-nbitq), 
to_sfixed(1646.0/65536.0,1,-nbitq), 
to_sfixed(-4672.0/65536.0,1,-nbitq), 
to_sfixed(3805.0/65536.0,1,-nbitq), 
to_sfixed(-5298.0/65536.0,1,-nbitq), 
to_sfixed(-609.0/65536.0,1,-nbitq), 
to_sfixed(-2005.0/65536.0,1,-nbitq), 
to_sfixed(-3396.0/65536.0,1,-nbitq), 
to_sfixed(4116.0/65536.0,1,-nbitq), 
to_sfixed(-2398.0/65536.0,1,-nbitq), 
to_sfixed(-1839.0/65536.0,1,-nbitq), 
to_sfixed(-1437.0/65536.0,1,-nbitq), 
to_sfixed(-1242.0/65536.0,1,-nbitq), 
to_sfixed(2966.0/65536.0,1,-nbitq), 
to_sfixed(909.0/65536.0,1,-nbitq), 
to_sfixed(261.0/65536.0,1,-nbitq), 
to_sfixed(-1543.0/65536.0,1,-nbitq), 
to_sfixed(2328.0/65536.0,1,-nbitq), 
to_sfixed(-4320.0/65536.0,1,-nbitq), 
to_sfixed(-2005.0/65536.0,1,-nbitq), 
to_sfixed(-831.0/65536.0,1,-nbitq), 
to_sfixed(-7561.0/65536.0,1,-nbitq), 
to_sfixed(-12393.0/65536.0,1,-nbitq), 
to_sfixed(1758.0/65536.0,1,-nbitq), 
to_sfixed(-4864.0/65536.0,1,-nbitq), 
to_sfixed(610.0/65536.0,1,-nbitq), 
to_sfixed(-1994.0/65536.0,1,-nbitq), 
to_sfixed(-4175.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(555.0/65536.0,1,-nbitq), 
to_sfixed(-533.0/65536.0,1,-nbitq), 
to_sfixed(3228.0/65536.0,1,-nbitq), 
to_sfixed(-6070.0/65536.0,1,-nbitq), 
to_sfixed(550.0/65536.0,1,-nbitq), 
to_sfixed(-7331.0/65536.0,1,-nbitq), 
to_sfixed(2880.0/65536.0,1,-nbitq), 
to_sfixed(-2488.0/65536.0,1,-nbitq), 
to_sfixed(-1300.0/65536.0,1,-nbitq), 
to_sfixed(-7993.0/65536.0,1,-nbitq), 
to_sfixed(8265.0/65536.0,1,-nbitq), 
to_sfixed(2128.0/65536.0,1,-nbitq), 
to_sfixed(-5315.0/65536.0,1,-nbitq), 
to_sfixed(-2279.0/65536.0,1,-nbitq), 
to_sfixed(12082.0/65536.0,1,-nbitq), 
to_sfixed(504.0/65536.0,1,-nbitq), 
to_sfixed(-1683.0/65536.0,1,-nbitq), 
to_sfixed(2074.0/65536.0,1,-nbitq), 
to_sfixed(-2754.0/65536.0,1,-nbitq), 
to_sfixed(841.0/65536.0,1,-nbitq), 
to_sfixed(-9974.0/65536.0,1,-nbitq), 
to_sfixed(-5428.0/65536.0,1,-nbitq), 
to_sfixed(-3576.0/65536.0,1,-nbitq), 
to_sfixed(-1770.0/65536.0,1,-nbitq), 
to_sfixed(715.0/65536.0,1,-nbitq), 
to_sfixed(394.0/65536.0,1,-nbitq), 
to_sfixed(7959.0/65536.0,1,-nbitq), 
to_sfixed(59.0/65536.0,1,-nbitq), 
to_sfixed(-1101.0/65536.0,1,-nbitq), 
to_sfixed(-808.0/65536.0,1,-nbitq), 
to_sfixed(-3092.0/65536.0,1,-nbitq), 
to_sfixed(14074.0/65536.0,1,-nbitq), 
to_sfixed(20387.0/65536.0,1,-nbitq), 
to_sfixed(-269.0/65536.0,1,-nbitq), 
to_sfixed(7672.0/65536.0,1,-nbitq), 
to_sfixed(2284.0/65536.0,1,-nbitq), 
to_sfixed(6489.0/65536.0,1,-nbitq), 
to_sfixed(571.0/65536.0,1,-nbitq), 
to_sfixed(199.0/65536.0,1,-nbitq), 
to_sfixed(-8332.0/65536.0,1,-nbitq), 
to_sfixed(-1725.0/65536.0,1,-nbitq), 
to_sfixed(1598.0/65536.0,1,-nbitq), 
to_sfixed(-7714.0/65536.0,1,-nbitq), 
to_sfixed(-818.0/65536.0,1,-nbitq), 
to_sfixed(-3751.0/65536.0,1,-nbitq), 
to_sfixed(2331.0/65536.0,1,-nbitq), 
to_sfixed(-7952.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-509.0/65536.0,1,-nbitq), 
to_sfixed(-5591.0/65536.0,1,-nbitq), 
to_sfixed(-6952.0/65536.0,1,-nbitq), 
to_sfixed(-1949.0/65536.0,1,-nbitq), 
to_sfixed(-12877.0/65536.0,1,-nbitq), 
to_sfixed(5067.0/65536.0,1,-nbitq), 
to_sfixed(841.0/65536.0,1,-nbitq), 
to_sfixed(4770.0/65536.0,1,-nbitq), 
to_sfixed(-339.0/65536.0,1,-nbitq), 
to_sfixed(2119.0/65536.0,1,-nbitq), 
to_sfixed(-915.0/65536.0,1,-nbitq), 
to_sfixed(-4482.0/65536.0,1,-nbitq), 
to_sfixed(1477.0/65536.0,1,-nbitq), 
to_sfixed(-5941.0/65536.0,1,-nbitq), 
to_sfixed(-643.0/65536.0,1,-nbitq), 
to_sfixed(1883.0/65536.0,1,-nbitq), 
to_sfixed(787.0/65536.0,1,-nbitq), 
to_sfixed(-14496.0/65536.0,1,-nbitq), 
to_sfixed(6108.0/65536.0,1,-nbitq), 
to_sfixed(2926.0/65536.0,1,-nbitq), 
to_sfixed(-5525.0/65536.0,1,-nbitq), 
to_sfixed(2359.0/65536.0,1,-nbitq), 
to_sfixed(-8999.0/65536.0,1,-nbitq), 
to_sfixed(4073.0/65536.0,1,-nbitq), 
to_sfixed(-31.0/65536.0,1,-nbitq), 
to_sfixed(-10759.0/65536.0,1,-nbitq), 
to_sfixed(-2301.0/65536.0,1,-nbitq), 
to_sfixed(-1518.0/65536.0,1,-nbitq), 
to_sfixed(689.0/65536.0,1,-nbitq), 
to_sfixed(3810.0/65536.0,1,-nbitq), 
to_sfixed(-4249.0/65536.0,1,-nbitq), 
to_sfixed(-3294.0/65536.0,1,-nbitq), 
to_sfixed(3958.0/65536.0,1,-nbitq), 
to_sfixed(10411.0/65536.0,1,-nbitq), 
to_sfixed(2952.0/65536.0,1,-nbitq), 
to_sfixed(-1483.0/65536.0,1,-nbitq), 
to_sfixed(-7572.0/65536.0,1,-nbitq), 
to_sfixed(3251.0/65536.0,1,-nbitq), 
to_sfixed(-10362.0/65536.0,1,-nbitq), 
to_sfixed(89.0/65536.0,1,-nbitq), 
to_sfixed(8305.0/65536.0,1,-nbitq), 
to_sfixed(2176.0/65536.0,1,-nbitq), 
to_sfixed(-8169.0/65536.0,1,-nbitq), 
to_sfixed(3128.0/65536.0,1,-nbitq), 
to_sfixed(2934.0/65536.0,1,-nbitq), 
to_sfixed(-2274.0/65536.0,1,-nbitq), 
to_sfixed(-2954.0/65536.0,1,-nbitq), 
to_sfixed(7211.0/65536.0,1,-nbitq), 
to_sfixed(2630.0/65536.0,1,-nbitq), 
to_sfixed(2278.0/65536.0,1,-nbitq), 
to_sfixed(-2544.0/65536.0,1,-nbitq), 
to_sfixed(-7311.0/65536.0,1,-nbitq), 
to_sfixed(1402.0/65536.0,1,-nbitq), 
to_sfixed(-9713.0/65536.0,1,-nbitq), 
to_sfixed(-549.0/65536.0,1,-nbitq), 
to_sfixed(-4391.0/65536.0,1,-nbitq), 
to_sfixed(-1344.0/65536.0,1,-nbitq), 
to_sfixed(2588.0/65536.0,1,-nbitq), 
to_sfixed(-2212.0/65536.0,1,-nbitq), 
to_sfixed(5691.0/65536.0,1,-nbitq), 
to_sfixed(-13850.0/65536.0,1,-nbitq), 
to_sfixed(-85.0/65536.0,1,-nbitq), 
to_sfixed(-1227.0/65536.0,1,-nbitq), 
to_sfixed(-48.0/65536.0,1,-nbitq), 
to_sfixed(16198.0/65536.0,1,-nbitq), 
to_sfixed(-2659.0/65536.0,1,-nbitq), 
to_sfixed(4798.0/65536.0,1,-nbitq), 
to_sfixed(9330.0/65536.0,1,-nbitq), 
to_sfixed(3486.0/65536.0,1,-nbitq), 
to_sfixed(3748.0/65536.0,1,-nbitq), 
to_sfixed(-5454.0/65536.0,1,-nbitq), 
to_sfixed(1488.0/65536.0,1,-nbitq), 
to_sfixed(-9866.0/65536.0,1,-nbitq), 
to_sfixed(2985.0/65536.0,1,-nbitq), 
to_sfixed(-137.0/65536.0,1,-nbitq), 
to_sfixed(-13376.0/65536.0,1,-nbitq), 
to_sfixed(1149.0/65536.0,1,-nbitq), 
to_sfixed(11628.0/65536.0,1,-nbitq), 
to_sfixed(-2598.0/65536.0,1,-nbitq), 
to_sfixed(-6191.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4670.0/65536.0,1,-nbitq), 
to_sfixed(-5402.0/65536.0,1,-nbitq), 
to_sfixed(-6742.0/65536.0,1,-nbitq), 
to_sfixed(-5916.0/65536.0,1,-nbitq), 
to_sfixed(-8143.0/65536.0,1,-nbitq), 
to_sfixed(1154.0/65536.0,1,-nbitq), 
to_sfixed(672.0/65536.0,1,-nbitq), 
to_sfixed(-7156.0/65536.0,1,-nbitq), 
to_sfixed(3500.0/65536.0,1,-nbitq), 
to_sfixed(1567.0/65536.0,1,-nbitq), 
to_sfixed(-4008.0/65536.0,1,-nbitq), 
to_sfixed(-1552.0/65536.0,1,-nbitq), 
to_sfixed(3974.0/65536.0,1,-nbitq), 
to_sfixed(-4084.0/65536.0,1,-nbitq), 
to_sfixed(-4490.0/65536.0,1,-nbitq), 
to_sfixed(576.0/65536.0,1,-nbitq), 
to_sfixed(1798.0/65536.0,1,-nbitq), 
to_sfixed(-7782.0/65536.0,1,-nbitq), 
to_sfixed(4938.0/65536.0,1,-nbitq), 
to_sfixed(267.0/65536.0,1,-nbitq), 
to_sfixed(-3798.0/65536.0,1,-nbitq), 
to_sfixed(9023.0/65536.0,1,-nbitq), 
to_sfixed(-1972.0/65536.0,1,-nbitq), 
to_sfixed(2375.0/65536.0,1,-nbitq), 
to_sfixed(-1634.0/65536.0,1,-nbitq), 
to_sfixed(-3162.0/65536.0,1,-nbitq), 
to_sfixed(2846.0/65536.0,1,-nbitq), 
to_sfixed(-2340.0/65536.0,1,-nbitq), 
to_sfixed(5201.0/65536.0,1,-nbitq), 
to_sfixed(2228.0/65536.0,1,-nbitq), 
to_sfixed(-2025.0/65536.0,1,-nbitq), 
to_sfixed(2001.0/65536.0,1,-nbitq), 
to_sfixed(5377.0/65536.0,1,-nbitq), 
to_sfixed(10030.0/65536.0,1,-nbitq), 
to_sfixed(2551.0/65536.0,1,-nbitq), 
to_sfixed(2921.0/65536.0,1,-nbitq), 
to_sfixed(-10784.0/65536.0,1,-nbitq), 
to_sfixed(6388.0/65536.0,1,-nbitq), 
to_sfixed(5746.0/65536.0,1,-nbitq), 
to_sfixed(-1362.0/65536.0,1,-nbitq), 
to_sfixed(12829.0/65536.0,1,-nbitq), 
to_sfixed(-337.0/65536.0,1,-nbitq), 
to_sfixed(2897.0/65536.0,1,-nbitq), 
to_sfixed(8108.0/65536.0,1,-nbitq), 
to_sfixed(107.0/65536.0,1,-nbitq), 
to_sfixed(-4282.0/65536.0,1,-nbitq), 
to_sfixed(-5784.0/65536.0,1,-nbitq), 
to_sfixed(6190.0/65536.0,1,-nbitq), 
to_sfixed(3329.0/65536.0,1,-nbitq), 
to_sfixed(2683.0/65536.0,1,-nbitq), 
to_sfixed(723.0/65536.0,1,-nbitq), 
to_sfixed(1116.0/65536.0,1,-nbitq), 
to_sfixed(5070.0/65536.0,1,-nbitq), 
to_sfixed(5537.0/65536.0,1,-nbitq), 
to_sfixed(-2975.0/65536.0,1,-nbitq), 
to_sfixed(-654.0/65536.0,1,-nbitq), 
to_sfixed(-2372.0/65536.0,1,-nbitq), 
to_sfixed(4597.0/65536.0,1,-nbitq), 
to_sfixed(-2776.0/65536.0,1,-nbitq), 
to_sfixed(10771.0/65536.0,1,-nbitq), 
to_sfixed(-15691.0/65536.0,1,-nbitq), 
to_sfixed(-1820.0/65536.0,1,-nbitq), 
to_sfixed(-2698.0/65536.0,1,-nbitq), 
to_sfixed(-775.0/65536.0,1,-nbitq), 
to_sfixed(9659.0/65536.0,1,-nbitq), 
to_sfixed(-15464.0/65536.0,1,-nbitq), 
to_sfixed(-241.0/65536.0,1,-nbitq), 
to_sfixed(3486.0/65536.0,1,-nbitq), 
to_sfixed(8508.0/65536.0,1,-nbitq), 
to_sfixed(6758.0/65536.0,1,-nbitq), 
to_sfixed(-3961.0/65536.0,1,-nbitq), 
to_sfixed(-4566.0/65536.0,1,-nbitq), 
to_sfixed(-9590.0/65536.0,1,-nbitq), 
to_sfixed(-1063.0/65536.0,1,-nbitq), 
to_sfixed(2790.0/65536.0,1,-nbitq), 
to_sfixed(-11586.0/65536.0,1,-nbitq), 
to_sfixed(-936.0/65536.0,1,-nbitq), 
to_sfixed(3798.0/65536.0,1,-nbitq), 
to_sfixed(80.0/65536.0,1,-nbitq), 
to_sfixed(2026.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-6616.0/65536.0,1,-nbitq), 
to_sfixed(-317.0/65536.0,1,-nbitq), 
to_sfixed(-10038.0/65536.0,1,-nbitq), 
to_sfixed(-3525.0/65536.0,1,-nbitq), 
to_sfixed(-6493.0/65536.0,1,-nbitq), 
to_sfixed(2899.0/65536.0,1,-nbitq), 
to_sfixed(3887.0/65536.0,1,-nbitq), 
to_sfixed(-7850.0/65536.0,1,-nbitq), 
to_sfixed(350.0/65536.0,1,-nbitq), 
to_sfixed(-2521.0/65536.0,1,-nbitq), 
to_sfixed(-8551.0/65536.0,1,-nbitq), 
to_sfixed(-370.0/65536.0,1,-nbitq), 
to_sfixed(4738.0/65536.0,1,-nbitq), 
to_sfixed(-8667.0/65536.0,1,-nbitq), 
to_sfixed(-3238.0/65536.0,1,-nbitq), 
to_sfixed(-1112.0/65536.0,1,-nbitq), 
to_sfixed(922.0/65536.0,1,-nbitq), 
to_sfixed(-3763.0/65536.0,1,-nbitq), 
to_sfixed(603.0/65536.0,1,-nbitq), 
to_sfixed(-1098.0/65536.0,1,-nbitq), 
to_sfixed(298.0/65536.0,1,-nbitq), 
to_sfixed(8941.0/65536.0,1,-nbitq), 
to_sfixed(-4247.0/65536.0,1,-nbitq), 
to_sfixed(3142.0/65536.0,1,-nbitq), 
to_sfixed(-3660.0/65536.0,1,-nbitq), 
to_sfixed(-6055.0/65536.0,1,-nbitq), 
to_sfixed(781.0/65536.0,1,-nbitq), 
to_sfixed(-1305.0/65536.0,1,-nbitq), 
to_sfixed(19855.0/65536.0,1,-nbitq), 
to_sfixed(-1853.0/65536.0,1,-nbitq), 
to_sfixed(3794.0/65536.0,1,-nbitq), 
to_sfixed(635.0/65536.0,1,-nbitq), 
to_sfixed(-2572.0/65536.0,1,-nbitq), 
to_sfixed(12702.0/65536.0,1,-nbitq), 
to_sfixed(1543.0/65536.0,1,-nbitq), 
to_sfixed(768.0/65536.0,1,-nbitq), 
to_sfixed(-6165.0/65536.0,1,-nbitq), 
to_sfixed(11915.0/65536.0,1,-nbitq), 
to_sfixed(22391.0/65536.0,1,-nbitq), 
to_sfixed(-3642.0/65536.0,1,-nbitq), 
to_sfixed(16196.0/65536.0,1,-nbitq), 
to_sfixed(-1270.0/65536.0,1,-nbitq), 
to_sfixed(3504.0/65536.0,1,-nbitq), 
to_sfixed(6836.0/65536.0,1,-nbitq), 
to_sfixed(1769.0/65536.0,1,-nbitq), 
to_sfixed(906.0/65536.0,1,-nbitq), 
to_sfixed(-3899.0/65536.0,1,-nbitq), 
to_sfixed(3694.0/65536.0,1,-nbitq), 
to_sfixed(2711.0/65536.0,1,-nbitq), 
to_sfixed(319.0/65536.0,1,-nbitq), 
to_sfixed(1441.0/65536.0,1,-nbitq), 
to_sfixed(3405.0/65536.0,1,-nbitq), 
to_sfixed(9083.0/65536.0,1,-nbitq), 
to_sfixed(-2173.0/65536.0,1,-nbitq), 
to_sfixed(6625.0/65536.0,1,-nbitq), 
to_sfixed(-14896.0/65536.0,1,-nbitq), 
to_sfixed(-2641.0/65536.0,1,-nbitq), 
to_sfixed(2949.0/65536.0,1,-nbitq), 
to_sfixed(1743.0/65536.0,1,-nbitq), 
to_sfixed(5461.0/65536.0,1,-nbitq), 
to_sfixed(-11314.0/65536.0,1,-nbitq), 
to_sfixed(2400.0/65536.0,1,-nbitq), 
to_sfixed(834.0/65536.0,1,-nbitq), 
to_sfixed(-3071.0/65536.0,1,-nbitq), 
to_sfixed(1051.0/65536.0,1,-nbitq), 
to_sfixed(-12173.0/65536.0,1,-nbitq), 
to_sfixed(-8984.0/65536.0,1,-nbitq), 
to_sfixed(-220.0/65536.0,1,-nbitq), 
to_sfixed(4410.0/65536.0,1,-nbitq), 
to_sfixed(-3966.0/65536.0,1,-nbitq), 
to_sfixed(-5404.0/65536.0,1,-nbitq), 
to_sfixed(-6914.0/65536.0,1,-nbitq), 
to_sfixed(-17756.0/65536.0,1,-nbitq), 
to_sfixed(-910.0/65536.0,1,-nbitq), 
to_sfixed(-887.0/65536.0,1,-nbitq), 
to_sfixed(-7518.0/65536.0,1,-nbitq), 
to_sfixed(2823.0/65536.0,1,-nbitq), 
to_sfixed(3862.0/65536.0,1,-nbitq), 
to_sfixed(-1936.0/65536.0,1,-nbitq), 
to_sfixed(-468.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-7971.0/65536.0,1,-nbitq), 
to_sfixed(2406.0/65536.0,1,-nbitq), 
to_sfixed(-786.0/65536.0,1,-nbitq), 
to_sfixed(-7150.0/65536.0,1,-nbitq), 
to_sfixed(6116.0/65536.0,1,-nbitq), 
to_sfixed(7300.0/65536.0,1,-nbitq), 
to_sfixed(6.0/65536.0,1,-nbitq), 
to_sfixed(-350.0/65536.0,1,-nbitq), 
to_sfixed(2546.0/65536.0,1,-nbitq), 
to_sfixed(1060.0/65536.0,1,-nbitq), 
to_sfixed(-2980.0/65536.0,1,-nbitq), 
to_sfixed(3237.0/65536.0,1,-nbitq), 
to_sfixed(469.0/65536.0,1,-nbitq), 
to_sfixed(-2105.0/65536.0,1,-nbitq), 
to_sfixed(-2270.0/65536.0,1,-nbitq), 
to_sfixed(-3170.0/65536.0,1,-nbitq), 
to_sfixed(-845.0/65536.0,1,-nbitq), 
to_sfixed(-1265.0/65536.0,1,-nbitq), 
to_sfixed(361.0/65536.0,1,-nbitq), 
to_sfixed(2309.0/65536.0,1,-nbitq), 
to_sfixed(5445.0/65536.0,1,-nbitq), 
to_sfixed(3762.0/65536.0,1,-nbitq), 
to_sfixed(228.0/65536.0,1,-nbitq), 
to_sfixed(-286.0/65536.0,1,-nbitq), 
to_sfixed(-12054.0/65536.0,1,-nbitq), 
to_sfixed(-5842.0/65536.0,1,-nbitq), 
to_sfixed(7334.0/65536.0,1,-nbitq), 
to_sfixed(1739.0/65536.0,1,-nbitq), 
to_sfixed(17306.0/65536.0,1,-nbitq), 
to_sfixed(-6.0/65536.0,1,-nbitq), 
to_sfixed(8294.0/65536.0,1,-nbitq), 
to_sfixed(10153.0/65536.0,1,-nbitq), 
to_sfixed(-3945.0/65536.0,1,-nbitq), 
to_sfixed(473.0/65536.0,1,-nbitq), 
to_sfixed(-1478.0/65536.0,1,-nbitq), 
to_sfixed(1263.0/65536.0,1,-nbitq), 
to_sfixed(-11420.0/65536.0,1,-nbitq), 
to_sfixed(18527.0/65536.0,1,-nbitq), 
to_sfixed(7787.0/65536.0,1,-nbitq), 
to_sfixed(481.0/65536.0,1,-nbitq), 
to_sfixed(18162.0/65536.0,1,-nbitq), 
to_sfixed(-3241.0/65536.0,1,-nbitq), 
to_sfixed(-1923.0/65536.0,1,-nbitq), 
to_sfixed(9634.0/65536.0,1,-nbitq), 
to_sfixed(1969.0/65536.0,1,-nbitq), 
to_sfixed(4366.0/65536.0,1,-nbitq), 
to_sfixed(-2005.0/65536.0,1,-nbitq), 
to_sfixed(-124.0/65536.0,1,-nbitq), 
to_sfixed(-2306.0/65536.0,1,-nbitq), 
to_sfixed(-1025.0/65536.0,1,-nbitq), 
to_sfixed(-1464.0/65536.0,1,-nbitq), 
to_sfixed(3272.0/65536.0,1,-nbitq), 
to_sfixed(8037.0/65536.0,1,-nbitq), 
to_sfixed(-1263.0/65536.0,1,-nbitq), 
to_sfixed(9294.0/65536.0,1,-nbitq), 
to_sfixed(-10480.0/65536.0,1,-nbitq), 
to_sfixed(-1480.0/65536.0,1,-nbitq), 
to_sfixed(-1532.0/65536.0,1,-nbitq), 
to_sfixed(-3145.0/65536.0,1,-nbitq), 
to_sfixed(9291.0/65536.0,1,-nbitq), 
to_sfixed(-798.0/65536.0,1,-nbitq), 
to_sfixed(465.0/65536.0,1,-nbitq), 
to_sfixed(1928.0/65536.0,1,-nbitq), 
to_sfixed(2316.0/65536.0,1,-nbitq), 
to_sfixed(-1866.0/65536.0,1,-nbitq), 
to_sfixed(-11471.0/65536.0,1,-nbitq), 
to_sfixed(-10283.0/65536.0,1,-nbitq), 
to_sfixed(-1369.0/65536.0,1,-nbitq), 
to_sfixed(2568.0/65536.0,1,-nbitq), 
to_sfixed(-12205.0/65536.0,1,-nbitq), 
to_sfixed(1064.0/65536.0,1,-nbitq), 
to_sfixed(-9093.0/65536.0,1,-nbitq), 
to_sfixed(-3774.0/65536.0,1,-nbitq), 
to_sfixed(-402.0/65536.0,1,-nbitq), 
to_sfixed(314.0/65536.0,1,-nbitq), 
to_sfixed(3527.0/65536.0,1,-nbitq), 
to_sfixed(3368.0/65536.0,1,-nbitq), 
to_sfixed(783.0/65536.0,1,-nbitq), 
to_sfixed(-2309.0/65536.0,1,-nbitq), 
to_sfixed(1648.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-6484.0/65536.0,1,-nbitq), 
to_sfixed(1823.0/65536.0,1,-nbitq), 
to_sfixed(1412.0/65536.0,1,-nbitq), 
to_sfixed(-3271.0/65536.0,1,-nbitq), 
to_sfixed(-2073.0/65536.0,1,-nbitq), 
to_sfixed(-2182.0/65536.0,1,-nbitq), 
to_sfixed(1160.0/65536.0,1,-nbitq), 
to_sfixed(8801.0/65536.0,1,-nbitq), 
to_sfixed(-4118.0/65536.0,1,-nbitq), 
to_sfixed(2802.0/65536.0,1,-nbitq), 
to_sfixed(-3347.0/65536.0,1,-nbitq), 
to_sfixed(-6149.0/65536.0,1,-nbitq), 
to_sfixed(869.0/65536.0,1,-nbitq), 
to_sfixed(1948.0/65536.0,1,-nbitq), 
to_sfixed(-665.0/65536.0,1,-nbitq), 
to_sfixed(-2778.0/65536.0,1,-nbitq), 
to_sfixed(781.0/65536.0,1,-nbitq), 
to_sfixed(-2650.0/65536.0,1,-nbitq), 
to_sfixed(1480.0/65536.0,1,-nbitq), 
to_sfixed(1900.0/65536.0,1,-nbitq), 
to_sfixed(-2960.0/65536.0,1,-nbitq), 
to_sfixed(11080.0/65536.0,1,-nbitq), 
to_sfixed(8754.0/65536.0,1,-nbitq), 
to_sfixed(-3608.0/65536.0,1,-nbitq), 
to_sfixed(-12900.0/65536.0,1,-nbitq), 
to_sfixed(-3208.0/65536.0,1,-nbitq), 
to_sfixed(8341.0/65536.0,1,-nbitq), 
to_sfixed(3979.0/65536.0,1,-nbitq), 
to_sfixed(16473.0/65536.0,1,-nbitq), 
to_sfixed(4080.0/65536.0,1,-nbitq), 
to_sfixed(4651.0/65536.0,1,-nbitq), 
to_sfixed(13055.0/65536.0,1,-nbitq), 
to_sfixed(2175.0/65536.0,1,-nbitq), 
to_sfixed(-9199.0/65536.0,1,-nbitq), 
to_sfixed(-2758.0/65536.0,1,-nbitq), 
to_sfixed(509.0/65536.0,1,-nbitq), 
to_sfixed(-7581.0/65536.0,1,-nbitq), 
to_sfixed(6051.0/65536.0,1,-nbitq), 
to_sfixed(-5346.0/65536.0,1,-nbitq), 
to_sfixed(4369.0/65536.0,1,-nbitq), 
to_sfixed(11082.0/65536.0,1,-nbitq), 
to_sfixed(1027.0/65536.0,1,-nbitq), 
to_sfixed(-603.0/65536.0,1,-nbitq), 
to_sfixed(5414.0/65536.0,1,-nbitq), 
to_sfixed(-2425.0/65536.0,1,-nbitq), 
to_sfixed(697.0/65536.0,1,-nbitq), 
to_sfixed(-1127.0/65536.0,1,-nbitq), 
to_sfixed(683.0/65536.0,1,-nbitq), 
to_sfixed(-2777.0/65536.0,1,-nbitq), 
to_sfixed(2478.0/65536.0,1,-nbitq), 
to_sfixed(-762.0/65536.0,1,-nbitq), 
to_sfixed(-479.0/65536.0,1,-nbitq), 
to_sfixed(3417.0/65536.0,1,-nbitq), 
to_sfixed(2606.0/65536.0,1,-nbitq), 
to_sfixed(13352.0/65536.0,1,-nbitq), 
to_sfixed(-9485.0/65536.0,1,-nbitq), 
to_sfixed(-125.0/65536.0,1,-nbitq), 
to_sfixed(-5907.0/65536.0,1,-nbitq), 
to_sfixed(-1270.0/65536.0,1,-nbitq), 
to_sfixed(2284.0/65536.0,1,-nbitq), 
to_sfixed(3473.0/65536.0,1,-nbitq), 
to_sfixed(-1409.0/65536.0,1,-nbitq), 
to_sfixed(1204.0/65536.0,1,-nbitq), 
to_sfixed(-1842.0/65536.0,1,-nbitq), 
to_sfixed(-6020.0/65536.0,1,-nbitq), 
to_sfixed(-11126.0/65536.0,1,-nbitq), 
to_sfixed(-5970.0/65536.0,1,-nbitq), 
to_sfixed(-431.0/65536.0,1,-nbitq), 
to_sfixed(-2569.0/65536.0,1,-nbitq), 
to_sfixed(-11191.0/65536.0,1,-nbitq), 
to_sfixed(4693.0/65536.0,1,-nbitq), 
to_sfixed(-319.0/65536.0,1,-nbitq), 
to_sfixed(1008.0/65536.0,1,-nbitq), 
to_sfixed(-649.0/65536.0,1,-nbitq), 
to_sfixed(-230.0/65536.0,1,-nbitq), 
to_sfixed(11814.0/65536.0,1,-nbitq), 
to_sfixed(935.0/65536.0,1,-nbitq), 
to_sfixed(-3819.0/65536.0,1,-nbitq), 
to_sfixed(-259.0/65536.0,1,-nbitq), 
to_sfixed(3722.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3784.0/65536.0,1,-nbitq), 
to_sfixed(-2071.0/65536.0,1,-nbitq), 
to_sfixed(-2309.0/65536.0,1,-nbitq), 
to_sfixed(-5029.0/65536.0,1,-nbitq), 
to_sfixed(-4875.0/65536.0,1,-nbitq), 
to_sfixed(-1517.0/65536.0,1,-nbitq), 
to_sfixed(4838.0/65536.0,1,-nbitq), 
to_sfixed(4629.0/65536.0,1,-nbitq), 
to_sfixed(-4060.0/65536.0,1,-nbitq), 
to_sfixed(753.0/65536.0,1,-nbitq), 
to_sfixed(-613.0/65536.0,1,-nbitq), 
to_sfixed(-3170.0/65536.0,1,-nbitq), 
to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(4966.0/65536.0,1,-nbitq), 
to_sfixed(-193.0/65536.0,1,-nbitq), 
to_sfixed(-1259.0/65536.0,1,-nbitq), 
to_sfixed(3033.0/65536.0,1,-nbitq), 
to_sfixed(-7657.0/65536.0,1,-nbitq), 
to_sfixed(-2135.0/65536.0,1,-nbitq), 
to_sfixed(2409.0/65536.0,1,-nbitq), 
to_sfixed(-2460.0/65536.0,1,-nbitq), 
to_sfixed(11624.0/65536.0,1,-nbitq), 
to_sfixed(6272.0/65536.0,1,-nbitq), 
to_sfixed(-8942.0/65536.0,1,-nbitq), 
to_sfixed(-10847.0/65536.0,1,-nbitq), 
to_sfixed(-11272.0/65536.0,1,-nbitq), 
to_sfixed(-1144.0/65536.0,1,-nbitq), 
to_sfixed(2783.0/65536.0,1,-nbitq), 
to_sfixed(15925.0/65536.0,1,-nbitq), 
to_sfixed(1128.0/65536.0,1,-nbitq), 
to_sfixed(1270.0/65536.0,1,-nbitq), 
to_sfixed(16567.0/65536.0,1,-nbitq), 
to_sfixed(1761.0/65536.0,1,-nbitq), 
to_sfixed(-9533.0/65536.0,1,-nbitq), 
to_sfixed(-3165.0/65536.0,1,-nbitq), 
to_sfixed(1318.0/65536.0,1,-nbitq), 
to_sfixed(1639.0/65536.0,1,-nbitq), 
to_sfixed(4406.0/65536.0,1,-nbitq), 
to_sfixed(-9103.0/65536.0,1,-nbitq), 
to_sfixed(4342.0/65536.0,1,-nbitq), 
to_sfixed(2070.0/65536.0,1,-nbitq), 
to_sfixed(-1885.0/65536.0,1,-nbitq), 
to_sfixed(9046.0/65536.0,1,-nbitq), 
to_sfixed(5559.0/65536.0,1,-nbitq), 
to_sfixed(2981.0/65536.0,1,-nbitq), 
to_sfixed(-5524.0/65536.0,1,-nbitq), 
to_sfixed(1605.0/65536.0,1,-nbitq), 
to_sfixed(2939.0/65536.0,1,-nbitq), 
to_sfixed(2417.0/65536.0,1,-nbitq), 
to_sfixed(2722.0/65536.0,1,-nbitq), 
to_sfixed(-2215.0/65536.0,1,-nbitq), 
to_sfixed(1844.0/65536.0,1,-nbitq), 
to_sfixed(2688.0/65536.0,1,-nbitq), 
to_sfixed(-229.0/65536.0,1,-nbitq), 
to_sfixed(4297.0/65536.0,1,-nbitq), 
to_sfixed(-8227.0/65536.0,1,-nbitq), 
to_sfixed(-1600.0/65536.0,1,-nbitq), 
to_sfixed(-3510.0/65536.0,1,-nbitq), 
to_sfixed(-3114.0/65536.0,1,-nbitq), 
to_sfixed(-3135.0/65536.0,1,-nbitq), 
to_sfixed(6891.0/65536.0,1,-nbitq), 
to_sfixed(-2962.0/65536.0,1,-nbitq), 
to_sfixed(225.0/65536.0,1,-nbitq), 
to_sfixed(-2107.0/65536.0,1,-nbitq), 
to_sfixed(-6067.0/65536.0,1,-nbitq), 
to_sfixed(-19303.0/65536.0,1,-nbitq), 
to_sfixed(1765.0/65536.0,1,-nbitq), 
to_sfixed(-5206.0/65536.0,1,-nbitq), 
to_sfixed(902.0/65536.0,1,-nbitq), 
to_sfixed(-3014.0/65536.0,1,-nbitq), 
to_sfixed(6675.0/65536.0,1,-nbitq), 
to_sfixed(-3836.0/65536.0,1,-nbitq), 
to_sfixed(8423.0/65536.0,1,-nbitq), 
to_sfixed(-329.0/65536.0,1,-nbitq), 
to_sfixed(1603.0/65536.0,1,-nbitq), 
to_sfixed(824.0/65536.0,1,-nbitq), 
to_sfixed(1718.0/65536.0,1,-nbitq), 
to_sfixed(-3495.0/65536.0,1,-nbitq), 
to_sfixed(-1351.0/65536.0,1,-nbitq), 
to_sfixed(1396.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2341.0/65536.0,1,-nbitq), 
to_sfixed(-4901.0/65536.0,1,-nbitq), 
to_sfixed(1343.0/65536.0,1,-nbitq), 
to_sfixed(-1883.0/65536.0,1,-nbitq), 
to_sfixed(-2578.0/65536.0,1,-nbitq), 
to_sfixed(343.0/65536.0,1,-nbitq), 
to_sfixed(205.0/65536.0,1,-nbitq), 
to_sfixed(-3372.0/65536.0,1,-nbitq), 
to_sfixed(2054.0/65536.0,1,-nbitq), 
to_sfixed(174.0/65536.0,1,-nbitq), 
to_sfixed(-861.0/65536.0,1,-nbitq), 
to_sfixed(-1646.0/65536.0,1,-nbitq), 
to_sfixed(2897.0/65536.0,1,-nbitq), 
to_sfixed(7111.0/65536.0,1,-nbitq), 
to_sfixed(1248.0/65536.0,1,-nbitq), 
to_sfixed(1360.0/65536.0,1,-nbitq), 
to_sfixed(3084.0/65536.0,1,-nbitq), 
to_sfixed(-7244.0/65536.0,1,-nbitq), 
to_sfixed(-5609.0/65536.0,1,-nbitq), 
to_sfixed(309.0/65536.0,1,-nbitq), 
to_sfixed(1529.0/65536.0,1,-nbitq), 
to_sfixed(10124.0/65536.0,1,-nbitq), 
to_sfixed(9870.0/65536.0,1,-nbitq), 
to_sfixed(-3450.0/65536.0,1,-nbitq), 
to_sfixed(-10429.0/65536.0,1,-nbitq), 
to_sfixed(-9441.0/65536.0,1,-nbitq), 
to_sfixed(-1220.0/65536.0,1,-nbitq), 
to_sfixed(1742.0/65536.0,1,-nbitq), 
to_sfixed(19087.0/65536.0,1,-nbitq), 
to_sfixed(2988.0/65536.0,1,-nbitq), 
to_sfixed(-1190.0/65536.0,1,-nbitq), 
to_sfixed(6715.0/65536.0,1,-nbitq), 
to_sfixed(-4483.0/65536.0,1,-nbitq), 
to_sfixed(-7209.0/65536.0,1,-nbitq), 
to_sfixed(988.0/65536.0,1,-nbitq), 
to_sfixed(-3925.0/65536.0,1,-nbitq), 
to_sfixed(-6131.0/65536.0,1,-nbitq), 
to_sfixed(-317.0/65536.0,1,-nbitq), 
to_sfixed(-8258.0/65536.0,1,-nbitq), 
to_sfixed(-1800.0/65536.0,1,-nbitq), 
to_sfixed(-907.0/65536.0,1,-nbitq), 
to_sfixed(2758.0/65536.0,1,-nbitq), 
to_sfixed(433.0/65536.0,1,-nbitq), 
to_sfixed(5159.0/65536.0,1,-nbitq), 
to_sfixed(1441.0/65536.0,1,-nbitq), 
to_sfixed(-7470.0/65536.0,1,-nbitq), 
to_sfixed(-1206.0/65536.0,1,-nbitq), 
to_sfixed(7094.0/65536.0,1,-nbitq), 
to_sfixed(2480.0/65536.0,1,-nbitq), 
to_sfixed(-621.0/65536.0,1,-nbitq), 
to_sfixed(1074.0/65536.0,1,-nbitq), 
to_sfixed(688.0/65536.0,1,-nbitq), 
to_sfixed(2912.0/65536.0,1,-nbitq), 
to_sfixed(-411.0/65536.0,1,-nbitq), 
to_sfixed(6446.0/65536.0,1,-nbitq), 
to_sfixed(-4873.0/65536.0,1,-nbitq), 
to_sfixed(-1403.0/65536.0,1,-nbitq), 
to_sfixed(-4766.0/65536.0,1,-nbitq), 
to_sfixed(270.0/65536.0,1,-nbitq), 
to_sfixed(-7173.0/65536.0,1,-nbitq), 
to_sfixed(6390.0/65536.0,1,-nbitq), 
to_sfixed(2626.0/65536.0,1,-nbitq), 
to_sfixed(2506.0/65536.0,1,-nbitq), 
to_sfixed(-3016.0/65536.0,1,-nbitq), 
to_sfixed(-8203.0/65536.0,1,-nbitq), 
to_sfixed(-10618.0/65536.0,1,-nbitq), 
to_sfixed(-1545.0/65536.0,1,-nbitq), 
to_sfixed(-3252.0/65536.0,1,-nbitq), 
to_sfixed(2517.0/65536.0,1,-nbitq), 
to_sfixed(1229.0/65536.0,1,-nbitq), 
to_sfixed(3313.0/65536.0,1,-nbitq), 
to_sfixed(1730.0/65536.0,1,-nbitq), 
to_sfixed(1638.0/65536.0,1,-nbitq), 
to_sfixed(-520.0/65536.0,1,-nbitq), 
to_sfixed(1944.0/65536.0,1,-nbitq), 
to_sfixed(434.0/65536.0,1,-nbitq), 
to_sfixed(129.0/65536.0,1,-nbitq), 
to_sfixed(-3595.0/65536.0,1,-nbitq), 
to_sfixed(1012.0/65536.0,1,-nbitq), 
to_sfixed(-748.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1474.0/65536.0,1,-nbitq), 
to_sfixed(-3000.0/65536.0,1,-nbitq), 
to_sfixed(4347.0/65536.0,1,-nbitq), 
to_sfixed(2350.0/65536.0,1,-nbitq), 
to_sfixed(-6696.0/65536.0,1,-nbitq), 
to_sfixed(-1049.0/65536.0,1,-nbitq), 
to_sfixed(2428.0/65536.0,1,-nbitq), 
to_sfixed(-1353.0/65536.0,1,-nbitq), 
to_sfixed(3807.0/65536.0,1,-nbitq), 
to_sfixed(-832.0/65536.0,1,-nbitq), 
to_sfixed(-177.0/65536.0,1,-nbitq), 
to_sfixed(-82.0/65536.0,1,-nbitq), 
to_sfixed(146.0/65536.0,1,-nbitq), 
to_sfixed(-2815.0/65536.0,1,-nbitq), 
to_sfixed(-1553.0/65536.0,1,-nbitq), 
to_sfixed(1559.0/65536.0,1,-nbitq), 
to_sfixed(-1309.0/65536.0,1,-nbitq), 
to_sfixed(-7764.0/65536.0,1,-nbitq), 
to_sfixed(-6862.0/65536.0,1,-nbitq), 
to_sfixed(2684.0/65536.0,1,-nbitq), 
to_sfixed(719.0/65536.0,1,-nbitq), 
to_sfixed(10167.0/65536.0,1,-nbitq), 
to_sfixed(6033.0/65536.0,1,-nbitq), 
to_sfixed(-8270.0/65536.0,1,-nbitq), 
to_sfixed(-9634.0/65536.0,1,-nbitq), 
to_sfixed(-10815.0/65536.0,1,-nbitq), 
to_sfixed(384.0/65536.0,1,-nbitq), 
to_sfixed(-1846.0/65536.0,1,-nbitq), 
to_sfixed(15550.0/65536.0,1,-nbitq), 
to_sfixed(4600.0/65536.0,1,-nbitq), 
to_sfixed(-2439.0/65536.0,1,-nbitq), 
to_sfixed(950.0/65536.0,1,-nbitq), 
to_sfixed(-1245.0/65536.0,1,-nbitq), 
to_sfixed(-10800.0/65536.0,1,-nbitq), 
to_sfixed(359.0/65536.0,1,-nbitq), 
to_sfixed(-417.0/65536.0,1,-nbitq), 
to_sfixed(-3866.0/65536.0,1,-nbitq), 
to_sfixed(-4472.0/65536.0,1,-nbitq), 
to_sfixed(-5831.0/65536.0,1,-nbitq), 
to_sfixed(-886.0/65536.0,1,-nbitq), 
to_sfixed(5100.0/65536.0,1,-nbitq), 
to_sfixed(-2276.0/65536.0,1,-nbitq), 
to_sfixed(815.0/65536.0,1,-nbitq), 
to_sfixed(4145.0/65536.0,1,-nbitq), 
to_sfixed(-2113.0/65536.0,1,-nbitq), 
to_sfixed(-4390.0/65536.0,1,-nbitq), 
to_sfixed(1274.0/65536.0,1,-nbitq), 
to_sfixed(10539.0/65536.0,1,-nbitq), 
to_sfixed(-652.0/65536.0,1,-nbitq), 
to_sfixed(-821.0/65536.0,1,-nbitq), 
to_sfixed(-1718.0/65536.0,1,-nbitq), 
to_sfixed(3439.0/65536.0,1,-nbitq), 
to_sfixed(-4625.0/65536.0,1,-nbitq), 
to_sfixed(-2432.0/65536.0,1,-nbitq), 
to_sfixed(1476.0/65536.0,1,-nbitq), 
to_sfixed(-9607.0/65536.0,1,-nbitq), 
to_sfixed(-1650.0/65536.0,1,-nbitq), 
to_sfixed(-6553.0/65536.0,1,-nbitq), 
to_sfixed(168.0/65536.0,1,-nbitq), 
to_sfixed(-5054.0/65536.0,1,-nbitq), 
to_sfixed(4007.0/65536.0,1,-nbitq), 
to_sfixed(-3104.0/65536.0,1,-nbitq), 
to_sfixed(94.0/65536.0,1,-nbitq), 
to_sfixed(2484.0/65536.0,1,-nbitq), 
to_sfixed(-2164.0/65536.0,1,-nbitq), 
to_sfixed(-8457.0/65536.0,1,-nbitq), 
to_sfixed(-1029.0/65536.0,1,-nbitq), 
to_sfixed(-9723.0/65536.0,1,-nbitq), 
to_sfixed(8037.0/65536.0,1,-nbitq), 
to_sfixed(5196.0/65536.0,1,-nbitq), 
to_sfixed(905.0/65536.0,1,-nbitq), 
to_sfixed(2888.0/65536.0,1,-nbitq), 
to_sfixed(859.0/65536.0,1,-nbitq), 
to_sfixed(-2214.0/65536.0,1,-nbitq), 
to_sfixed(-747.0/65536.0,1,-nbitq), 
to_sfixed(-553.0/65536.0,1,-nbitq), 
to_sfixed(-10638.0/65536.0,1,-nbitq), 
to_sfixed(201.0/65536.0,1,-nbitq), 
to_sfixed(-1372.0/65536.0,1,-nbitq), 
to_sfixed(-3406.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2077.0/65536.0,1,-nbitq), 
to_sfixed(-3166.0/65536.0,1,-nbitq), 
to_sfixed(5908.0/65536.0,1,-nbitq), 
to_sfixed(-67.0/65536.0,1,-nbitq), 
to_sfixed(-3528.0/65536.0,1,-nbitq), 
to_sfixed(-315.0/65536.0,1,-nbitq), 
to_sfixed(4159.0/65536.0,1,-nbitq), 
to_sfixed(-836.0/65536.0,1,-nbitq), 
to_sfixed(900.0/65536.0,1,-nbitq), 
to_sfixed(-521.0/65536.0,1,-nbitq), 
to_sfixed(1961.0/65536.0,1,-nbitq), 
to_sfixed(-1677.0/65536.0,1,-nbitq), 
to_sfixed(121.0/65536.0,1,-nbitq), 
to_sfixed(-8221.0/65536.0,1,-nbitq), 
to_sfixed(164.0/65536.0,1,-nbitq), 
to_sfixed(3377.0/65536.0,1,-nbitq), 
to_sfixed(707.0/65536.0,1,-nbitq), 
to_sfixed(-6915.0/65536.0,1,-nbitq), 
to_sfixed(-5998.0/65536.0,1,-nbitq), 
to_sfixed(219.0/65536.0,1,-nbitq), 
to_sfixed(840.0/65536.0,1,-nbitq), 
to_sfixed(10669.0/65536.0,1,-nbitq), 
to_sfixed(3017.0/65536.0,1,-nbitq), 
to_sfixed(-10446.0/65536.0,1,-nbitq), 
to_sfixed(-4220.0/65536.0,1,-nbitq), 
to_sfixed(-8129.0/65536.0,1,-nbitq), 
to_sfixed(-2511.0/65536.0,1,-nbitq), 
to_sfixed(1661.0/65536.0,1,-nbitq), 
to_sfixed(14155.0/65536.0,1,-nbitq), 
to_sfixed(1237.0/65536.0,1,-nbitq), 
to_sfixed(1525.0/65536.0,1,-nbitq), 
to_sfixed(3697.0/65536.0,1,-nbitq), 
to_sfixed(1993.0/65536.0,1,-nbitq), 
to_sfixed(-4449.0/65536.0,1,-nbitq), 
to_sfixed(2986.0/65536.0,1,-nbitq), 
to_sfixed(842.0/65536.0,1,-nbitq), 
to_sfixed(-4192.0/65536.0,1,-nbitq), 
to_sfixed(-6610.0/65536.0,1,-nbitq), 
to_sfixed(-1218.0/65536.0,1,-nbitq), 
to_sfixed(-47.0/65536.0,1,-nbitq), 
to_sfixed(2853.0/65536.0,1,-nbitq), 
to_sfixed(114.0/65536.0,1,-nbitq), 
to_sfixed(-2446.0/65536.0,1,-nbitq), 
to_sfixed(3196.0/65536.0,1,-nbitq), 
to_sfixed(-2506.0/65536.0,1,-nbitq), 
to_sfixed(-2903.0/65536.0,1,-nbitq), 
to_sfixed(2303.0/65536.0,1,-nbitq), 
to_sfixed(8468.0/65536.0,1,-nbitq), 
to_sfixed(-1647.0/65536.0,1,-nbitq), 
to_sfixed(-605.0/65536.0,1,-nbitq), 
to_sfixed(2689.0/65536.0,1,-nbitq), 
to_sfixed(5342.0/65536.0,1,-nbitq), 
to_sfixed(-3745.0/65536.0,1,-nbitq), 
to_sfixed(3767.0/65536.0,1,-nbitq), 
to_sfixed(-1172.0/65536.0,1,-nbitq), 
to_sfixed(-4958.0/65536.0,1,-nbitq), 
to_sfixed(-2409.0/65536.0,1,-nbitq), 
to_sfixed(-3820.0/65536.0,1,-nbitq), 
to_sfixed(1300.0/65536.0,1,-nbitq), 
to_sfixed(-6588.0/65536.0,1,-nbitq), 
to_sfixed(3265.0/65536.0,1,-nbitq), 
to_sfixed(2525.0/65536.0,1,-nbitq), 
to_sfixed(-2804.0/65536.0,1,-nbitq), 
to_sfixed(1749.0/65536.0,1,-nbitq), 
to_sfixed(1957.0/65536.0,1,-nbitq), 
to_sfixed(-7615.0/65536.0,1,-nbitq), 
to_sfixed(1699.0/65536.0,1,-nbitq), 
to_sfixed(-6956.0/65536.0,1,-nbitq), 
to_sfixed(8030.0/65536.0,1,-nbitq), 
to_sfixed(12739.0/65536.0,1,-nbitq), 
to_sfixed(1969.0/65536.0,1,-nbitq), 
to_sfixed(9341.0/65536.0,1,-nbitq), 
to_sfixed(3234.0/65536.0,1,-nbitq), 
to_sfixed(1167.0/65536.0,1,-nbitq), 
to_sfixed(2612.0/65536.0,1,-nbitq), 
to_sfixed(-1989.0/65536.0,1,-nbitq), 
to_sfixed(-11703.0/65536.0,1,-nbitq), 
to_sfixed(-233.0/65536.0,1,-nbitq), 
to_sfixed(-497.0/65536.0,1,-nbitq), 
to_sfixed(-3287.0/65536.0,1,-nbitq)  ), 
( to_sfixed(812.0/65536.0,1,-nbitq), 
to_sfixed(-2046.0/65536.0,1,-nbitq), 
to_sfixed(7578.0/65536.0,1,-nbitq), 
to_sfixed(1758.0/65536.0,1,-nbitq), 
to_sfixed(-3460.0/65536.0,1,-nbitq), 
to_sfixed(-3879.0/65536.0,1,-nbitq), 
to_sfixed(889.0/65536.0,1,-nbitq), 
to_sfixed(1239.0/65536.0,1,-nbitq), 
to_sfixed(-1974.0/65536.0,1,-nbitq), 
to_sfixed(2338.0/65536.0,1,-nbitq), 
to_sfixed(781.0/65536.0,1,-nbitq), 
to_sfixed(-2678.0/65536.0,1,-nbitq), 
to_sfixed(1546.0/65536.0,1,-nbitq), 
to_sfixed(-12779.0/65536.0,1,-nbitq), 
to_sfixed(1642.0/65536.0,1,-nbitq), 
to_sfixed(313.0/65536.0,1,-nbitq), 
to_sfixed(-2649.0/65536.0,1,-nbitq), 
to_sfixed(-5003.0/65536.0,1,-nbitq), 
to_sfixed(-7250.0/65536.0,1,-nbitq), 
to_sfixed(3054.0/65536.0,1,-nbitq), 
to_sfixed(4003.0/65536.0,1,-nbitq), 
to_sfixed(4062.0/65536.0,1,-nbitq), 
to_sfixed(2885.0/65536.0,1,-nbitq), 
to_sfixed(-5967.0/65536.0,1,-nbitq), 
to_sfixed(-3788.0/65536.0,1,-nbitq), 
to_sfixed(-6875.0/65536.0,1,-nbitq), 
to_sfixed(-1061.0/65536.0,1,-nbitq), 
to_sfixed(984.0/65536.0,1,-nbitq), 
to_sfixed(8996.0/65536.0,1,-nbitq), 
to_sfixed(-2847.0/65536.0,1,-nbitq), 
to_sfixed(-4433.0/65536.0,1,-nbitq), 
to_sfixed(1207.0/65536.0,1,-nbitq), 
to_sfixed(1865.0/65536.0,1,-nbitq), 
to_sfixed(3452.0/65536.0,1,-nbitq), 
to_sfixed(-1801.0/65536.0,1,-nbitq), 
to_sfixed(-1420.0/65536.0,1,-nbitq), 
to_sfixed(834.0/65536.0,1,-nbitq), 
to_sfixed(-3499.0/65536.0,1,-nbitq), 
to_sfixed(3697.0/65536.0,1,-nbitq), 
to_sfixed(2187.0/65536.0,1,-nbitq), 
to_sfixed(3021.0/65536.0,1,-nbitq), 
to_sfixed(-2112.0/65536.0,1,-nbitq), 
to_sfixed(70.0/65536.0,1,-nbitq), 
to_sfixed(-2101.0/65536.0,1,-nbitq), 
to_sfixed(-486.0/65536.0,1,-nbitq), 
to_sfixed(2608.0/65536.0,1,-nbitq), 
to_sfixed(2410.0/65536.0,1,-nbitq), 
to_sfixed(6555.0/65536.0,1,-nbitq), 
to_sfixed(1248.0/65536.0,1,-nbitq), 
to_sfixed(-1649.0/65536.0,1,-nbitq), 
to_sfixed(1005.0/65536.0,1,-nbitq), 
to_sfixed(-1948.0/65536.0,1,-nbitq), 
to_sfixed(-3577.0/65536.0,1,-nbitq), 
to_sfixed(11830.0/65536.0,1,-nbitq), 
to_sfixed(2885.0/65536.0,1,-nbitq), 
to_sfixed(-5674.0/65536.0,1,-nbitq), 
to_sfixed(378.0/65536.0,1,-nbitq), 
to_sfixed(4806.0/65536.0,1,-nbitq), 
to_sfixed(-2543.0/65536.0,1,-nbitq), 
to_sfixed(-3804.0/65536.0,1,-nbitq), 
to_sfixed(3897.0/65536.0,1,-nbitq), 
to_sfixed(-1205.0/65536.0,1,-nbitq), 
to_sfixed(2273.0/65536.0,1,-nbitq), 
to_sfixed(-2910.0/65536.0,1,-nbitq), 
to_sfixed(1153.0/65536.0,1,-nbitq), 
to_sfixed(-5093.0/65536.0,1,-nbitq), 
to_sfixed(5834.0/65536.0,1,-nbitq), 
to_sfixed(3090.0/65536.0,1,-nbitq), 
to_sfixed(4646.0/65536.0,1,-nbitq), 
to_sfixed(9056.0/65536.0,1,-nbitq), 
to_sfixed(-2369.0/65536.0,1,-nbitq), 
to_sfixed(3264.0/65536.0,1,-nbitq), 
to_sfixed(2819.0/65536.0,1,-nbitq), 
to_sfixed(-316.0/65536.0,1,-nbitq), 
to_sfixed(1618.0/65536.0,1,-nbitq), 
to_sfixed(4204.0/65536.0,1,-nbitq), 
to_sfixed(-7667.0/65536.0,1,-nbitq), 
to_sfixed(6091.0/65536.0,1,-nbitq), 
to_sfixed(-2018.0/65536.0,1,-nbitq), 
to_sfixed(-5231.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2766.0/65536.0,1,-nbitq), 
to_sfixed(-1798.0/65536.0,1,-nbitq), 
to_sfixed(5286.0/65536.0,1,-nbitq), 
to_sfixed(5396.0/65536.0,1,-nbitq), 
to_sfixed(-2351.0/65536.0,1,-nbitq), 
to_sfixed(-2066.0/65536.0,1,-nbitq), 
to_sfixed(2940.0/65536.0,1,-nbitq), 
to_sfixed(2034.0/65536.0,1,-nbitq), 
to_sfixed(2427.0/65536.0,1,-nbitq), 
to_sfixed(1562.0/65536.0,1,-nbitq), 
to_sfixed(646.0/65536.0,1,-nbitq), 
to_sfixed(-7105.0/65536.0,1,-nbitq), 
to_sfixed(-866.0/65536.0,1,-nbitq), 
to_sfixed(-9161.0/65536.0,1,-nbitq), 
to_sfixed(168.0/65536.0,1,-nbitq), 
to_sfixed(-681.0/65536.0,1,-nbitq), 
to_sfixed(-1001.0/65536.0,1,-nbitq), 
to_sfixed(-40.0/65536.0,1,-nbitq), 
to_sfixed(-1744.0/65536.0,1,-nbitq), 
to_sfixed(1214.0/65536.0,1,-nbitq), 
to_sfixed(1338.0/65536.0,1,-nbitq), 
to_sfixed(-2784.0/65536.0,1,-nbitq), 
to_sfixed(-463.0/65536.0,1,-nbitq), 
to_sfixed(-9187.0/65536.0,1,-nbitq), 
to_sfixed(-4306.0/65536.0,1,-nbitq), 
to_sfixed(-4104.0/65536.0,1,-nbitq), 
to_sfixed(-2444.0/65536.0,1,-nbitq), 
to_sfixed(-135.0/65536.0,1,-nbitq), 
to_sfixed(7832.0/65536.0,1,-nbitq), 
to_sfixed(285.0/65536.0,1,-nbitq), 
to_sfixed(-2326.0/65536.0,1,-nbitq), 
to_sfixed(-5333.0/65536.0,1,-nbitq), 
to_sfixed(11.0/65536.0,1,-nbitq), 
to_sfixed(-368.0/65536.0,1,-nbitq), 
to_sfixed(-1438.0/65536.0,1,-nbitq), 
to_sfixed(-851.0/65536.0,1,-nbitq), 
to_sfixed(-1325.0/65536.0,1,-nbitq), 
to_sfixed(815.0/65536.0,1,-nbitq), 
to_sfixed(630.0/65536.0,1,-nbitq), 
to_sfixed(2756.0/65536.0,1,-nbitq), 
to_sfixed(2399.0/65536.0,1,-nbitq), 
to_sfixed(1737.0/65536.0,1,-nbitq), 
to_sfixed(-78.0/65536.0,1,-nbitq), 
to_sfixed(-1812.0/65536.0,1,-nbitq), 
to_sfixed(386.0/65536.0,1,-nbitq), 
to_sfixed(117.0/65536.0,1,-nbitq), 
to_sfixed(2509.0/65536.0,1,-nbitq), 
to_sfixed(1886.0/65536.0,1,-nbitq), 
to_sfixed(2035.0/65536.0,1,-nbitq), 
to_sfixed(2737.0/65536.0,1,-nbitq), 
to_sfixed(1315.0/65536.0,1,-nbitq), 
to_sfixed(458.0/65536.0,1,-nbitq), 
to_sfixed(-3801.0/65536.0,1,-nbitq), 
to_sfixed(8709.0/65536.0,1,-nbitq), 
to_sfixed(-3836.0/65536.0,1,-nbitq), 
to_sfixed(-7208.0/65536.0,1,-nbitq), 
to_sfixed(2573.0/65536.0,1,-nbitq), 
to_sfixed(2877.0/65536.0,1,-nbitq), 
to_sfixed(-1581.0/65536.0,1,-nbitq), 
to_sfixed(-4249.0/65536.0,1,-nbitq), 
to_sfixed(4125.0/65536.0,1,-nbitq), 
to_sfixed(1800.0/65536.0,1,-nbitq), 
to_sfixed(1755.0/65536.0,1,-nbitq), 
to_sfixed(1795.0/65536.0,1,-nbitq), 
to_sfixed(2658.0/65536.0,1,-nbitq), 
to_sfixed(484.0/65536.0,1,-nbitq), 
to_sfixed(1020.0/65536.0,1,-nbitq), 
to_sfixed(3503.0/65536.0,1,-nbitq), 
to_sfixed(3505.0/65536.0,1,-nbitq), 
to_sfixed(5431.0/65536.0,1,-nbitq), 
to_sfixed(-2821.0/65536.0,1,-nbitq), 
to_sfixed(1981.0/65536.0,1,-nbitq), 
to_sfixed(3823.0/65536.0,1,-nbitq), 
to_sfixed(1965.0/65536.0,1,-nbitq), 
to_sfixed(-1494.0/65536.0,1,-nbitq), 
to_sfixed(-2388.0/65536.0,1,-nbitq), 
to_sfixed(-7629.0/65536.0,1,-nbitq), 
to_sfixed(2242.0/65536.0,1,-nbitq), 
to_sfixed(-3226.0/65536.0,1,-nbitq), 
to_sfixed(-3557.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3018.0/65536.0,1,-nbitq), 
to_sfixed(-270.0/65536.0,1,-nbitq), 
to_sfixed(2848.0/65536.0,1,-nbitq), 
to_sfixed(2218.0/65536.0,1,-nbitq), 
to_sfixed(-1225.0/65536.0,1,-nbitq), 
to_sfixed(4009.0/65536.0,1,-nbitq), 
to_sfixed(1671.0/65536.0,1,-nbitq), 
to_sfixed(2480.0/65536.0,1,-nbitq), 
to_sfixed(188.0/65536.0,1,-nbitq), 
to_sfixed(2727.0/65536.0,1,-nbitq), 
to_sfixed(232.0/65536.0,1,-nbitq), 
to_sfixed(-7614.0/65536.0,1,-nbitq), 
to_sfixed(105.0/65536.0,1,-nbitq), 
to_sfixed(-8233.0/65536.0,1,-nbitq), 
to_sfixed(-506.0/65536.0,1,-nbitq), 
to_sfixed(-963.0/65536.0,1,-nbitq), 
to_sfixed(-1559.0/65536.0,1,-nbitq), 
to_sfixed(-1985.0/65536.0,1,-nbitq), 
to_sfixed(-3479.0/65536.0,1,-nbitq), 
to_sfixed(1580.0/65536.0,1,-nbitq), 
to_sfixed(2410.0/65536.0,1,-nbitq), 
to_sfixed(2220.0/65536.0,1,-nbitq), 
to_sfixed(-3378.0/65536.0,1,-nbitq), 
to_sfixed(-6348.0/65536.0,1,-nbitq), 
to_sfixed(-2509.0/65536.0,1,-nbitq), 
to_sfixed(1686.0/65536.0,1,-nbitq), 
to_sfixed(1316.0/65536.0,1,-nbitq), 
to_sfixed(-3931.0/65536.0,1,-nbitq), 
to_sfixed(7545.0/65536.0,1,-nbitq), 
to_sfixed(678.0/65536.0,1,-nbitq), 
to_sfixed(-2801.0/65536.0,1,-nbitq), 
to_sfixed(-1554.0/65536.0,1,-nbitq), 
to_sfixed(5121.0/65536.0,1,-nbitq), 
to_sfixed(-1188.0/65536.0,1,-nbitq), 
to_sfixed(-532.0/65536.0,1,-nbitq), 
to_sfixed(2394.0/65536.0,1,-nbitq), 
to_sfixed(3081.0/65536.0,1,-nbitq), 
to_sfixed(-3463.0/65536.0,1,-nbitq), 
to_sfixed(-1526.0/65536.0,1,-nbitq), 
to_sfixed(-201.0/65536.0,1,-nbitq), 
to_sfixed(-2129.0/65536.0,1,-nbitq), 
to_sfixed(1314.0/65536.0,1,-nbitq), 
to_sfixed(3267.0/65536.0,1,-nbitq), 
to_sfixed(-2639.0/65536.0,1,-nbitq), 
to_sfixed(1432.0/65536.0,1,-nbitq), 
to_sfixed(674.0/65536.0,1,-nbitq), 
to_sfixed(-2328.0/65536.0,1,-nbitq), 
to_sfixed(5150.0/65536.0,1,-nbitq), 
to_sfixed(-2635.0/65536.0,1,-nbitq), 
to_sfixed(2153.0/65536.0,1,-nbitq), 
to_sfixed(3173.0/65536.0,1,-nbitq), 
to_sfixed(-281.0/65536.0,1,-nbitq), 
to_sfixed(-757.0/65536.0,1,-nbitq), 
to_sfixed(11972.0/65536.0,1,-nbitq), 
to_sfixed(-1410.0/65536.0,1,-nbitq), 
to_sfixed(-1524.0/65536.0,1,-nbitq), 
to_sfixed(1073.0/65536.0,1,-nbitq), 
to_sfixed(4235.0/65536.0,1,-nbitq), 
to_sfixed(-1003.0/65536.0,1,-nbitq), 
to_sfixed(-1325.0/65536.0,1,-nbitq), 
to_sfixed(5426.0/65536.0,1,-nbitq), 
to_sfixed(1715.0/65536.0,1,-nbitq), 
to_sfixed(90.0/65536.0,1,-nbitq), 
to_sfixed(257.0/65536.0,1,-nbitq), 
to_sfixed(4741.0/65536.0,1,-nbitq), 
to_sfixed(5424.0/65536.0,1,-nbitq), 
to_sfixed(1440.0/65536.0,1,-nbitq), 
to_sfixed(1506.0/65536.0,1,-nbitq), 
to_sfixed(2580.0/65536.0,1,-nbitq), 
to_sfixed(9145.0/65536.0,1,-nbitq), 
to_sfixed(759.0/65536.0,1,-nbitq), 
to_sfixed(1016.0/65536.0,1,-nbitq), 
to_sfixed(8338.0/65536.0,1,-nbitq), 
to_sfixed(2620.0/65536.0,1,-nbitq), 
to_sfixed(-640.0/65536.0,1,-nbitq), 
to_sfixed(2305.0/65536.0,1,-nbitq), 
to_sfixed(-4956.0/65536.0,1,-nbitq), 
to_sfixed(4135.0/65536.0,1,-nbitq), 
to_sfixed(-2850.0/65536.0,1,-nbitq), 
to_sfixed(-1198.0/65536.0,1,-nbitq)  ), 
( to_sfixed(550.0/65536.0,1,-nbitq), 
to_sfixed(-2603.0/65536.0,1,-nbitq), 
to_sfixed(-1456.0/65536.0,1,-nbitq), 
to_sfixed(6159.0/65536.0,1,-nbitq), 
to_sfixed(1251.0/65536.0,1,-nbitq), 
to_sfixed(1551.0/65536.0,1,-nbitq), 
to_sfixed(2984.0/65536.0,1,-nbitq), 
to_sfixed(4694.0/65536.0,1,-nbitq), 
to_sfixed(-4906.0/65536.0,1,-nbitq), 
to_sfixed(341.0/65536.0,1,-nbitq), 
to_sfixed(-141.0/65536.0,1,-nbitq), 
to_sfixed(-4169.0/65536.0,1,-nbitq), 
to_sfixed(2558.0/65536.0,1,-nbitq), 
to_sfixed(-4466.0/65536.0,1,-nbitq), 
to_sfixed(-3707.0/65536.0,1,-nbitq), 
to_sfixed(2719.0/65536.0,1,-nbitq), 
to_sfixed(478.0/65536.0,1,-nbitq), 
to_sfixed(-3636.0/65536.0,1,-nbitq), 
to_sfixed(-1120.0/65536.0,1,-nbitq), 
to_sfixed(1601.0/65536.0,1,-nbitq), 
to_sfixed(6051.0/65536.0,1,-nbitq), 
to_sfixed(1729.0/65536.0,1,-nbitq), 
to_sfixed(-4398.0/65536.0,1,-nbitq), 
to_sfixed(-5138.0/65536.0,1,-nbitq), 
to_sfixed(-4413.0/65536.0,1,-nbitq), 
to_sfixed(-1692.0/65536.0,1,-nbitq), 
to_sfixed(-2527.0/65536.0,1,-nbitq), 
to_sfixed(-3692.0/65536.0,1,-nbitq), 
to_sfixed(4861.0/65536.0,1,-nbitq), 
to_sfixed(-161.0/65536.0,1,-nbitq), 
to_sfixed(-3152.0/65536.0,1,-nbitq), 
to_sfixed(-2774.0/65536.0,1,-nbitq), 
to_sfixed(5203.0/65536.0,1,-nbitq), 
to_sfixed(765.0/65536.0,1,-nbitq), 
to_sfixed(32.0/65536.0,1,-nbitq), 
to_sfixed(-1073.0/65536.0,1,-nbitq), 
to_sfixed(-1962.0/65536.0,1,-nbitq), 
to_sfixed(-4871.0/65536.0,1,-nbitq), 
to_sfixed(-3354.0/65536.0,1,-nbitq), 
to_sfixed(2839.0/65536.0,1,-nbitq), 
to_sfixed(-1678.0/65536.0,1,-nbitq), 
to_sfixed(-2747.0/65536.0,1,-nbitq), 
to_sfixed(769.0/65536.0,1,-nbitq), 
to_sfixed(-5339.0/65536.0,1,-nbitq), 
to_sfixed(-1667.0/65536.0,1,-nbitq), 
to_sfixed(4877.0/65536.0,1,-nbitq), 
to_sfixed(-331.0/65536.0,1,-nbitq), 
to_sfixed(4070.0/65536.0,1,-nbitq), 
to_sfixed(3116.0/65536.0,1,-nbitq), 
to_sfixed(-538.0/65536.0,1,-nbitq), 
to_sfixed(-2609.0/65536.0,1,-nbitq), 
to_sfixed(-2935.0/65536.0,1,-nbitq), 
to_sfixed(-50.0/65536.0,1,-nbitq), 
to_sfixed(8070.0/65536.0,1,-nbitq), 
to_sfixed(-2577.0/65536.0,1,-nbitq), 
to_sfixed(-2931.0/65536.0,1,-nbitq), 
to_sfixed(-1726.0/65536.0,1,-nbitq), 
to_sfixed(3164.0/65536.0,1,-nbitq), 
to_sfixed(1030.0/65536.0,1,-nbitq), 
to_sfixed(-3315.0/65536.0,1,-nbitq), 
to_sfixed(1307.0/65536.0,1,-nbitq), 
to_sfixed(-1772.0/65536.0,1,-nbitq), 
to_sfixed(2347.0/65536.0,1,-nbitq), 
to_sfixed(2371.0/65536.0,1,-nbitq), 
to_sfixed(-71.0/65536.0,1,-nbitq), 
to_sfixed(1326.0/65536.0,1,-nbitq), 
to_sfixed(5042.0/65536.0,1,-nbitq), 
to_sfixed(1730.0/65536.0,1,-nbitq), 
to_sfixed(5615.0/65536.0,1,-nbitq), 
to_sfixed(9432.0/65536.0,1,-nbitq), 
to_sfixed(-2076.0/65536.0,1,-nbitq), 
to_sfixed(-3965.0/65536.0,1,-nbitq), 
to_sfixed(8136.0/65536.0,1,-nbitq), 
to_sfixed(-1774.0/65536.0,1,-nbitq), 
to_sfixed(-2532.0/65536.0,1,-nbitq), 
to_sfixed(895.0/65536.0,1,-nbitq), 
to_sfixed(-6682.0/65536.0,1,-nbitq), 
to_sfixed(2019.0/65536.0,1,-nbitq), 
to_sfixed(-1262.0/65536.0,1,-nbitq), 
to_sfixed(750.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-407.0/65536.0,1,-nbitq), 
to_sfixed(2514.0/65536.0,1,-nbitq), 
to_sfixed(-2546.0/65536.0,1,-nbitq), 
to_sfixed(4587.0/65536.0,1,-nbitq), 
to_sfixed(-2214.0/65536.0,1,-nbitq), 
to_sfixed(-2046.0/65536.0,1,-nbitq), 
to_sfixed(1219.0/65536.0,1,-nbitq), 
to_sfixed(4271.0/65536.0,1,-nbitq), 
to_sfixed(-386.0/65536.0,1,-nbitq), 
to_sfixed(1715.0/65536.0,1,-nbitq), 
to_sfixed(2882.0/65536.0,1,-nbitq), 
to_sfixed(-1750.0/65536.0,1,-nbitq), 
to_sfixed(1710.0/65536.0,1,-nbitq), 
to_sfixed(-3788.0/65536.0,1,-nbitq), 
to_sfixed(2038.0/65536.0,1,-nbitq), 
to_sfixed(2881.0/65536.0,1,-nbitq), 
to_sfixed(-1773.0/65536.0,1,-nbitq), 
to_sfixed(1526.0/65536.0,1,-nbitq), 
to_sfixed(3132.0/65536.0,1,-nbitq), 
to_sfixed(1148.0/65536.0,1,-nbitq), 
to_sfixed(-1455.0/65536.0,1,-nbitq), 
to_sfixed(7617.0/65536.0,1,-nbitq), 
to_sfixed(-4835.0/65536.0,1,-nbitq), 
to_sfixed(-288.0/65536.0,1,-nbitq), 
to_sfixed(-1106.0/65536.0,1,-nbitq), 
to_sfixed(2577.0/65536.0,1,-nbitq), 
to_sfixed(1094.0/65536.0,1,-nbitq), 
to_sfixed(-1246.0/65536.0,1,-nbitq), 
to_sfixed(951.0/65536.0,1,-nbitq), 
to_sfixed(-997.0/65536.0,1,-nbitq), 
to_sfixed(-511.0/65536.0,1,-nbitq), 
to_sfixed(-1436.0/65536.0,1,-nbitq), 
to_sfixed(1947.0/65536.0,1,-nbitq), 
to_sfixed(-363.0/65536.0,1,-nbitq), 
to_sfixed(-1166.0/65536.0,1,-nbitq), 
to_sfixed(-2544.0/65536.0,1,-nbitq), 
to_sfixed(-5885.0/65536.0,1,-nbitq), 
to_sfixed(1737.0/65536.0,1,-nbitq), 
to_sfixed(-3747.0/65536.0,1,-nbitq), 
to_sfixed(-2327.0/65536.0,1,-nbitq), 
to_sfixed(3072.0/65536.0,1,-nbitq), 
to_sfixed(-1175.0/65536.0,1,-nbitq), 
to_sfixed(650.0/65536.0,1,-nbitq), 
to_sfixed(-260.0/65536.0,1,-nbitq), 
to_sfixed(-2490.0/65536.0,1,-nbitq), 
to_sfixed(5243.0/65536.0,1,-nbitq), 
to_sfixed(1719.0/65536.0,1,-nbitq), 
to_sfixed(3892.0/65536.0,1,-nbitq), 
to_sfixed(2832.0/65536.0,1,-nbitq), 
to_sfixed(3919.0/65536.0,1,-nbitq), 
to_sfixed(2355.0/65536.0,1,-nbitq), 
to_sfixed(1968.0/65536.0,1,-nbitq), 
to_sfixed(-4070.0/65536.0,1,-nbitq), 
to_sfixed(7322.0/65536.0,1,-nbitq), 
to_sfixed(-4103.0/65536.0,1,-nbitq), 
to_sfixed(-13.0/65536.0,1,-nbitq), 
to_sfixed(-500.0/65536.0,1,-nbitq), 
to_sfixed(2824.0/65536.0,1,-nbitq), 
to_sfixed(2864.0/65536.0,1,-nbitq), 
to_sfixed(-3474.0/65536.0,1,-nbitq), 
to_sfixed(-2134.0/65536.0,1,-nbitq), 
to_sfixed(-2997.0/65536.0,1,-nbitq), 
to_sfixed(268.0/65536.0,1,-nbitq), 
to_sfixed(344.0/65536.0,1,-nbitq), 
to_sfixed(-1725.0/65536.0,1,-nbitq), 
to_sfixed(-2600.0/65536.0,1,-nbitq), 
to_sfixed(5715.0/65536.0,1,-nbitq), 
to_sfixed(1557.0/65536.0,1,-nbitq), 
to_sfixed(4965.0/65536.0,1,-nbitq), 
to_sfixed(971.0/65536.0,1,-nbitq), 
to_sfixed(-3713.0/65536.0,1,-nbitq), 
to_sfixed(-706.0/65536.0,1,-nbitq), 
to_sfixed(1346.0/65536.0,1,-nbitq), 
to_sfixed(2216.0/65536.0,1,-nbitq), 
to_sfixed(2414.0/65536.0,1,-nbitq), 
to_sfixed(-1644.0/65536.0,1,-nbitq), 
to_sfixed(-2779.0/65536.0,1,-nbitq), 
to_sfixed(1749.0/65536.0,1,-nbitq), 
to_sfixed(-2302.0/65536.0,1,-nbitq), 
to_sfixed(3099.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2243.0/65536.0,1,-nbitq), 
to_sfixed(10.0/65536.0,1,-nbitq), 
to_sfixed(1365.0/65536.0,1,-nbitq), 
to_sfixed(2806.0/65536.0,1,-nbitq), 
to_sfixed(689.0/65536.0,1,-nbitq), 
to_sfixed(-2564.0/65536.0,1,-nbitq), 
to_sfixed(2093.0/65536.0,1,-nbitq), 
to_sfixed(2323.0/65536.0,1,-nbitq), 
to_sfixed(-156.0/65536.0,1,-nbitq), 
to_sfixed(772.0/65536.0,1,-nbitq), 
to_sfixed(-3618.0/65536.0,1,-nbitq), 
to_sfixed(-777.0/65536.0,1,-nbitq), 
to_sfixed(2344.0/65536.0,1,-nbitq), 
to_sfixed(1206.0/65536.0,1,-nbitq), 
to_sfixed(-291.0/65536.0,1,-nbitq), 
to_sfixed(-893.0/65536.0,1,-nbitq), 
to_sfixed(-2463.0/65536.0,1,-nbitq), 
to_sfixed(3736.0/65536.0,1,-nbitq), 
to_sfixed(164.0/65536.0,1,-nbitq), 
to_sfixed(-2371.0/65536.0,1,-nbitq), 
to_sfixed(441.0/65536.0,1,-nbitq), 
to_sfixed(2325.0/65536.0,1,-nbitq), 
to_sfixed(-1056.0/65536.0,1,-nbitq), 
to_sfixed(978.0/65536.0,1,-nbitq), 
to_sfixed(2428.0/65536.0,1,-nbitq), 
to_sfixed(3421.0/65536.0,1,-nbitq), 
to_sfixed(-2066.0/65536.0,1,-nbitq), 
to_sfixed(-1835.0/65536.0,1,-nbitq), 
to_sfixed(-1698.0/65536.0,1,-nbitq), 
to_sfixed(-1443.0/65536.0,1,-nbitq), 
to_sfixed(1799.0/65536.0,1,-nbitq), 
to_sfixed(349.0/65536.0,1,-nbitq), 
to_sfixed(-3050.0/65536.0,1,-nbitq), 
to_sfixed(-4137.0/65536.0,1,-nbitq), 
to_sfixed(-2098.0/65536.0,1,-nbitq), 
to_sfixed(-1036.0/65536.0,1,-nbitq), 
to_sfixed(-3384.0/65536.0,1,-nbitq), 
to_sfixed(-1300.0/65536.0,1,-nbitq), 
to_sfixed(-3707.0/65536.0,1,-nbitq), 
to_sfixed(-198.0/65536.0,1,-nbitq), 
to_sfixed(-3169.0/65536.0,1,-nbitq), 
to_sfixed(-1739.0/65536.0,1,-nbitq), 
to_sfixed(-1988.0/65536.0,1,-nbitq), 
to_sfixed(694.0/65536.0,1,-nbitq), 
to_sfixed(-2520.0/65536.0,1,-nbitq), 
to_sfixed(1150.0/65536.0,1,-nbitq), 
to_sfixed(1028.0/65536.0,1,-nbitq), 
to_sfixed(728.0/65536.0,1,-nbitq), 
to_sfixed(-1415.0/65536.0,1,-nbitq), 
to_sfixed(753.0/65536.0,1,-nbitq), 
to_sfixed(1153.0/65536.0,1,-nbitq), 
to_sfixed(365.0/65536.0,1,-nbitq), 
to_sfixed(1093.0/65536.0,1,-nbitq), 
to_sfixed(-1143.0/65536.0,1,-nbitq), 
to_sfixed(3179.0/65536.0,1,-nbitq), 
to_sfixed(-2685.0/65536.0,1,-nbitq), 
to_sfixed(1436.0/65536.0,1,-nbitq), 
to_sfixed(3730.0/65536.0,1,-nbitq), 
to_sfixed(-283.0/65536.0,1,-nbitq), 
to_sfixed(902.0/65536.0,1,-nbitq), 
to_sfixed(-788.0/65536.0,1,-nbitq), 
to_sfixed(2501.0/65536.0,1,-nbitq), 
to_sfixed(-1152.0/65536.0,1,-nbitq), 
to_sfixed(2240.0/65536.0,1,-nbitq), 
to_sfixed(-1088.0/65536.0,1,-nbitq), 
to_sfixed(2442.0/65536.0,1,-nbitq), 
to_sfixed(351.0/65536.0,1,-nbitq), 
to_sfixed(-2515.0/65536.0,1,-nbitq), 
to_sfixed(174.0/65536.0,1,-nbitq), 
to_sfixed(3714.0/65536.0,1,-nbitq), 
to_sfixed(-2870.0/65536.0,1,-nbitq), 
to_sfixed(1294.0/65536.0,1,-nbitq), 
to_sfixed(473.0/65536.0,1,-nbitq), 
to_sfixed(800.0/65536.0,1,-nbitq), 
to_sfixed(686.0/65536.0,1,-nbitq), 
to_sfixed(-1466.0/65536.0,1,-nbitq), 
to_sfixed(-2402.0/65536.0,1,-nbitq), 
to_sfixed(1048.0/65536.0,1,-nbitq), 
to_sfixed(-2411.0/65536.0,1,-nbitq), 
to_sfixed(2429.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1449.0/65536.0,1,-nbitq), 
to_sfixed(-2839.0/65536.0,1,-nbitq), 
to_sfixed(-971.0/65536.0,1,-nbitq), 
to_sfixed(-901.0/65536.0,1,-nbitq), 
to_sfixed(-56.0/65536.0,1,-nbitq), 
to_sfixed(515.0/65536.0,1,-nbitq), 
to_sfixed(-1019.0/65536.0,1,-nbitq), 
to_sfixed(1526.0/65536.0,1,-nbitq), 
to_sfixed(-968.0/65536.0,1,-nbitq), 
to_sfixed(-1560.0/65536.0,1,-nbitq), 
to_sfixed(284.0/65536.0,1,-nbitq), 
to_sfixed(-1797.0/65536.0,1,-nbitq), 
to_sfixed(2275.0/65536.0,1,-nbitq), 
to_sfixed(-248.0/65536.0,1,-nbitq), 
to_sfixed(-61.0/65536.0,1,-nbitq), 
to_sfixed(-687.0/65536.0,1,-nbitq), 
to_sfixed(-2193.0/65536.0,1,-nbitq), 
to_sfixed(2228.0/65536.0,1,-nbitq), 
to_sfixed(2506.0/65536.0,1,-nbitq), 
to_sfixed(1128.0/65536.0,1,-nbitq), 
to_sfixed(1429.0/65536.0,1,-nbitq), 
to_sfixed(1919.0/65536.0,1,-nbitq), 
to_sfixed(-1881.0/65536.0,1,-nbitq), 
to_sfixed(2305.0/65536.0,1,-nbitq), 
to_sfixed(1222.0/65536.0,1,-nbitq), 
to_sfixed(3373.0/65536.0,1,-nbitq), 
to_sfixed(-759.0/65536.0,1,-nbitq), 
to_sfixed(2330.0/65536.0,1,-nbitq), 
to_sfixed(692.0/65536.0,1,-nbitq), 
to_sfixed(-2995.0/65536.0,1,-nbitq), 
to_sfixed(2479.0/65536.0,1,-nbitq), 
to_sfixed(-3167.0/65536.0,1,-nbitq), 
to_sfixed(-4510.0/65536.0,1,-nbitq), 
to_sfixed(-2252.0/65536.0,1,-nbitq), 
to_sfixed(-1875.0/65536.0,1,-nbitq), 
to_sfixed(778.0/65536.0,1,-nbitq), 
to_sfixed(-686.0/65536.0,1,-nbitq), 
to_sfixed(521.0/65536.0,1,-nbitq), 
to_sfixed(-2913.0/65536.0,1,-nbitq), 
to_sfixed(-1446.0/65536.0,1,-nbitq), 
to_sfixed(1761.0/65536.0,1,-nbitq), 
to_sfixed(-2415.0/65536.0,1,-nbitq), 
to_sfixed(-3702.0/65536.0,1,-nbitq), 
to_sfixed(1597.0/65536.0,1,-nbitq), 
to_sfixed(1366.0/65536.0,1,-nbitq), 
to_sfixed(2018.0/65536.0,1,-nbitq), 
to_sfixed(278.0/65536.0,1,-nbitq), 
to_sfixed(-1374.0/65536.0,1,-nbitq), 
to_sfixed(925.0/65536.0,1,-nbitq), 
to_sfixed(909.0/65536.0,1,-nbitq), 
to_sfixed(344.0/65536.0,1,-nbitq), 
to_sfixed(-227.0/65536.0,1,-nbitq), 
to_sfixed(2530.0/65536.0,1,-nbitq), 
to_sfixed(2833.0/65536.0,1,-nbitq), 
to_sfixed(3144.0/65536.0,1,-nbitq), 
to_sfixed(-2011.0/65536.0,1,-nbitq), 
to_sfixed(2029.0/65536.0,1,-nbitq), 
to_sfixed(-928.0/65536.0,1,-nbitq), 
to_sfixed(58.0/65536.0,1,-nbitq), 
to_sfixed(-282.0/65536.0,1,-nbitq), 
to_sfixed(-1769.0/65536.0,1,-nbitq), 
to_sfixed(-1356.0/65536.0,1,-nbitq), 
to_sfixed(869.0/65536.0,1,-nbitq), 
to_sfixed(-1258.0/65536.0,1,-nbitq), 
to_sfixed(1252.0/65536.0,1,-nbitq), 
to_sfixed(3356.0/65536.0,1,-nbitq), 
to_sfixed(2740.0/65536.0,1,-nbitq), 
to_sfixed(-598.0/65536.0,1,-nbitq), 
to_sfixed(1331.0/65536.0,1,-nbitq), 
to_sfixed(-869.0/65536.0,1,-nbitq), 
to_sfixed(-2299.0/65536.0,1,-nbitq), 
to_sfixed(-2398.0/65536.0,1,-nbitq), 
to_sfixed(2063.0/65536.0,1,-nbitq), 
to_sfixed(-417.0/65536.0,1,-nbitq), 
to_sfixed(-2892.0/65536.0,1,-nbitq), 
to_sfixed(1412.0/65536.0,1,-nbitq), 
to_sfixed(-1766.0/65536.0,1,-nbitq), 
to_sfixed(-392.0/65536.0,1,-nbitq), 
to_sfixed(687.0/65536.0,1,-nbitq), 
to_sfixed(2392.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-935.0/65536.0,1,-nbitq), 
to_sfixed(1628.0/65536.0,1,-nbitq), 
to_sfixed(179.0/65536.0,1,-nbitq), 
to_sfixed(1065.0/65536.0,1,-nbitq), 
to_sfixed(-904.0/65536.0,1,-nbitq), 
to_sfixed(-1859.0/65536.0,1,-nbitq), 
to_sfixed(214.0/65536.0,1,-nbitq), 
to_sfixed(2851.0/65536.0,1,-nbitq), 
to_sfixed(2802.0/65536.0,1,-nbitq), 
to_sfixed(2923.0/65536.0,1,-nbitq), 
to_sfixed(-858.0/65536.0,1,-nbitq), 
to_sfixed(128.0/65536.0,1,-nbitq), 
to_sfixed(1888.0/65536.0,1,-nbitq), 
to_sfixed(-1387.0/65536.0,1,-nbitq), 
to_sfixed(1947.0/65536.0,1,-nbitq), 
to_sfixed(317.0/65536.0,1,-nbitq), 
to_sfixed(-1764.0/65536.0,1,-nbitq), 
to_sfixed(926.0/65536.0,1,-nbitq), 
to_sfixed(2270.0/65536.0,1,-nbitq), 
to_sfixed(1378.0/65536.0,1,-nbitq), 
to_sfixed(145.0/65536.0,1,-nbitq), 
to_sfixed(1918.0/65536.0,1,-nbitq), 
to_sfixed(447.0/65536.0,1,-nbitq), 
to_sfixed(-1150.0/65536.0,1,-nbitq), 
to_sfixed(-554.0/65536.0,1,-nbitq), 
to_sfixed(2536.0/65536.0,1,-nbitq), 
to_sfixed(-1669.0/65536.0,1,-nbitq), 
to_sfixed(-1002.0/65536.0,1,-nbitq), 
to_sfixed(-66.0/65536.0,1,-nbitq), 
to_sfixed(-569.0/65536.0,1,-nbitq), 
to_sfixed(-734.0/65536.0,1,-nbitq), 
to_sfixed(552.0/65536.0,1,-nbitq), 
to_sfixed(-4848.0/65536.0,1,-nbitq), 
to_sfixed(-4481.0/65536.0,1,-nbitq), 
to_sfixed(-6.0/65536.0,1,-nbitq), 
to_sfixed(22.0/65536.0,1,-nbitq), 
to_sfixed(-1137.0/65536.0,1,-nbitq), 
to_sfixed(-1109.0/65536.0,1,-nbitq), 
to_sfixed(-2212.0/65536.0,1,-nbitq), 
to_sfixed(-2328.0/65536.0,1,-nbitq), 
to_sfixed(1461.0/65536.0,1,-nbitq), 
to_sfixed(-1171.0/65536.0,1,-nbitq), 
to_sfixed(-851.0/65536.0,1,-nbitq), 
to_sfixed(2201.0/65536.0,1,-nbitq), 
to_sfixed(1132.0/65536.0,1,-nbitq), 
to_sfixed(3319.0/65536.0,1,-nbitq), 
to_sfixed(1379.0/65536.0,1,-nbitq), 
to_sfixed(1698.0/65536.0,1,-nbitq), 
to_sfixed(50.0/65536.0,1,-nbitq), 
to_sfixed(-220.0/65536.0,1,-nbitq), 
to_sfixed(-2425.0/65536.0,1,-nbitq), 
to_sfixed(259.0/65536.0,1,-nbitq), 
to_sfixed(2743.0/65536.0,1,-nbitq), 
to_sfixed(1378.0/65536.0,1,-nbitq), 
to_sfixed(2967.0/65536.0,1,-nbitq), 
to_sfixed(567.0/65536.0,1,-nbitq), 
to_sfixed(1279.0/65536.0,1,-nbitq), 
to_sfixed(1418.0/65536.0,1,-nbitq), 
to_sfixed(1730.0/65536.0,1,-nbitq), 
to_sfixed(829.0/65536.0,1,-nbitq), 
to_sfixed(-3084.0/65536.0,1,-nbitq), 
to_sfixed(978.0/65536.0,1,-nbitq), 
to_sfixed(-732.0/65536.0,1,-nbitq), 
to_sfixed(387.0/65536.0,1,-nbitq), 
to_sfixed(2682.0/65536.0,1,-nbitq), 
to_sfixed(63.0/65536.0,1,-nbitq), 
to_sfixed(2025.0/65536.0,1,-nbitq), 
to_sfixed(2136.0/65536.0,1,-nbitq), 
to_sfixed(361.0/65536.0,1,-nbitq), 
to_sfixed(-857.0/65536.0,1,-nbitq), 
to_sfixed(-1735.0/65536.0,1,-nbitq), 
to_sfixed(2009.0/65536.0,1,-nbitq), 
to_sfixed(3223.0/65536.0,1,-nbitq), 
to_sfixed(810.0/65536.0,1,-nbitq), 
to_sfixed(-1828.0/65536.0,1,-nbitq), 
to_sfixed(107.0/65536.0,1,-nbitq), 
to_sfixed(-3204.0/65536.0,1,-nbitq), 
to_sfixed(-200.0/65536.0,1,-nbitq), 
to_sfixed(-840.0/65536.0,1,-nbitq), 
to_sfixed(4679.0/65536.0,1,-nbitq)  ), 
( to_sfixed(904.0/65536.0,1,-nbitq), 
to_sfixed(-1242.0/65536.0,1,-nbitq), 
to_sfixed(4015.0/65536.0,1,-nbitq), 
to_sfixed(-2431.0/65536.0,1,-nbitq), 
to_sfixed(2916.0/65536.0,1,-nbitq), 
to_sfixed(-2653.0/65536.0,1,-nbitq), 
to_sfixed(207.0/65536.0,1,-nbitq), 
to_sfixed(1391.0/65536.0,1,-nbitq), 
to_sfixed(-3896.0/65536.0,1,-nbitq), 
to_sfixed(2221.0/65536.0,1,-nbitq), 
to_sfixed(1874.0/65536.0,1,-nbitq), 
to_sfixed(-532.0/65536.0,1,-nbitq), 
to_sfixed(-726.0/65536.0,1,-nbitq), 
to_sfixed(190.0/65536.0,1,-nbitq), 
to_sfixed(5268.0/65536.0,1,-nbitq), 
to_sfixed(176.0/65536.0,1,-nbitq), 
to_sfixed(-2167.0/65536.0,1,-nbitq), 
to_sfixed(976.0/65536.0,1,-nbitq), 
to_sfixed(-2550.0/65536.0,1,-nbitq), 
to_sfixed(2909.0/65536.0,1,-nbitq), 
to_sfixed(536.0/65536.0,1,-nbitq), 
to_sfixed(-882.0/65536.0,1,-nbitq), 
to_sfixed(-869.0/65536.0,1,-nbitq), 
to_sfixed(3703.0/65536.0,1,-nbitq), 
to_sfixed(1590.0/65536.0,1,-nbitq), 
to_sfixed(3852.0/65536.0,1,-nbitq), 
to_sfixed(-2156.0/65536.0,1,-nbitq), 
to_sfixed(-1256.0/65536.0,1,-nbitq), 
to_sfixed(3180.0/65536.0,1,-nbitq), 
to_sfixed(81.0/65536.0,1,-nbitq), 
to_sfixed(-526.0/65536.0,1,-nbitq), 
to_sfixed(1296.0/65536.0,1,-nbitq), 
to_sfixed(-1180.0/65536.0,1,-nbitq), 
to_sfixed(-5011.0/65536.0,1,-nbitq), 
to_sfixed(-2996.0/65536.0,1,-nbitq), 
to_sfixed(-3111.0/65536.0,1,-nbitq), 
to_sfixed(-3234.0/65536.0,1,-nbitq), 
to_sfixed(388.0/65536.0,1,-nbitq), 
to_sfixed(-3728.0/65536.0,1,-nbitq), 
to_sfixed(-476.0/65536.0,1,-nbitq), 
to_sfixed(282.0/65536.0,1,-nbitq), 
to_sfixed(-1101.0/65536.0,1,-nbitq), 
to_sfixed(-934.0/65536.0,1,-nbitq), 
to_sfixed(-903.0/65536.0,1,-nbitq), 
to_sfixed(817.0/65536.0,1,-nbitq), 
to_sfixed(3966.0/65536.0,1,-nbitq), 
to_sfixed(1527.0/65536.0,1,-nbitq), 
to_sfixed(-2069.0/65536.0,1,-nbitq), 
to_sfixed(3399.0/65536.0,1,-nbitq), 
to_sfixed(1118.0/65536.0,1,-nbitq), 
to_sfixed(2147.0/65536.0,1,-nbitq), 
to_sfixed(-534.0/65536.0,1,-nbitq), 
to_sfixed(2540.0/65536.0,1,-nbitq), 
to_sfixed(-1135.0/65536.0,1,-nbitq), 
to_sfixed(1136.0/65536.0,1,-nbitq), 
to_sfixed(-2597.0/65536.0,1,-nbitq), 
to_sfixed(769.0/65536.0,1,-nbitq), 
to_sfixed(-699.0/65536.0,1,-nbitq), 
to_sfixed(1240.0/65536.0,1,-nbitq), 
to_sfixed(2180.0/65536.0,1,-nbitq), 
to_sfixed(-3107.0/65536.0,1,-nbitq), 
to_sfixed(1783.0/65536.0,1,-nbitq), 
to_sfixed(-2270.0/65536.0,1,-nbitq), 
to_sfixed(-1793.0/65536.0,1,-nbitq), 
to_sfixed(331.0/65536.0,1,-nbitq), 
to_sfixed(2812.0/65536.0,1,-nbitq), 
to_sfixed(-2229.0/65536.0,1,-nbitq), 
to_sfixed(-3236.0/65536.0,1,-nbitq), 
to_sfixed(-2841.0/65536.0,1,-nbitq), 
to_sfixed(-787.0/65536.0,1,-nbitq), 
to_sfixed(-797.0/65536.0,1,-nbitq), 
to_sfixed(-1028.0/65536.0,1,-nbitq), 
to_sfixed(2271.0/65536.0,1,-nbitq), 
to_sfixed(1277.0/65536.0,1,-nbitq), 
to_sfixed(2284.0/65536.0,1,-nbitq), 
to_sfixed(1244.0/65536.0,1,-nbitq), 
to_sfixed(1698.0/65536.0,1,-nbitq), 
to_sfixed(-752.0/65536.0,1,-nbitq), 
to_sfixed(851.0/65536.0,1,-nbitq), 
to_sfixed(3602.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-756.0/65536.0,1,-nbitq), 
to_sfixed(373.0/65536.0,1,-nbitq), 
to_sfixed(-1415.0/65536.0,1,-nbitq), 
to_sfixed(-422.0/65536.0,1,-nbitq), 
to_sfixed(960.0/65536.0,1,-nbitq), 
to_sfixed(-3612.0/65536.0,1,-nbitq), 
to_sfixed(-666.0/65536.0,1,-nbitq), 
to_sfixed(-597.0/65536.0,1,-nbitq), 
to_sfixed(-2238.0/65536.0,1,-nbitq), 
to_sfixed(-572.0/65536.0,1,-nbitq), 
to_sfixed(-114.0/65536.0,1,-nbitq), 
to_sfixed(-1515.0/65536.0,1,-nbitq), 
to_sfixed(764.0/65536.0,1,-nbitq), 
to_sfixed(-3579.0/65536.0,1,-nbitq), 
to_sfixed(4909.0/65536.0,1,-nbitq), 
to_sfixed(2470.0/65536.0,1,-nbitq), 
to_sfixed(-1689.0/65536.0,1,-nbitq), 
to_sfixed(1770.0/65536.0,1,-nbitq), 
to_sfixed(-3677.0/65536.0,1,-nbitq), 
to_sfixed(-2428.0/65536.0,1,-nbitq), 
to_sfixed(192.0/65536.0,1,-nbitq), 
to_sfixed(2079.0/65536.0,1,-nbitq), 
to_sfixed(-414.0/65536.0,1,-nbitq), 
to_sfixed(3463.0/65536.0,1,-nbitq), 
to_sfixed(1469.0/65536.0,1,-nbitq), 
to_sfixed(3539.0/65536.0,1,-nbitq), 
to_sfixed(1996.0/65536.0,1,-nbitq), 
to_sfixed(-1862.0/65536.0,1,-nbitq), 
to_sfixed(4996.0/65536.0,1,-nbitq), 
to_sfixed(-5473.0/65536.0,1,-nbitq), 
to_sfixed(-2114.0/65536.0,1,-nbitq), 
to_sfixed(970.0/65536.0,1,-nbitq), 
to_sfixed(-2629.0/65536.0,1,-nbitq), 
to_sfixed(-1035.0/65536.0,1,-nbitq), 
to_sfixed(2544.0/65536.0,1,-nbitq), 
to_sfixed(-160.0/65536.0,1,-nbitq), 
to_sfixed(-1577.0/65536.0,1,-nbitq), 
to_sfixed(-1004.0/65536.0,1,-nbitq), 
to_sfixed(-896.0/65536.0,1,-nbitq), 
to_sfixed(96.0/65536.0,1,-nbitq), 
to_sfixed(-5431.0/65536.0,1,-nbitq), 
to_sfixed(597.0/65536.0,1,-nbitq), 
to_sfixed(-1588.0/65536.0,1,-nbitq), 
to_sfixed(180.0/65536.0,1,-nbitq), 
to_sfixed(-2048.0/65536.0,1,-nbitq), 
to_sfixed(2972.0/65536.0,1,-nbitq), 
to_sfixed(2713.0/65536.0,1,-nbitq), 
to_sfixed(1103.0/65536.0,1,-nbitq), 
to_sfixed(-914.0/65536.0,1,-nbitq), 
to_sfixed(-71.0/65536.0,1,-nbitq), 
to_sfixed(343.0/65536.0,1,-nbitq), 
to_sfixed(1238.0/65536.0,1,-nbitq), 
to_sfixed(-755.0/65536.0,1,-nbitq), 
to_sfixed(148.0/65536.0,1,-nbitq), 
to_sfixed(3051.0/65536.0,1,-nbitq), 
to_sfixed(-1458.0/65536.0,1,-nbitq), 
to_sfixed(-144.0/65536.0,1,-nbitq), 
to_sfixed(1769.0/65536.0,1,-nbitq), 
to_sfixed(2327.0/65536.0,1,-nbitq), 
to_sfixed(-779.0/65536.0,1,-nbitq), 
to_sfixed(-4220.0/65536.0,1,-nbitq), 
to_sfixed(2320.0/65536.0,1,-nbitq), 
to_sfixed(1877.0/65536.0,1,-nbitq), 
to_sfixed(-2487.0/65536.0,1,-nbitq), 
to_sfixed(1101.0/65536.0,1,-nbitq), 
to_sfixed(-432.0/65536.0,1,-nbitq), 
to_sfixed(-1150.0/65536.0,1,-nbitq), 
to_sfixed(1533.0/65536.0,1,-nbitq), 
to_sfixed(-995.0/65536.0,1,-nbitq), 
to_sfixed(1478.0/65536.0,1,-nbitq), 
to_sfixed(2426.0/65536.0,1,-nbitq), 
to_sfixed(-1257.0/65536.0,1,-nbitq), 
to_sfixed(-495.0/65536.0,1,-nbitq), 
to_sfixed(341.0/65536.0,1,-nbitq), 
to_sfixed(2395.0/65536.0,1,-nbitq), 
to_sfixed(3598.0/65536.0,1,-nbitq), 
to_sfixed(-5280.0/65536.0,1,-nbitq), 
to_sfixed(3047.0/65536.0,1,-nbitq), 
to_sfixed(-1514.0/65536.0,1,-nbitq), 
to_sfixed(-630.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-587.0/65536.0,1,-nbitq), 
to_sfixed(-2450.0/65536.0,1,-nbitq), 
to_sfixed(-1460.0/65536.0,1,-nbitq), 
to_sfixed(1994.0/65536.0,1,-nbitq), 
to_sfixed(-210.0/65536.0,1,-nbitq), 
to_sfixed(895.0/65536.0,1,-nbitq), 
to_sfixed(-2535.0/65536.0,1,-nbitq), 
to_sfixed(-1016.0/65536.0,1,-nbitq), 
to_sfixed(1048.0/65536.0,1,-nbitq), 
to_sfixed(2349.0/65536.0,1,-nbitq), 
to_sfixed(2128.0/65536.0,1,-nbitq), 
to_sfixed(-9063.0/65536.0,1,-nbitq), 
to_sfixed(996.0/65536.0,1,-nbitq), 
to_sfixed(3492.0/65536.0,1,-nbitq), 
to_sfixed(3752.0/65536.0,1,-nbitq), 
to_sfixed(946.0/65536.0,1,-nbitq), 
to_sfixed(-707.0/65536.0,1,-nbitq), 
to_sfixed(1064.0/65536.0,1,-nbitq), 
to_sfixed(1347.0/65536.0,1,-nbitq), 
to_sfixed(454.0/65536.0,1,-nbitq), 
to_sfixed(1527.0/65536.0,1,-nbitq), 
to_sfixed(3134.0/65536.0,1,-nbitq), 
to_sfixed(3558.0/65536.0,1,-nbitq), 
to_sfixed(2954.0/65536.0,1,-nbitq), 
to_sfixed(2606.0/65536.0,1,-nbitq), 
to_sfixed(7448.0/65536.0,1,-nbitq), 
to_sfixed(1738.0/65536.0,1,-nbitq), 
to_sfixed(-502.0/65536.0,1,-nbitq), 
to_sfixed(6582.0/65536.0,1,-nbitq), 
to_sfixed(-2386.0/65536.0,1,-nbitq), 
to_sfixed(-991.0/65536.0,1,-nbitq), 
to_sfixed(-345.0/65536.0,1,-nbitq), 
to_sfixed(3313.0/65536.0,1,-nbitq), 
to_sfixed(-6432.0/65536.0,1,-nbitq), 
to_sfixed(-3.0/65536.0,1,-nbitq), 
to_sfixed(1708.0/65536.0,1,-nbitq), 
to_sfixed(-7901.0/65536.0,1,-nbitq), 
to_sfixed(1164.0/65536.0,1,-nbitq), 
to_sfixed(-8407.0/65536.0,1,-nbitq), 
to_sfixed(-2547.0/65536.0,1,-nbitq), 
to_sfixed(-33.0/65536.0,1,-nbitq), 
to_sfixed(-545.0/65536.0,1,-nbitq), 
to_sfixed(1364.0/65536.0,1,-nbitq), 
to_sfixed(1839.0/65536.0,1,-nbitq), 
to_sfixed(185.0/65536.0,1,-nbitq), 
to_sfixed(3064.0/65536.0,1,-nbitq), 
to_sfixed(37.0/65536.0,1,-nbitq), 
to_sfixed(-580.0/65536.0,1,-nbitq), 
to_sfixed(-1170.0/65536.0,1,-nbitq), 
to_sfixed(-1755.0/65536.0,1,-nbitq), 
to_sfixed(1537.0/65536.0,1,-nbitq), 
to_sfixed(1128.0/65536.0,1,-nbitq), 
to_sfixed(-2082.0/65536.0,1,-nbitq), 
to_sfixed(1103.0/65536.0,1,-nbitq), 
to_sfixed(447.0/65536.0,1,-nbitq), 
to_sfixed(2283.0/65536.0,1,-nbitq), 
to_sfixed(1768.0/65536.0,1,-nbitq), 
to_sfixed(3298.0/65536.0,1,-nbitq), 
to_sfixed(-2147.0/65536.0,1,-nbitq), 
to_sfixed(-2143.0/65536.0,1,-nbitq), 
to_sfixed(-7991.0/65536.0,1,-nbitq), 
to_sfixed(1008.0/65536.0,1,-nbitq), 
to_sfixed(1161.0/65536.0,1,-nbitq), 
to_sfixed(726.0/65536.0,1,-nbitq), 
to_sfixed(2120.0/65536.0,1,-nbitq), 
to_sfixed(1572.0/65536.0,1,-nbitq), 
to_sfixed(568.0/65536.0,1,-nbitq), 
to_sfixed(2525.0/65536.0,1,-nbitq), 
to_sfixed(3477.0/65536.0,1,-nbitq), 
to_sfixed(-4511.0/65536.0,1,-nbitq), 
to_sfixed(1663.0/65536.0,1,-nbitq), 
to_sfixed(2013.0/65536.0,1,-nbitq), 
to_sfixed(2742.0/65536.0,1,-nbitq), 
to_sfixed(1157.0/65536.0,1,-nbitq), 
to_sfixed(-780.0/65536.0,1,-nbitq), 
to_sfixed(4703.0/65536.0,1,-nbitq), 
to_sfixed(-3220.0/65536.0,1,-nbitq), 
to_sfixed(-3630.0/65536.0,1,-nbitq), 
to_sfixed(68.0/65536.0,1,-nbitq), 
to_sfixed(368.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3822.0/65536.0,1,-nbitq), 
to_sfixed(-2813.0/65536.0,1,-nbitq), 
to_sfixed(-388.0/65536.0,1,-nbitq), 
to_sfixed(-695.0/65536.0,1,-nbitq), 
to_sfixed(402.0/65536.0,1,-nbitq), 
to_sfixed(-4232.0/65536.0,1,-nbitq), 
to_sfixed(-995.0/65536.0,1,-nbitq), 
to_sfixed(-6248.0/65536.0,1,-nbitq), 
to_sfixed(-2361.0/65536.0,1,-nbitq), 
to_sfixed(695.0/65536.0,1,-nbitq), 
to_sfixed(1089.0/65536.0,1,-nbitq), 
to_sfixed(-893.0/65536.0,1,-nbitq), 
to_sfixed(-342.0/65536.0,1,-nbitq), 
to_sfixed(3032.0/65536.0,1,-nbitq), 
to_sfixed(-901.0/65536.0,1,-nbitq), 
to_sfixed(-61.0/65536.0,1,-nbitq), 
to_sfixed(2745.0/65536.0,1,-nbitq), 
to_sfixed(-2704.0/65536.0,1,-nbitq), 
to_sfixed(639.0/65536.0,1,-nbitq), 
to_sfixed(2266.0/65536.0,1,-nbitq), 
to_sfixed(4575.0/65536.0,1,-nbitq), 
to_sfixed(3988.0/65536.0,1,-nbitq), 
to_sfixed(6281.0/65536.0,1,-nbitq), 
to_sfixed(-2006.0/65536.0,1,-nbitq), 
to_sfixed(2386.0/65536.0,1,-nbitq), 
to_sfixed(-378.0/65536.0,1,-nbitq), 
to_sfixed(2644.0/65536.0,1,-nbitq), 
to_sfixed(-1482.0/65536.0,1,-nbitq), 
to_sfixed(355.0/65536.0,1,-nbitq), 
to_sfixed(-1430.0/65536.0,1,-nbitq), 
to_sfixed(-1962.0/65536.0,1,-nbitq), 
to_sfixed(2491.0/65536.0,1,-nbitq), 
to_sfixed(-58.0/65536.0,1,-nbitq), 
to_sfixed(-15820.0/65536.0,1,-nbitq), 
to_sfixed(-1472.0/65536.0,1,-nbitq), 
to_sfixed(2537.0/65536.0,1,-nbitq), 
to_sfixed(-11042.0/65536.0,1,-nbitq), 
to_sfixed(3969.0/65536.0,1,-nbitq), 
to_sfixed(-12121.0/65536.0,1,-nbitq), 
to_sfixed(-2505.0/65536.0,1,-nbitq), 
to_sfixed(7367.0/65536.0,1,-nbitq), 
to_sfixed(-2736.0/65536.0,1,-nbitq), 
to_sfixed(244.0/65536.0,1,-nbitq), 
to_sfixed(1390.0/65536.0,1,-nbitq), 
to_sfixed(2626.0/65536.0,1,-nbitq), 
to_sfixed(4357.0/65536.0,1,-nbitq), 
to_sfixed(1318.0/65536.0,1,-nbitq), 
to_sfixed(468.0/65536.0,1,-nbitq), 
to_sfixed(2952.0/65536.0,1,-nbitq), 
to_sfixed(1277.0/65536.0,1,-nbitq), 
to_sfixed(1160.0/65536.0,1,-nbitq), 
to_sfixed(5179.0/65536.0,1,-nbitq), 
to_sfixed(2361.0/65536.0,1,-nbitq), 
to_sfixed(2152.0/65536.0,1,-nbitq), 
to_sfixed(-1973.0/65536.0,1,-nbitq), 
to_sfixed(6908.0/65536.0,1,-nbitq), 
to_sfixed(-1007.0/65536.0,1,-nbitq), 
to_sfixed(4415.0/65536.0,1,-nbitq), 
to_sfixed(2654.0/65536.0,1,-nbitq), 
to_sfixed(-13786.0/65536.0,1,-nbitq), 
to_sfixed(-9920.0/65536.0,1,-nbitq), 
to_sfixed(-2965.0/65536.0,1,-nbitq), 
to_sfixed(-424.0/65536.0,1,-nbitq), 
to_sfixed(194.0/65536.0,1,-nbitq), 
to_sfixed(3417.0/65536.0,1,-nbitq), 
to_sfixed(3553.0/65536.0,1,-nbitq), 
to_sfixed(-1985.0/65536.0,1,-nbitq), 
to_sfixed(2511.0/65536.0,1,-nbitq), 
to_sfixed(4682.0/65536.0,1,-nbitq), 
to_sfixed(-2937.0/65536.0,1,-nbitq), 
to_sfixed(-688.0/65536.0,1,-nbitq), 
to_sfixed(1997.0/65536.0,1,-nbitq), 
to_sfixed(-1222.0/65536.0,1,-nbitq), 
to_sfixed(-1478.0/65536.0,1,-nbitq), 
to_sfixed(-2043.0/65536.0,1,-nbitq), 
to_sfixed(-3816.0/65536.0,1,-nbitq), 
to_sfixed(-4510.0/65536.0,1,-nbitq), 
to_sfixed(-980.0/65536.0,1,-nbitq), 
to_sfixed(2642.0/65536.0,1,-nbitq), 
to_sfixed(2401.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-432.0/65536.0,1,-nbitq), 
to_sfixed(-3065.0/65536.0,1,-nbitq), 
to_sfixed(-2274.0/65536.0,1,-nbitq), 
to_sfixed(901.0/65536.0,1,-nbitq), 
to_sfixed(624.0/65536.0,1,-nbitq), 
to_sfixed(-4132.0/65536.0,1,-nbitq), 
to_sfixed(-4892.0/65536.0,1,-nbitq), 
to_sfixed(-4964.0/65536.0,1,-nbitq), 
to_sfixed(-1136.0/65536.0,1,-nbitq), 
to_sfixed(-2452.0/65536.0,1,-nbitq), 
to_sfixed(3664.0/65536.0,1,-nbitq), 
to_sfixed(4726.0/65536.0,1,-nbitq), 
to_sfixed(1839.0/65536.0,1,-nbitq), 
to_sfixed(-3119.0/65536.0,1,-nbitq), 
to_sfixed(-576.0/65536.0,1,-nbitq), 
to_sfixed(-1336.0/65536.0,1,-nbitq), 
to_sfixed(993.0/65536.0,1,-nbitq), 
to_sfixed(-1070.0/65536.0,1,-nbitq), 
to_sfixed(3697.0/65536.0,1,-nbitq), 
to_sfixed(-821.0/65536.0,1,-nbitq), 
to_sfixed(1237.0/65536.0,1,-nbitq), 
to_sfixed(-1585.0/65536.0,1,-nbitq), 
to_sfixed(4171.0/65536.0,1,-nbitq), 
to_sfixed(-5243.0/65536.0,1,-nbitq), 
to_sfixed(2778.0/65536.0,1,-nbitq), 
to_sfixed(-9086.0/65536.0,1,-nbitq), 
to_sfixed(-282.0/65536.0,1,-nbitq), 
to_sfixed(4263.0/65536.0,1,-nbitq), 
to_sfixed(-125.0/65536.0,1,-nbitq), 
to_sfixed(-4757.0/65536.0,1,-nbitq), 
to_sfixed(3186.0/65536.0,1,-nbitq), 
to_sfixed(-3941.0/65536.0,1,-nbitq), 
to_sfixed(-2105.0/65536.0,1,-nbitq), 
to_sfixed(-15154.0/65536.0,1,-nbitq), 
to_sfixed(1183.0/65536.0,1,-nbitq), 
to_sfixed(1788.0/65536.0,1,-nbitq), 
to_sfixed(-10976.0/65536.0,1,-nbitq), 
to_sfixed(6023.0/65536.0,1,-nbitq), 
to_sfixed(-9221.0/65536.0,1,-nbitq), 
to_sfixed(-9231.0/65536.0,1,-nbitq), 
to_sfixed(9669.0/65536.0,1,-nbitq), 
to_sfixed(506.0/65536.0,1,-nbitq), 
to_sfixed(6307.0/65536.0,1,-nbitq), 
to_sfixed(-795.0/65536.0,1,-nbitq), 
to_sfixed(-2275.0/65536.0,1,-nbitq), 
to_sfixed(1137.0/65536.0,1,-nbitq), 
to_sfixed(274.0/65536.0,1,-nbitq), 
to_sfixed(1148.0/65536.0,1,-nbitq), 
to_sfixed(-1205.0/65536.0,1,-nbitq), 
to_sfixed(276.0/65536.0,1,-nbitq), 
to_sfixed(1058.0/65536.0,1,-nbitq), 
to_sfixed(6762.0/65536.0,1,-nbitq), 
to_sfixed(-1150.0/65536.0,1,-nbitq), 
to_sfixed(-3933.0/65536.0,1,-nbitq), 
to_sfixed(-5883.0/65536.0,1,-nbitq), 
to_sfixed(10587.0/65536.0,1,-nbitq), 
to_sfixed(2643.0/65536.0,1,-nbitq), 
to_sfixed(-365.0/65536.0,1,-nbitq), 
to_sfixed(-2378.0/65536.0,1,-nbitq), 
to_sfixed(-9018.0/65536.0,1,-nbitq), 
to_sfixed(-8825.0/65536.0,1,-nbitq), 
to_sfixed(2637.0/65536.0,1,-nbitq), 
to_sfixed(241.0/65536.0,1,-nbitq), 
to_sfixed(-1350.0/65536.0,1,-nbitq), 
to_sfixed(7562.0/65536.0,1,-nbitq), 
to_sfixed(5933.0/65536.0,1,-nbitq), 
to_sfixed(5036.0/65536.0,1,-nbitq), 
to_sfixed(3248.0/65536.0,1,-nbitq), 
to_sfixed(-20.0/65536.0,1,-nbitq), 
to_sfixed(-403.0/65536.0,1,-nbitq), 
to_sfixed(-1231.0/65536.0,1,-nbitq), 
to_sfixed(-2588.0/65536.0,1,-nbitq), 
to_sfixed(3342.0/65536.0,1,-nbitq), 
to_sfixed(889.0/65536.0,1,-nbitq), 
to_sfixed(-253.0/65536.0,1,-nbitq), 
to_sfixed(-3809.0/65536.0,1,-nbitq), 
to_sfixed(-3002.0/65536.0,1,-nbitq), 
to_sfixed(-4107.0/65536.0,1,-nbitq), 
to_sfixed(332.0/65536.0,1,-nbitq), 
to_sfixed(1070.0/65536.0,1,-nbitq)  ), 
( to_sfixed(375.0/65536.0,1,-nbitq), 
to_sfixed(-323.0/65536.0,1,-nbitq), 
to_sfixed(6277.0/65536.0,1,-nbitq), 
to_sfixed(3065.0/65536.0,1,-nbitq), 
to_sfixed(-2219.0/65536.0,1,-nbitq), 
to_sfixed(-4056.0/65536.0,1,-nbitq), 
to_sfixed(-6254.0/65536.0,1,-nbitq), 
to_sfixed(-8572.0/65536.0,1,-nbitq), 
to_sfixed(2272.0/65536.0,1,-nbitq), 
to_sfixed(1698.0/65536.0,1,-nbitq), 
to_sfixed(2751.0/65536.0,1,-nbitq), 
to_sfixed(13722.0/65536.0,1,-nbitq), 
to_sfixed(383.0/65536.0,1,-nbitq), 
to_sfixed(-1350.0/65536.0,1,-nbitq), 
to_sfixed(-3439.0/65536.0,1,-nbitq), 
to_sfixed(622.0/65536.0,1,-nbitq), 
to_sfixed(-840.0/65536.0,1,-nbitq), 
to_sfixed(1455.0/65536.0,1,-nbitq), 
to_sfixed(-1538.0/65536.0,1,-nbitq), 
to_sfixed(3226.0/65536.0,1,-nbitq), 
to_sfixed(-7911.0/65536.0,1,-nbitq), 
to_sfixed(-8476.0/65536.0,1,-nbitq), 
to_sfixed(-4569.0/65536.0,1,-nbitq), 
to_sfixed(1955.0/65536.0,1,-nbitq), 
to_sfixed(2263.0/65536.0,1,-nbitq), 
to_sfixed(-9154.0/65536.0,1,-nbitq), 
to_sfixed(-5287.0/65536.0,1,-nbitq), 
to_sfixed(5797.0/65536.0,1,-nbitq), 
to_sfixed(-1902.0/65536.0,1,-nbitq), 
to_sfixed(-5045.0/65536.0,1,-nbitq), 
to_sfixed(-897.0/65536.0,1,-nbitq), 
to_sfixed(-368.0/65536.0,1,-nbitq), 
to_sfixed(-2361.0/65536.0,1,-nbitq), 
to_sfixed(-12794.0/65536.0,1,-nbitq), 
to_sfixed(-479.0/65536.0,1,-nbitq), 
to_sfixed(-2474.0/65536.0,1,-nbitq), 
to_sfixed(-16763.0/65536.0,1,-nbitq), 
to_sfixed(2245.0/65536.0,1,-nbitq), 
to_sfixed(-14201.0/65536.0,1,-nbitq), 
to_sfixed(-9678.0/65536.0,1,-nbitq), 
to_sfixed(6355.0/65536.0,1,-nbitq), 
to_sfixed(1088.0/65536.0,1,-nbitq), 
to_sfixed(-1800.0/65536.0,1,-nbitq), 
to_sfixed(204.0/65536.0,1,-nbitq), 
to_sfixed(688.0/65536.0,1,-nbitq), 
to_sfixed(618.0/65536.0,1,-nbitq), 
to_sfixed(507.0/65536.0,1,-nbitq), 
to_sfixed(1693.0/65536.0,1,-nbitq), 
to_sfixed(3354.0/65536.0,1,-nbitq), 
to_sfixed(3494.0/65536.0,1,-nbitq), 
to_sfixed(2515.0/65536.0,1,-nbitq), 
to_sfixed(7277.0/65536.0,1,-nbitq), 
to_sfixed(-2032.0/65536.0,1,-nbitq), 
to_sfixed(266.0/65536.0,1,-nbitq), 
to_sfixed(-6085.0/65536.0,1,-nbitq), 
to_sfixed(2066.0/65536.0,1,-nbitq), 
to_sfixed(1743.0/65536.0,1,-nbitq), 
to_sfixed(-5461.0/65536.0,1,-nbitq), 
to_sfixed(543.0/65536.0,1,-nbitq), 
to_sfixed(-4635.0/65536.0,1,-nbitq), 
to_sfixed(-2137.0/65536.0,1,-nbitq), 
to_sfixed(3056.0/65536.0,1,-nbitq), 
to_sfixed(1241.0/65536.0,1,-nbitq), 
to_sfixed(-1128.0/65536.0,1,-nbitq), 
to_sfixed(2932.0/65536.0,1,-nbitq), 
to_sfixed(4581.0/65536.0,1,-nbitq), 
to_sfixed(96.0/65536.0,1,-nbitq), 
to_sfixed(3934.0/65536.0,1,-nbitq), 
to_sfixed(88.0/65536.0,1,-nbitq), 
to_sfixed(9671.0/65536.0,1,-nbitq), 
to_sfixed(-3294.0/65536.0,1,-nbitq), 
to_sfixed(2423.0/65536.0,1,-nbitq), 
to_sfixed(2474.0/65536.0,1,-nbitq), 
to_sfixed(-2732.0/65536.0,1,-nbitq), 
to_sfixed(1501.0/65536.0,1,-nbitq), 
to_sfixed(1059.0/65536.0,1,-nbitq), 
to_sfixed(-6106.0/65536.0,1,-nbitq), 
to_sfixed(-6203.0/65536.0,1,-nbitq), 
to_sfixed(866.0/65536.0,1,-nbitq), 
to_sfixed(3168.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4465.0/65536.0,1,-nbitq), 
to_sfixed(-233.0/65536.0,1,-nbitq), 
to_sfixed(6037.0/65536.0,1,-nbitq), 
to_sfixed(5618.0/65536.0,1,-nbitq), 
to_sfixed(-3280.0/65536.0,1,-nbitq), 
to_sfixed(-1024.0/65536.0,1,-nbitq), 
to_sfixed(-5226.0/65536.0,1,-nbitq), 
to_sfixed(1791.0/65536.0,1,-nbitq), 
to_sfixed(5682.0/65536.0,1,-nbitq), 
to_sfixed(-214.0/65536.0,1,-nbitq), 
to_sfixed(2345.0/65536.0,1,-nbitq), 
to_sfixed(1729.0/65536.0,1,-nbitq), 
to_sfixed(516.0/65536.0,1,-nbitq), 
to_sfixed(-721.0/65536.0,1,-nbitq), 
to_sfixed(1362.0/65536.0,1,-nbitq), 
to_sfixed(2394.0/65536.0,1,-nbitq), 
to_sfixed(-2651.0/65536.0,1,-nbitq), 
to_sfixed(6103.0/65536.0,1,-nbitq), 
to_sfixed(1665.0/65536.0,1,-nbitq), 
to_sfixed(29.0/65536.0,1,-nbitq), 
to_sfixed(-3667.0/65536.0,1,-nbitq), 
to_sfixed(-1885.0/65536.0,1,-nbitq), 
to_sfixed(-3864.0/65536.0,1,-nbitq), 
to_sfixed(13228.0/65536.0,1,-nbitq), 
to_sfixed(-2722.0/65536.0,1,-nbitq), 
to_sfixed(-12315.0/65536.0,1,-nbitq), 
to_sfixed(-1148.0/65536.0,1,-nbitq), 
to_sfixed(2213.0/65536.0,1,-nbitq), 
to_sfixed(-139.0/65536.0,1,-nbitq), 
to_sfixed(-2063.0/65536.0,1,-nbitq), 
to_sfixed(2181.0/65536.0,1,-nbitq), 
to_sfixed(5869.0/65536.0,1,-nbitq), 
to_sfixed(2740.0/65536.0,1,-nbitq), 
to_sfixed(-13510.0/65536.0,1,-nbitq), 
to_sfixed(-3617.0/65536.0,1,-nbitq), 
to_sfixed(358.0/65536.0,1,-nbitq), 
to_sfixed(-10894.0/65536.0,1,-nbitq), 
to_sfixed(4086.0/65536.0,1,-nbitq), 
to_sfixed(-4328.0/65536.0,1,-nbitq), 
to_sfixed(-5499.0/65536.0,1,-nbitq), 
to_sfixed(6410.0/65536.0,1,-nbitq), 
to_sfixed(-1451.0/65536.0,1,-nbitq), 
to_sfixed(-2227.0/65536.0,1,-nbitq), 
to_sfixed(6352.0/65536.0,1,-nbitq), 
to_sfixed(-1554.0/65536.0,1,-nbitq), 
to_sfixed(-1818.0/65536.0,1,-nbitq), 
to_sfixed(3896.0/65536.0,1,-nbitq), 
to_sfixed(3753.0/65536.0,1,-nbitq), 
to_sfixed(1276.0/65536.0,1,-nbitq), 
to_sfixed(3479.0/65536.0,1,-nbitq), 
to_sfixed(178.0/65536.0,1,-nbitq), 
to_sfixed(4206.0/65536.0,1,-nbitq), 
to_sfixed(-884.0/65536.0,1,-nbitq), 
to_sfixed(727.0/65536.0,1,-nbitq), 
to_sfixed(-4758.0/65536.0,1,-nbitq), 
to_sfixed(5813.0/65536.0,1,-nbitq), 
to_sfixed(-301.0/65536.0,1,-nbitq), 
to_sfixed(-3068.0/65536.0,1,-nbitq), 
to_sfixed(767.0/65536.0,1,-nbitq), 
to_sfixed(-4480.0/65536.0,1,-nbitq), 
to_sfixed(7256.0/65536.0,1,-nbitq), 
to_sfixed(2497.0/65536.0,1,-nbitq), 
to_sfixed(1678.0/65536.0,1,-nbitq), 
to_sfixed(1336.0/65536.0,1,-nbitq), 
to_sfixed(6967.0/65536.0,1,-nbitq), 
to_sfixed(5109.0/65536.0,1,-nbitq), 
to_sfixed(4575.0/65536.0,1,-nbitq), 
to_sfixed(15406.0/65536.0,1,-nbitq), 
to_sfixed(-2055.0/65536.0,1,-nbitq), 
to_sfixed(5014.0/65536.0,1,-nbitq), 
to_sfixed(396.0/65536.0,1,-nbitq), 
to_sfixed(1469.0/65536.0,1,-nbitq), 
to_sfixed(-1107.0/65536.0,1,-nbitq), 
to_sfixed(-781.0/65536.0,1,-nbitq), 
to_sfixed(1250.0/65536.0,1,-nbitq), 
to_sfixed(1123.0/65536.0,1,-nbitq), 
to_sfixed(-7207.0/65536.0,1,-nbitq), 
to_sfixed(-6125.0/65536.0,1,-nbitq), 
to_sfixed(-45.0/65536.0,1,-nbitq), 
to_sfixed(535.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3342.0/65536.0,1,-nbitq), 
to_sfixed(5518.0/65536.0,1,-nbitq), 
to_sfixed(-1618.0/65536.0,1,-nbitq), 
to_sfixed(3962.0/65536.0,1,-nbitq), 
to_sfixed(3613.0/65536.0,1,-nbitq), 
to_sfixed(3012.0/65536.0,1,-nbitq), 
to_sfixed(-8265.0/65536.0,1,-nbitq), 
to_sfixed(6777.0/65536.0,1,-nbitq), 
to_sfixed(2924.0/65536.0,1,-nbitq), 
to_sfixed(400.0/65536.0,1,-nbitq), 
to_sfixed(2734.0/65536.0,1,-nbitq), 
to_sfixed(1975.0/65536.0,1,-nbitq), 
to_sfixed(-2530.0/65536.0,1,-nbitq), 
to_sfixed(2578.0/65536.0,1,-nbitq), 
to_sfixed(2737.0/65536.0,1,-nbitq), 
to_sfixed(3886.0/65536.0,1,-nbitq), 
to_sfixed(-597.0/65536.0,1,-nbitq), 
to_sfixed(7975.0/65536.0,1,-nbitq), 
to_sfixed(-142.0/65536.0,1,-nbitq), 
to_sfixed(87.0/65536.0,1,-nbitq), 
to_sfixed(-3248.0/65536.0,1,-nbitq), 
to_sfixed(-6961.0/65536.0,1,-nbitq), 
to_sfixed(-2911.0/65536.0,1,-nbitq), 
to_sfixed(18728.0/65536.0,1,-nbitq), 
to_sfixed(-3813.0/65536.0,1,-nbitq), 
to_sfixed(-11815.0/65536.0,1,-nbitq), 
to_sfixed(-10927.0/65536.0,1,-nbitq), 
to_sfixed(1783.0/65536.0,1,-nbitq), 
to_sfixed(-1215.0/65536.0,1,-nbitq), 
to_sfixed(520.0/65536.0,1,-nbitq), 
to_sfixed(3923.0/65536.0,1,-nbitq), 
to_sfixed(4814.0/65536.0,1,-nbitq), 
to_sfixed(5178.0/65536.0,1,-nbitq), 
to_sfixed(-15922.0/65536.0,1,-nbitq), 
to_sfixed(-2489.0/65536.0,1,-nbitq), 
to_sfixed(2551.0/65536.0,1,-nbitq), 
to_sfixed(-3085.0/65536.0,1,-nbitq), 
to_sfixed(6339.0/65536.0,1,-nbitq), 
to_sfixed(614.0/65536.0,1,-nbitq), 
to_sfixed(-111.0/65536.0,1,-nbitq), 
to_sfixed(7094.0/65536.0,1,-nbitq), 
to_sfixed(1750.0/65536.0,1,-nbitq), 
to_sfixed(6263.0/65536.0,1,-nbitq), 
to_sfixed(7419.0/65536.0,1,-nbitq), 
to_sfixed(-2432.0/65536.0,1,-nbitq), 
to_sfixed(-11807.0/65536.0,1,-nbitq), 
to_sfixed(4562.0/65536.0,1,-nbitq), 
to_sfixed(3707.0/65536.0,1,-nbitq), 
to_sfixed(5340.0/65536.0,1,-nbitq), 
to_sfixed(3497.0/65536.0,1,-nbitq), 
to_sfixed(2654.0/65536.0,1,-nbitq), 
to_sfixed(-435.0/65536.0,1,-nbitq), 
to_sfixed(3976.0/65536.0,1,-nbitq), 
to_sfixed(5871.0/65536.0,1,-nbitq), 
to_sfixed(-4610.0/65536.0,1,-nbitq), 
to_sfixed(-3064.0/65536.0,1,-nbitq), 
to_sfixed(-2347.0/65536.0,1,-nbitq), 
to_sfixed(-3793.0/65536.0,1,-nbitq), 
to_sfixed(235.0/65536.0,1,-nbitq), 
to_sfixed(4138.0/65536.0,1,-nbitq), 
to_sfixed(16132.0/65536.0,1,-nbitq), 
to_sfixed(2712.0/65536.0,1,-nbitq), 
to_sfixed(-2212.0/65536.0,1,-nbitq), 
to_sfixed(-2454.0/65536.0,1,-nbitq), 
to_sfixed(12403.0/65536.0,1,-nbitq), 
to_sfixed(2700.0/65536.0,1,-nbitq), 
to_sfixed(-4310.0/65536.0,1,-nbitq), 
to_sfixed(7251.0/65536.0,1,-nbitq), 
to_sfixed(4052.0/65536.0,1,-nbitq), 
to_sfixed(6557.0/65536.0,1,-nbitq), 
to_sfixed(-3574.0/65536.0,1,-nbitq), 
to_sfixed(-4318.0/65536.0,1,-nbitq), 
to_sfixed(-5018.0/65536.0,1,-nbitq), 
to_sfixed(1975.0/65536.0,1,-nbitq), 
to_sfixed(618.0/65536.0,1,-nbitq), 
to_sfixed(5607.0/65536.0,1,-nbitq), 
to_sfixed(-7949.0/65536.0,1,-nbitq), 
to_sfixed(-12851.0/65536.0,1,-nbitq), 
to_sfixed(-1724.0/65536.0,1,-nbitq), 
to_sfixed(322.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1684.0/65536.0,1,-nbitq), 
to_sfixed(-2159.0/65536.0,1,-nbitq), 
to_sfixed(-1716.0/65536.0,1,-nbitq), 
to_sfixed(3441.0/65536.0,1,-nbitq), 
to_sfixed(951.0/65536.0,1,-nbitq), 
to_sfixed(3709.0/65536.0,1,-nbitq), 
to_sfixed(-4252.0/65536.0,1,-nbitq), 
to_sfixed(6823.0/65536.0,1,-nbitq), 
to_sfixed(-3416.0/65536.0,1,-nbitq), 
to_sfixed(1217.0/65536.0,1,-nbitq), 
to_sfixed(2246.0/65536.0,1,-nbitq), 
to_sfixed(-12364.0/65536.0,1,-nbitq), 
to_sfixed(-1676.0/65536.0,1,-nbitq), 
to_sfixed(-539.0/65536.0,1,-nbitq), 
to_sfixed(221.0/65536.0,1,-nbitq), 
to_sfixed(-871.0/65536.0,1,-nbitq), 
to_sfixed(-2164.0/65536.0,1,-nbitq), 
to_sfixed(16491.0/65536.0,1,-nbitq), 
to_sfixed(-873.0/65536.0,1,-nbitq), 
to_sfixed(2571.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(-15548.0/65536.0,1,-nbitq), 
to_sfixed(-7282.0/65536.0,1,-nbitq), 
to_sfixed(9213.0/65536.0,1,-nbitq), 
to_sfixed(-3146.0/65536.0,1,-nbitq), 
to_sfixed(2554.0/65536.0,1,-nbitq), 
to_sfixed(-7614.0/65536.0,1,-nbitq), 
to_sfixed(2975.0/65536.0,1,-nbitq), 
to_sfixed(6523.0/65536.0,1,-nbitq), 
to_sfixed(1776.0/65536.0,1,-nbitq), 
to_sfixed(1203.0/65536.0,1,-nbitq), 
to_sfixed(2671.0/65536.0,1,-nbitq), 
to_sfixed(5024.0/65536.0,1,-nbitq), 
to_sfixed(-7484.0/65536.0,1,-nbitq), 
to_sfixed(-265.0/65536.0,1,-nbitq), 
to_sfixed(2629.0/65536.0,1,-nbitq), 
to_sfixed(-3677.0/65536.0,1,-nbitq), 
to_sfixed(1267.0/65536.0,1,-nbitq), 
to_sfixed(-6458.0/65536.0,1,-nbitq), 
to_sfixed(-305.0/65536.0,1,-nbitq), 
to_sfixed(2296.0/65536.0,1,-nbitq), 
to_sfixed(2874.0/65536.0,1,-nbitq), 
to_sfixed(5513.0/65536.0,1,-nbitq), 
to_sfixed(5151.0/65536.0,1,-nbitq), 
to_sfixed(-1881.0/65536.0,1,-nbitq), 
to_sfixed(-10250.0/65536.0,1,-nbitq), 
to_sfixed(2047.0/65536.0,1,-nbitq), 
to_sfixed(3744.0/65536.0,1,-nbitq), 
to_sfixed(2893.0/65536.0,1,-nbitq), 
to_sfixed(-1570.0/65536.0,1,-nbitq), 
to_sfixed(583.0/65536.0,1,-nbitq), 
to_sfixed(-1725.0/65536.0,1,-nbitq), 
to_sfixed(1268.0/65536.0,1,-nbitq), 
to_sfixed(-2105.0/65536.0,1,-nbitq), 
to_sfixed(-5090.0/65536.0,1,-nbitq), 
to_sfixed(-6611.0/65536.0,1,-nbitq), 
to_sfixed(1481.0/65536.0,1,-nbitq), 
to_sfixed(1244.0/65536.0,1,-nbitq), 
to_sfixed(-341.0/65536.0,1,-nbitq), 
to_sfixed(8005.0/65536.0,1,-nbitq), 
to_sfixed(18230.0/65536.0,1,-nbitq), 
to_sfixed(-1883.0/65536.0,1,-nbitq), 
to_sfixed(9.0/65536.0,1,-nbitq), 
to_sfixed(2003.0/65536.0,1,-nbitq), 
to_sfixed(12493.0/65536.0,1,-nbitq), 
to_sfixed(11623.0/65536.0,1,-nbitq), 
to_sfixed(2434.0/65536.0,1,-nbitq), 
to_sfixed(6080.0/65536.0,1,-nbitq), 
to_sfixed(5496.0/65536.0,1,-nbitq), 
to_sfixed(7833.0/65536.0,1,-nbitq), 
to_sfixed(-3559.0/65536.0,1,-nbitq), 
to_sfixed(-1334.0/65536.0,1,-nbitq), 
to_sfixed(-2447.0/65536.0,1,-nbitq), 
to_sfixed(-868.0/65536.0,1,-nbitq), 
to_sfixed(-896.0/65536.0,1,-nbitq), 
to_sfixed(-1058.0/65536.0,1,-nbitq), 
to_sfixed(-6069.0/65536.0,1,-nbitq), 
to_sfixed(-10221.0/65536.0,1,-nbitq), 
to_sfixed(1403.0/65536.0,1,-nbitq), 
to_sfixed(-3596.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5144.0/65536.0,1,-nbitq), 
to_sfixed(-5389.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(-2779.0/65536.0,1,-nbitq), 
to_sfixed(-13035.0/65536.0,1,-nbitq), 
to_sfixed(1833.0/65536.0,1,-nbitq), 
to_sfixed(-6955.0/65536.0,1,-nbitq), 
to_sfixed(3092.0/65536.0,1,-nbitq), 
to_sfixed(3443.0/65536.0,1,-nbitq), 
to_sfixed(-2927.0/65536.0,1,-nbitq), 
to_sfixed(-1247.0/65536.0,1,-nbitq), 
to_sfixed(-5090.0/65536.0,1,-nbitq), 
to_sfixed(-1739.0/65536.0,1,-nbitq), 
to_sfixed(1857.0/65536.0,1,-nbitq), 
to_sfixed(439.0/65536.0,1,-nbitq), 
to_sfixed(871.0/65536.0,1,-nbitq), 
to_sfixed(847.0/65536.0,1,-nbitq), 
to_sfixed(17196.0/65536.0,1,-nbitq), 
to_sfixed(-3361.0/65536.0,1,-nbitq), 
to_sfixed(1871.0/65536.0,1,-nbitq), 
to_sfixed(-3661.0/65536.0,1,-nbitq), 
to_sfixed(-8256.0/65536.0,1,-nbitq), 
to_sfixed(-373.0/65536.0,1,-nbitq), 
to_sfixed(15423.0/65536.0,1,-nbitq), 
to_sfixed(1671.0/65536.0,1,-nbitq), 
to_sfixed(8859.0/65536.0,1,-nbitq), 
to_sfixed(-676.0/65536.0,1,-nbitq), 
to_sfixed(-536.0/65536.0,1,-nbitq), 
to_sfixed(4192.0/65536.0,1,-nbitq), 
to_sfixed(-365.0/65536.0,1,-nbitq), 
to_sfixed(-2001.0/65536.0,1,-nbitq), 
to_sfixed(-4067.0/65536.0,1,-nbitq), 
to_sfixed(4777.0/65536.0,1,-nbitq), 
to_sfixed(8189.0/65536.0,1,-nbitq), 
to_sfixed(-3087.0/65536.0,1,-nbitq), 
to_sfixed(3071.0/65536.0,1,-nbitq), 
to_sfixed(-2898.0/65536.0,1,-nbitq), 
to_sfixed(1039.0/65536.0,1,-nbitq), 
to_sfixed(-5070.0/65536.0,1,-nbitq), 
to_sfixed(-1775.0/65536.0,1,-nbitq), 
to_sfixed(-5103.0/65536.0,1,-nbitq), 
to_sfixed(-2590.0/65536.0,1,-nbitq), 
to_sfixed(-7839.0/65536.0,1,-nbitq), 
to_sfixed(6575.0/65536.0,1,-nbitq), 
to_sfixed(1554.0/65536.0,1,-nbitq), 
to_sfixed(-7699.0/65536.0,1,-nbitq), 
to_sfixed(-1561.0/65536.0,1,-nbitq), 
to_sfixed(4915.0/65536.0,1,-nbitq), 
to_sfixed(-43.0/65536.0,1,-nbitq), 
to_sfixed(2989.0/65536.0,1,-nbitq), 
to_sfixed(1136.0/65536.0,1,-nbitq), 
to_sfixed(-8110.0/65536.0,1,-nbitq), 
to_sfixed(-2454.0/65536.0,1,-nbitq), 
to_sfixed(-8783.0/65536.0,1,-nbitq), 
to_sfixed(-7817.0/65536.0,1,-nbitq), 
to_sfixed(-933.0/65536.0,1,-nbitq), 
to_sfixed(-3016.0/65536.0,1,-nbitq), 
to_sfixed(2421.0/65536.0,1,-nbitq), 
to_sfixed(2472.0/65536.0,1,-nbitq), 
to_sfixed(12280.0/65536.0,1,-nbitq), 
to_sfixed(6135.0/65536.0,1,-nbitq), 
to_sfixed(-1767.0/65536.0,1,-nbitq), 
to_sfixed(764.0/65536.0,1,-nbitq), 
to_sfixed(1777.0/65536.0,1,-nbitq), 
to_sfixed(11180.0/65536.0,1,-nbitq), 
to_sfixed(15159.0/65536.0,1,-nbitq), 
to_sfixed(-416.0/65536.0,1,-nbitq), 
to_sfixed(3749.0/65536.0,1,-nbitq), 
to_sfixed(2680.0/65536.0,1,-nbitq), 
to_sfixed(7944.0/65536.0,1,-nbitq), 
to_sfixed(-3647.0/65536.0,1,-nbitq), 
to_sfixed(-8170.0/65536.0,1,-nbitq), 
to_sfixed(-7543.0/65536.0,1,-nbitq), 
to_sfixed(1144.0/65536.0,1,-nbitq), 
to_sfixed(-721.0/65536.0,1,-nbitq), 
to_sfixed(-6182.0/65536.0,1,-nbitq), 
to_sfixed(-80.0/65536.0,1,-nbitq), 
to_sfixed(-477.0/65536.0,1,-nbitq), 
to_sfixed(-3028.0/65536.0,1,-nbitq), 
to_sfixed(-5436.0/65536.0,1,-nbitq)  ), 
( to_sfixed(207.0/65536.0,1,-nbitq), 
to_sfixed(-8916.0/65536.0,1,-nbitq), 
to_sfixed(-405.0/65536.0,1,-nbitq), 
to_sfixed(-6455.0/65536.0,1,-nbitq), 
to_sfixed(-13446.0/65536.0,1,-nbitq), 
to_sfixed(-1217.0/65536.0,1,-nbitq), 
to_sfixed(-1796.0/65536.0,1,-nbitq), 
to_sfixed(6018.0/65536.0,1,-nbitq), 
to_sfixed(-1540.0/65536.0,1,-nbitq), 
to_sfixed(-250.0/65536.0,1,-nbitq), 
to_sfixed(-19.0/65536.0,1,-nbitq), 
to_sfixed(-6709.0/65536.0,1,-nbitq), 
to_sfixed(4725.0/65536.0,1,-nbitq), 
to_sfixed(-672.0/65536.0,1,-nbitq), 
to_sfixed(-4071.0/65536.0,1,-nbitq), 
to_sfixed(2651.0/65536.0,1,-nbitq), 
to_sfixed(218.0/65536.0,1,-nbitq), 
to_sfixed(-15584.0/65536.0,1,-nbitq), 
to_sfixed(4734.0/65536.0,1,-nbitq), 
to_sfixed(1993.0/65536.0,1,-nbitq), 
to_sfixed(-11148.0/65536.0,1,-nbitq), 
to_sfixed(1578.0/65536.0,1,-nbitq), 
to_sfixed(-621.0/65536.0,1,-nbitq), 
to_sfixed(6286.0/65536.0,1,-nbitq), 
to_sfixed(3741.0/65536.0,1,-nbitq), 
to_sfixed(4168.0/65536.0,1,-nbitq), 
to_sfixed(-899.0/65536.0,1,-nbitq), 
to_sfixed(-1802.0/65536.0,1,-nbitq), 
to_sfixed(10747.0/65536.0,1,-nbitq), 
to_sfixed(-528.0/65536.0,1,-nbitq), 
to_sfixed(-3542.0/65536.0,1,-nbitq), 
to_sfixed(-9109.0/65536.0,1,-nbitq), 
to_sfixed(7236.0/65536.0,1,-nbitq), 
to_sfixed(15432.0/65536.0,1,-nbitq), 
to_sfixed(2040.0/65536.0,1,-nbitq), 
to_sfixed(2067.0/65536.0,1,-nbitq), 
to_sfixed(-6369.0/65536.0,1,-nbitq), 
to_sfixed(1037.0/65536.0,1,-nbitq), 
to_sfixed(-8996.0/65536.0,1,-nbitq), 
to_sfixed(-3407.0/65536.0,1,-nbitq), 
to_sfixed(-2658.0/65536.0,1,-nbitq), 
to_sfixed(901.0/65536.0,1,-nbitq), 
to_sfixed(-12689.0/65536.0,1,-nbitq), 
to_sfixed(4539.0/65536.0,1,-nbitq), 
to_sfixed(2009.0/65536.0,1,-nbitq), 
to_sfixed(-1004.0/65536.0,1,-nbitq), 
to_sfixed(-2376.0/65536.0,1,-nbitq), 
to_sfixed(4098.0/65536.0,1,-nbitq), 
to_sfixed(2848.0/65536.0,1,-nbitq), 
to_sfixed(-1134.0/65536.0,1,-nbitq), 
to_sfixed(2254.0/65536.0,1,-nbitq), 
to_sfixed(-9766.0/65536.0,1,-nbitq), 
to_sfixed(7423.0/65536.0,1,-nbitq), 
to_sfixed(-14696.0/65536.0,1,-nbitq), 
to_sfixed(-4081.0/65536.0,1,-nbitq), 
to_sfixed(-5546.0/65536.0,1,-nbitq), 
to_sfixed(-2149.0/65536.0,1,-nbitq), 
to_sfixed(-762.0/65536.0,1,-nbitq), 
to_sfixed(-1361.0/65536.0,1,-nbitq), 
to_sfixed(15466.0/65536.0,1,-nbitq), 
to_sfixed(-10019.0/65536.0,1,-nbitq), 
to_sfixed(1742.0/65536.0,1,-nbitq), 
to_sfixed(403.0/65536.0,1,-nbitq), 
to_sfixed(-2182.0/65536.0,1,-nbitq), 
to_sfixed(9284.0/65536.0,1,-nbitq), 
to_sfixed(-18372.0/65536.0,1,-nbitq), 
to_sfixed(-757.0/65536.0,1,-nbitq), 
to_sfixed(8618.0/65536.0,1,-nbitq), 
to_sfixed(4169.0/65536.0,1,-nbitq), 
to_sfixed(11243.0/65536.0,1,-nbitq), 
to_sfixed(-6055.0/65536.0,1,-nbitq), 
to_sfixed(-2607.0/65536.0,1,-nbitq), 
to_sfixed(-8353.0/65536.0,1,-nbitq), 
to_sfixed(-2233.0/65536.0,1,-nbitq), 
to_sfixed(-1003.0/65536.0,1,-nbitq), 
to_sfixed(-14376.0/65536.0,1,-nbitq), 
to_sfixed(-26.0/65536.0,1,-nbitq), 
to_sfixed(11504.0/65536.0,1,-nbitq), 
to_sfixed(3.0/65536.0,1,-nbitq), 
to_sfixed(-7763.0/65536.0,1,-nbitq)  ), 
( to_sfixed(370.0/65536.0,1,-nbitq), 
to_sfixed(-5078.0/65536.0,1,-nbitq), 
to_sfixed(-8649.0/65536.0,1,-nbitq), 
to_sfixed(-12103.0/65536.0,1,-nbitq), 
to_sfixed(-3609.0/65536.0,1,-nbitq), 
to_sfixed(2959.0/65536.0,1,-nbitq), 
to_sfixed(-3522.0/65536.0,1,-nbitq), 
to_sfixed(4611.0/65536.0,1,-nbitq), 
to_sfixed(-1431.0/65536.0,1,-nbitq), 
to_sfixed(-1502.0/65536.0,1,-nbitq), 
to_sfixed(-4743.0/65536.0,1,-nbitq), 
to_sfixed(-8454.0/65536.0,1,-nbitq), 
to_sfixed(6748.0/65536.0,1,-nbitq), 
to_sfixed(-3197.0/65536.0,1,-nbitq), 
to_sfixed(-7331.0/65536.0,1,-nbitq), 
to_sfixed(2863.0/65536.0,1,-nbitq), 
to_sfixed(2341.0/65536.0,1,-nbitq), 
to_sfixed(-12498.0/65536.0,1,-nbitq), 
to_sfixed(2305.0/65536.0,1,-nbitq), 
to_sfixed(860.0/65536.0,1,-nbitq), 
to_sfixed(-5147.0/65536.0,1,-nbitq), 
to_sfixed(2106.0/65536.0,1,-nbitq), 
to_sfixed(-13045.0/65536.0,1,-nbitq), 
to_sfixed(4948.0/65536.0,1,-nbitq), 
to_sfixed(7322.0/65536.0,1,-nbitq), 
to_sfixed(12716.0/65536.0,1,-nbitq), 
to_sfixed(-3195.0/65536.0,1,-nbitq), 
to_sfixed(-276.0/65536.0,1,-nbitq), 
to_sfixed(12559.0/65536.0,1,-nbitq), 
to_sfixed(-1774.0/65536.0,1,-nbitq), 
to_sfixed(-763.0/65536.0,1,-nbitq), 
to_sfixed(-6035.0/65536.0,1,-nbitq), 
to_sfixed(9851.0/65536.0,1,-nbitq), 
to_sfixed(13270.0/65536.0,1,-nbitq), 
to_sfixed(-599.0/65536.0,1,-nbitq), 
to_sfixed(3691.0/65536.0,1,-nbitq), 
to_sfixed(-7533.0/65536.0,1,-nbitq), 
to_sfixed(3034.0/65536.0,1,-nbitq), 
to_sfixed(-4276.0/65536.0,1,-nbitq), 
to_sfixed(-4459.0/65536.0,1,-nbitq), 
to_sfixed(4248.0/65536.0,1,-nbitq), 
to_sfixed(-761.0/65536.0,1,-nbitq), 
to_sfixed(-1221.0/65536.0,1,-nbitq), 
to_sfixed(11.0/65536.0,1,-nbitq), 
to_sfixed(-894.0/65536.0,1,-nbitq), 
to_sfixed(2433.0/65536.0,1,-nbitq), 
to_sfixed(-1992.0/65536.0,1,-nbitq), 
to_sfixed(-1223.0/65536.0,1,-nbitq), 
to_sfixed(3491.0/65536.0,1,-nbitq), 
to_sfixed(-794.0/65536.0,1,-nbitq), 
to_sfixed(1271.0/65536.0,1,-nbitq), 
to_sfixed(-6354.0/65536.0,1,-nbitq), 
to_sfixed(5479.0/65536.0,1,-nbitq), 
to_sfixed(-15464.0/65536.0,1,-nbitq), 
to_sfixed(-5255.0/65536.0,1,-nbitq), 
to_sfixed(1018.0/65536.0,1,-nbitq), 
to_sfixed(-3055.0/65536.0,1,-nbitq), 
to_sfixed(5856.0/65536.0,1,-nbitq), 
to_sfixed(-1707.0/65536.0,1,-nbitq), 
to_sfixed(21342.0/65536.0,1,-nbitq), 
to_sfixed(-19469.0/65536.0,1,-nbitq), 
to_sfixed(-1921.0/65536.0,1,-nbitq), 
to_sfixed(-2878.0/65536.0,1,-nbitq), 
to_sfixed(-63.0/65536.0,1,-nbitq), 
to_sfixed(8753.0/65536.0,1,-nbitq), 
to_sfixed(-20294.0/65536.0,1,-nbitq), 
to_sfixed(-5639.0/65536.0,1,-nbitq), 
to_sfixed(6750.0/65536.0,1,-nbitq), 
to_sfixed(4932.0/65536.0,1,-nbitq), 
to_sfixed(4003.0/65536.0,1,-nbitq), 
to_sfixed(-9502.0/65536.0,1,-nbitq), 
to_sfixed(-9471.0/65536.0,1,-nbitq), 
to_sfixed(-8218.0/65536.0,1,-nbitq), 
to_sfixed(2239.0/65536.0,1,-nbitq), 
to_sfixed(-2797.0/65536.0,1,-nbitq), 
to_sfixed(-17451.0/65536.0,1,-nbitq), 
to_sfixed(2136.0/65536.0,1,-nbitq), 
to_sfixed(6051.0/65536.0,1,-nbitq), 
to_sfixed(-505.0/65536.0,1,-nbitq), 
to_sfixed(-547.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-563.0/65536.0,1,-nbitq), 
to_sfixed(-5949.0/65536.0,1,-nbitq), 
to_sfixed(-12025.0/65536.0,1,-nbitq), 
to_sfixed(-13625.0/65536.0,1,-nbitq), 
to_sfixed(-3025.0/65536.0,1,-nbitq), 
to_sfixed(1538.0/65536.0,1,-nbitq), 
to_sfixed(-2358.0/65536.0,1,-nbitq), 
to_sfixed(-7363.0/65536.0,1,-nbitq), 
to_sfixed(-928.0/65536.0,1,-nbitq), 
to_sfixed(224.0/65536.0,1,-nbitq), 
to_sfixed(-4504.0/65536.0,1,-nbitq), 
to_sfixed(493.0/65536.0,1,-nbitq), 
to_sfixed(2828.0/65536.0,1,-nbitq), 
to_sfixed(-1629.0/65536.0,1,-nbitq), 
to_sfixed(-4816.0/65536.0,1,-nbitq), 
to_sfixed(431.0/65536.0,1,-nbitq), 
to_sfixed(2725.0/65536.0,1,-nbitq), 
to_sfixed(-1297.0/65536.0,1,-nbitq), 
to_sfixed(5194.0/65536.0,1,-nbitq), 
to_sfixed(2393.0/65536.0,1,-nbitq), 
to_sfixed(-3263.0/65536.0,1,-nbitq), 
to_sfixed(3598.0/65536.0,1,-nbitq), 
to_sfixed(-9045.0/65536.0,1,-nbitq), 
to_sfixed(4732.0/65536.0,1,-nbitq), 
to_sfixed(12649.0/65536.0,1,-nbitq), 
to_sfixed(3491.0/65536.0,1,-nbitq), 
to_sfixed(-1236.0/65536.0,1,-nbitq), 
to_sfixed(1647.0/65536.0,1,-nbitq), 
to_sfixed(8744.0/65536.0,1,-nbitq), 
to_sfixed(-470.0/65536.0,1,-nbitq), 
to_sfixed(5413.0/65536.0,1,-nbitq), 
to_sfixed(2093.0/65536.0,1,-nbitq), 
to_sfixed(-4500.0/65536.0,1,-nbitq), 
to_sfixed(3894.0/65536.0,1,-nbitq), 
to_sfixed(-906.0/65536.0,1,-nbitq), 
to_sfixed(2320.0/65536.0,1,-nbitq), 
to_sfixed(-8636.0/65536.0,1,-nbitq), 
to_sfixed(6370.0/65536.0,1,-nbitq), 
to_sfixed(21869.0/65536.0,1,-nbitq), 
to_sfixed(284.0/65536.0,1,-nbitq), 
to_sfixed(8128.0/65536.0,1,-nbitq), 
to_sfixed(-1697.0/65536.0,1,-nbitq), 
to_sfixed(-154.0/65536.0,1,-nbitq), 
to_sfixed(472.0/65536.0,1,-nbitq), 
to_sfixed(-2610.0/65536.0,1,-nbitq), 
to_sfixed(4723.0/65536.0,1,-nbitq), 
to_sfixed(-985.0/65536.0,1,-nbitq), 
to_sfixed(-3455.0/65536.0,1,-nbitq), 
to_sfixed(-10.0/65536.0,1,-nbitq), 
to_sfixed(-911.0/65536.0,1,-nbitq), 
to_sfixed(2413.0/65536.0,1,-nbitq), 
to_sfixed(-3889.0/65536.0,1,-nbitq), 
to_sfixed(9619.0/65536.0,1,-nbitq), 
to_sfixed(-10634.0/65536.0,1,-nbitq), 
to_sfixed(1468.0/65536.0,1,-nbitq), 
to_sfixed(-10059.0/65536.0,1,-nbitq), 
to_sfixed(919.0/65536.0,1,-nbitq), 
to_sfixed(5276.0/65536.0,1,-nbitq), 
to_sfixed(-2407.0/65536.0,1,-nbitq), 
to_sfixed(10561.0/65536.0,1,-nbitq), 
to_sfixed(-11071.0/65536.0,1,-nbitq), 
to_sfixed(2112.0/65536.0,1,-nbitq), 
to_sfixed(-2531.0/65536.0,1,-nbitq), 
to_sfixed(340.0/65536.0,1,-nbitq), 
to_sfixed(-735.0/65536.0,1,-nbitq), 
to_sfixed(-13013.0/65536.0,1,-nbitq), 
to_sfixed(-6455.0/65536.0,1,-nbitq), 
to_sfixed(-4291.0/65536.0,1,-nbitq), 
to_sfixed(-4400.0/65536.0,1,-nbitq), 
to_sfixed(104.0/65536.0,1,-nbitq), 
to_sfixed(-3525.0/65536.0,1,-nbitq), 
to_sfixed(-4139.0/65536.0,1,-nbitq), 
to_sfixed(-15144.0/65536.0,1,-nbitq), 
to_sfixed(2389.0/65536.0,1,-nbitq), 
to_sfixed(2590.0/65536.0,1,-nbitq), 
to_sfixed(-16957.0/65536.0,1,-nbitq), 
to_sfixed(-128.0/65536.0,1,-nbitq), 
to_sfixed(2134.0/65536.0,1,-nbitq), 
to_sfixed(-292.0/65536.0,1,-nbitq), 
to_sfixed(2341.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-928.0/65536.0,1,-nbitq), 
to_sfixed(-4666.0/65536.0,1,-nbitq), 
to_sfixed(-4283.0/65536.0,1,-nbitq), 
to_sfixed(-8532.0/65536.0,1,-nbitq), 
to_sfixed(-979.0/65536.0,1,-nbitq), 
to_sfixed(4574.0/65536.0,1,-nbitq), 
to_sfixed(-916.0/65536.0,1,-nbitq), 
to_sfixed(-9445.0/65536.0,1,-nbitq), 
to_sfixed(4413.0/65536.0,1,-nbitq), 
to_sfixed(1094.0/65536.0,1,-nbitq), 
to_sfixed(-5266.0/65536.0,1,-nbitq), 
to_sfixed(15399.0/65536.0,1,-nbitq), 
to_sfixed(4273.0/65536.0,1,-nbitq), 
to_sfixed(6160.0/65536.0,1,-nbitq), 
to_sfixed(-934.0/65536.0,1,-nbitq), 
to_sfixed(-1430.0/65536.0,1,-nbitq), 
to_sfixed(75.0/65536.0,1,-nbitq), 
to_sfixed(4573.0/65536.0,1,-nbitq), 
to_sfixed(5151.0/65536.0,1,-nbitq), 
to_sfixed(-118.0/65536.0,1,-nbitq), 
to_sfixed(26.0/65536.0,1,-nbitq), 
to_sfixed(7299.0/65536.0,1,-nbitq), 
to_sfixed(-4836.0/65536.0,1,-nbitq), 
to_sfixed(2048.0/65536.0,1,-nbitq), 
to_sfixed(8413.0/65536.0,1,-nbitq), 
to_sfixed(-5191.0/65536.0,1,-nbitq), 
to_sfixed(4955.0/65536.0,1,-nbitq), 
to_sfixed(-2211.0/65536.0,1,-nbitq), 
to_sfixed(9662.0/65536.0,1,-nbitq), 
to_sfixed(-6246.0/65536.0,1,-nbitq), 
to_sfixed(8822.0/65536.0,1,-nbitq), 
to_sfixed(8414.0/65536.0,1,-nbitq), 
to_sfixed(1702.0/65536.0,1,-nbitq), 
to_sfixed(-14906.0/65536.0,1,-nbitq), 
to_sfixed(-1283.0/65536.0,1,-nbitq), 
to_sfixed(-1143.0/65536.0,1,-nbitq), 
to_sfixed(-18634.0/65536.0,1,-nbitq), 
to_sfixed(11331.0/65536.0,1,-nbitq), 
to_sfixed(4714.0/65536.0,1,-nbitq), 
to_sfixed(-1551.0/65536.0,1,-nbitq), 
to_sfixed(15276.0/65536.0,1,-nbitq), 
to_sfixed(297.0/65536.0,1,-nbitq), 
to_sfixed(-317.0/65536.0,1,-nbitq), 
to_sfixed(4504.0/65536.0,1,-nbitq), 
to_sfixed(292.0/65536.0,1,-nbitq), 
to_sfixed(5438.0/65536.0,1,-nbitq), 
to_sfixed(-2570.0/65536.0,1,-nbitq), 
to_sfixed(-81.0/65536.0,1,-nbitq), 
to_sfixed(-3043.0/65536.0,1,-nbitq), 
to_sfixed(-913.0/65536.0,1,-nbitq), 
to_sfixed(382.0/65536.0,1,-nbitq), 
to_sfixed(-4701.0/65536.0,1,-nbitq), 
to_sfixed(5665.0/65536.0,1,-nbitq), 
to_sfixed(-5232.0/65536.0,1,-nbitq), 
to_sfixed(7098.0/65536.0,1,-nbitq), 
to_sfixed(-15159.0/65536.0,1,-nbitq), 
to_sfixed(887.0/65536.0,1,-nbitq), 
to_sfixed(177.0/65536.0,1,-nbitq), 
to_sfixed(1920.0/65536.0,1,-nbitq), 
to_sfixed(1627.0/65536.0,1,-nbitq), 
to_sfixed(-4094.0/65536.0,1,-nbitq), 
to_sfixed(-913.0/65536.0,1,-nbitq), 
to_sfixed(2480.0/65536.0,1,-nbitq), 
to_sfixed(-542.0/65536.0,1,-nbitq), 
to_sfixed(-10024.0/65536.0,1,-nbitq), 
to_sfixed(-12551.0/65536.0,1,-nbitq), 
to_sfixed(-4143.0/65536.0,1,-nbitq), 
to_sfixed(-1880.0/65536.0,1,-nbitq), 
to_sfixed(-1553.0/65536.0,1,-nbitq), 
to_sfixed(-2292.0/65536.0,1,-nbitq), 
to_sfixed(1979.0/65536.0,1,-nbitq), 
to_sfixed(-10138.0/65536.0,1,-nbitq), 
to_sfixed(-15499.0/65536.0,1,-nbitq), 
to_sfixed(2000.0/65536.0,1,-nbitq), 
to_sfixed(1580.0/65536.0,1,-nbitq), 
to_sfixed(5350.0/65536.0,1,-nbitq), 
to_sfixed(-6416.0/65536.0,1,-nbitq), 
to_sfixed(-1595.0/65536.0,1,-nbitq), 
to_sfixed(-1427.0/65536.0,1,-nbitq), 
to_sfixed(9234.0/65536.0,1,-nbitq)  ), 
( to_sfixed(550.0/65536.0,1,-nbitq), 
to_sfixed(184.0/65536.0,1,-nbitq), 
to_sfixed(-3153.0/65536.0,1,-nbitq), 
to_sfixed(-4706.0/65536.0,1,-nbitq), 
to_sfixed(-3421.0/65536.0,1,-nbitq), 
to_sfixed(4749.0/65536.0,1,-nbitq), 
to_sfixed(2034.0/65536.0,1,-nbitq), 
to_sfixed(1076.0/65536.0,1,-nbitq), 
to_sfixed(-5038.0/65536.0,1,-nbitq), 
to_sfixed(-2652.0/65536.0,1,-nbitq), 
to_sfixed(-3158.0/65536.0,1,-nbitq), 
to_sfixed(9093.0/65536.0,1,-nbitq), 
to_sfixed(4127.0/65536.0,1,-nbitq), 
to_sfixed(11277.0/65536.0,1,-nbitq), 
to_sfixed(1040.0/65536.0,1,-nbitq), 
to_sfixed(1327.0/65536.0,1,-nbitq), 
to_sfixed(-945.0/65536.0,1,-nbitq), 
to_sfixed(2653.0/65536.0,1,-nbitq), 
to_sfixed(3829.0/65536.0,1,-nbitq), 
to_sfixed(-1420.0/65536.0,1,-nbitq), 
to_sfixed(-506.0/65536.0,1,-nbitq), 
to_sfixed(2654.0/65536.0,1,-nbitq), 
to_sfixed(-4110.0/65536.0,1,-nbitq), 
to_sfixed(-2587.0/65536.0,1,-nbitq), 
to_sfixed(2311.0/65536.0,1,-nbitq), 
to_sfixed(-8171.0/65536.0,1,-nbitq), 
to_sfixed(1901.0/65536.0,1,-nbitq), 
to_sfixed(2575.0/65536.0,1,-nbitq), 
to_sfixed(6024.0/65536.0,1,-nbitq), 
to_sfixed(547.0/65536.0,1,-nbitq), 
to_sfixed(2826.0/65536.0,1,-nbitq), 
to_sfixed(13950.0/65536.0,1,-nbitq), 
to_sfixed(-312.0/65536.0,1,-nbitq), 
to_sfixed(-13966.0/65536.0,1,-nbitq), 
to_sfixed(2138.0/65536.0,1,-nbitq), 
to_sfixed(-2058.0/65536.0,1,-nbitq), 
to_sfixed(-9851.0/65536.0,1,-nbitq), 
to_sfixed(7519.0/65536.0,1,-nbitq), 
to_sfixed(-1839.0/65536.0,1,-nbitq), 
to_sfixed(615.0/65536.0,1,-nbitq), 
to_sfixed(16397.0/65536.0,1,-nbitq), 
to_sfixed(2339.0/65536.0,1,-nbitq), 
to_sfixed(-2010.0/65536.0,1,-nbitq), 
to_sfixed(9163.0/65536.0,1,-nbitq), 
to_sfixed(-1447.0/65536.0,1,-nbitq), 
to_sfixed(2239.0/65536.0,1,-nbitq), 
to_sfixed(-2600.0/65536.0,1,-nbitq), 
to_sfixed(291.0/65536.0,1,-nbitq), 
to_sfixed(1095.0/65536.0,1,-nbitq), 
to_sfixed(19.0/65536.0,1,-nbitq), 
to_sfixed(-1018.0/65536.0,1,-nbitq), 
to_sfixed(-6227.0/65536.0,1,-nbitq), 
to_sfixed(3465.0/65536.0,1,-nbitq), 
to_sfixed(6294.0/65536.0,1,-nbitq), 
to_sfixed(15046.0/65536.0,1,-nbitq), 
to_sfixed(-16089.0/65536.0,1,-nbitq), 
to_sfixed(-1744.0/65536.0,1,-nbitq), 
to_sfixed(-2787.0/65536.0,1,-nbitq), 
to_sfixed(-3555.0/65536.0,1,-nbitq), 
to_sfixed(-3462.0/65536.0,1,-nbitq), 
to_sfixed(-7100.0/65536.0,1,-nbitq), 
to_sfixed(-1165.0/65536.0,1,-nbitq), 
to_sfixed(498.0/65536.0,1,-nbitq), 
to_sfixed(-2450.0/65536.0,1,-nbitq), 
to_sfixed(-6680.0/65536.0,1,-nbitq), 
to_sfixed(-8725.0/65536.0,1,-nbitq), 
to_sfixed(1599.0/65536.0,1,-nbitq), 
to_sfixed(-4479.0/65536.0,1,-nbitq), 
to_sfixed(7284.0/65536.0,1,-nbitq), 
to_sfixed(-1324.0/65536.0,1,-nbitq), 
to_sfixed(54.0/65536.0,1,-nbitq), 
to_sfixed(1533.0/65536.0,1,-nbitq), 
to_sfixed(7911.0/65536.0,1,-nbitq), 
to_sfixed(-456.0/65536.0,1,-nbitq), 
to_sfixed(-1864.0/65536.0,1,-nbitq), 
to_sfixed(12077.0/65536.0,1,-nbitq), 
to_sfixed(-2138.0/65536.0,1,-nbitq), 
to_sfixed(-4528.0/65536.0,1,-nbitq), 
to_sfixed(1134.0/65536.0,1,-nbitq), 
to_sfixed(8664.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4011.0/65536.0,1,-nbitq), 
to_sfixed(1970.0/65536.0,1,-nbitq), 
to_sfixed(-3161.0/65536.0,1,-nbitq), 
to_sfixed(559.0/65536.0,1,-nbitq), 
to_sfixed(-4762.0/65536.0,1,-nbitq), 
to_sfixed(7684.0/65536.0,1,-nbitq), 
to_sfixed(3793.0/65536.0,1,-nbitq), 
to_sfixed(4981.0/65536.0,1,-nbitq), 
to_sfixed(-4084.0/65536.0,1,-nbitq), 
to_sfixed(2325.0/65536.0,1,-nbitq), 
to_sfixed(-1022.0/65536.0,1,-nbitq), 
to_sfixed(-787.0/65536.0,1,-nbitq), 
to_sfixed(434.0/65536.0,1,-nbitq), 
to_sfixed(7218.0/65536.0,1,-nbitq), 
to_sfixed(-65.0/65536.0,1,-nbitq), 
to_sfixed(-773.0/65536.0,1,-nbitq), 
to_sfixed(2536.0/65536.0,1,-nbitq), 
to_sfixed(-4830.0/65536.0,1,-nbitq), 
to_sfixed(4479.0/65536.0,1,-nbitq), 
to_sfixed(-296.0/65536.0,1,-nbitq), 
to_sfixed(-3865.0/65536.0,1,-nbitq), 
to_sfixed(6891.0/65536.0,1,-nbitq), 
to_sfixed(-1579.0/65536.0,1,-nbitq), 
to_sfixed(-6823.0/65536.0,1,-nbitq), 
to_sfixed(-873.0/65536.0,1,-nbitq), 
to_sfixed(-10721.0/65536.0,1,-nbitq), 
to_sfixed(-5516.0/65536.0,1,-nbitq), 
to_sfixed(595.0/65536.0,1,-nbitq), 
to_sfixed(3295.0/65536.0,1,-nbitq), 
to_sfixed(4520.0/65536.0,1,-nbitq), 
to_sfixed(-374.0/65536.0,1,-nbitq), 
to_sfixed(10183.0/65536.0,1,-nbitq), 
to_sfixed(-450.0/65536.0,1,-nbitq), 
to_sfixed(-11911.0/65536.0,1,-nbitq), 
to_sfixed(-3236.0/65536.0,1,-nbitq), 
to_sfixed(-2449.0/65536.0,1,-nbitq), 
to_sfixed(-4607.0/65536.0,1,-nbitq), 
to_sfixed(7865.0/65536.0,1,-nbitq), 
to_sfixed(-5525.0/65536.0,1,-nbitq), 
to_sfixed(-2635.0/65536.0,1,-nbitq), 
to_sfixed(8215.0/65536.0,1,-nbitq), 
to_sfixed(2077.0/65536.0,1,-nbitq), 
to_sfixed(5641.0/65536.0,1,-nbitq), 
to_sfixed(7395.0/65536.0,1,-nbitq), 
to_sfixed(2403.0/65536.0,1,-nbitq), 
to_sfixed(-8603.0/65536.0,1,-nbitq), 
to_sfixed(1789.0/65536.0,1,-nbitq), 
to_sfixed(-204.0/65536.0,1,-nbitq), 
to_sfixed(1771.0/65536.0,1,-nbitq), 
to_sfixed(-46.0/65536.0,1,-nbitq), 
to_sfixed(2303.0/65536.0,1,-nbitq), 
to_sfixed(-1606.0/65536.0,1,-nbitq), 
to_sfixed(6325.0/65536.0,1,-nbitq), 
to_sfixed(1885.0/65536.0,1,-nbitq), 
to_sfixed(4202.0/65536.0,1,-nbitq), 
to_sfixed(-11711.0/65536.0,1,-nbitq), 
to_sfixed(1736.0/65536.0,1,-nbitq), 
to_sfixed(-5123.0/65536.0,1,-nbitq), 
to_sfixed(1602.0/65536.0,1,-nbitq), 
to_sfixed(-7292.0/65536.0,1,-nbitq), 
to_sfixed(3306.0/65536.0,1,-nbitq), 
to_sfixed(1264.0/65536.0,1,-nbitq), 
to_sfixed(-2443.0/65536.0,1,-nbitq), 
to_sfixed(-101.0/65536.0,1,-nbitq), 
to_sfixed(-4721.0/65536.0,1,-nbitq), 
to_sfixed(-13015.0/65536.0,1,-nbitq), 
to_sfixed(-796.0/65536.0,1,-nbitq), 
to_sfixed(-5703.0/65536.0,1,-nbitq), 
to_sfixed(8397.0/65536.0,1,-nbitq), 
to_sfixed(163.0/65536.0,1,-nbitq), 
to_sfixed(-1036.0/65536.0,1,-nbitq), 
to_sfixed(937.0/65536.0,1,-nbitq), 
to_sfixed(8510.0/65536.0,1,-nbitq), 
to_sfixed(-968.0/65536.0,1,-nbitq), 
to_sfixed(1574.0/65536.0,1,-nbitq), 
to_sfixed(-162.0/65536.0,1,-nbitq), 
to_sfixed(-8071.0/65536.0,1,-nbitq), 
to_sfixed(-10168.0/65536.0,1,-nbitq), 
to_sfixed(1740.0/65536.0,1,-nbitq), 
to_sfixed(2131.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2082.0/65536.0,1,-nbitq), 
to_sfixed(1976.0/65536.0,1,-nbitq), 
to_sfixed(-2644.0/65536.0,1,-nbitq), 
to_sfixed(5152.0/65536.0,1,-nbitq), 
to_sfixed(-4792.0/65536.0,1,-nbitq), 
to_sfixed(9544.0/65536.0,1,-nbitq), 
to_sfixed(-1264.0/65536.0,1,-nbitq), 
to_sfixed(-6418.0/65536.0,1,-nbitq), 
to_sfixed(1806.0/65536.0,1,-nbitq), 
to_sfixed(1307.0/65536.0,1,-nbitq), 
to_sfixed(862.0/65536.0,1,-nbitq), 
to_sfixed(-4581.0/65536.0,1,-nbitq), 
to_sfixed(2238.0/65536.0,1,-nbitq), 
to_sfixed(7532.0/65536.0,1,-nbitq), 
to_sfixed(3591.0/65536.0,1,-nbitq), 
to_sfixed(-2882.0/65536.0,1,-nbitq), 
to_sfixed(-1838.0/65536.0,1,-nbitq), 
to_sfixed(-1329.0/65536.0,1,-nbitq), 
to_sfixed(-1920.0/65536.0,1,-nbitq), 
to_sfixed(2001.0/65536.0,1,-nbitq), 
to_sfixed(-822.0/65536.0,1,-nbitq), 
to_sfixed(11514.0/65536.0,1,-nbitq), 
to_sfixed(2434.0/65536.0,1,-nbitq), 
to_sfixed(-2307.0/65536.0,1,-nbitq), 
to_sfixed(1063.0/65536.0,1,-nbitq), 
to_sfixed(-4755.0/65536.0,1,-nbitq), 
to_sfixed(-4990.0/65536.0,1,-nbitq), 
to_sfixed(1577.0/65536.0,1,-nbitq), 
to_sfixed(14856.0/65536.0,1,-nbitq), 
to_sfixed(1221.0/65536.0,1,-nbitq), 
to_sfixed(-4546.0/65536.0,1,-nbitq), 
to_sfixed(3075.0/65536.0,1,-nbitq), 
to_sfixed(-4970.0/65536.0,1,-nbitq), 
to_sfixed(-12634.0/65536.0,1,-nbitq), 
to_sfixed(-2465.0/65536.0,1,-nbitq), 
to_sfixed(1627.0/65536.0,1,-nbitq), 
to_sfixed(-4872.0/65536.0,1,-nbitq), 
to_sfixed(1878.0/65536.0,1,-nbitq), 
to_sfixed(-9488.0/65536.0,1,-nbitq), 
to_sfixed(-675.0/65536.0,1,-nbitq), 
to_sfixed(4349.0/65536.0,1,-nbitq), 
to_sfixed(-1359.0/65536.0,1,-nbitq), 
to_sfixed(2514.0/65536.0,1,-nbitq), 
to_sfixed(7659.0/65536.0,1,-nbitq), 
to_sfixed(1405.0/65536.0,1,-nbitq), 
to_sfixed(-10319.0/65536.0,1,-nbitq), 
to_sfixed(-3049.0/65536.0,1,-nbitq), 
to_sfixed(6435.0/65536.0,1,-nbitq), 
to_sfixed(1382.0/65536.0,1,-nbitq), 
to_sfixed(-2553.0/65536.0,1,-nbitq), 
to_sfixed(-1592.0/65536.0,1,-nbitq), 
to_sfixed(-1969.0/65536.0,1,-nbitq), 
to_sfixed(2487.0/65536.0,1,-nbitq), 
to_sfixed(2539.0/65536.0,1,-nbitq), 
to_sfixed(-1413.0/65536.0,1,-nbitq), 
to_sfixed(-8393.0/65536.0,1,-nbitq), 
to_sfixed(-3085.0/65536.0,1,-nbitq), 
to_sfixed(-5718.0/65536.0,1,-nbitq), 
to_sfixed(-156.0/65536.0,1,-nbitq), 
to_sfixed(-7683.0/65536.0,1,-nbitq), 
to_sfixed(2329.0/65536.0,1,-nbitq), 
to_sfixed(-2165.0/65536.0,1,-nbitq), 
to_sfixed(-2298.0/65536.0,1,-nbitq), 
to_sfixed(-931.0/65536.0,1,-nbitq), 
to_sfixed(-6286.0/65536.0,1,-nbitq), 
to_sfixed(-3015.0/65536.0,1,-nbitq), 
to_sfixed(-3996.0/65536.0,1,-nbitq), 
to_sfixed(-3580.0/65536.0,1,-nbitq), 
to_sfixed(7809.0/65536.0,1,-nbitq), 
to_sfixed(12582.0/65536.0,1,-nbitq), 
to_sfixed(953.0/65536.0,1,-nbitq), 
to_sfixed(2330.0/65536.0,1,-nbitq), 
to_sfixed(692.0/65536.0,1,-nbitq), 
to_sfixed(-775.0/65536.0,1,-nbitq), 
to_sfixed(-2861.0/65536.0,1,-nbitq), 
to_sfixed(-3741.0/65536.0,1,-nbitq), 
to_sfixed(-4874.0/65536.0,1,-nbitq), 
to_sfixed(-9686.0/65536.0,1,-nbitq), 
to_sfixed(-2796.0/65536.0,1,-nbitq), 
to_sfixed(-1096.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3705.0/65536.0,1,-nbitq), 
to_sfixed(-3552.0/65536.0,1,-nbitq), 
to_sfixed(-4227.0/65536.0,1,-nbitq), 
to_sfixed(2681.0/65536.0,1,-nbitq), 
to_sfixed(-2018.0/65536.0,1,-nbitq), 
to_sfixed(5271.0/65536.0,1,-nbitq), 
to_sfixed(1390.0/65536.0,1,-nbitq), 
to_sfixed(-2747.0/65536.0,1,-nbitq), 
to_sfixed(3748.0/65536.0,1,-nbitq), 
to_sfixed(995.0/65536.0,1,-nbitq), 
to_sfixed(2288.0/65536.0,1,-nbitq), 
to_sfixed(-8625.0/65536.0,1,-nbitq), 
to_sfixed(-1224.0/65536.0,1,-nbitq), 
to_sfixed(1647.0/65536.0,1,-nbitq), 
to_sfixed(-1445.0/65536.0,1,-nbitq), 
to_sfixed(310.0/65536.0,1,-nbitq), 
to_sfixed(-645.0/65536.0,1,-nbitq), 
to_sfixed(-5470.0/65536.0,1,-nbitq), 
to_sfixed(479.0/65536.0,1,-nbitq), 
to_sfixed(1697.0/65536.0,1,-nbitq), 
to_sfixed(1808.0/65536.0,1,-nbitq), 
to_sfixed(13119.0/65536.0,1,-nbitq), 
to_sfixed(3816.0/65536.0,1,-nbitq), 
to_sfixed(-8775.0/65536.0,1,-nbitq), 
to_sfixed(-2273.0/65536.0,1,-nbitq), 
to_sfixed(-4948.0/65536.0,1,-nbitq), 
to_sfixed(-3580.0/65536.0,1,-nbitq), 
to_sfixed(890.0/65536.0,1,-nbitq), 
to_sfixed(21461.0/65536.0,1,-nbitq), 
to_sfixed(2760.0/65536.0,1,-nbitq), 
to_sfixed(-4067.0/65536.0,1,-nbitq), 
to_sfixed(-5893.0/65536.0,1,-nbitq), 
to_sfixed(-5997.0/65536.0,1,-nbitq), 
to_sfixed(-8948.0/65536.0,1,-nbitq), 
to_sfixed(1587.0/65536.0,1,-nbitq), 
to_sfixed(1108.0/65536.0,1,-nbitq), 
to_sfixed(-5802.0/65536.0,1,-nbitq), 
to_sfixed(-4990.0/65536.0,1,-nbitq), 
to_sfixed(-4496.0/65536.0,1,-nbitq), 
to_sfixed(2482.0/65536.0,1,-nbitq), 
to_sfixed(5372.0/65536.0,1,-nbitq), 
to_sfixed(-128.0/65536.0,1,-nbitq), 
to_sfixed(672.0/65536.0,1,-nbitq), 
to_sfixed(4454.0/65536.0,1,-nbitq), 
to_sfixed(191.0/65536.0,1,-nbitq), 
to_sfixed(-7710.0/65536.0,1,-nbitq), 
to_sfixed(1579.0/65536.0,1,-nbitq), 
to_sfixed(9977.0/65536.0,1,-nbitq), 
to_sfixed(-2333.0/65536.0,1,-nbitq), 
to_sfixed(426.0/65536.0,1,-nbitq), 
to_sfixed(2507.0/65536.0,1,-nbitq), 
to_sfixed(-2330.0/65536.0,1,-nbitq), 
to_sfixed(-2262.0/65536.0,1,-nbitq), 
to_sfixed(3714.0/65536.0,1,-nbitq), 
to_sfixed(-1413.0/65536.0,1,-nbitq), 
to_sfixed(-8955.0/65536.0,1,-nbitq), 
to_sfixed(-3343.0/65536.0,1,-nbitq), 
to_sfixed(-2064.0/65536.0,1,-nbitq), 
to_sfixed(-1108.0/65536.0,1,-nbitq), 
to_sfixed(-4526.0/65536.0,1,-nbitq), 
to_sfixed(5348.0/65536.0,1,-nbitq), 
to_sfixed(841.0/65536.0,1,-nbitq), 
to_sfixed(2926.0/65536.0,1,-nbitq), 
to_sfixed(-97.0/65536.0,1,-nbitq), 
to_sfixed(-1549.0/65536.0,1,-nbitq), 
to_sfixed(-108.0/65536.0,1,-nbitq), 
to_sfixed(106.0/65536.0,1,-nbitq), 
to_sfixed(-6891.0/65536.0,1,-nbitq), 
to_sfixed(9196.0/65536.0,1,-nbitq), 
to_sfixed(9819.0/65536.0,1,-nbitq), 
to_sfixed(1199.0/65536.0,1,-nbitq), 
to_sfixed(7978.0/65536.0,1,-nbitq), 
to_sfixed(-200.0/65536.0,1,-nbitq), 
to_sfixed(1343.0/65536.0,1,-nbitq), 
to_sfixed(-2794.0/65536.0,1,-nbitq), 
to_sfixed(-862.0/65536.0,1,-nbitq), 
to_sfixed(-9094.0/65536.0,1,-nbitq), 
to_sfixed(-5373.0/65536.0,1,-nbitq), 
to_sfixed(1296.0/65536.0,1,-nbitq), 
to_sfixed(-4587.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1846.0/65536.0,1,-nbitq), 
to_sfixed(-2117.0/65536.0,1,-nbitq), 
to_sfixed(1667.0/65536.0,1,-nbitq), 
to_sfixed(4230.0/65536.0,1,-nbitq), 
to_sfixed(6303.0/65536.0,1,-nbitq), 
to_sfixed(-2388.0/65536.0,1,-nbitq), 
to_sfixed(4015.0/65536.0,1,-nbitq), 
to_sfixed(-4305.0/65536.0,1,-nbitq), 
to_sfixed(2448.0/65536.0,1,-nbitq), 
to_sfixed(-1790.0/65536.0,1,-nbitq), 
to_sfixed(3282.0/65536.0,1,-nbitq), 
to_sfixed(3703.0/65536.0,1,-nbitq), 
to_sfixed(-2164.0/65536.0,1,-nbitq), 
to_sfixed(-4717.0/65536.0,1,-nbitq), 
to_sfixed(-1854.0/65536.0,1,-nbitq), 
to_sfixed(1439.0/65536.0,1,-nbitq), 
to_sfixed(-2715.0/65536.0,1,-nbitq), 
to_sfixed(-7756.0/65536.0,1,-nbitq), 
to_sfixed(-1451.0/65536.0,1,-nbitq), 
to_sfixed(-2228.0/65536.0,1,-nbitq), 
to_sfixed(3624.0/65536.0,1,-nbitq), 
to_sfixed(2386.0/65536.0,1,-nbitq), 
to_sfixed(6462.0/65536.0,1,-nbitq), 
to_sfixed(-8374.0/65536.0,1,-nbitq), 
to_sfixed(-212.0/65536.0,1,-nbitq), 
to_sfixed(-3841.0/65536.0,1,-nbitq), 
to_sfixed(-773.0/65536.0,1,-nbitq), 
to_sfixed(3337.0/65536.0,1,-nbitq), 
to_sfixed(20137.0/65536.0,1,-nbitq), 
to_sfixed(2011.0/65536.0,1,-nbitq), 
to_sfixed(1147.0/65536.0,1,-nbitq), 
to_sfixed(-2756.0/65536.0,1,-nbitq), 
to_sfixed(4080.0/65536.0,1,-nbitq), 
to_sfixed(-4743.0/65536.0,1,-nbitq), 
to_sfixed(1002.0/65536.0,1,-nbitq), 
to_sfixed(-2922.0/65536.0,1,-nbitq), 
to_sfixed(-8720.0/65536.0,1,-nbitq), 
to_sfixed(-8444.0/65536.0,1,-nbitq), 
to_sfixed(-4536.0/65536.0,1,-nbitq), 
to_sfixed(2130.0/65536.0,1,-nbitq), 
to_sfixed(4744.0/65536.0,1,-nbitq), 
to_sfixed(-2333.0/65536.0,1,-nbitq), 
to_sfixed(1234.0/65536.0,1,-nbitq), 
to_sfixed(2911.0/65536.0,1,-nbitq), 
to_sfixed(2252.0/65536.0,1,-nbitq), 
to_sfixed(-23.0/65536.0,1,-nbitq), 
to_sfixed(-1504.0/65536.0,1,-nbitq), 
to_sfixed(10299.0/65536.0,1,-nbitq), 
to_sfixed(2029.0/65536.0,1,-nbitq), 
to_sfixed(-1847.0/65536.0,1,-nbitq), 
to_sfixed(-1930.0/65536.0,1,-nbitq), 
to_sfixed(155.0/65536.0,1,-nbitq), 
to_sfixed(1060.0/65536.0,1,-nbitq), 
to_sfixed(12751.0/65536.0,1,-nbitq), 
to_sfixed(-837.0/65536.0,1,-nbitq), 
to_sfixed(-2275.0/65536.0,1,-nbitq), 
to_sfixed(431.0/65536.0,1,-nbitq), 
to_sfixed(-4085.0/65536.0,1,-nbitq), 
to_sfixed(-498.0/65536.0,1,-nbitq), 
to_sfixed(682.0/65536.0,1,-nbitq), 
to_sfixed(7367.0/65536.0,1,-nbitq), 
to_sfixed(532.0/65536.0,1,-nbitq), 
to_sfixed(-1082.0/65536.0,1,-nbitq), 
to_sfixed(1968.0/65536.0,1,-nbitq), 
to_sfixed(3856.0/65536.0,1,-nbitq), 
to_sfixed(-5708.0/65536.0,1,-nbitq), 
to_sfixed(-2702.0/65536.0,1,-nbitq), 
to_sfixed(-4565.0/65536.0,1,-nbitq), 
to_sfixed(8051.0/65536.0,1,-nbitq), 
to_sfixed(9582.0/65536.0,1,-nbitq), 
to_sfixed(590.0/65536.0,1,-nbitq), 
to_sfixed(5102.0/65536.0,1,-nbitq), 
to_sfixed(4945.0/65536.0,1,-nbitq), 
to_sfixed(-304.0/65536.0,1,-nbitq), 
to_sfixed(139.0/65536.0,1,-nbitq), 
to_sfixed(-2644.0/65536.0,1,-nbitq), 
to_sfixed(-17880.0/65536.0,1,-nbitq), 
to_sfixed(-7561.0/65536.0,1,-nbitq), 
to_sfixed(996.0/65536.0,1,-nbitq), 
to_sfixed(-5576.0/65536.0,1,-nbitq)  ), 
( to_sfixed(660.0/65536.0,1,-nbitq), 
to_sfixed(-2062.0/65536.0,1,-nbitq), 
to_sfixed(5457.0/65536.0,1,-nbitq), 
to_sfixed(8648.0/65536.0,1,-nbitq), 
to_sfixed(5838.0/65536.0,1,-nbitq), 
to_sfixed(3015.0/65536.0,1,-nbitq), 
to_sfixed(2552.0/65536.0,1,-nbitq), 
to_sfixed(-900.0/65536.0,1,-nbitq), 
to_sfixed(-3971.0/65536.0,1,-nbitq), 
to_sfixed(-906.0/65536.0,1,-nbitq), 
to_sfixed(-1222.0/65536.0,1,-nbitq), 
to_sfixed(-6638.0/65536.0,1,-nbitq), 
to_sfixed(-388.0/65536.0,1,-nbitq), 
to_sfixed(-4430.0/65536.0,1,-nbitq), 
to_sfixed(1529.0/65536.0,1,-nbitq), 
to_sfixed(-2267.0/65536.0,1,-nbitq), 
to_sfixed(-2215.0/65536.0,1,-nbitq), 
to_sfixed(-1550.0/65536.0,1,-nbitq), 
to_sfixed(-2221.0/65536.0,1,-nbitq), 
to_sfixed(-145.0/65536.0,1,-nbitq), 
to_sfixed(2836.0/65536.0,1,-nbitq), 
to_sfixed(1204.0/65536.0,1,-nbitq), 
to_sfixed(-1630.0/65536.0,1,-nbitq), 
to_sfixed(-5456.0/65536.0,1,-nbitq), 
to_sfixed(-2381.0/65536.0,1,-nbitq), 
to_sfixed(3422.0/65536.0,1,-nbitq), 
to_sfixed(321.0/65536.0,1,-nbitq), 
to_sfixed(259.0/65536.0,1,-nbitq), 
to_sfixed(13459.0/65536.0,1,-nbitq), 
to_sfixed(-1497.0/65536.0,1,-nbitq), 
to_sfixed(-12.0/65536.0,1,-nbitq), 
to_sfixed(-4414.0/65536.0,1,-nbitq), 
to_sfixed(3962.0/65536.0,1,-nbitq), 
to_sfixed(-2111.0/65536.0,1,-nbitq), 
to_sfixed(-274.0/65536.0,1,-nbitq), 
to_sfixed(-3062.0/65536.0,1,-nbitq), 
to_sfixed(-6648.0/65536.0,1,-nbitq), 
to_sfixed(-2415.0/65536.0,1,-nbitq), 
to_sfixed(-3071.0/65536.0,1,-nbitq), 
to_sfixed(-1603.0/65536.0,1,-nbitq), 
to_sfixed(7393.0/65536.0,1,-nbitq), 
to_sfixed(312.0/65536.0,1,-nbitq), 
to_sfixed(3426.0/65536.0,1,-nbitq), 
to_sfixed(1522.0/65536.0,1,-nbitq), 
to_sfixed(-2472.0/65536.0,1,-nbitq), 
to_sfixed(4216.0/65536.0,1,-nbitq), 
to_sfixed(-1041.0/65536.0,1,-nbitq), 
to_sfixed(6645.0/65536.0,1,-nbitq), 
to_sfixed(-2670.0/65536.0,1,-nbitq), 
to_sfixed(-1354.0/65536.0,1,-nbitq), 
to_sfixed(1161.0/65536.0,1,-nbitq), 
to_sfixed(-743.0/65536.0,1,-nbitq), 
to_sfixed(-2623.0/65536.0,1,-nbitq), 
to_sfixed(11716.0/65536.0,1,-nbitq), 
to_sfixed(-1517.0/65536.0,1,-nbitq), 
to_sfixed(-98.0/65536.0,1,-nbitq), 
to_sfixed(2718.0/65536.0,1,-nbitq), 
to_sfixed(1114.0/65536.0,1,-nbitq), 
to_sfixed(-601.0/65536.0,1,-nbitq), 
to_sfixed(-4293.0/65536.0,1,-nbitq), 
to_sfixed(4147.0/65536.0,1,-nbitq), 
to_sfixed(2207.0/65536.0,1,-nbitq), 
to_sfixed(2564.0/65536.0,1,-nbitq), 
to_sfixed(-2675.0/65536.0,1,-nbitq), 
to_sfixed(4156.0/65536.0,1,-nbitq), 
to_sfixed(-1397.0/65536.0,1,-nbitq), 
to_sfixed(2003.0/65536.0,1,-nbitq), 
to_sfixed(5417.0/65536.0,1,-nbitq), 
to_sfixed(5674.0/65536.0,1,-nbitq), 
to_sfixed(14895.0/65536.0,1,-nbitq), 
to_sfixed(783.0/65536.0,1,-nbitq), 
to_sfixed(4467.0/65536.0,1,-nbitq), 
to_sfixed(3897.0/65536.0,1,-nbitq), 
to_sfixed(2351.0/65536.0,1,-nbitq), 
to_sfixed(-1059.0/65536.0,1,-nbitq), 
to_sfixed(11.0/65536.0,1,-nbitq), 
to_sfixed(-8981.0/65536.0,1,-nbitq), 
to_sfixed(27.0/65536.0,1,-nbitq), 
to_sfixed(-2076.0/65536.0,1,-nbitq), 
to_sfixed(-4927.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2251.0/65536.0,1,-nbitq), 
to_sfixed(303.0/65536.0,1,-nbitq), 
to_sfixed(4962.0/65536.0,1,-nbitq), 
to_sfixed(4979.0/65536.0,1,-nbitq), 
to_sfixed(193.0/65536.0,1,-nbitq), 
to_sfixed(4848.0/65536.0,1,-nbitq), 
to_sfixed(634.0/65536.0,1,-nbitq), 
to_sfixed(2076.0/65536.0,1,-nbitq), 
to_sfixed(-3906.0/65536.0,1,-nbitq), 
to_sfixed(1241.0/65536.0,1,-nbitq), 
to_sfixed(2572.0/65536.0,1,-nbitq), 
to_sfixed(-4671.0/65536.0,1,-nbitq), 
to_sfixed(3727.0/65536.0,1,-nbitq), 
to_sfixed(-8861.0/65536.0,1,-nbitq), 
to_sfixed(1410.0/65536.0,1,-nbitq), 
to_sfixed(2711.0/65536.0,1,-nbitq), 
to_sfixed(-332.0/65536.0,1,-nbitq), 
to_sfixed(-1466.0/65536.0,1,-nbitq), 
to_sfixed(-6406.0/65536.0,1,-nbitq), 
to_sfixed(-1991.0/65536.0,1,-nbitq), 
to_sfixed(4663.0/65536.0,1,-nbitq), 
to_sfixed(178.0/65536.0,1,-nbitq), 
to_sfixed(-4775.0/65536.0,1,-nbitq), 
to_sfixed(-8072.0/65536.0,1,-nbitq), 
to_sfixed(-1900.0/65536.0,1,-nbitq), 
to_sfixed(3329.0/65536.0,1,-nbitq), 
to_sfixed(-161.0/65536.0,1,-nbitq), 
to_sfixed(-2373.0/65536.0,1,-nbitq), 
to_sfixed(8422.0/65536.0,1,-nbitq), 
to_sfixed(-3770.0/65536.0,1,-nbitq), 
to_sfixed(-591.0/65536.0,1,-nbitq), 
to_sfixed(-2134.0/65536.0,1,-nbitq), 
to_sfixed(6594.0/65536.0,1,-nbitq), 
to_sfixed(2190.0/65536.0,1,-nbitq), 
to_sfixed(-1348.0/65536.0,1,-nbitq), 
to_sfixed(1957.0/65536.0,1,-nbitq), 
to_sfixed(1636.0/65536.0,1,-nbitq), 
to_sfixed(2787.0/65536.0,1,-nbitq), 
to_sfixed(-2031.0/65536.0,1,-nbitq), 
to_sfixed(1653.0/65536.0,1,-nbitq), 
to_sfixed(2208.0/65536.0,1,-nbitq), 
to_sfixed(2660.0/65536.0,1,-nbitq), 
to_sfixed(-451.0/65536.0,1,-nbitq), 
to_sfixed(129.0/65536.0,1,-nbitq), 
to_sfixed(1352.0/65536.0,1,-nbitq), 
to_sfixed(782.0/65536.0,1,-nbitq), 
to_sfixed(-694.0/65536.0,1,-nbitq), 
to_sfixed(3201.0/65536.0,1,-nbitq), 
to_sfixed(-2026.0/65536.0,1,-nbitq), 
to_sfixed(3044.0/65536.0,1,-nbitq), 
to_sfixed(-647.0/65536.0,1,-nbitq), 
to_sfixed(3565.0/65536.0,1,-nbitq), 
to_sfixed(3927.0/65536.0,1,-nbitq), 
to_sfixed(13259.0/65536.0,1,-nbitq), 
to_sfixed(-4856.0/65536.0,1,-nbitq), 
to_sfixed(-6793.0/65536.0,1,-nbitq), 
to_sfixed(-3101.0/65536.0,1,-nbitq), 
to_sfixed(703.0/65536.0,1,-nbitq), 
to_sfixed(2039.0/65536.0,1,-nbitq), 
to_sfixed(-6495.0/65536.0,1,-nbitq), 
to_sfixed(10750.0/65536.0,1,-nbitq), 
to_sfixed(1917.0/65536.0,1,-nbitq), 
to_sfixed(2532.0/65536.0,1,-nbitq), 
to_sfixed(-3010.0/65536.0,1,-nbitq), 
to_sfixed(6404.0/65536.0,1,-nbitq), 
to_sfixed(-2473.0/65536.0,1,-nbitq), 
to_sfixed(1425.0/65536.0,1,-nbitq), 
to_sfixed(2297.0/65536.0,1,-nbitq), 
to_sfixed(3557.0/65536.0,1,-nbitq), 
to_sfixed(8061.0/65536.0,1,-nbitq), 
to_sfixed(1072.0/65536.0,1,-nbitq), 
to_sfixed(-3347.0/65536.0,1,-nbitq), 
to_sfixed(6401.0/65536.0,1,-nbitq), 
to_sfixed(-1350.0/65536.0,1,-nbitq), 
to_sfixed(587.0/65536.0,1,-nbitq), 
to_sfixed(1208.0/65536.0,1,-nbitq), 
to_sfixed(-9412.0/65536.0,1,-nbitq), 
to_sfixed(2849.0/65536.0,1,-nbitq), 
to_sfixed(284.0/65536.0,1,-nbitq), 
to_sfixed(-2718.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3621.0/65536.0,1,-nbitq), 
to_sfixed(-3029.0/65536.0,1,-nbitq), 
to_sfixed(1072.0/65536.0,1,-nbitq), 
to_sfixed(7284.0/65536.0,1,-nbitq), 
to_sfixed(-360.0/65536.0,1,-nbitq), 
to_sfixed(1262.0/65536.0,1,-nbitq), 
to_sfixed(-990.0/65536.0,1,-nbitq), 
to_sfixed(6901.0/65536.0,1,-nbitq), 
to_sfixed(-3985.0/65536.0,1,-nbitq), 
to_sfixed(-77.0/65536.0,1,-nbitq), 
to_sfixed(4111.0/65536.0,1,-nbitq), 
to_sfixed(-4648.0/65536.0,1,-nbitq), 
to_sfixed(1047.0/65536.0,1,-nbitq), 
to_sfixed(-5928.0/65536.0,1,-nbitq), 
to_sfixed(-119.0/65536.0,1,-nbitq), 
to_sfixed(1115.0/65536.0,1,-nbitq), 
to_sfixed(-1969.0/65536.0,1,-nbitq), 
to_sfixed(-727.0/65536.0,1,-nbitq), 
to_sfixed(159.0/65536.0,1,-nbitq), 
to_sfixed(1856.0/65536.0,1,-nbitq), 
to_sfixed(6868.0/65536.0,1,-nbitq), 
to_sfixed(-1884.0/65536.0,1,-nbitq), 
to_sfixed(-1265.0/65536.0,1,-nbitq), 
to_sfixed(-4839.0/65536.0,1,-nbitq), 
to_sfixed(-3208.0/65536.0,1,-nbitq), 
to_sfixed(6330.0/65536.0,1,-nbitq), 
to_sfixed(4721.0/65536.0,1,-nbitq), 
to_sfixed(-1247.0/65536.0,1,-nbitq), 
to_sfixed(7297.0/65536.0,1,-nbitq), 
to_sfixed(-1583.0/65536.0,1,-nbitq), 
to_sfixed(-1387.0/65536.0,1,-nbitq), 
to_sfixed(-1779.0/65536.0,1,-nbitq), 
to_sfixed(3354.0/65536.0,1,-nbitq), 
to_sfixed(-1431.0/65536.0,1,-nbitq), 
to_sfixed(1773.0/65536.0,1,-nbitq), 
to_sfixed(3046.0/65536.0,1,-nbitq), 
to_sfixed(111.0/65536.0,1,-nbitq), 
to_sfixed(-3451.0/65536.0,1,-nbitq), 
to_sfixed(-2983.0/65536.0,1,-nbitq), 
to_sfixed(1990.0/65536.0,1,-nbitq), 
to_sfixed(-2959.0/65536.0,1,-nbitq), 
to_sfixed(-1779.0/65536.0,1,-nbitq), 
to_sfixed(701.0/65536.0,1,-nbitq), 
to_sfixed(-857.0/65536.0,1,-nbitq), 
to_sfixed(-35.0/65536.0,1,-nbitq), 
to_sfixed(2110.0/65536.0,1,-nbitq), 
to_sfixed(-3196.0/65536.0,1,-nbitq), 
to_sfixed(596.0/65536.0,1,-nbitq), 
to_sfixed(2120.0/65536.0,1,-nbitq), 
to_sfixed(4025.0/65536.0,1,-nbitq), 
to_sfixed(1905.0/65536.0,1,-nbitq), 
to_sfixed(-956.0/65536.0,1,-nbitq), 
to_sfixed(-1498.0/65536.0,1,-nbitq), 
to_sfixed(16457.0/65536.0,1,-nbitq), 
to_sfixed(-4012.0/65536.0,1,-nbitq), 
to_sfixed(-6413.0/65536.0,1,-nbitq), 
to_sfixed(1487.0/65536.0,1,-nbitq), 
to_sfixed(4757.0/65536.0,1,-nbitq), 
to_sfixed(-2578.0/65536.0,1,-nbitq), 
to_sfixed(-2534.0/65536.0,1,-nbitq), 
to_sfixed(5505.0/65536.0,1,-nbitq), 
to_sfixed(-854.0/65536.0,1,-nbitq), 
to_sfixed(2631.0/65536.0,1,-nbitq), 
to_sfixed(-2382.0/65536.0,1,-nbitq), 
to_sfixed(1754.0/65536.0,1,-nbitq), 
to_sfixed(4132.0/65536.0,1,-nbitq), 
to_sfixed(4172.0/65536.0,1,-nbitq), 
to_sfixed(613.0/65536.0,1,-nbitq), 
to_sfixed(-2069.0/65536.0,1,-nbitq), 
to_sfixed(-1153.0/65536.0,1,-nbitq), 
to_sfixed(618.0/65536.0,1,-nbitq), 
to_sfixed(-2011.0/65536.0,1,-nbitq), 
to_sfixed(7303.0/65536.0,1,-nbitq), 
to_sfixed(2367.0/65536.0,1,-nbitq), 
to_sfixed(-1965.0/65536.0,1,-nbitq), 
to_sfixed(-1663.0/65536.0,1,-nbitq), 
to_sfixed(-2122.0/65536.0,1,-nbitq), 
to_sfixed(1675.0/65536.0,1,-nbitq), 
to_sfixed(-1471.0/65536.0,1,-nbitq), 
to_sfixed(-3336.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4276.0/65536.0,1,-nbitq), 
to_sfixed(195.0/65536.0,1,-nbitq), 
to_sfixed(-4222.0/65536.0,1,-nbitq), 
to_sfixed(5765.0/65536.0,1,-nbitq), 
to_sfixed(2977.0/65536.0,1,-nbitq), 
to_sfixed(1500.0/65536.0,1,-nbitq), 
to_sfixed(-870.0/65536.0,1,-nbitq), 
to_sfixed(7292.0/65536.0,1,-nbitq), 
to_sfixed(-3220.0/65536.0,1,-nbitq), 
to_sfixed(659.0/65536.0,1,-nbitq), 
to_sfixed(-1243.0/65536.0,1,-nbitq), 
to_sfixed(-7279.0/65536.0,1,-nbitq), 
to_sfixed(1459.0/65536.0,1,-nbitq), 
to_sfixed(-1667.0/65536.0,1,-nbitq), 
to_sfixed(-2759.0/65536.0,1,-nbitq), 
to_sfixed(107.0/65536.0,1,-nbitq), 
to_sfixed(2559.0/65536.0,1,-nbitq), 
to_sfixed(-2356.0/65536.0,1,-nbitq), 
to_sfixed(-516.0/65536.0,1,-nbitq), 
to_sfixed(2115.0/65536.0,1,-nbitq), 
to_sfixed(2030.0/65536.0,1,-nbitq), 
to_sfixed(1887.0/65536.0,1,-nbitq), 
to_sfixed(-2808.0/65536.0,1,-nbitq), 
to_sfixed(-868.0/65536.0,1,-nbitq), 
to_sfixed(-2241.0/65536.0,1,-nbitq), 
to_sfixed(3390.0/65536.0,1,-nbitq), 
to_sfixed(-4083.0/65536.0,1,-nbitq), 
to_sfixed(-2366.0/65536.0,1,-nbitq), 
to_sfixed(6645.0/65536.0,1,-nbitq), 
to_sfixed(-1128.0/65536.0,1,-nbitq), 
to_sfixed(-1407.0/65536.0,1,-nbitq), 
to_sfixed(-6795.0/65536.0,1,-nbitq), 
to_sfixed(4334.0/65536.0,1,-nbitq), 
to_sfixed(-3560.0/65536.0,1,-nbitq), 
to_sfixed(-1292.0/65536.0,1,-nbitq), 
to_sfixed(830.0/65536.0,1,-nbitq), 
to_sfixed(-3904.0/65536.0,1,-nbitq), 
to_sfixed(-1490.0/65536.0,1,-nbitq), 
to_sfixed(-1870.0/65536.0,1,-nbitq), 
to_sfixed(1609.0/65536.0,1,-nbitq), 
to_sfixed(-2480.0/65536.0,1,-nbitq), 
to_sfixed(-920.0/65536.0,1,-nbitq), 
to_sfixed(-1513.0/65536.0,1,-nbitq), 
to_sfixed(-893.0/65536.0,1,-nbitq), 
to_sfixed(-1047.0/65536.0,1,-nbitq), 
to_sfixed(194.0/65536.0,1,-nbitq), 
to_sfixed(-2209.0/65536.0,1,-nbitq), 
to_sfixed(2891.0/65536.0,1,-nbitq), 
to_sfixed(1733.0/65536.0,1,-nbitq), 
to_sfixed(1038.0/65536.0,1,-nbitq), 
to_sfixed(896.0/65536.0,1,-nbitq), 
to_sfixed(-670.0/65536.0,1,-nbitq), 
to_sfixed(-4509.0/65536.0,1,-nbitq), 
to_sfixed(8761.0/65536.0,1,-nbitq), 
to_sfixed(-4090.0/65536.0,1,-nbitq), 
to_sfixed(-5885.0/65536.0,1,-nbitq), 
to_sfixed(-2579.0/65536.0,1,-nbitq), 
to_sfixed(2063.0/65536.0,1,-nbitq), 
to_sfixed(-1919.0/65536.0,1,-nbitq), 
to_sfixed(-2709.0/65536.0,1,-nbitq), 
to_sfixed(-415.0/65536.0,1,-nbitq), 
to_sfixed(-2725.0/65536.0,1,-nbitq), 
to_sfixed(-473.0/65536.0,1,-nbitq), 
to_sfixed(-1734.0/65536.0,1,-nbitq), 
to_sfixed(2358.0/65536.0,1,-nbitq), 
to_sfixed(1416.0/65536.0,1,-nbitq), 
to_sfixed(6159.0/65536.0,1,-nbitq), 
to_sfixed(-2313.0/65536.0,1,-nbitq), 
to_sfixed(2736.0/65536.0,1,-nbitq), 
to_sfixed(2533.0/65536.0,1,-nbitq), 
to_sfixed(1638.0/65536.0,1,-nbitq), 
to_sfixed(-4146.0/65536.0,1,-nbitq), 
to_sfixed(6779.0/65536.0,1,-nbitq), 
to_sfixed(2490.0/65536.0,1,-nbitq), 
to_sfixed(-894.0/65536.0,1,-nbitq), 
to_sfixed(-328.0/65536.0,1,-nbitq), 
to_sfixed(-5328.0/65536.0,1,-nbitq), 
to_sfixed(1193.0/65536.0,1,-nbitq), 
to_sfixed(-1708.0/65536.0,1,-nbitq), 
to_sfixed(-2360.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3362.0/65536.0,1,-nbitq), 
to_sfixed(-2454.0/65536.0,1,-nbitq), 
to_sfixed(-5084.0/65536.0,1,-nbitq), 
to_sfixed(2170.0/65536.0,1,-nbitq), 
to_sfixed(-2315.0/65536.0,1,-nbitq), 
to_sfixed(-1329.0/65536.0,1,-nbitq), 
to_sfixed(-1638.0/65536.0,1,-nbitq), 
to_sfixed(3492.0/65536.0,1,-nbitq), 
to_sfixed(-5245.0/65536.0,1,-nbitq), 
to_sfixed(2868.0/65536.0,1,-nbitq), 
to_sfixed(-2650.0/65536.0,1,-nbitq), 
to_sfixed(-5295.0/65536.0,1,-nbitq), 
to_sfixed(-1234.0/65536.0,1,-nbitq), 
to_sfixed(-3448.0/65536.0,1,-nbitq), 
to_sfixed(-1630.0/65536.0,1,-nbitq), 
to_sfixed(-555.0/65536.0,1,-nbitq), 
to_sfixed(-637.0/65536.0,1,-nbitq), 
to_sfixed(5997.0/65536.0,1,-nbitq), 
to_sfixed(3171.0/65536.0,1,-nbitq), 
to_sfixed(3155.0/65536.0,1,-nbitq), 
to_sfixed(-479.0/65536.0,1,-nbitq), 
to_sfixed(662.0/65536.0,1,-nbitq), 
to_sfixed(-4663.0/65536.0,1,-nbitq), 
to_sfixed(-3466.0/65536.0,1,-nbitq), 
to_sfixed(-2780.0/65536.0,1,-nbitq), 
to_sfixed(-132.0/65536.0,1,-nbitq), 
to_sfixed(-4445.0/65536.0,1,-nbitq), 
to_sfixed(-1124.0/65536.0,1,-nbitq), 
to_sfixed(4444.0/65536.0,1,-nbitq), 
to_sfixed(2077.0/65536.0,1,-nbitq), 
to_sfixed(-704.0/65536.0,1,-nbitq), 
to_sfixed(-1416.0/65536.0,1,-nbitq), 
to_sfixed(-2017.0/65536.0,1,-nbitq), 
to_sfixed(-5558.0/65536.0,1,-nbitq), 
to_sfixed(-142.0/65536.0,1,-nbitq), 
to_sfixed(2730.0/65536.0,1,-nbitq), 
to_sfixed(-6782.0/65536.0,1,-nbitq), 
to_sfixed(-3619.0/65536.0,1,-nbitq), 
to_sfixed(-251.0/65536.0,1,-nbitq), 
to_sfixed(1717.0/65536.0,1,-nbitq), 
to_sfixed(3376.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(2063.0/65536.0,1,-nbitq), 
to_sfixed(-1759.0/65536.0,1,-nbitq), 
to_sfixed(-145.0/65536.0,1,-nbitq), 
to_sfixed(1497.0/65536.0,1,-nbitq), 
to_sfixed(-406.0/65536.0,1,-nbitq), 
to_sfixed(-2562.0/65536.0,1,-nbitq), 
to_sfixed(2179.0/65536.0,1,-nbitq), 
to_sfixed(604.0/65536.0,1,-nbitq), 
to_sfixed(-1438.0/65536.0,1,-nbitq), 
to_sfixed(-636.0/65536.0,1,-nbitq), 
to_sfixed(-2448.0/65536.0,1,-nbitq), 
to_sfixed(6694.0/65536.0,1,-nbitq), 
to_sfixed(-4588.0/65536.0,1,-nbitq), 
to_sfixed(-3611.0/65536.0,1,-nbitq), 
to_sfixed(-438.0/65536.0,1,-nbitq), 
to_sfixed(5238.0/65536.0,1,-nbitq), 
to_sfixed(-1236.0/65536.0,1,-nbitq), 
to_sfixed(-3259.0/65536.0,1,-nbitq), 
to_sfixed(-732.0/65536.0,1,-nbitq), 
to_sfixed(762.0/65536.0,1,-nbitq), 
to_sfixed(-2809.0/65536.0,1,-nbitq), 
to_sfixed(-2840.0/65536.0,1,-nbitq), 
to_sfixed(-1843.0/65536.0,1,-nbitq), 
to_sfixed(-2033.0/65536.0,1,-nbitq), 
to_sfixed(1930.0/65536.0,1,-nbitq), 
to_sfixed(-1301.0/65536.0,1,-nbitq), 
to_sfixed(3177.0/65536.0,1,-nbitq), 
to_sfixed(3855.0/65536.0,1,-nbitq), 
to_sfixed(1923.0/65536.0,1,-nbitq), 
to_sfixed(-4385.0/65536.0,1,-nbitq), 
to_sfixed(1647.0/65536.0,1,-nbitq), 
to_sfixed(1478.0/65536.0,1,-nbitq), 
to_sfixed(-122.0/65536.0,1,-nbitq), 
to_sfixed(-947.0/65536.0,1,-nbitq), 
to_sfixed(-7328.0/65536.0,1,-nbitq), 
to_sfixed(3356.0/65536.0,1,-nbitq), 
to_sfixed(-1595.0/65536.0,1,-nbitq), 
to_sfixed(1057.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2242.0/65536.0,1,-nbitq), 
to_sfixed(2861.0/65536.0,1,-nbitq), 
to_sfixed(2021.0/65536.0,1,-nbitq), 
to_sfixed(732.0/65536.0,1,-nbitq), 
to_sfixed(-642.0/65536.0,1,-nbitq), 
to_sfixed(711.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(-563.0/65536.0,1,-nbitq), 
to_sfixed(-3641.0/65536.0,1,-nbitq), 
to_sfixed(-1673.0/65536.0,1,-nbitq), 
to_sfixed(-635.0/65536.0,1,-nbitq), 
to_sfixed(-1905.0/65536.0,1,-nbitq), 
to_sfixed(-1867.0/65536.0,1,-nbitq), 
to_sfixed(-2662.0/65536.0,1,-nbitq), 
to_sfixed(1702.0/65536.0,1,-nbitq), 
to_sfixed(-377.0/65536.0,1,-nbitq), 
to_sfixed(-51.0/65536.0,1,-nbitq), 
to_sfixed(4354.0/65536.0,1,-nbitq), 
to_sfixed(4305.0/65536.0,1,-nbitq), 
to_sfixed(-1606.0/65536.0,1,-nbitq), 
to_sfixed(-884.0/65536.0,1,-nbitq), 
to_sfixed(618.0/65536.0,1,-nbitq), 
to_sfixed(-1577.0/65536.0,1,-nbitq), 
to_sfixed(-922.0/65536.0,1,-nbitq), 
to_sfixed(3007.0/65536.0,1,-nbitq), 
to_sfixed(-1830.0/65536.0,1,-nbitq), 
to_sfixed(-4893.0/65536.0,1,-nbitq), 
to_sfixed(2509.0/65536.0,1,-nbitq), 
to_sfixed(3301.0/65536.0,1,-nbitq), 
to_sfixed(571.0/65536.0,1,-nbitq), 
to_sfixed(-2851.0/65536.0,1,-nbitq), 
to_sfixed(-1672.0/65536.0,1,-nbitq), 
to_sfixed(-2442.0/65536.0,1,-nbitq), 
to_sfixed(-1200.0/65536.0,1,-nbitq), 
to_sfixed(2426.0/65536.0,1,-nbitq), 
to_sfixed(-3098.0/65536.0,1,-nbitq), 
to_sfixed(-2626.0/65536.0,1,-nbitq), 
to_sfixed(1843.0/65536.0,1,-nbitq), 
to_sfixed(-4258.0/65536.0,1,-nbitq), 
to_sfixed(-1471.0/65536.0,1,-nbitq), 
to_sfixed(-2697.0/65536.0,1,-nbitq), 
to_sfixed(950.0/65536.0,1,-nbitq), 
to_sfixed(-2749.0/65536.0,1,-nbitq), 
to_sfixed(-1406.0/65536.0,1,-nbitq), 
to_sfixed(-1317.0/65536.0,1,-nbitq), 
to_sfixed(5237.0/65536.0,1,-nbitq), 
to_sfixed(1769.0/65536.0,1,-nbitq), 
to_sfixed(-1864.0/65536.0,1,-nbitq), 
to_sfixed(-262.0/65536.0,1,-nbitq), 
to_sfixed(195.0/65536.0,1,-nbitq), 
to_sfixed(983.0/65536.0,1,-nbitq), 
to_sfixed(2098.0/65536.0,1,-nbitq), 
to_sfixed(-3787.0/65536.0,1,-nbitq), 
to_sfixed(892.0/65536.0,1,-nbitq), 
to_sfixed(-1497.0/65536.0,1,-nbitq), 
to_sfixed(1748.0/65536.0,1,-nbitq), 
to_sfixed(-824.0/65536.0,1,-nbitq), 
to_sfixed(-477.0/65536.0,1,-nbitq), 
to_sfixed(-2616.0/65536.0,1,-nbitq), 
to_sfixed(1691.0/65536.0,1,-nbitq), 
to_sfixed(-1799.0/65536.0,1,-nbitq), 
to_sfixed(-1553.0/65536.0,1,-nbitq), 
to_sfixed(1577.0/65536.0,1,-nbitq), 
to_sfixed(2345.0/65536.0,1,-nbitq), 
to_sfixed(2772.0/65536.0,1,-nbitq), 
to_sfixed(2670.0/65536.0,1,-nbitq), 
to_sfixed(50.0/65536.0,1,-nbitq), 
to_sfixed(480.0/65536.0,1,-nbitq), 
to_sfixed(2133.0/65536.0,1,-nbitq), 
to_sfixed(-846.0/65536.0,1,-nbitq), 
to_sfixed(-914.0/65536.0,1,-nbitq), 
to_sfixed(-2859.0/65536.0,1,-nbitq), 
to_sfixed(4438.0/65536.0,1,-nbitq), 
to_sfixed(2518.0/65536.0,1,-nbitq), 
to_sfixed(1006.0/65536.0,1,-nbitq), 
to_sfixed(-839.0/65536.0,1,-nbitq), 
to_sfixed(-1282.0/65536.0,1,-nbitq), 
to_sfixed(-71.0/65536.0,1,-nbitq), 
to_sfixed(2638.0/65536.0,1,-nbitq), 
to_sfixed(2880.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2782.0/65536.0,1,-nbitq), 
to_sfixed(-2722.0/65536.0,1,-nbitq), 
to_sfixed(-1278.0/65536.0,1,-nbitq), 
to_sfixed(147.0/65536.0,1,-nbitq), 
to_sfixed(545.0/65536.0,1,-nbitq), 
to_sfixed(71.0/65536.0,1,-nbitq), 
to_sfixed(2490.0/65536.0,1,-nbitq), 
to_sfixed(1018.0/65536.0,1,-nbitq), 
to_sfixed(-1360.0/65536.0,1,-nbitq), 
to_sfixed(-2742.0/65536.0,1,-nbitq), 
to_sfixed(-2590.0/65536.0,1,-nbitq), 
to_sfixed(-162.0/65536.0,1,-nbitq), 
to_sfixed(-614.0/65536.0,1,-nbitq), 
to_sfixed(-3000.0/65536.0,1,-nbitq), 
to_sfixed(971.0/65536.0,1,-nbitq), 
to_sfixed(735.0/65536.0,1,-nbitq), 
to_sfixed(1783.0/65536.0,1,-nbitq), 
to_sfixed(1680.0/65536.0,1,-nbitq), 
to_sfixed(3903.0/65536.0,1,-nbitq), 
to_sfixed(2676.0/65536.0,1,-nbitq), 
to_sfixed(-1120.0/65536.0,1,-nbitq), 
to_sfixed(548.0/65536.0,1,-nbitq), 
to_sfixed(949.0/65536.0,1,-nbitq), 
to_sfixed(2734.0/65536.0,1,-nbitq), 
to_sfixed(-1866.0/65536.0,1,-nbitq), 
to_sfixed(1152.0/65536.0,1,-nbitq), 
to_sfixed(130.0/65536.0,1,-nbitq), 
to_sfixed(2701.0/65536.0,1,-nbitq), 
to_sfixed(-2339.0/65536.0,1,-nbitq), 
to_sfixed(1316.0/65536.0,1,-nbitq), 
to_sfixed(-1532.0/65536.0,1,-nbitq), 
to_sfixed(319.0/65536.0,1,-nbitq), 
to_sfixed(-4634.0/65536.0,1,-nbitq), 
to_sfixed(-3006.0/65536.0,1,-nbitq), 
to_sfixed(-2645.0/65536.0,1,-nbitq), 
to_sfixed(-1040.0/65536.0,1,-nbitq), 
to_sfixed(21.0/65536.0,1,-nbitq), 
to_sfixed(-4027.0/65536.0,1,-nbitq), 
to_sfixed(-640.0/65536.0,1,-nbitq), 
to_sfixed(2554.0/65536.0,1,-nbitq), 
to_sfixed(-1199.0/65536.0,1,-nbitq), 
to_sfixed(1949.0/65536.0,1,-nbitq), 
to_sfixed(-480.0/65536.0,1,-nbitq), 
to_sfixed(864.0/65536.0,1,-nbitq), 
to_sfixed(993.0/65536.0,1,-nbitq), 
to_sfixed(4534.0/65536.0,1,-nbitq), 
to_sfixed(-1464.0/65536.0,1,-nbitq), 
to_sfixed(81.0/65536.0,1,-nbitq), 
to_sfixed(-2166.0/65536.0,1,-nbitq), 
to_sfixed(2384.0/65536.0,1,-nbitq), 
to_sfixed(-2457.0/65536.0,1,-nbitq), 
to_sfixed(894.0/65536.0,1,-nbitq), 
to_sfixed(-1851.0/65536.0,1,-nbitq), 
to_sfixed(188.0/65536.0,1,-nbitq), 
to_sfixed(913.0/65536.0,1,-nbitq), 
to_sfixed(1582.0/65536.0,1,-nbitq), 
to_sfixed(1204.0/65536.0,1,-nbitq), 
to_sfixed(1818.0/65536.0,1,-nbitq), 
to_sfixed(-448.0/65536.0,1,-nbitq), 
to_sfixed(1041.0/65536.0,1,-nbitq), 
to_sfixed(-1241.0/65536.0,1,-nbitq), 
to_sfixed(1902.0/65536.0,1,-nbitq), 
to_sfixed(2674.0/65536.0,1,-nbitq), 
to_sfixed(366.0/65536.0,1,-nbitq), 
to_sfixed(690.0/65536.0,1,-nbitq), 
to_sfixed(1452.0/65536.0,1,-nbitq), 
to_sfixed(-1244.0/65536.0,1,-nbitq), 
to_sfixed(-3025.0/65536.0,1,-nbitq), 
to_sfixed(989.0/65536.0,1,-nbitq), 
to_sfixed(866.0/65536.0,1,-nbitq), 
to_sfixed(1105.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(-1509.0/65536.0,1,-nbitq), 
to_sfixed(313.0/65536.0,1,-nbitq), 
to_sfixed(-728.0/65536.0,1,-nbitq), 
to_sfixed(701.0/65536.0,1,-nbitq), 
to_sfixed(-3441.0/65536.0,1,-nbitq), 
to_sfixed(1898.0/65536.0,1,-nbitq), 
to_sfixed(-2512.0/65536.0,1,-nbitq), 
to_sfixed(5174.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(846.0/65536.0,1,-nbitq), 
to_sfixed(-423.0/65536.0,1,-nbitq), 
to_sfixed(-404.0/65536.0,1,-nbitq), 
to_sfixed(948.0/65536.0,1,-nbitq), 
to_sfixed(2079.0/65536.0,1,-nbitq), 
to_sfixed(767.0/65536.0,1,-nbitq), 
to_sfixed(2102.0/65536.0,1,-nbitq), 
to_sfixed(-1779.0/65536.0,1,-nbitq), 
to_sfixed(-2344.0/65536.0,1,-nbitq), 
to_sfixed(2145.0/65536.0,1,-nbitq), 
to_sfixed(-1229.0/65536.0,1,-nbitq), 
to_sfixed(1192.0/65536.0,1,-nbitq), 
to_sfixed(-1474.0/65536.0,1,-nbitq), 
to_sfixed(-2959.0/65536.0,1,-nbitq), 
to_sfixed(3448.0/65536.0,1,-nbitq), 
to_sfixed(482.0/65536.0,1,-nbitq), 
to_sfixed(288.0/65536.0,1,-nbitq), 
to_sfixed(-878.0/65536.0,1,-nbitq), 
to_sfixed(-1152.0/65536.0,1,-nbitq), 
to_sfixed(-1370.0/65536.0,1,-nbitq), 
to_sfixed(1624.0/65536.0,1,-nbitq), 
to_sfixed(1309.0/65536.0,1,-nbitq), 
to_sfixed(534.0/65536.0,1,-nbitq), 
to_sfixed(-803.0/65536.0,1,-nbitq), 
to_sfixed(817.0/65536.0,1,-nbitq), 
to_sfixed(908.0/65536.0,1,-nbitq), 
to_sfixed(-1968.0/65536.0,1,-nbitq), 
to_sfixed(1633.0/65536.0,1,-nbitq), 
to_sfixed(3659.0/65536.0,1,-nbitq), 
to_sfixed(-4123.0/65536.0,1,-nbitq), 
to_sfixed(123.0/65536.0,1,-nbitq), 
to_sfixed(-2269.0/65536.0,1,-nbitq), 
to_sfixed(142.0/65536.0,1,-nbitq), 
to_sfixed(-2797.0/65536.0,1,-nbitq), 
to_sfixed(163.0/65536.0,1,-nbitq), 
to_sfixed(941.0/65536.0,1,-nbitq), 
to_sfixed(1386.0/65536.0,1,-nbitq), 
to_sfixed(466.0/65536.0,1,-nbitq), 
to_sfixed(-737.0/65536.0,1,-nbitq), 
to_sfixed(-2984.0/65536.0,1,-nbitq), 
to_sfixed(-2540.0/65536.0,1,-nbitq), 
to_sfixed(-3005.0/65536.0,1,-nbitq), 
to_sfixed(-1693.0/65536.0,1,-nbitq), 
to_sfixed(1720.0/65536.0,1,-nbitq), 
to_sfixed(830.0/65536.0,1,-nbitq), 
to_sfixed(5132.0/65536.0,1,-nbitq), 
to_sfixed(-2011.0/65536.0,1,-nbitq), 
to_sfixed(1912.0/65536.0,1,-nbitq), 
to_sfixed(-744.0/65536.0,1,-nbitq), 
to_sfixed(3892.0/65536.0,1,-nbitq), 
to_sfixed(2191.0/65536.0,1,-nbitq), 
to_sfixed(-469.0/65536.0,1,-nbitq), 
to_sfixed(3198.0/65536.0,1,-nbitq), 
to_sfixed(-308.0/65536.0,1,-nbitq), 
to_sfixed(-580.0/65536.0,1,-nbitq), 
to_sfixed(-1531.0/65536.0,1,-nbitq), 
to_sfixed(-2721.0/65536.0,1,-nbitq), 
to_sfixed(-139.0/65536.0,1,-nbitq), 
to_sfixed(2131.0/65536.0,1,-nbitq), 
to_sfixed(466.0/65536.0,1,-nbitq), 
to_sfixed(-199.0/65536.0,1,-nbitq), 
to_sfixed(-2135.0/65536.0,1,-nbitq), 
to_sfixed(-1076.0/65536.0,1,-nbitq), 
to_sfixed(-1185.0/65536.0,1,-nbitq), 
to_sfixed(1711.0/65536.0,1,-nbitq), 
to_sfixed(2558.0/65536.0,1,-nbitq), 
to_sfixed(516.0/65536.0,1,-nbitq), 
to_sfixed(-4021.0/65536.0,1,-nbitq), 
to_sfixed(1877.0/65536.0,1,-nbitq), 
to_sfixed(-2806.0/65536.0,1,-nbitq), 
to_sfixed(1352.0/65536.0,1,-nbitq), 
to_sfixed(2771.0/65536.0,1,-nbitq), 
to_sfixed(541.0/65536.0,1,-nbitq), 
to_sfixed(431.0/65536.0,1,-nbitq), 
to_sfixed(977.0/65536.0,1,-nbitq), 
to_sfixed(2876.0/65536.0,1,-nbitq), 
to_sfixed(256.0/65536.0,1,-nbitq), 
to_sfixed(3470.0/65536.0,1,-nbitq), 
to_sfixed(1638.0/65536.0,1,-nbitq), 
to_sfixed(1467.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3184.0/65536.0,1,-nbitq), 
to_sfixed(-2638.0/65536.0,1,-nbitq), 
to_sfixed(2765.0/65536.0,1,-nbitq), 
to_sfixed(1470.0/65536.0,1,-nbitq), 
to_sfixed(-465.0/65536.0,1,-nbitq), 
to_sfixed(1119.0/65536.0,1,-nbitq), 
to_sfixed(-2836.0/65536.0,1,-nbitq), 
to_sfixed(2189.0/65536.0,1,-nbitq), 
to_sfixed(1502.0/65536.0,1,-nbitq), 
to_sfixed(2245.0/65536.0,1,-nbitq), 
to_sfixed(-3479.0/65536.0,1,-nbitq), 
to_sfixed(-2789.0/65536.0,1,-nbitq), 
to_sfixed(-1656.0/65536.0,1,-nbitq), 
to_sfixed(512.0/65536.0,1,-nbitq), 
to_sfixed(255.0/65536.0,1,-nbitq), 
to_sfixed(2532.0/65536.0,1,-nbitq), 
to_sfixed(-2072.0/65536.0,1,-nbitq), 
to_sfixed(3824.0/65536.0,1,-nbitq), 
to_sfixed(-197.0/65536.0,1,-nbitq), 
to_sfixed(1437.0/65536.0,1,-nbitq), 
to_sfixed(-2134.0/65536.0,1,-nbitq), 
to_sfixed(-2139.0/65536.0,1,-nbitq), 
to_sfixed(-294.0/65536.0,1,-nbitq), 
to_sfixed(772.0/65536.0,1,-nbitq), 
to_sfixed(1322.0/65536.0,1,-nbitq), 
to_sfixed(2044.0/65536.0,1,-nbitq), 
to_sfixed(1740.0/65536.0,1,-nbitq), 
to_sfixed(-1511.0/65536.0,1,-nbitq), 
to_sfixed(-1508.0/65536.0,1,-nbitq), 
to_sfixed(-4310.0/65536.0,1,-nbitq), 
to_sfixed(2438.0/65536.0,1,-nbitq), 
to_sfixed(-2687.0/65536.0,1,-nbitq), 
to_sfixed(-2226.0/65536.0,1,-nbitq), 
to_sfixed(-5198.0/65536.0,1,-nbitq), 
to_sfixed(-2087.0/65536.0,1,-nbitq), 
to_sfixed(836.0/65536.0,1,-nbitq), 
to_sfixed(113.0/65536.0,1,-nbitq), 
to_sfixed(-175.0/65536.0,1,-nbitq), 
to_sfixed(-1319.0/65536.0,1,-nbitq), 
to_sfixed(1850.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(-190.0/65536.0,1,-nbitq), 
to_sfixed(-1749.0/65536.0,1,-nbitq), 
to_sfixed(125.0/65536.0,1,-nbitq), 
to_sfixed(311.0/65536.0,1,-nbitq), 
to_sfixed(4732.0/65536.0,1,-nbitq), 
to_sfixed(2266.0/65536.0,1,-nbitq), 
to_sfixed(1550.0/65536.0,1,-nbitq), 
to_sfixed(-2148.0/65536.0,1,-nbitq), 
to_sfixed(4056.0/65536.0,1,-nbitq), 
to_sfixed(-1060.0/65536.0,1,-nbitq), 
to_sfixed(116.0/65536.0,1,-nbitq), 
to_sfixed(1111.0/65536.0,1,-nbitq), 
to_sfixed(1490.0/65536.0,1,-nbitq), 
to_sfixed(1220.0/65536.0,1,-nbitq), 
to_sfixed(-2361.0/65536.0,1,-nbitq), 
to_sfixed(2155.0/65536.0,1,-nbitq), 
to_sfixed(3770.0/65536.0,1,-nbitq), 
to_sfixed(2092.0/65536.0,1,-nbitq), 
to_sfixed(1301.0/65536.0,1,-nbitq), 
to_sfixed(-1267.0/65536.0,1,-nbitq), 
to_sfixed(693.0/65536.0,1,-nbitq), 
to_sfixed(1353.0/65536.0,1,-nbitq), 
to_sfixed(1299.0/65536.0,1,-nbitq), 
to_sfixed(3143.0/65536.0,1,-nbitq), 
to_sfixed(850.0/65536.0,1,-nbitq), 
to_sfixed(1897.0/65536.0,1,-nbitq), 
to_sfixed(664.0/65536.0,1,-nbitq), 
to_sfixed(3160.0/65536.0,1,-nbitq), 
to_sfixed(-2675.0/65536.0,1,-nbitq), 
to_sfixed(1501.0/65536.0,1,-nbitq), 
to_sfixed(1420.0/65536.0,1,-nbitq), 
to_sfixed(-668.0/65536.0,1,-nbitq), 
to_sfixed(-1171.0/65536.0,1,-nbitq), 
to_sfixed(-831.0/65536.0,1,-nbitq), 
to_sfixed(1558.0/65536.0,1,-nbitq), 
to_sfixed(-2646.0/65536.0,1,-nbitq), 
to_sfixed(-111.0/65536.0,1,-nbitq), 
to_sfixed(2319.0/65536.0,1,-nbitq), 
to_sfixed(1253.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3106.0/65536.0,1,-nbitq), 
to_sfixed(-2409.0/65536.0,1,-nbitq), 
to_sfixed(2936.0/65536.0,1,-nbitq), 
to_sfixed(-251.0/65536.0,1,-nbitq), 
to_sfixed(1252.0/65536.0,1,-nbitq), 
to_sfixed(-991.0/65536.0,1,-nbitq), 
to_sfixed(-3624.0/65536.0,1,-nbitq), 
to_sfixed(-2732.0/65536.0,1,-nbitq), 
to_sfixed(-283.0/65536.0,1,-nbitq), 
to_sfixed(1093.0/65536.0,1,-nbitq), 
to_sfixed(1650.0/65536.0,1,-nbitq), 
to_sfixed(-1804.0/65536.0,1,-nbitq), 
to_sfixed(-2375.0/65536.0,1,-nbitq), 
to_sfixed(299.0/65536.0,1,-nbitq), 
to_sfixed(4770.0/65536.0,1,-nbitq), 
to_sfixed(-1932.0/65536.0,1,-nbitq), 
to_sfixed(-2057.0/65536.0,1,-nbitq), 
to_sfixed(3704.0/65536.0,1,-nbitq), 
to_sfixed(216.0/65536.0,1,-nbitq), 
to_sfixed(-995.0/65536.0,1,-nbitq), 
to_sfixed(-77.0/65536.0,1,-nbitq), 
to_sfixed(3471.0/65536.0,1,-nbitq), 
to_sfixed(623.0/65536.0,1,-nbitq), 
to_sfixed(5014.0/65536.0,1,-nbitq), 
to_sfixed(1388.0/65536.0,1,-nbitq), 
to_sfixed(9007.0/65536.0,1,-nbitq), 
to_sfixed(3345.0/65536.0,1,-nbitq), 
to_sfixed(3188.0/65536.0,1,-nbitq), 
to_sfixed(70.0/65536.0,1,-nbitq), 
to_sfixed(1124.0/65536.0,1,-nbitq), 
to_sfixed(1678.0/65536.0,1,-nbitq), 
to_sfixed(870.0/65536.0,1,-nbitq), 
to_sfixed(-2532.0/65536.0,1,-nbitq), 
to_sfixed(-3583.0/65536.0,1,-nbitq), 
to_sfixed(-1781.0/65536.0,1,-nbitq), 
to_sfixed(2097.0/65536.0,1,-nbitq), 
to_sfixed(-4983.0/65536.0,1,-nbitq), 
to_sfixed(-4882.0/65536.0,1,-nbitq), 
to_sfixed(-3251.0/65536.0,1,-nbitq), 
to_sfixed(-342.0/65536.0,1,-nbitq), 
to_sfixed(-4257.0/65536.0,1,-nbitq), 
to_sfixed(9.0/65536.0,1,-nbitq), 
to_sfixed(1160.0/65536.0,1,-nbitq), 
to_sfixed(-440.0/65536.0,1,-nbitq), 
to_sfixed(-134.0/65536.0,1,-nbitq), 
to_sfixed(4651.0/65536.0,1,-nbitq), 
to_sfixed(831.0/65536.0,1,-nbitq), 
to_sfixed(2224.0/65536.0,1,-nbitq), 
to_sfixed(2855.0/65536.0,1,-nbitq), 
to_sfixed(785.0/65536.0,1,-nbitq), 
to_sfixed(-1098.0/65536.0,1,-nbitq), 
to_sfixed(-2603.0/65536.0,1,-nbitq), 
to_sfixed(1231.0/65536.0,1,-nbitq), 
to_sfixed(2613.0/65536.0,1,-nbitq), 
to_sfixed(2153.0/65536.0,1,-nbitq), 
to_sfixed(724.0/65536.0,1,-nbitq), 
to_sfixed(530.0/65536.0,1,-nbitq), 
to_sfixed(2663.0/65536.0,1,-nbitq), 
to_sfixed(1909.0/65536.0,1,-nbitq), 
to_sfixed(3222.0/65536.0,1,-nbitq), 
to_sfixed(51.0/65536.0,1,-nbitq), 
to_sfixed(-760.0/65536.0,1,-nbitq), 
to_sfixed(2195.0/65536.0,1,-nbitq), 
to_sfixed(349.0/65536.0,1,-nbitq), 
to_sfixed(-781.0/65536.0,1,-nbitq), 
to_sfixed(2290.0/65536.0,1,-nbitq), 
to_sfixed(854.0/65536.0,1,-nbitq), 
to_sfixed(-2474.0/65536.0,1,-nbitq), 
to_sfixed(-430.0/65536.0,1,-nbitq), 
to_sfixed(-1192.0/65536.0,1,-nbitq), 
to_sfixed(-2527.0/65536.0,1,-nbitq), 
to_sfixed(-966.0/65536.0,1,-nbitq), 
to_sfixed(1014.0/65536.0,1,-nbitq), 
to_sfixed(-1362.0/65536.0,1,-nbitq), 
to_sfixed(2237.0/65536.0,1,-nbitq), 
to_sfixed(2713.0/65536.0,1,-nbitq), 
to_sfixed(-4068.0/65536.0,1,-nbitq), 
to_sfixed(2455.0/65536.0,1,-nbitq), 
to_sfixed(2379.0/65536.0,1,-nbitq), 
to_sfixed(3071.0/65536.0,1,-nbitq)  ), 
( to_sfixed(675.0/65536.0,1,-nbitq), 
to_sfixed(2752.0/65536.0,1,-nbitq), 
to_sfixed(-148.0/65536.0,1,-nbitq), 
to_sfixed(5996.0/65536.0,1,-nbitq), 
to_sfixed(-1118.0/65536.0,1,-nbitq), 
to_sfixed(2525.0/65536.0,1,-nbitq), 
to_sfixed(-2439.0/65536.0,1,-nbitq), 
to_sfixed(1053.0/65536.0,1,-nbitq), 
to_sfixed(-2590.0/65536.0,1,-nbitq), 
to_sfixed(368.0/65536.0,1,-nbitq), 
to_sfixed(1860.0/65536.0,1,-nbitq), 
to_sfixed(876.0/65536.0,1,-nbitq), 
to_sfixed(-681.0/65536.0,1,-nbitq), 
to_sfixed(2172.0/65536.0,1,-nbitq), 
to_sfixed(37.0/65536.0,1,-nbitq), 
to_sfixed(-569.0/65536.0,1,-nbitq), 
to_sfixed(-564.0/65536.0,1,-nbitq), 
to_sfixed(977.0/65536.0,1,-nbitq), 
to_sfixed(-382.0/65536.0,1,-nbitq), 
to_sfixed(2619.0/65536.0,1,-nbitq), 
to_sfixed(-1511.0/65536.0,1,-nbitq), 
to_sfixed(2266.0/65536.0,1,-nbitq), 
to_sfixed(3571.0/65536.0,1,-nbitq), 
to_sfixed(7884.0/65536.0,1,-nbitq), 
to_sfixed(-352.0/65536.0,1,-nbitq), 
to_sfixed(9384.0/65536.0,1,-nbitq), 
to_sfixed(4162.0/65536.0,1,-nbitq), 
to_sfixed(3917.0/65536.0,1,-nbitq), 
to_sfixed(5158.0/65536.0,1,-nbitq), 
to_sfixed(2443.0/65536.0,1,-nbitq), 
to_sfixed(-2530.0/65536.0,1,-nbitq), 
to_sfixed(558.0/65536.0,1,-nbitq), 
to_sfixed(312.0/65536.0,1,-nbitq), 
to_sfixed(-3528.0/65536.0,1,-nbitq), 
to_sfixed(3496.0/65536.0,1,-nbitq), 
to_sfixed(-1809.0/65536.0,1,-nbitq), 
to_sfixed(-5458.0/65536.0,1,-nbitq), 
to_sfixed(2909.0/65536.0,1,-nbitq), 
to_sfixed(-6622.0/65536.0,1,-nbitq), 
to_sfixed(-3711.0/65536.0,1,-nbitq), 
to_sfixed(3815.0/65536.0,1,-nbitq), 
to_sfixed(-1496.0/65536.0,1,-nbitq), 
to_sfixed(-1879.0/65536.0,1,-nbitq), 
to_sfixed(1904.0/65536.0,1,-nbitq), 
to_sfixed(869.0/65536.0,1,-nbitq), 
to_sfixed(4378.0/65536.0,1,-nbitq), 
to_sfixed(-256.0/65536.0,1,-nbitq), 
to_sfixed(-1548.0/65536.0,1,-nbitq), 
to_sfixed(-2237.0/65536.0,1,-nbitq), 
to_sfixed(2685.0/65536.0,1,-nbitq), 
to_sfixed(-1686.0/65536.0,1,-nbitq), 
to_sfixed(2858.0/65536.0,1,-nbitq), 
to_sfixed(468.0/65536.0,1,-nbitq), 
to_sfixed(2102.0/65536.0,1,-nbitq), 
to_sfixed(-4432.0/65536.0,1,-nbitq), 
to_sfixed(6836.0/65536.0,1,-nbitq), 
to_sfixed(1939.0/65536.0,1,-nbitq), 
to_sfixed(-1654.0/65536.0,1,-nbitq), 
to_sfixed(-1686.0/65536.0,1,-nbitq), 
to_sfixed(-2132.0/65536.0,1,-nbitq), 
to_sfixed(-4284.0/65536.0,1,-nbitq), 
to_sfixed(-927.0/65536.0,1,-nbitq), 
to_sfixed(-2360.0/65536.0,1,-nbitq), 
to_sfixed(-928.0/65536.0,1,-nbitq), 
to_sfixed(4026.0/65536.0,1,-nbitq), 
to_sfixed(2519.0/65536.0,1,-nbitq), 
to_sfixed(93.0/65536.0,1,-nbitq), 
to_sfixed(2493.0/65536.0,1,-nbitq), 
to_sfixed(1909.0/65536.0,1,-nbitq), 
to_sfixed(-2973.0/65536.0,1,-nbitq), 
to_sfixed(505.0/65536.0,1,-nbitq), 
to_sfixed(5.0/65536.0,1,-nbitq), 
to_sfixed(1086.0/65536.0,1,-nbitq), 
to_sfixed(2271.0/65536.0,1,-nbitq), 
to_sfixed(-1911.0/65536.0,1,-nbitq), 
to_sfixed(2973.0/65536.0,1,-nbitq), 
to_sfixed(-1387.0/65536.0,1,-nbitq), 
to_sfixed(-1888.0/65536.0,1,-nbitq), 
to_sfixed(-1076.0/65536.0,1,-nbitq), 
to_sfixed(672.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1337.0/65536.0,1,-nbitq), 
to_sfixed(2394.0/65536.0,1,-nbitq), 
to_sfixed(-1658.0/65536.0,1,-nbitq), 
to_sfixed(3842.0/65536.0,1,-nbitq), 
to_sfixed(-1164.0/65536.0,1,-nbitq), 
to_sfixed(190.0/65536.0,1,-nbitq), 
to_sfixed(-4142.0/65536.0,1,-nbitq), 
to_sfixed(-2479.0/65536.0,1,-nbitq), 
to_sfixed(-3294.0/65536.0,1,-nbitq), 
to_sfixed(-308.0/65536.0,1,-nbitq), 
to_sfixed(5391.0/65536.0,1,-nbitq), 
to_sfixed(2629.0/65536.0,1,-nbitq), 
to_sfixed(71.0/65536.0,1,-nbitq), 
to_sfixed(3163.0/65536.0,1,-nbitq), 
to_sfixed(-2051.0/65536.0,1,-nbitq), 
to_sfixed(1288.0/65536.0,1,-nbitq), 
to_sfixed(1575.0/65536.0,1,-nbitq), 
to_sfixed(-1296.0/65536.0,1,-nbitq), 
to_sfixed(-4129.0/65536.0,1,-nbitq), 
to_sfixed(3014.0/65536.0,1,-nbitq), 
to_sfixed(1381.0/65536.0,1,-nbitq), 
to_sfixed(6781.0/65536.0,1,-nbitq), 
to_sfixed(5232.0/65536.0,1,-nbitq), 
to_sfixed(4330.0/65536.0,1,-nbitq), 
to_sfixed(1885.0/65536.0,1,-nbitq), 
to_sfixed(1106.0/65536.0,1,-nbitq), 
to_sfixed(4150.0/65536.0,1,-nbitq), 
to_sfixed(2082.0/65536.0,1,-nbitq), 
to_sfixed(1510.0/65536.0,1,-nbitq), 
to_sfixed(-2731.0/65536.0,1,-nbitq), 
to_sfixed(-2924.0/65536.0,1,-nbitq), 
to_sfixed(-1319.0/65536.0,1,-nbitq), 
to_sfixed(470.0/65536.0,1,-nbitq), 
to_sfixed(-11297.0/65536.0,1,-nbitq), 
to_sfixed(1886.0/65536.0,1,-nbitq), 
to_sfixed(-352.0/65536.0,1,-nbitq), 
to_sfixed(-8903.0/65536.0,1,-nbitq), 
to_sfixed(3511.0/65536.0,1,-nbitq), 
to_sfixed(-6043.0/65536.0,1,-nbitq), 
to_sfixed(-5327.0/65536.0,1,-nbitq), 
to_sfixed(7081.0/65536.0,1,-nbitq), 
to_sfixed(-2653.0/65536.0,1,-nbitq), 
to_sfixed(-777.0/65536.0,1,-nbitq), 
to_sfixed(388.0/65536.0,1,-nbitq), 
to_sfixed(-392.0/65536.0,1,-nbitq), 
to_sfixed(4526.0/65536.0,1,-nbitq), 
to_sfixed(797.0/65536.0,1,-nbitq), 
to_sfixed(-2805.0/65536.0,1,-nbitq), 
to_sfixed(2711.0/65536.0,1,-nbitq), 
to_sfixed(832.0/65536.0,1,-nbitq), 
to_sfixed(-1484.0/65536.0,1,-nbitq), 
to_sfixed(4799.0/65536.0,1,-nbitq), 
to_sfixed(-954.0/65536.0,1,-nbitq), 
to_sfixed(3807.0/65536.0,1,-nbitq), 
to_sfixed(-6490.0/65536.0,1,-nbitq), 
to_sfixed(11982.0/65536.0,1,-nbitq), 
to_sfixed(424.0/65536.0,1,-nbitq), 
to_sfixed(-2471.0/65536.0,1,-nbitq), 
to_sfixed(-1570.0/65536.0,1,-nbitq), 
to_sfixed(-6436.0/65536.0,1,-nbitq), 
to_sfixed(-6469.0/65536.0,1,-nbitq), 
to_sfixed(215.0/65536.0,1,-nbitq), 
to_sfixed(2637.0/65536.0,1,-nbitq), 
to_sfixed(2283.0/65536.0,1,-nbitq), 
to_sfixed(4160.0/65536.0,1,-nbitq), 
to_sfixed(6401.0/65536.0,1,-nbitq), 
to_sfixed(-1465.0/65536.0,1,-nbitq), 
to_sfixed(3825.0/65536.0,1,-nbitq), 
to_sfixed(1395.0/65536.0,1,-nbitq), 
to_sfixed(-136.0/65536.0,1,-nbitq), 
to_sfixed(-3297.0/65536.0,1,-nbitq), 
to_sfixed(-809.0/65536.0,1,-nbitq), 
to_sfixed(1259.0/65536.0,1,-nbitq), 
to_sfixed(1375.0/65536.0,1,-nbitq), 
to_sfixed(-896.0/65536.0,1,-nbitq), 
to_sfixed(-4105.0/65536.0,1,-nbitq), 
to_sfixed(-4095.0/65536.0,1,-nbitq), 
to_sfixed(-2675.0/65536.0,1,-nbitq), 
to_sfixed(864.0/65536.0,1,-nbitq), 
to_sfixed(685.0/65536.0,1,-nbitq)  ), 
( to_sfixed(640.0/65536.0,1,-nbitq), 
to_sfixed(-4611.0/65536.0,1,-nbitq), 
to_sfixed(5711.0/65536.0,1,-nbitq), 
to_sfixed(1876.0/65536.0,1,-nbitq), 
to_sfixed(3225.0/65536.0,1,-nbitq), 
to_sfixed(-2386.0/65536.0,1,-nbitq), 
to_sfixed(-4959.0/65536.0,1,-nbitq), 
to_sfixed(-6922.0/65536.0,1,-nbitq), 
to_sfixed(-76.0/65536.0,1,-nbitq), 
to_sfixed(-1586.0/65536.0,1,-nbitq), 
to_sfixed(3944.0/65536.0,1,-nbitq), 
to_sfixed(7891.0/65536.0,1,-nbitq), 
to_sfixed(-1526.0/65536.0,1,-nbitq), 
to_sfixed(10236.0/65536.0,1,-nbitq), 
to_sfixed(-7740.0/65536.0,1,-nbitq), 
to_sfixed(-302.0/65536.0,1,-nbitq), 
to_sfixed(-2870.0/65536.0,1,-nbitq), 
to_sfixed(4585.0/65536.0,1,-nbitq), 
to_sfixed(-1636.0/65536.0,1,-nbitq), 
to_sfixed(-146.0/65536.0,1,-nbitq), 
to_sfixed(820.0/65536.0,1,-nbitq), 
to_sfixed(-10534.0/65536.0,1,-nbitq), 
to_sfixed(-2344.0/65536.0,1,-nbitq), 
to_sfixed(-4365.0/65536.0,1,-nbitq), 
to_sfixed(2615.0/65536.0,1,-nbitq), 
to_sfixed(1166.0/65536.0,1,-nbitq), 
to_sfixed(2728.0/65536.0,1,-nbitq), 
to_sfixed(2751.0/65536.0,1,-nbitq), 
to_sfixed(1268.0/65536.0,1,-nbitq), 
to_sfixed(-3676.0/65536.0,1,-nbitq), 
to_sfixed(715.0/65536.0,1,-nbitq), 
to_sfixed(-2553.0/65536.0,1,-nbitq), 
to_sfixed(-3988.0/65536.0,1,-nbitq), 
to_sfixed(-11815.0/65536.0,1,-nbitq), 
to_sfixed(-1636.0/65536.0,1,-nbitq), 
to_sfixed(-1396.0/65536.0,1,-nbitq), 
to_sfixed(-7788.0/65536.0,1,-nbitq), 
to_sfixed(11162.0/65536.0,1,-nbitq), 
to_sfixed(-14748.0/65536.0,1,-nbitq), 
to_sfixed(-10809.0/65536.0,1,-nbitq), 
to_sfixed(9334.0/65536.0,1,-nbitq), 
to_sfixed(2680.0/65536.0,1,-nbitq), 
to_sfixed(-3783.0/65536.0,1,-nbitq), 
to_sfixed(-4231.0/65536.0,1,-nbitq), 
to_sfixed(-113.0/65536.0,1,-nbitq), 
to_sfixed(602.0/65536.0,1,-nbitq), 
to_sfixed(248.0/65536.0,1,-nbitq), 
to_sfixed(-1128.0/65536.0,1,-nbitq), 
to_sfixed(987.0/65536.0,1,-nbitq), 
to_sfixed(1645.0/65536.0,1,-nbitq), 
to_sfixed(-1655.0/65536.0,1,-nbitq), 
to_sfixed(2785.0/65536.0,1,-nbitq), 
to_sfixed(-602.0/65536.0,1,-nbitq), 
to_sfixed(1276.0/65536.0,1,-nbitq), 
to_sfixed(-6736.0/65536.0,1,-nbitq), 
to_sfixed(15306.0/65536.0,1,-nbitq), 
to_sfixed(818.0/65536.0,1,-nbitq), 
to_sfixed(-1246.0/65536.0,1,-nbitq), 
to_sfixed(1044.0/65536.0,1,-nbitq), 
to_sfixed(-1969.0/65536.0,1,-nbitq), 
to_sfixed(-9496.0/65536.0,1,-nbitq), 
to_sfixed(-2227.0/65536.0,1,-nbitq), 
to_sfixed(513.0/65536.0,1,-nbitq), 
to_sfixed(-126.0/65536.0,1,-nbitq), 
to_sfixed(9474.0/65536.0,1,-nbitq), 
to_sfixed(6233.0/65536.0,1,-nbitq), 
to_sfixed(3030.0/65536.0,1,-nbitq), 
to_sfixed(-402.0/65536.0,1,-nbitq), 
to_sfixed(-5307.0/65536.0,1,-nbitq), 
to_sfixed(1409.0/65536.0,1,-nbitq), 
to_sfixed(-309.0/65536.0,1,-nbitq), 
to_sfixed(762.0/65536.0,1,-nbitq), 
to_sfixed(2861.0/65536.0,1,-nbitq), 
to_sfixed(-1708.0/65536.0,1,-nbitq), 
to_sfixed(-2471.0/65536.0,1,-nbitq), 
to_sfixed(-4800.0/65536.0,1,-nbitq), 
to_sfixed(-2824.0/65536.0,1,-nbitq), 
to_sfixed(-4612.0/65536.0,1,-nbitq), 
to_sfixed(936.0/65536.0,1,-nbitq), 
to_sfixed(-3787.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1836.0/65536.0,1,-nbitq), 
to_sfixed(-711.0/65536.0,1,-nbitq), 
to_sfixed(3784.0/65536.0,1,-nbitq), 
to_sfixed(2844.0/65536.0,1,-nbitq), 
to_sfixed(-2552.0/65536.0,1,-nbitq), 
to_sfixed(221.0/65536.0,1,-nbitq), 
to_sfixed(-1349.0/65536.0,1,-nbitq), 
to_sfixed(-10406.0/65536.0,1,-nbitq), 
to_sfixed(2505.0/65536.0,1,-nbitq), 
to_sfixed(-469.0/65536.0,1,-nbitq), 
to_sfixed(5180.0/65536.0,1,-nbitq), 
to_sfixed(16958.0/65536.0,1,-nbitq), 
to_sfixed(1057.0/65536.0,1,-nbitq), 
to_sfixed(8132.0/65536.0,1,-nbitq), 
to_sfixed(-2772.0/65536.0,1,-nbitq), 
to_sfixed(2439.0/65536.0,1,-nbitq), 
to_sfixed(-899.0/65536.0,1,-nbitq), 
to_sfixed(7888.0/65536.0,1,-nbitq), 
to_sfixed(1922.0/65536.0,1,-nbitq), 
to_sfixed(-1627.0/65536.0,1,-nbitq), 
to_sfixed(-6319.0/65536.0,1,-nbitq), 
to_sfixed(-9073.0/65536.0,1,-nbitq), 
to_sfixed(-7608.0/65536.0,1,-nbitq), 
to_sfixed(101.0/65536.0,1,-nbitq), 
to_sfixed(3155.0/65536.0,1,-nbitq), 
to_sfixed(5202.0/65536.0,1,-nbitq), 
to_sfixed(-2839.0/65536.0,1,-nbitq), 
to_sfixed(6581.0/65536.0,1,-nbitq), 
to_sfixed(-2178.0/65536.0,1,-nbitq), 
to_sfixed(-4999.0/65536.0,1,-nbitq), 
to_sfixed(-1475.0/65536.0,1,-nbitq), 
to_sfixed(-4858.0/65536.0,1,-nbitq), 
to_sfixed(-4823.0/65536.0,1,-nbitq), 
to_sfixed(-6795.0/65536.0,1,-nbitq), 
to_sfixed(-3122.0/65536.0,1,-nbitq), 
to_sfixed(-1721.0/65536.0,1,-nbitq), 
to_sfixed(-12973.0/65536.0,1,-nbitq), 
to_sfixed(5712.0/65536.0,1,-nbitq), 
to_sfixed(-13956.0/65536.0,1,-nbitq), 
to_sfixed(-10418.0/65536.0,1,-nbitq), 
to_sfixed(8327.0/65536.0,1,-nbitq), 
to_sfixed(2024.0/65536.0,1,-nbitq), 
to_sfixed(-9695.0/65536.0,1,-nbitq), 
to_sfixed(-920.0/65536.0,1,-nbitq), 
to_sfixed(2924.0/65536.0,1,-nbitq), 
to_sfixed(-192.0/65536.0,1,-nbitq), 
to_sfixed(-2044.0/65536.0,1,-nbitq), 
to_sfixed(4466.0/65536.0,1,-nbitq), 
to_sfixed(3512.0/65536.0,1,-nbitq), 
to_sfixed(-627.0/65536.0,1,-nbitq), 
to_sfixed(305.0/65536.0,1,-nbitq), 
to_sfixed(543.0/65536.0,1,-nbitq), 
to_sfixed(-169.0/65536.0,1,-nbitq), 
to_sfixed(-1741.0/65536.0,1,-nbitq), 
to_sfixed(-6154.0/65536.0,1,-nbitq), 
to_sfixed(10964.0/65536.0,1,-nbitq), 
to_sfixed(-1898.0/65536.0,1,-nbitq), 
to_sfixed(-7132.0/65536.0,1,-nbitq), 
to_sfixed(2205.0/65536.0,1,-nbitq), 
to_sfixed(2608.0/65536.0,1,-nbitq), 
to_sfixed(-734.0/65536.0,1,-nbitq), 
to_sfixed(2122.0/65536.0,1,-nbitq), 
to_sfixed(-542.0/65536.0,1,-nbitq), 
to_sfixed(-1596.0/65536.0,1,-nbitq), 
to_sfixed(9189.0/65536.0,1,-nbitq), 
to_sfixed(4793.0/65536.0,1,-nbitq), 
to_sfixed(4846.0/65536.0,1,-nbitq), 
to_sfixed(11149.0/65536.0,1,-nbitq), 
to_sfixed(-5550.0/65536.0,1,-nbitq), 
to_sfixed(1029.0/65536.0,1,-nbitq), 
to_sfixed(-3180.0/65536.0,1,-nbitq), 
to_sfixed(2477.0/65536.0,1,-nbitq), 
to_sfixed(667.0/65536.0,1,-nbitq), 
to_sfixed(2246.0/65536.0,1,-nbitq), 
to_sfixed(-2504.0/65536.0,1,-nbitq), 
to_sfixed(-4421.0/65536.0,1,-nbitq), 
to_sfixed(3875.0/65536.0,1,-nbitq), 
to_sfixed(-2510.0/65536.0,1,-nbitq), 
to_sfixed(-2116.0/65536.0,1,-nbitq), 
to_sfixed(-1426.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3354.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(4904.0/65536.0,1,-nbitq), 
to_sfixed(7800.0/65536.0,1,-nbitq), 
to_sfixed(-1736.0/65536.0,1,-nbitq), 
to_sfixed(-3033.0/65536.0,1,-nbitq), 
to_sfixed(-3881.0/65536.0,1,-nbitq), 
to_sfixed(-6105.0/65536.0,1,-nbitq), 
to_sfixed(55.0/65536.0,1,-nbitq), 
to_sfixed(-182.0/65536.0,1,-nbitq), 
to_sfixed(3704.0/65536.0,1,-nbitq), 
to_sfixed(3162.0/65536.0,1,-nbitq), 
to_sfixed(1699.0/65536.0,1,-nbitq), 
to_sfixed(3754.0/65536.0,1,-nbitq), 
to_sfixed(-3915.0/65536.0,1,-nbitq), 
to_sfixed(-2559.0/65536.0,1,-nbitq), 
to_sfixed(-939.0/65536.0,1,-nbitq), 
to_sfixed(5504.0/65536.0,1,-nbitq), 
to_sfixed(3867.0/65536.0,1,-nbitq), 
to_sfixed(2096.0/65536.0,1,-nbitq), 
to_sfixed(-9341.0/65536.0,1,-nbitq), 
to_sfixed(-3269.0/65536.0,1,-nbitq), 
to_sfixed(-9996.0/65536.0,1,-nbitq), 
to_sfixed(14791.0/65536.0,1,-nbitq), 
to_sfixed(-5742.0/65536.0,1,-nbitq), 
to_sfixed(4318.0/65536.0,1,-nbitq), 
to_sfixed(-4756.0/65536.0,1,-nbitq), 
to_sfixed(2488.0/65536.0,1,-nbitq), 
to_sfixed(4902.0/65536.0,1,-nbitq), 
to_sfixed(-11042.0/65536.0,1,-nbitq), 
to_sfixed(-1052.0/65536.0,1,-nbitq), 
to_sfixed(1608.0/65536.0,1,-nbitq), 
to_sfixed(-2822.0/65536.0,1,-nbitq), 
to_sfixed(-9677.0/65536.0,1,-nbitq), 
to_sfixed(-2085.0/65536.0,1,-nbitq), 
to_sfixed(1458.0/65536.0,1,-nbitq), 
to_sfixed(-13650.0/65536.0,1,-nbitq), 
to_sfixed(7595.0/65536.0,1,-nbitq), 
to_sfixed(-4981.0/65536.0,1,-nbitq), 
to_sfixed(-3565.0/65536.0,1,-nbitq), 
to_sfixed(13043.0/65536.0,1,-nbitq), 
to_sfixed(-1947.0/65536.0,1,-nbitq), 
to_sfixed(-3015.0/65536.0,1,-nbitq), 
to_sfixed(-1468.0/65536.0,1,-nbitq), 
to_sfixed(2529.0/65536.0,1,-nbitq), 
to_sfixed(-1211.0/65536.0,1,-nbitq), 
to_sfixed(-1525.0/65536.0,1,-nbitq), 
to_sfixed(7092.0/65536.0,1,-nbitq), 
to_sfixed(4595.0/65536.0,1,-nbitq), 
to_sfixed(453.0/65536.0,1,-nbitq), 
to_sfixed(784.0/65536.0,1,-nbitq), 
to_sfixed(2703.0/65536.0,1,-nbitq), 
to_sfixed(-2452.0/65536.0,1,-nbitq), 
to_sfixed(-6903.0/65536.0,1,-nbitq), 
to_sfixed(-3967.0/65536.0,1,-nbitq), 
to_sfixed(3115.0/65536.0,1,-nbitq), 
to_sfixed(2360.0/65536.0,1,-nbitq), 
to_sfixed(-2525.0/65536.0,1,-nbitq), 
to_sfixed(2411.0/65536.0,1,-nbitq), 
to_sfixed(-2571.0/65536.0,1,-nbitq), 
to_sfixed(10820.0/65536.0,1,-nbitq), 
to_sfixed(1209.0/65536.0,1,-nbitq), 
to_sfixed(164.0/65536.0,1,-nbitq), 
to_sfixed(53.0/65536.0,1,-nbitq), 
to_sfixed(6845.0/65536.0,1,-nbitq), 
to_sfixed(2854.0/65536.0,1,-nbitq), 
to_sfixed(2424.0/65536.0,1,-nbitq), 
to_sfixed(15877.0/65536.0,1,-nbitq), 
to_sfixed(1576.0/65536.0,1,-nbitq), 
to_sfixed(2551.0/65536.0,1,-nbitq), 
to_sfixed(-2465.0/65536.0,1,-nbitq), 
to_sfixed(-6743.0/65536.0,1,-nbitq), 
to_sfixed(1106.0/65536.0,1,-nbitq), 
to_sfixed(-531.0/65536.0,1,-nbitq), 
to_sfixed(1654.0/65536.0,1,-nbitq), 
to_sfixed(2784.0/65536.0,1,-nbitq), 
to_sfixed(-2680.0/65536.0,1,-nbitq), 
to_sfixed(-365.0/65536.0,1,-nbitq), 
to_sfixed(-1201.0/65536.0,1,-nbitq), 
to_sfixed(-1505.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3278.0/65536.0,1,-nbitq), 
to_sfixed(5210.0/65536.0,1,-nbitq), 
to_sfixed(-325.0/65536.0,1,-nbitq), 
to_sfixed(5563.0/65536.0,1,-nbitq), 
to_sfixed(-3652.0/65536.0,1,-nbitq), 
to_sfixed(8515.0/65536.0,1,-nbitq), 
to_sfixed(-6148.0/65536.0,1,-nbitq), 
to_sfixed(3250.0/65536.0,1,-nbitq), 
to_sfixed(-1670.0/65536.0,1,-nbitq), 
to_sfixed(-1258.0/65536.0,1,-nbitq), 
to_sfixed(3987.0/65536.0,1,-nbitq), 
to_sfixed(-2667.0/65536.0,1,-nbitq), 
to_sfixed(-2339.0/65536.0,1,-nbitq), 
to_sfixed(2336.0/65536.0,1,-nbitq), 
to_sfixed(128.0/65536.0,1,-nbitq), 
to_sfixed(2127.0/65536.0,1,-nbitq), 
to_sfixed(-1771.0/65536.0,1,-nbitq), 
to_sfixed(6408.0/65536.0,1,-nbitq), 
to_sfixed(1506.0/65536.0,1,-nbitq), 
to_sfixed(-2753.0/65536.0,1,-nbitq), 
to_sfixed(-6456.0/65536.0,1,-nbitq), 
to_sfixed(-3567.0/65536.0,1,-nbitq), 
to_sfixed(-9865.0/65536.0,1,-nbitq), 
to_sfixed(17772.0/65536.0,1,-nbitq), 
to_sfixed(-2086.0/65536.0,1,-nbitq), 
to_sfixed(9706.0/65536.0,1,-nbitq), 
to_sfixed(-2886.0/65536.0,1,-nbitq), 
to_sfixed(6319.0/65536.0,1,-nbitq), 
to_sfixed(6994.0/65536.0,1,-nbitq), 
to_sfixed(-1645.0/65536.0,1,-nbitq), 
to_sfixed(3432.0/65536.0,1,-nbitq), 
to_sfixed(2280.0/65536.0,1,-nbitq), 
to_sfixed(1642.0/65536.0,1,-nbitq), 
to_sfixed(-14186.0/65536.0,1,-nbitq), 
to_sfixed(-415.0/65536.0,1,-nbitq), 
to_sfixed(-231.0/65536.0,1,-nbitq), 
to_sfixed(-3121.0/65536.0,1,-nbitq), 
to_sfixed(2771.0/65536.0,1,-nbitq), 
to_sfixed(-12312.0/65536.0,1,-nbitq), 
to_sfixed(-3485.0/65536.0,1,-nbitq), 
to_sfixed(-3470.0/65536.0,1,-nbitq), 
to_sfixed(-408.0/65536.0,1,-nbitq), 
to_sfixed(850.0/65536.0,1,-nbitq), 
to_sfixed(-860.0/65536.0,1,-nbitq), 
to_sfixed(-2520.0/65536.0,1,-nbitq), 
to_sfixed(-11573.0/65536.0,1,-nbitq), 
to_sfixed(929.0/65536.0,1,-nbitq), 
to_sfixed(9881.0/65536.0,1,-nbitq), 
to_sfixed(4334.0/65536.0,1,-nbitq), 
to_sfixed(2545.0/65536.0,1,-nbitq), 
to_sfixed(-1704.0/65536.0,1,-nbitq), 
to_sfixed(-3051.0/65536.0,1,-nbitq), 
to_sfixed(-2149.0/65536.0,1,-nbitq), 
to_sfixed(-7234.0/65536.0,1,-nbitq), 
to_sfixed(-6197.0/65536.0,1,-nbitq), 
to_sfixed(6570.0/65536.0,1,-nbitq), 
to_sfixed(-1640.0/65536.0,1,-nbitq), 
to_sfixed(15.0/65536.0,1,-nbitq), 
to_sfixed(2209.0/65536.0,1,-nbitq), 
to_sfixed(5279.0/65536.0,1,-nbitq), 
to_sfixed(17152.0/65536.0,1,-nbitq), 
to_sfixed(1290.0/65536.0,1,-nbitq), 
to_sfixed(-2127.0/65536.0,1,-nbitq), 
to_sfixed(-1316.0/65536.0,1,-nbitq), 
to_sfixed(7762.0/65536.0,1,-nbitq), 
to_sfixed(2532.0/65536.0,1,-nbitq), 
to_sfixed(258.0/65536.0,1,-nbitq), 
to_sfixed(5551.0/65536.0,1,-nbitq), 
to_sfixed(-482.0/65536.0,1,-nbitq), 
to_sfixed(1129.0/65536.0,1,-nbitq), 
to_sfixed(474.0/65536.0,1,-nbitq), 
to_sfixed(-9756.0/65536.0,1,-nbitq), 
to_sfixed(1581.0/65536.0,1,-nbitq), 
to_sfixed(-2476.0/65536.0,1,-nbitq), 
to_sfixed(-614.0/65536.0,1,-nbitq), 
to_sfixed(3044.0/65536.0,1,-nbitq), 
to_sfixed(-8762.0/65536.0,1,-nbitq), 
to_sfixed(-8374.0/65536.0,1,-nbitq), 
to_sfixed(-2156.0/65536.0,1,-nbitq), 
to_sfixed(1587.0/65536.0,1,-nbitq)  ), 
( to_sfixed(852.0/65536.0,1,-nbitq), 
to_sfixed(7239.0/65536.0,1,-nbitq), 
to_sfixed(2685.0/65536.0,1,-nbitq), 
to_sfixed(4166.0/65536.0,1,-nbitq), 
to_sfixed(-779.0/65536.0,1,-nbitq), 
to_sfixed(-1952.0/65536.0,1,-nbitq), 
to_sfixed(-2836.0/65536.0,1,-nbitq), 
to_sfixed(9615.0/65536.0,1,-nbitq), 
to_sfixed(-5889.0/65536.0,1,-nbitq), 
to_sfixed(1175.0/65536.0,1,-nbitq), 
to_sfixed(985.0/65536.0,1,-nbitq), 
to_sfixed(-3866.0/65536.0,1,-nbitq), 
to_sfixed(-2423.0/65536.0,1,-nbitq), 
to_sfixed(-662.0/65536.0,1,-nbitq), 
to_sfixed(779.0/65536.0,1,-nbitq), 
to_sfixed(1436.0/65536.0,1,-nbitq), 
to_sfixed(-381.0/65536.0,1,-nbitq), 
to_sfixed(13863.0/65536.0,1,-nbitq), 
to_sfixed(-5771.0/65536.0,1,-nbitq), 
to_sfixed(2228.0/65536.0,1,-nbitq), 
to_sfixed(-2562.0/65536.0,1,-nbitq), 
to_sfixed(-20547.0/65536.0,1,-nbitq), 
to_sfixed(2713.0/65536.0,1,-nbitq), 
to_sfixed(7923.0/65536.0,1,-nbitq), 
to_sfixed(-24.0/65536.0,1,-nbitq), 
to_sfixed(11024.0/65536.0,1,-nbitq), 
to_sfixed(-2337.0/65536.0,1,-nbitq), 
to_sfixed(197.0/65536.0,1,-nbitq), 
to_sfixed(10087.0/65536.0,1,-nbitq), 
to_sfixed(4583.0/65536.0,1,-nbitq), 
to_sfixed(-1073.0/65536.0,1,-nbitq), 
to_sfixed(-2440.0/65536.0,1,-nbitq), 
to_sfixed(1901.0/65536.0,1,-nbitq), 
to_sfixed(-500.0/65536.0,1,-nbitq), 
to_sfixed(-189.0/65536.0,1,-nbitq), 
to_sfixed(390.0/65536.0,1,-nbitq), 
to_sfixed(4398.0/65536.0,1,-nbitq), 
to_sfixed(-3077.0/65536.0,1,-nbitq), 
to_sfixed(-11133.0/65536.0,1,-nbitq), 
to_sfixed(2071.0/65536.0,1,-nbitq), 
to_sfixed(-8857.0/65536.0,1,-nbitq), 
to_sfixed(-2313.0/65536.0,1,-nbitq), 
to_sfixed(4036.0/65536.0,1,-nbitq), 
to_sfixed(-5681.0/65536.0,1,-nbitq), 
to_sfixed(-2993.0/65536.0,1,-nbitq), 
to_sfixed(-13083.0/65536.0,1,-nbitq), 
to_sfixed(1022.0/65536.0,1,-nbitq), 
to_sfixed(6238.0/65536.0,1,-nbitq), 
to_sfixed(1610.0/65536.0,1,-nbitq), 
to_sfixed(709.0/65536.0,1,-nbitq), 
to_sfixed(2761.0/65536.0,1,-nbitq), 
to_sfixed(363.0/65536.0,1,-nbitq), 
to_sfixed(-1261.0/65536.0,1,-nbitq), 
to_sfixed(-2971.0/65536.0,1,-nbitq), 
to_sfixed(-7762.0/65536.0,1,-nbitq), 
to_sfixed(4001.0/65536.0,1,-nbitq), 
to_sfixed(3009.0/65536.0,1,-nbitq), 
to_sfixed(-645.0/65536.0,1,-nbitq), 
to_sfixed(828.0/65536.0,1,-nbitq), 
to_sfixed(5982.0/65536.0,1,-nbitq), 
to_sfixed(17053.0/65536.0,1,-nbitq), 
to_sfixed(2827.0/65536.0,1,-nbitq), 
to_sfixed(-2272.0/65536.0,1,-nbitq), 
to_sfixed(-1145.0/65536.0,1,-nbitq), 
to_sfixed(14842.0/65536.0,1,-nbitq), 
to_sfixed(10692.0/65536.0,1,-nbitq), 
to_sfixed(-3113.0/65536.0,1,-nbitq), 
to_sfixed(717.0/65536.0,1,-nbitq), 
to_sfixed(6929.0/65536.0,1,-nbitq), 
to_sfixed(4490.0/65536.0,1,-nbitq), 
to_sfixed(798.0/65536.0,1,-nbitq), 
to_sfixed(-8485.0/65536.0,1,-nbitq), 
to_sfixed(-3987.0/65536.0,1,-nbitq), 
to_sfixed(-1371.0/65536.0,1,-nbitq), 
to_sfixed(195.0/65536.0,1,-nbitq), 
to_sfixed(2693.0/65536.0,1,-nbitq), 
to_sfixed(-6596.0/65536.0,1,-nbitq), 
to_sfixed(-9563.0/65536.0,1,-nbitq), 
to_sfixed(-1726.0/65536.0,1,-nbitq), 
to_sfixed(-2579.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1032.0/65536.0,1,-nbitq), 
to_sfixed(7159.0/65536.0,1,-nbitq), 
to_sfixed(7217.0/65536.0,1,-nbitq), 
to_sfixed(3155.0/65536.0,1,-nbitq), 
to_sfixed(-5988.0/65536.0,1,-nbitq), 
to_sfixed(-1003.0/65536.0,1,-nbitq), 
to_sfixed(-2011.0/65536.0,1,-nbitq), 
to_sfixed(9811.0/65536.0,1,-nbitq), 
to_sfixed(1513.0/65536.0,1,-nbitq), 
to_sfixed(-1892.0/65536.0,1,-nbitq), 
to_sfixed(4899.0/65536.0,1,-nbitq), 
to_sfixed(-157.0/65536.0,1,-nbitq), 
to_sfixed(-832.0/65536.0,1,-nbitq), 
to_sfixed(-1611.0/65536.0,1,-nbitq), 
to_sfixed(-1419.0/65536.0,1,-nbitq), 
to_sfixed(1455.0/65536.0,1,-nbitq), 
to_sfixed(965.0/65536.0,1,-nbitq), 
to_sfixed(18606.0/65536.0,1,-nbitq), 
to_sfixed(-8619.0/65536.0,1,-nbitq), 
to_sfixed(-25.0/65536.0,1,-nbitq), 
to_sfixed(-5550.0/65536.0,1,-nbitq), 
to_sfixed(-22406.0/65536.0,1,-nbitq), 
to_sfixed(2038.0/65536.0,1,-nbitq), 
to_sfixed(8372.0/65536.0,1,-nbitq), 
to_sfixed(-2997.0/65536.0,1,-nbitq), 
to_sfixed(16486.0/65536.0,1,-nbitq), 
to_sfixed(-2635.0/65536.0,1,-nbitq), 
to_sfixed(516.0/65536.0,1,-nbitq), 
to_sfixed(9814.0/65536.0,1,-nbitq), 
to_sfixed(2753.0/65536.0,1,-nbitq), 
to_sfixed(-2212.0/65536.0,1,-nbitq), 
to_sfixed(120.0/65536.0,1,-nbitq), 
to_sfixed(5012.0/65536.0,1,-nbitq), 
to_sfixed(10544.0/65536.0,1,-nbitq), 
to_sfixed(463.0/65536.0,1,-nbitq), 
to_sfixed(3577.0/65536.0,1,-nbitq), 
to_sfixed(4984.0/65536.0,1,-nbitq), 
to_sfixed(-2057.0/65536.0,1,-nbitq), 
to_sfixed(-3701.0/65536.0,1,-nbitq), 
to_sfixed(587.0/65536.0,1,-nbitq), 
to_sfixed(-1956.0/65536.0,1,-nbitq), 
to_sfixed(1728.0/65536.0,1,-nbitq), 
to_sfixed(2364.0/65536.0,1,-nbitq), 
to_sfixed(-2851.0/65536.0,1,-nbitq), 
to_sfixed(-1844.0/65536.0,1,-nbitq), 
to_sfixed(-9801.0/65536.0,1,-nbitq), 
to_sfixed(-782.0/65536.0,1,-nbitq), 
to_sfixed(-3134.0/65536.0,1,-nbitq), 
to_sfixed(2037.0/65536.0,1,-nbitq), 
to_sfixed(-1706.0/65536.0,1,-nbitq), 
to_sfixed(-1698.0/65536.0,1,-nbitq), 
to_sfixed(-1765.0/65536.0,1,-nbitq), 
to_sfixed(1874.0/65536.0,1,-nbitq), 
to_sfixed(-10422.0/65536.0,1,-nbitq), 
to_sfixed(-5821.0/65536.0,1,-nbitq), 
to_sfixed(5085.0/65536.0,1,-nbitq), 
to_sfixed(304.0/65536.0,1,-nbitq), 
to_sfixed(-1953.0/65536.0,1,-nbitq), 
to_sfixed(-375.0/65536.0,1,-nbitq), 
to_sfixed(8058.0/65536.0,1,-nbitq), 
to_sfixed(12152.0/65536.0,1,-nbitq), 
to_sfixed(2286.0/65536.0,1,-nbitq), 
to_sfixed(-309.0/65536.0,1,-nbitq), 
to_sfixed(-2067.0/65536.0,1,-nbitq), 
to_sfixed(16841.0/65536.0,1,-nbitq), 
to_sfixed(-5966.0/65536.0,1,-nbitq), 
to_sfixed(-4712.0/65536.0,1,-nbitq), 
to_sfixed(728.0/65536.0,1,-nbitq), 
to_sfixed(8124.0/65536.0,1,-nbitq), 
to_sfixed(5618.0/65536.0,1,-nbitq), 
to_sfixed(-4304.0/65536.0,1,-nbitq), 
to_sfixed(-15657.0/65536.0,1,-nbitq), 
to_sfixed(-2764.0/65536.0,1,-nbitq), 
to_sfixed(-2413.0/65536.0,1,-nbitq), 
to_sfixed(-28.0/65536.0,1,-nbitq), 
to_sfixed(-3556.0/65536.0,1,-nbitq), 
to_sfixed(-986.0/65536.0,1,-nbitq), 
to_sfixed(-2140.0/65536.0,1,-nbitq), 
to_sfixed(-1255.0/65536.0,1,-nbitq), 
to_sfixed(-6646.0/65536.0,1,-nbitq)  ), 
( to_sfixed(385.0/65536.0,1,-nbitq), 
to_sfixed(2022.0/65536.0,1,-nbitq), 
to_sfixed(869.0/65536.0,1,-nbitq), 
to_sfixed(-344.0/65536.0,1,-nbitq), 
to_sfixed(-8615.0/65536.0,1,-nbitq), 
to_sfixed(-2227.0/65536.0,1,-nbitq), 
to_sfixed(1880.0/65536.0,1,-nbitq), 
to_sfixed(6875.0/65536.0,1,-nbitq), 
to_sfixed(-3783.0/65536.0,1,-nbitq), 
to_sfixed(483.0/65536.0,1,-nbitq), 
to_sfixed(5303.0/65536.0,1,-nbitq), 
to_sfixed(313.0/65536.0,1,-nbitq), 
to_sfixed(4429.0/65536.0,1,-nbitq), 
to_sfixed(-7565.0/65536.0,1,-nbitq), 
to_sfixed(-7872.0/65536.0,1,-nbitq), 
to_sfixed(-1009.0/65536.0,1,-nbitq), 
to_sfixed(725.0/65536.0,1,-nbitq), 
to_sfixed(-19529.0/65536.0,1,-nbitq), 
to_sfixed(-7699.0/65536.0,1,-nbitq), 
to_sfixed(-2959.0/65536.0,1,-nbitq), 
to_sfixed(-6535.0/65536.0,1,-nbitq), 
to_sfixed(-10197.0/65536.0,1,-nbitq), 
to_sfixed(-10831.0/65536.0,1,-nbitq), 
to_sfixed(10151.0/65536.0,1,-nbitq), 
to_sfixed(2902.0/65536.0,1,-nbitq), 
to_sfixed(4758.0/65536.0,1,-nbitq), 
to_sfixed(-1266.0/65536.0,1,-nbitq), 
to_sfixed(-1063.0/65536.0,1,-nbitq), 
to_sfixed(18924.0/65536.0,1,-nbitq), 
to_sfixed(-324.0/65536.0,1,-nbitq), 
to_sfixed(-2983.0/65536.0,1,-nbitq), 
to_sfixed(-4835.0/65536.0,1,-nbitq), 
to_sfixed(9265.0/65536.0,1,-nbitq), 
to_sfixed(14444.0/65536.0,1,-nbitq), 
to_sfixed(-3083.0/65536.0,1,-nbitq), 
to_sfixed(3413.0/65536.0,1,-nbitq), 
to_sfixed(-883.0/65536.0,1,-nbitq), 
to_sfixed(-2171.0/65536.0,1,-nbitq), 
to_sfixed(-6281.0/65536.0,1,-nbitq), 
to_sfixed(-2085.0/65536.0,1,-nbitq), 
to_sfixed(-737.0/65536.0,1,-nbitq), 
to_sfixed(-1364.0/65536.0,1,-nbitq), 
to_sfixed(2263.0/65536.0,1,-nbitq), 
to_sfixed(-10829.0/65536.0,1,-nbitq), 
to_sfixed(1549.0/65536.0,1,-nbitq), 
to_sfixed(141.0/65536.0,1,-nbitq), 
to_sfixed(-121.0/65536.0,1,-nbitq), 
to_sfixed(-5120.0/65536.0,1,-nbitq), 
to_sfixed(158.0/65536.0,1,-nbitq), 
to_sfixed(-1428.0/65536.0,1,-nbitq), 
to_sfixed(96.0/65536.0,1,-nbitq), 
to_sfixed(-6827.0/65536.0,1,-nbitq), 
to_sfixed(2115.0/65536.0,1,-nbitq), 
to_sfixed(1261.0/65536.0,1,-nbitq), 
to_sfixed(-1861.0/65536.0,1,-nbitq), 
to_sfixed(129.0/65536.0,1,-nbitq), 
to_sfixed(1328.0/65536.0,1,-nbitq), 
to_sfixed(970.0/65536.0,1,-nbitq), 
to_sfixed(-1635.0/65536.0,1,-nbitq), 
to_sfixed(16353.0/65536.0,1,-nbitq), 
to_sfixed(188.0/65536.0,1,-nbitq), 
to_sfixed(1325.0/65536.0,1,-nbitq), 
to_sfixed(-1062.0/65536.0,1,-nbitq), 
to_sfixed(-2041.0/65536.0,1,-nbitq), 
to_sfixed(12612.0/65536.0,1,-nbitq), 
to_sfixed(-26394.0/65536.0,1,-nbitq), 
to_sfixed(-5760.0/65536.0,1,-nbitq), 
to_sfixed(2441.0/65536.0,1,-nbitq), 
to_sfixed(3504.0/65536.0,1,-nbitq), 
to_sfixed(1531.0/65536.0,1,-nbitq), 
to_sfixed(-8128.0/65536.0,1,-nbitq), 
to_sfixed(-14823.0/65536.0,1,-nbitq), 
to_sfixed(1618.0/65536.0,1,-nbitq), 
to_sfixed(-1774.0/65536.0,1,-nbitq), 
to_sfixed(782.0/65536.0,1,-nbitq), 
to_sfixed(-8994.0/65536.0,1,-nbitq), 
to_sfixed(-9847.0/65536.0,1,-nbitq), 
to_sfixed(11370.0/65536.0,1,-nbitq), 
to_sfixed(1097.0/65536.0,1,-nbitq), 
to_sfixed(-5330.0/65536.0,1,-nbitq)  ), 
( to_sfixed(526.0/65536.0,1,-nbitq), 
to_sfixed(-3604.0/65536.0,1,-nbitq), 
to_sfixed(1081.0/65536.0,1,-nbitq), 
to_sfixed(-294.0/65536.0,1,-nbitq), 
to_sfixed(-5497.0/65536.0,1,-nbitq), 
to_sfixed(-2930.0/65536.0,1,-nbitq), 
to_sfixed(-123.0/65536.0,1,-nbitq), 
to_sfixed(7060.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(-36.0/65536.0,1,-nbitq), 
to_sfixed(4833.0/65536.0,1,-nbitq), 
to_sfixed(86.0/65536.0,1,-nbitq), 
to_sfixed(2632.0/65536.0,1,-nbitq), 
to_sfixed(-4199.0/65536.0,1,-nbitq), 
to_sfixed(-10352.0/65536.0,1,-nbitq), 
to_sfixed(433.0/65536.0,1,-nbitq), 
to_sfixed(-736.0/65536.0,1,-nbitq), 
to_sfixed(-16909.0/65536.0,1,-nbitq), 
to_sfixed(-5990.0/65536.0,1,-nbitq), 
to_sfixed(2330.0/65536.0,1,-nbitq), 
to_sfixed(-3007.0/65536.0,1,-nbitq), 
to_sfixed(-3694.0/65536.0,1,-nbitq), 
to_sfixed(-15487.0/65536.0,1,-nbitq), 
to_sfixed(518.0/65536.0,1,-nbitq), 
to_sfixed(7048.0/65536.0,1,-nbitq), 
to_sfixed(12174.0/65536.0,1,-nbitq), 
to_sfixed(-4386.0/65536.0,1,-nbitq), 
to_sfixed(168.0/65536.0,1,-nbitq), 
to_sfixed(2859.0/65536.0,1,-nbitq), 
to_sfixed(-2070.0/65536.0,1,-nbitq), 
to_sfixed(-6320.0/65536.0,1,-nbitq), 
to_sfixed(-1894.0/65536.0,1,-nbitq), 
to_sfixed(8965.0/65536.0,1,-nbitq), 
to_sfixed(3969.0/65536.0,1,-nbitq), 
to_sfixed(-772.0/65536.0,1,-nbitq), 
to_sfixed(4052.0/65536.0,1,-nbitq), 
to_sfixed(-4582.0/65536.0,1,-nbitq), 
to_sfixed(-1405.0/65536.0,1,-nbitq), 
to_sfixed(1417.0/65536.0,1,-nbitq), 
to_sfixed(-251.0/65536.0,1,-nbitq), 
to_sfixed(-184.0/65536.0,1,-nbitq), 
to_sfixed(-861.0/65536.0,1,-nbitq), 
to_sfixed(4853.0/65536.0,1,-nbitq), 
to_sfixed(-10012.0/65536.0,1,-nbitq), 
to_sfixed(-2547.0/65536.0,1,-nbitq), 
to_sfixed(11326.0/65536.0,1,-nbitq), 
to_sfixed(-253.0/65536.0,1,-nbitq), 
to_sfixed(-5283.0/65536.0,1,-nbitq), 
to_sfixed(1508.0/65536.0,1,-nbitq), 
to_sfixed(423.0/65536.0,1,-nbitq), 
to_sfixed(-2580.0/65536.0,1,-nbitq), 
to_sfixed(-4153.0/65536.0,1,-nbitq), 
to_sfixed(6918.0/65536.0,1,-nbitq), 
to_sfixed(-374.0/65536.0,1,-nbitq), 
to_sfixed(-1493.0/65536.0,1,-nbitq), 
to_sfixed(10794.0/65536.0,1,-nbitq), 
to_sfixed(-1609.0/65536.0,1,-nbitq), 
to_sfixed(3128.0/65536.0,1,-nbitq), 
to_sfixed(-2421.0/65536.0,1,-nbitq), 
to_sfixed(21029.0/65536.0,1,-nbitq), 
to_sfixed(-3519.0/65536.0,1,-nbitq), 
to_sfixed(-2089.0/65536.0,1,-nbitq), 
to_sfixed(-2495.0/65536.0,1,-nbitq), 
to_sfixed(-2662.0/65536.0,1,-nbitq), 
to_sfixed(8063.0/65536.0,1,-nbitq), 
to_sfixed(-24183.0/65536.0,1,-nbitq), 
to_sfixed(-210.0/65536.0,1,-nbitq), 
to_sfixed(-179.0/65536.0,1,-nbitq), 
to_sfixed(3921.0/65536.0,1,-nbitq), 
to_sfixed(3839.0/65536.0,1,-nbitq), 
to_sfixed(-6017.0/65536.0,1,-nbitq), 
to_sfixed(-2694.0/65536.0,1,-nbitq), 
to_sfixed(-849.0/65536.0,1,-nbitq), 
to_sfixed(-2841.0/65536.0,1,-nbitq), 
to_sfixed(971.0/65536.0,1,-nbitq), 
to_sfixed(-19472.0/65536.0,1,-nbitq), 
to_sfixed(-6436.0/65536.0,1,-nbitq), 
to_sfixed(4309.0/65536.0,1,-nbitq), 
to_sfixed(-2509.0/65536.0,1,-nbitq), 
to_sfixed(-1514.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-792.0/65536.0,1,-nbitq), 
to_sfixed(-7292.0/65536.0,1,-nbitq), 
to_sfixed(-5494.0/65536.0,1,-nbitq), 
to_sfixed(-139.0/65536.0,1,-nbitq), 
to_sfixed(-1981.0/65536.0,1,-nbitq), 
to_sfixed(-7153.0/65536.0,1,-nbitq), 
to_sfixed(-887.0/65536.0,1,-nbitq), 
to_sfixed(1605.0/65536.0,1,-nbitq), 
to_sfixed(-2687.0/65536.0,1,-nbitq), 
to_sfixed(1524.0/65536.0,1,-nbitq), 
to_sfixed(451.0/65536.0,1,-nbitq), 
to_sfixed(7712.0/65536.0,1,-nbitq), 
to_sfixed(3968.0/65536.0,1,-nbitq), 
to_sfixed(1581.0/65536.0,1,-nbitq), 
to_sfixed(-2156.0/65536.0,1,-nbitq), 
to_sfixed(-2251.0/65536.0,1,-nbitq), 
to_sfixed(495.0/65536.0,1,-nbitq), 
to_sfixed(-4150.0/65536.0,1,-nbitq), 
to_sfixed(-9514.0/65536.0,1,-nbitq), 
to_sfixed(-781.0/65536.0,1,-nbitq), 
to_sfixed(3843.0/65536.0,1,-nbitq), 
to_sfixed(-7932.0/65536.0,1,-nbitq), 
to_sfixed(-17050.0/65536.0,1,-nbitq), 
to_sfixed(3698.0/65536.0,1,-nbitq), 
to_sfixed(6698.0/65536.0,1,-nbitq), 
to_sfixed(9059.0/65536.0,1,-nbitq), 
to_sfixed(2145.0/65536.0,1,-nbitq), 
to_sfixed(-3863.0/65536.0,1,-nbitq), 
to_sfixed(-335.0/65536.0,1,-nbitq), 
to_sfixed(-6989.0/65536.0,1,-nbitq), 
to_sfixed(-3199.0/65536.0,1,-nbitq), 
to_sfixed(11060.0/65536.0,1,-nbitq), 
to_sfixed(2542.0/65536.0,1,-nbitq), 
to_sfixed(-6822.0/65536.0,1,-nbitq), 
to_sfixed(2362.0/65536.0,1,-nbitq), 
to_sfixed(-3221.0/65536.0,1,-nbitq), 
to_sfixed(-11223.0/65536.0,1,-nbitq), 
to_sfixed(2142.0/65536.0,1,-nbitq), 
to_sfixed(18566.0/65536.0,1,-nbitq), 
to_sfixed(1993.0/65536.0,1,-nbitq), 
to_sfixed(-3593.0/65536.0,1,-nbitq), 
to_sfixed(1277.0/65536.0,1,-nbitq), 
to_sfixed(9565.0/65536.0,1,-nbitq), 
to_sfixed(-8393.0/65536.0,1,-nbitq), 
to_sfixed(-1994.0/65536.0,1,-nbitq), 
to_sfixed(6857.0/65536.0,1,-nbitq), 
to_sfixed(-3434.0/65536.0,1,-nbitq), 
to_sfixed(-1655.0/65536.0,1,-nbitq), 
to_sfixed(1665.0/65536.0,1,-nbitq), 
to_sfixed(2431.0/65536.0,1,-nbitq), 
to_sfixed(2647.0/65536.0,1,-nbitq), 
to_sfixed(-1701.0/65536.0,1,-nbitq), 
to_sfixed(8330.0/65536.0,1,-nbitq), 
to_sfixed(-5797.0/65536.0,1,-nbitq), 
to_sfixed(-4072.0/65536.0,1,-nbitq), 
to_sfixed(696.0/65536.0,1,-nbitq), 
to_sfixed(127.0/65536.0,1,-nbitq), 
to_sfixed(3726.0/65536.0,1,-nbitq), 
to_sfixed(285.0/65536.0,1,-nbitq), 
to_sfixed(9500.0/65536.0,1,-nbitq), 
to_sfixed(-5887.0/65536.0,1,-nbitq), 
to_sfixed(2033.0/65536.0,1,-nbitq), 
to_sfixed(1476.0/65536.0,1,-nbitq), 
to_sfixed(298.0/65536.0,1,-nbitq), 
to_sfixed(1144.0/65536.0,1,-nbitq), 
to_sfixed(-9403.0/65536.0,1,-nbitq), 
to_sfixed(-3272.0/65536.0,1,-nbitq), 
to_sfixed(-2957.0/65536.0,1,-nbitq), 
to_sfixed(-4151.0/65536.0,1,-nbitq), 
to_sfixed(2724.0/65536.0,1,-nbitq), 
to_sfixed(-5163.0/65536.0,1,-nbitq), 
to_sfixed(677.0/65536.0,1,-nbitq), 
to_sfixed(-12447.0/65536.0,1,-nbitq), 
to_sfixed(2221.0/65536.0,1,-nbitq), 
to_sfixed(185.0/65536.0,1,-nbitq), 
to_sfixed(-12229.0/65536.0,1,-nbitq), 
to_sfixed(-6373.0/65536.0,1,-nbitq), 
to_sfixed(-1188.0/65536.0,1,-nbitq), 
to_sfixed(-2050.0/65536.0,1,-nbitq), 
to_sfixed(4251.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2434.0/65536.0,1,-nbitq), 
to_sfixed(-2952.0/65536.0,1,-nbitq), 
to_sfixed(-806.0/65536.0,1,-nbitq), 
to_sfixed(-1285.0/65536.0,1,-nbitq), 
to_sfixed(-4265.0/65536.0,1,-nbitq), 
to_sfixed(80.0/65536.0,1,-nbitq), 
to_sfixed(3335.0/65536.0,1,-nbitq), 
to_sfixed(-13609.0/65536.0,1,-nbitq), 
to_sfixed(-3284.0/65536.0,1,-nbitq), 
to_sfixed(1733.0/65536.0,1,-nbitq), 
to_sfixed(-3643.0/65536.0,1,-nbitq), 
to_sfixed(15787.0/65536.0,1,-nbitq), 
to_sfixed(5879.0/65536.0,1,-nbitq), 
to_sfixed(4064.0/65536.0,1,-nbitq), 
to_sfixed(1420.0/65536.0,1,-nbitq), 
to_sfixed(-1535.0/65536.0,1,-nbitq), 
to_sfixed(-1984.0/65536.0,1,-nbitq), 
to_sfixed(566.0/65536.0,1,-nbitq), 
to_sfixed(-1638.0/65536.0,1,-nbitq), 
to_sfixed(1678.0/65536.0,1,-nbitq), 
to_sfixed(897.0/65536.0,1,-nbitq), 
to_sfixed(-2565.0/65536.0,1,-nbitq), 
to_sfixed(-17393.0/65536.0,1,-nbitq), 
to_sfixed(-1635.0/65536.0,1,-nbitq), 
to_sfixed(8700.0/65536.0,1,-nbitq), 
to_sfixed(2580.0/65536.0,1,-nbitq), 
to_sfixed(-6401.0/65536.0,1,-nbitq), 
to_sfixed(-2653.0/65536.0,1,-nbitq), 
to_sfixed(5201.0/65536.0,1,-nbitq), 
to_sfixed(-7753.0/65536.0,1,-nbitq), 
to_sfixed(4236.0/65536.0,1,-nbitq), 
to_sfixed(9181.0/65536.0,1,-nbitq), 
to_sfixed(-3027.0/65536.0,1,-nbitq), 
to_sfixed(-17203.0/65536.0,1,-nbitq), 
to_sfixed(-701.0/65536.0,1,-nbitq), 
to_sfixed(-2528.0/65536.0,1,-nbitq), 
to_sfixed(-2711.0/65536.0,1,-nbitq), 
to_sfixed(9350.0/65536.0,1,-nbitq), 
to_sfixed(8991.0/65536.0,1,-nbitq), 
to_sfixed(-138.0/65536.0,1,-nbitq), 
to_sfixed(4207.0/65536.0,1,-nbitq), 
to_sfixed(-1223.0/65536.0,1,-nbitq), 
to_sfixed(4705.0/65536.0,1,-nbitq), 
to_sfixed(-5459.0/65536.0,1,-nbitq), 
to_sfixed(3281.0/65536.0,1,-nbitq), 
to_sfixed(7450.0/65536.0,1,-nbitq), 
to_sfixed(341.0/65536.0,1,-nbitq), 
to_sfixed(-8381.0/65536.0,1,-nbitq), 
to_sfixed(2461.0/65536.0,1,-nbitq), 
to_sfixed(1035.0/65536.0,1,-nbitq), 
to_sfixed(-985.0/65536.0,1,-nbitq), 
to_sfixed(-10351.0/65536.0,1,-nbitq), 
to_sfixed(11259.0/65536.0,1,-nbitq), 
to_sfixed(-2292.0/65536.0,1,-nbitq), 
to_sfixed(10145.0/65536.0,1,-nbitq), 
to_sfixed(-14668.0/65536.0,1,-nbitq), 
to_sfixed(1730.0/65536.0,1,-nbitq), 
to_sfixed(1899.0/65536.0,1,-nbitq), 
to_sfixed(428.0/65536.0,1,-nbitq), 
to_sfixed(-2918.0/65536.0,1,-nbitq), 
to_sfixed(-8811.0/65536.0,1,-nbitq), 
to_sfixed(2395.0/65536.0,1,-nbitq), 
to_sfixed(-2347.0/65536.0,1,-nbitq), 
to_sfixed(1238.0/65536.0,1,-nbitq), 
to_sfixed(-2217.0/65536.0,1,-nbitq), 
to_sfixed(-4394.0/65536.0,1,-nbitq), 
to_sfixed(-1909.0/65536.0,1,-nbitq), 
to_sfixed(-6081.0/65536.0,1,-nbitq), 
to_sfixed(-5326.0/65536.0,1,-nbitq), 
to_sfixed(2304.0/65536.0,1,-nbitq), 
to_sfixed(-977.0/65536.0,1,-nbitq), 
to_sfixed(-1687.0/65536.0,1,-nbitq), 
to_sfixed(-14248.0/65536.0,1,-nbitq), 
to_sfixed(-761.0/65536.0,1,-nbitq), 
to_sfixed(-1112.0/65536.0,1,-nbitq), 
to_sfixed(2272.0/65536.0,1,-nbitq), 
to_sfixed(-7608.0/65536.0,1,-nbitq), 
to_sfixed(2018.0/65536.0,1,-nbitq), 
to_sfixed(888.0/65536.0,1,-nbitq), 
to_sfixed(10027.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2085.0/65536.0,1,-nbitq), 
to_sfixed(-6472.0/65536.0,1,-nbitq), 
to_sfixed(5353.0/65536.0,1,-nbitq), 
to_sfixed(2440.0/65536.0,1,-nbitq), 
to_sfixed(-2800.0/65536.0,1,-nbitq), 
to_sfixed(14513.0/65536.0,1,-nbitq), 
to_sfixed(11.0/65536.0,1,-nbitq), 
to_sfixed(-17691.0/65536.0,1,-nbitq), 
to_sfixed(-4671.0/65536.0,1,-nbitq), 
to_sfixed(-1977.0/65536.0,1,-nbitq), 
to_sfixed(-1287.0/65536.0,1,-nbitq), 
to_sfixed(6398.0/65536.0,1,-nbitq), 
to_sfixed(5067.0/65536.0,1,-nbitq), 
to_sfixed(5236.0/65536.0,1,-nbitq), 
to_sfixed(1225.0/65536.0,1,-nbitq), 
to_sfixed(-253.0/65536.0,1,-nbitq), 
to_sfixed(161.0/65536.0,1,-nbitq), 
to_sfixed(1509.0/65536.0,1,-nbitq), 
to_sfixed(648.0/65536.0,1,-nbitq), 
to_sfixed(-1050.0/65536.0,1,-nbitq), 
to_sfixed(-500.0/65536.0,1,-nbitq), 
to_sfixed(-1670.0/65536.0,1,-nbitq), 
to_sfixed(-18340.0/65536.0,1,-nbitq), 
to_sfixed(-2474.0/65536.0,1,-nbitq), 
to_sfixed(9564.0/65536.0,1,-nbitq), 
to_sfixed(-5415.0/65536.0,1,-nbitq), 
to_sfixed(-737.0/65536.0,1,-nbitq), 
to_sfixed(4108.0/65536.0,1,-nbitq), 
to_sfixed(2939.0/65536.0,1,-nbitq), 
to_sfixed(-3501.0/65536.0,1,-nbitq), 
to_sfixed(2761.0/65536.0,1,-nbitq), 
to_sfixed(5985.0/65536.0,1,-nbitq), 
to_sfixed(-2642.0/65536.0,1,-nbitq), 
to_sfixed(-15174.0/65536.0,1,-nbitq), 
to_sfixed(635.0/65536.0,1,-nbitq), 
to_sfixed(-2974.0/65536.0,1,-nbitq), 
to_sfixed(-8290.0/65536.0,1,-nbitq), 
to_sfixed(5874.0/65536.0,1,-nbitq), 
to_sfixed(-2855.0/65536.0,1,-nbitq), 
to_sfixed(1137.0/65536.0,1,-nbitq), 
to_sfixed(14411.0/65536.0,1,-nbitq), 
to_sfixed(-1717.0/65536.0,1,-nbitq), 
to_sfixed(863.0/65536.0,1,-nbitq), 
to_sfixed(2046.0/65536.0,1,-nbitq), 
to_sfixed(-2250.0/65536.0,1,-nbitq), 
to_sfixed(1604.0/65536.0,1,-nbitq), 
to_sfixed(1505.0/65536.0,1,-nbitq), 
to_sfixed(440.0/65536.0,1,-nbitq), 
to_sfixed(-614.0/65536.0,1,-nbitq), 
to_sfixed(3896.0/65536.0,1,-nbitq), 
to_sfixed(2933.0/65536.0,1,-nbitq), 
to_sfixed(-10217.0/65536.0,1,-nbitq), 
to_sfixed(10673.0/65536.0,1,-nbitq), 
to_sfixed(10374.0/65536.0,1,-nbitq), 
to_sfixed(17196.0/65536.0,1,-nbitq), 
to_sfixed(-14636.0/65536.0,1,-nbitq), 
to_sfixed(1759.0/65536.0,1,-nbitq), 
to_sfixed(-2086.0/65536.0,1,-nbitq), 
to_sfixed(129.0/65536.0,1,-nbitq), 
to_sfixed(-3178.0/65536.0,1,-nbitq), 
to_sfixed(-5513.0/65536.0,1,-nbitq), 
to_sfixed(2573.0/65536.0,1,-nbitq), 
to_sfixed(-2222.0/65536.0,1,-nbitq), 
to_sfixed(-590.0/65536.0,1,-nbitq), 
to_sfixed(-5163.0/65536.0,1,-nbitq), 
to_sfixed(-9423.0/65536.0,1,-nbitq), 
to_sfixed(319.0/65536.0,1,-nbitq), 
to_sfixed(-4275.0/65536.0,1,-nbitq), 
to_sfixed(-674.0/65536.0,1,-nbitq), 
to_sfixed(3085.0/65536.0,1,-nbitq), 
to_sfixed(-3526.0/65536.0,1,-nbitq), 
to_sfixed(-1266.0/65536.0,1,-nbitq), 
to_sfixed(8228.0/65536.0,1,-nbitq), 
to_sfixed(-1614.0/65536.0,1,-nbitq), 
to_sfixed(-845.0/65536.0,1,-nbitq), 
to_sfixed(13709.0/65536.0,1,-nbitq), 
to_sfixed(-6995.0/65536.0,1,-nbitq), 
to_sfixed(-1385.0/65536.0,1,-nbitq), 
to_sfixed(249.0/65536.0,1,-nbitq), 
to_sfixed(13019.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1789.0/65536.0,1,-nbitq), 
to_sfixed(-1520.0/65536.0,1,-nbitq), 
to_sfixed(-1562.0/65536.0,1,-nbitq), 
to_sfixed(285.0/65536.0,1,-nbitq), 
to_sfixed(2334.0/65536.0,1,-nbitq), 
to_sfixed(14233.0/65536.0,1,-nbitq), 
to_sfixed(-886.0/65536.0,1,-nbitq), 
to_sfixed(-12629.0/65536.0,1,-nbitq), 
to_sfixed(2704.0/65536.0,1,-nbitq), 
to_sfixed(1089.0/65536.0,1,-nbitq), 
to_sfixed(-2681.0/65536.0,1,-nbitq), 
to_sfixed(3414.0/65536.0,1,-nbitq), 
to_sfixed(5645.0/65536.0,1,-nbitq), 
to_sfixed(8148.0/65536.0,1,-nbitq), 
to_sfixed(-3567.0/65536.0,1,-nbitq), 
to_sfixed(1965.0/65536.0,1,-nbitq), 
to_sfixed(3087.0/65536.0,1,-nbitq), 
to_sfixed(4591.0/65536.0,1,-nbitq), 
to_sfixed(1336.0/65536.0,1,-nbitq), 
to_sfixed(-646.0/65536.0,1,-nbitq), 
to_sfixed(-4248.0/65536.0,1,-nbitq), 
to_sfixed(2190.0/65536.0,1,-nbitq), 
to_sfixed(-17483.0/65536.0,1,-nbitq), 
to_sfixed(-1197.0/65536.0,1,-nbitq), 
to_sfixed(6994.0/65536.0,1,-nbitq), 
to_sfixed(-4749.0/65536.0,1,-nbitq), 
to_sfixed(-8148.0/65536.0,1,-nbitq), 
to_sfixed(2889.0/65536.0,1,-nbitq), 
to_sfixed(855.0/65536.0,1,-nbitq), 
to_sfixed(4447.0/65536.0,1,-nbitq), 
to_sfixed(2012.0/65536.0,1,-nbitq), 
to_sfixed(-654.0/65536.0,1,-nbitq), 
to_sfixed(-4858.0/65536.0,1,-nbitq), 
to_sfixed(-6419.0/65536.0,1,-nbitq), 
to_sfixed(-2946.0/65536.0,1,-nbitq), 
to_sfixed(-2999.0/65536.0,1,-nbitq), 
to_sfixed(2235.0/65536.0,1,-nbitq), 
to_sfixed(658.0/65536.0,1,-nbitq), 
to_sfixed(-4738.0/65536.0,1,-nbitq), 
to_sfixed(1314.0/65536.0,1,-nbitq), 
to_sfixed(12326.0/65536.0,1,-nbitq), 
to_sfixed(-990.0/65536.0,1,-nbitq), 
to_sfixed(3685.0/65536.0,1,-nbitq), 
to_sfixed(4241.0/65536.0,1,-nbitq), 
to_sfixed(-874.0/65536.0,1,-nbitq), 
to_sfixed(-7174.0/65536.0,1,-nbitq), 
to_sfixed(1214.0/65536.0,1,-nbitq), 
to_sfixed(5582.0/65536.0,1,-nbitq), 
to_sfixed(4824.0/65536.0,1,-nbitq), 
to_sfixed(2650.0/65536.0,1,-nbitq), 
to_sfixed(-2645.0/65536.0,1,-nbitq), 
to_sfixed(-8023.0/65536.0,1,-nbitq), 
to_sfixed(10839.0/65536.0,1,-nbitq), 
to_sfixed(13034.0/65536.0,1,-nbitq), 
to_sfixed(6662.0/65536.0,1,-nbitq), 
to_sfixed(-10397.0/65536.0,1,-nbitq), 
to_sfixed(2453.0/65536.0,1,-nbitq), 
to_sfixed(-5113.0/65536.0,1,-nbitq), 
to_sfixed(-841.0/65536.0,1,-nbitq), 
to_sfixed(-3367.0/65536.0,1,-nbitq), 
to_sfixed(-4761.0/65536.0,1,-nbitq), 
to_sfixed(-2202.0/65536.0,1,-nbitq), 
to_sfixed(-1691.0/65536.0,1,-nbitq), 
to_sfixed(1881.0/65536.0,1,-nbitq), 
to_sfixed(-4700.0/65536.0,1,-nbitq), 
to_sfixed(-1832.0/65536.0,1,-nbitq), 
to_sfixed(-1779.0/65536.0,1,-nbitq), 
to_sfixed(-1159.0/65536.0,1,-nbitq), 
to_sfixed(1343.0/65536.0,1,-nbitq), 
to_sfixed(14133.0/65536.0,1,-nbitq), 
to_sfixed(5115.0/65536.0,1,-nbitq), 
to_sfixed(5653.0/65536.0,1,-nbitq), 
to_sfixed(10761.0/65536.0,1,-nbitq), 
to_sfixed(1975.0/65536.0,1,-nbitq), 
to_sfixed(-2216.0/65536.0,1,-nbitq), 
to_sfixed(4307.0/65536.0,1,-nbitq), 
to_sfixed(-12419.0/65536.0,1,-nbitq), 
to_sfixed(-11750.0/65536.0,1,-nbitq), 
to_sfixed(1317.0/65536.0,1,-nbitq), 
to_sfixed(5475.0/65536.0,1,-nbitq)  ), 
( to_sfixed(6420.0/65536.0,1,-nbitq), 
to_sfixed(2245.0/65536.0,1,-nbitq), 
to_sfixed(2170.0/65536.0,1,-nbitq), 
to_sfixed(732.0/65536.0,1,-nbitq), 
to_sfixed(6112.0/65536.0,1,-nbitq), 
to_sfixed(14084.0/65536.0,1,-nbitq), 
to_sfixed(-1906.0/65536.0,1,-nbitq), 
to_sfixed(-13108.0/65536.0,1,-nbitq), 
to_sfixed(3776.0/65536.0,1,-nbitq), 
to_sfixed(2021.0/65536.0,1,-nbitq), 
to_sfixed(-429.0/65536.0,1,-nbitq), 
to_sfixed(-1644.0/65536.0,1,-nbitq), 
to_sfixed(2546.0/65536.0,1,-nbitq), 
to_sfixed(4429.0/65536.0,1,-nbitq), 
to_sfixed(1909.0/65536.0,1,-nbitq), 
to_sfixed(-956.0/65536.0,1,-nbitq), 
to_sfixed(-1127.0/65536.0,1,-nbitq), 
to_sfixed(4397.0/65536.0,1,-nbitq), 
to_sfixed(-2206.0/65536.0,1,-nbitq), 
to_sfixed(-800.0/65536.0,1,-nbitq), 
to_sfixed(238.0/65536.0,1,-nbitq), 
to_sfixed(5713.0/65536.0,1,-nbitq), 
to_sfixed(-4616.0/65536.0,1,-nbitq), 
to_sfixed(475.0/65536.0,1,-nbitq), 
to_sfixed(9102.0/65536.0,1,-nbitq), 
to_sfixed(-5471.0/65536.0,1,-nbitq), 
to_sfixed(-8668.0/65536.0,1,-nbitq), 
to_sfixed(408.0/65536.0,1,-nbitq), 
to_sfixed(2698.0/65536.0,1,-nbitq), 
to_sfixed(1194.0/65536.0,1,-nbitq), 
to_sfixed(-3853.0/65536.0,1,-nbitq), 
to_sfixed(-3205.0/65536.0,1,-nbitq), 
to_sfixed(-4019.0/65536.0,1,-nbitq), 
to_sfixed(-7322.0/65536.0,1,-nbitq), 
to_sfixed(-1770.0/65536.0,1,-nbitq), 
to_sfixed(-985.0/65536.0,1,-nbitq), 
to_sfixed(-6200.0/65536.0,1,-nbitq), 
to_sfixed(2460.0/65536.0,1,-nbitq), 
to_sfixed(-11119.0/65536.0,1,-nbitq), 
to_sfixed(633.0/65536.0,1,-nbitq), 
to_sfixed(10032.0/65536.0,1,-nbitq), 
to_sfixed(-550.0/65536.0,1,-nbitq), 
to_sfixed(-2393.0/65536.0,1,-nbitq), 
to_sfixed(4126.0/65536.0,1,-nbitq), 
to_sfixed(-1542.0/65536.0,1,-nbitq), 
to_sfixed(-9917.0/65536.0,1,-nbitq), 
to_sfixed(823.0/65536.0,1,-nbitq), 
to_sfixed(4523.0/65536.0,1,-nbitq), 
to_sfixed(1642.0/65536.0,1,-nbitq), 
to_sfixed(2268.0/65536.0,1,-nbitq), 
to_sfixed(1131.0/65536.0,1,-nbitq), 
to_sfixed(867.0/65536.0,1,-nbitq), 
to_sfixed(8478.0/65536.0,1,-nbitq), 
to_sfixed(19761.0/65536.0,1,-nbitq), 
to_sfixed(2067.0/65536.0,1,-nbitq), 
to_sfixed(-12796.0/65536.0,1,-nbitq), 
to_sfixed(-1608.0/65536.0,1,-nbitq), 
to_sfixed(-91.0/65536.0,1,-nbitq), 
to_sfixed(685.0/65536.0,1,-nbitq), 
to_sfixed(-5508.0/65536.0,1,-nbitq), 
to_sfixed(5258.0/65536.0,1,-nbitq), 
to_sfixed(493.0/65536.0,1,-nbitq), 
to_sfixed(-1969.0/65536.0,1,-nbitq), 
to_sfixed(912.0/65536.0,1,-nbitq), 
to_sfixed(-2578.0/65536.0,1,-nbitq), 
to_sfixed(-3067.0/65536.0,1,-nbitq), 
to_sfixed(-4109.0/65536.0,1,-nbitq), 
to_sfixed(-4880.0/65536.0,1,-nbitq), 
to_sfixed(980.0/65536.0,1,-nbitq), 
to_sfixed(13663.0/65536.0,1,-nbitq), 
to_sfixed(5645.0/65536.0,1,-nbitq), 
to_sfixed(9849.0/65536.0,1,-nbitq), 
to_sfixed(5129.0/65536.0,1,-nbitq), 
to_sfixed(-2203.0/65536.0,1,-nbitq), 
to_sfixed(-1108.0/65536.0,1,-nbitq), 
to_sfixed(-1713.0/65536.0,1,-nbitq), 
to_sfixed(-9266.0/65536.0,1,-nbitq), 
to_sfixed(-10558.0/65536.0,1,-nbitq), 
to_sfixed(-653.0/65536.0,1,-nbitq), 
to_sfixed(-2268.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3727.0/65536.0,1,-nbitq), 
to_sfixed(-179.0/65536.0,1,-nbitq), 
to_sfixed(-3378.0/65536.0,1,-nbitq), 
to_sfixed(4190.0/65536.0,1,-nbitq), 
to_sfixed(-3258.0/65536.0,1,-nbitq), 
to_sfixed(6131.0/65536.0,1,-nbitq), 
to_sfixed(1450.0/65536.0,1,-nbitq), 
to_sfixed(-5703.0/65536.0,1,-nbitq), 
to_sfixed(3941.0/65536.0,1,-nbitq), 
to_sfixed(1904.0/65536.0,1,-nbitq), 
to_sfixed(-3936.0/65536.0,1,-nbitq), 
to_sfixed(3768.0/65536.0,1,-nbitq), 
to_sfixed(3695.0/65536.0,1,-nbitq), 
to_sfixed(1232.0/65536.0,1,-nbitq), 
to_sfixed(-4608.0/65536.0,1,-nbitq), 
to_sfixed(-1450.0/65536.0,1,-nbitq), 
to_sfixed(-789.0/65536.0,1,-nbitq), 
to_sfixed(-542.0/65536.0,1,-nbitq), 
to_sfixed(399.0/65536.0,1,-nbitq), 
to_sfixed(1382.0/65536.0,1,-nbitq), 
to_sfixed(-600.0/65536.0,1,-nbitq), 
to_sfixed(12157.0/65536.0,1,-nbitq), 
to_sfixed(3663.0/65536.0,1,-nbitq), 
to_sfixed(-1378.0/65536.0,1,-nbitq), 
to_sfixed(2718.0/65536.0,1,-nbitq), 
to_sfixed(-3873.0/65536.0,1,-nbitq), 
to_sfixed(-5931.0/65536.0,1,-nbitq), 
to_sfixed(2069.0/65536.0,1,-nbitq), 
to_sfixed(9635.0/65536.0,1,-nbitq), 
to_sfixed(-1388.0/65536.0,1,-nbitq), 
to_sfixed(-3655.0/65536.0,1,-nbitq), 
to_sfixed(-6596.0/65536.0,1,-nbitq), 
to_sfixed(-2109.0/65536.0,1,-nbitq), 
to_sfixed(-227.0/65536.0,1,-nbitq), 
to_sfixed(-777.0/65536.0,1,-nbitq), 
to_sfixed(2091.0/65536.0,1,-nbitq), 
to_sfixed(-8677.0/65536.0,1,-nbitq), 
to_sfixed(-3672.0/65536.0,1,-nbitq), 
to_sfixed(-4867.0/65536.0,1,-nbitq), 
to_sfixed(1944.0/65536.0,1,-nbitq), 
to_sfixed(12124.0/65536.0,1,-nbitq), 
to_sfixed(2134.0/65536.0,1,-nbitq), 
to_sfixed(896.0/65536.0,1,-nbitq), 
to_sfixed(8760.0/65536.0,1,-nbitq), 
to_sfixed(771.0/65536.0,1,-nbitq), 
to_sfixed(-1998.0/65536.0,1,-nbitq), 
to_sfixed(-4464.0/65536.0,1,-nbitq), 
to_sfixed(8636.0/65536.0,1,-nbitq), 
to_sfixed(-1524.0/65536.0,1,-nbitq), 
to_sfixed(923.0/65536.0,1,-nbitq), 
to_sfixed(1890.0/65536.0,1,-nbitq), 
to_sfixed(-1422.0/65536.0,1,-nbitq), 
to_sfixed(11538.0/65536.0,1,-nbitq), 
to_sfixed(16553.0/65536.0,1,-nbitq), 
to_sfixed(6556.0/65536.0,1,-nbitq), 
to_sfixed(-11773.0/65536.0,1,-nbitq), 
to_sfixed(-2973.0/65536.0,1,-nbitq), 
to_sfixed(-1691.0/65536.0,1,-nbitq), 
to_sfixed(-2389.0/65536.0,1,-nbitq), 
to_sfixed(-2208.0/65536.0,1,-nbitq), 
to_sfixed(8019.0/65536.0,1,-nbitq), 
to_sfixed(1058.0/65536.0,1,-nbitq), 
to_sfixed(2430.0/65536.0,1,-nbitq), 
to_sfixed(-2341.0/65536.0,1,-nbitq), 
to_sfixed(6875.0/65536.0,1,-nbitq), 
to_sfixed(-2309.0/65536.0,1,-nbitq), 
to_sfixed(-906.0/65536.0,1,-nbitq), 
to_sfixed(-4852.0/65536.0,1,-nbitq), 
to_sfixed(701.0/65536.0,1,-nbitq), 
to_sfixed(1910.0/65536.0,1,-nbitq), 
to_sfixed(5233.0/65536.0,1,-nbitq), 
to_sfixed(3337.0/65536.0,1,-nbitq), 
to_sfixed(9632.0/65536.0,1,-nbitq), 
to_sfixed(2064.0/65536.0,1,-nbitq), 
to_sfixed(1361.0/65536.0,1,-nbitq), 
to_sfixed(-6797.0/65536.0,1,-nbitq), 
to_sfixed(-9825.0/65536.0,1,-nbitq), 
to_sfixed(-10173.0/65536.0,1,-nbitq), 
to_sfixed(-1878.0/65536.0,1,-nbitq), 
to_sfixed(-2334.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-624.0/65536.0,1,-nbitq), 
to_sfixed(-684.0/65536.0,1,-nbitq), 
to_sfixed(-2264.0/65536.0,1,-nbitq), 
to_sfixed(4053.0/65536.0,1,-nbitq), 
to_sfixed(7980.0/65536.0,1,-nbitq), 
to_sfixed(3309.0/65536.0,1,-nbitq), 
to_sfixed(1059.0/65536.0,1,-nbitq), 
to_sfixed(-2705.0/65536.0,1,-nbitq), 
to_sfixed(451.0/65536.0,1,-nbitq), 
to_sfixed(10.0/65536.0,1,-nbitq), 
to_sfixed(919.0/65536.0,1,-nbitq), 
to_sfixed(-4406.0/65536.0,1,-nbitq), 
to_sfixed(1976.0/65536.0,1,-nbitq), 
to_sfixed(883.0/65536.0,1,-nbitq), 
to_sfixed(-211.0/65536.0,1,-nbitq), 
to_sfixed(2719.0/65536.0,1,-nbitq), 
to_sfixed(1501.0/65536.0,1,-nbitq), 
to_sfixed(-2563.0/65536.0,1,-nbitq), 
to_sfixed(-1222.0/65536.0,1,-nbitq), 
to_sfixed(1360.0/65536.0,1,-nbitq), 
to_sfixed(-601.0/65536.0,1,-nbitq), 
to_sfixed(5361.0/65536.0,1,-nbitq), 
to_sfixed(-627.0/65536.0,1,-nbitq), 
to_sfixed(-7096.0/65536.0,1,-nbitq), 
to_sfixed(-1754.0/65536.0,1,-nbitq), 
to_sfixed(3706.0/65536.0,1,-nbitq), 
to_sfixed(-5658.0/65536.0,1,-nbitq), 
to_sfixed(955.0/65536.0,1,-nbitq), 
to_sfixed(14066.0/65536.0,1,-nbitq), 
to_sfixed(-2779.0/65536.0,1,-nbitq), 
to_sfixed(-25.0/65536.0,1,-nbitq), 
to_sfixed(-5748.0/65536.0,1,-nbitq), 
to_sfixed(5581.0/65536.0,1,-nbitq), 
to_sfixed(5064.0/65536.0,1,-nbitq), 
to_sfixed(-2104.0/65536.0,1,-nbitq), 
to_sfixed(207.0/65536.0,1,-nbitq), 
to_sfixed(-6301.0/65536.0,1,-nbitq), 
to_sfixed(-5869.0/65536.0,1,-nbitq), 
to_sfixed(-4681.0/65536.0,1,-nbitq), 
to_sfixed(-1005.0/65536.0,1,-nbitq), 
to_sfixed(9422.0/65536.0,1,-nbitq), 
to_sfixed(-1240.0/65536.0,1,-nbitq), 
to_sfixed(3138.0/65536.0,1,-nbitq), 
to_sfixed(3800.0/65536.0,1,-nbitq), 
to_sfixed(-2057.0/65536.0,1,-nbitq), 
to_sfixed(176.0/65536.0,1,-nbitq), 
to_sfixed(-1429.0/65536.0,1,-nbitq), 
to_sfixed(13975.0/65536.0,1,-nbitq), 
to_sfixed(-464.0/65536.0,1,-nbitq), 
to_sfixed(2202.0/65536.0,1,-nbitq), 
to_sfixed(-942.0/65536.0,1,-nbitq), 
to_sfixed(-2824.0/65536.0,1,-nbitq), 
to_sfixed(5084.0/65536.0,1,-nbitq), 
to_sfixed(18872.0/65536.0,1,-nbitq), 
to_sfixed(4188.0/65536.0,1,-nbitq), 
to_sfixed(-4901.0/65536.0,1,-nbitq), 
to_sfixed(1693.0/65536.0,1,-nbitq), 
to_sfixed(-5271.0/65536.0,1,-nbitq), 
to_sfixed(2849.0/65536.0,1,-nbitq), 
to_sfixed(-788.0/65536.0,1,-nbitq), 
to_sfixed(8055.0/65536.0,1,-nbitq), 
to_sfixed(-1538.0/65536.0,1,-nbitq), 
to_sfixed(1982.0/65536.0,1,-nbitq), 
to_sfixed(585.0/65536.0,1,-nbitq), 
to_sfixed(4801.0/65536.0,1,-nbitq), 
to_sfixed(-4539.0/65536.0,1,-nbitq), 
to_sfixed(2075.0/65536.0,1,-nbitq), 
to_sfixed(-5151.0/65536.0,1,-nbitq), 
to_sfixed(1136.0/65536.0,1,-nbitq), 
to_sfixed(9410.0/65536.0,1,-nbitq), 
to_sfixed(4124.0/65536.0,1,-nbitq), 
to_sfixed(5979.0/65536.0,1,-nbitq), 
to_sfixed(9810.0/65536.0,1,-nbitq), 
to_sfixed(-3146.0/65536.0,1,-nbitq), 
to_sfixed(-2441.0/65536.0,1,-nbitq), 
to_sfixed(-404.0/65536.0,1,-nbitq), 
to_sfixed(-10585.0/65536.0,1,-nbitq), 
to_sfixed(-6444.0/65536.0,1,-nbitq), 
to_sfixed(-2484.0/65536.0,1,-nbitq), 
to_sfixed(-5074.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2611.0/65536.0,1,-nbitq), 
to_sfixed(2576.0/65536.0,1,-nbitq), 
to_sfixed(-3317.0/65536.0,1,-nbitq), 
to_sfixed(4597.0/65536.0,1,-nbitq), 
to_sfixed(8850.0/65536.0,1,-nbitq), 
to_sfixed(7566.0/65536.0,1,-nbitq), 
to_sfixed(563.0/65536.0,1,-nbitq), 
to_sfixed(-1842.0/65536.0,1,-nbitq), 
to_sfixed(368.0/65536.0,1,-nbitq), 
to_sfixed(2756.0/65536.0,1,-nbitq), 
to_sfixed(-1039.0/65536.0,1,-nbitq), 
to_sfixed(-13843.0/65536.0,1,-nbitq), 
to_sfixed(-1.0/65536.0,1,-nbitq), 
to_sfixed(1918.0/65536.0,1,-nbitq), 
to_sfixed(-4021.0/65536.0,1,-nbitq), 
to_sfixed(2070.0/65536.0,1,-nbitq), 
to_sfixed(-1649.0/65536.0,1,-nbitq), 
to_sfixed(-4098.0/65536.0,1,-nbitq), 
to_sfixed(-214.0/65536.0,1,-nbitq), 
to_sfixed(2142.0/65536.0,1,-nbitq), 
to_sfixed(-467.0/65536.0,1,-nbitq), 
to_sfixed(2061.0/65536.0,1,-nbitq), 
to_sfixed(-3691.0/65536.0,1,-nbitq), 
to_sfixed(-9082.0/65536.0,1,-nbitq), 
to_sfixed(-1072.0/65536.0,1,-nbitq), 
to_sfixed(6629.0/65536.0,1,-nbitq), 
to_sfixed(-6211.0/65536.0,1,-nbitq), 
to_sfixed(3989.0/65536.0,1,-nbitq), 
to_sfixed(14573.0/65536.0,1,-nbitq), 
to_sfixed(794.0/65536.0,1,-nbitq), 
to_sfixed(-1205.0/65536.0,1,-nbitq), 
to_sfixed(-10141.0/65536.0,1,-nbitq), 
to_sfixed(7188.0/65536.0,1,-nbitq), 
to_sfixed(6621.0/65536.0,1,-nbitq), 
to_sfixed(-1194.0/65536.0,1,-nbitq), 
to_sfixed(-209.0/65536.0,1,-nbitq), 
to_sfixed(-8985.0/65536.0,1,-nbitq), 
to_sfixed(-432.0/65536.0,1,-nbitq), 
to_sfixed(-6983.0/65536.0,1,-nbitq), 
to_sfixed(-2551.0/65536.0,1,-nbitq), 
to_sfixed(6168.0/65536.0,1,-nbitq), 
to_sfixed(2829.0/65536.0,1,-nbitq), 
to_sfixed(7872.0/65536.0,1,-nbitq), 
to_sfixed(5596.0/65536.0,1,-nbitq), 
to_sfixed(-1896.0/65536.0,1,-nbitq), 
to_sfixed(2940.0/65536.0,1,-nbitq), 
to_sfixed(-3252.0/65536.0,1,-nbitq), 
to_sfixed(7573.0/65536.0,1,-nbitq), 
to_sfixed(441.0/65536.0,1,-nbitq), 
to_sfixed(-2147.0/65536.0,1,-nbitq), 
to_sfixed(554.0/65536.0,1,-nbitq), 
to_sfixed(-1883.0/65536.0,1,-nbitq), 
to_sfixed(5.0/65536.0,1,-nbitq), 
to_sfixed(15710.0/65536.0,1,-nbitq), 
to_sfixed(-1572.0/65536.0,1,-nbitq), 
to_sfixed(698.0/65536.0,1,-nbitq), 
to_sfixed(-1921.0/65536.0,1,-nbitq), 
to_sfixed(-1260.0/65536.0,1,-nbitq), 
to_sfixed(-1336.0/65536.0,1,-nbitq), 
to_sfixed(-7428.0/65536.0,1,-nbitq), 
to_sfixed(8259.0/65536.0,1,-nbitq), 
to_sfixed(938.0/65536.0,1,-nbitq), 
to_sfixed(-819.0/65536.0,1,-nbitq), 
to_sfixed(886.0/65536.0,1,-nbitq), 
to_sfixed(4231.0/65536.0,1,-nbitq), 
to_sfixed(888.0/65536.0,1,-nbitq), 
to_sfixed(-727.0/65536.0,1,-nbitq), 
to_sfixed(5396.0/65536.0,1,-nbitq), 
to_sfixed(5863.0/65536.0,1,-nbitq), 
to_sfixed(12291.0/65536.0,1,-nbitq), 
to_sfixed(-1119.0/65536.0,1,-nbitq), 
to_sfixed(-1430.0/65536.0,1,-nbitq), 
to_sfixed(10556.0/65536.0,1,-nbitq), 
to_sfixed(-2997.0/65536.0,1,-nbitq), 
to_sfixed(447.0/65536.0,1,-nbitq), 
to_sfixed(1593.0/65536.0,1,-nbitq), 
to_sfixed(-8484.0/65536.0,1,-nbitq), 
to_sfixed(1145.0/65536.0,1,-nbitq), 
to_sfixed(808.0/65536.0,1,-nbitq), 
to_sfixed(-6103.0/65536.0,1,-nbitq)  ), 
( to_sfixed(660.0/65536.0,1,-nbitq), 
to_sfixed(1867.0/65536.0,1,-nbitq), 
to_sfixed(1648.0/65536.0,1,-nbitq), 
to_sfixed(4112.0/65536.0,1,-nbitq), 
to_sfixed(1540.0/65536.0,1,-nbitq), 
to_sfixed(4469.0/65536.0,1,-nbitq), 
to_sfixed(-1477.0/65536.0,1,-nbitq), 
to_sfixed(1339.0/65536.0,1,-nbitq), 
to_sfixed(-2825.0/65536.0,1,-nbitq), 
to_sfixed(-241.0/65536.0,1,-nbitq), 
to_sfixed(2205.0/65536.0,1,-nbitq), 
to_sfixed(-6532.0/65536.0,1,-nbitq), 
to_sfixed(-864.0/65536.0,1,-nbitq), 
to_sfixed(291.0/65536.0,1,-nbitq), 
to_sfixed(4939.0/65536.0,1,-nbitq), 
to_sfixed(-1700.0/65536.0,1,-nbitq), 
to_sfixed(1524.0/65536.0,1,-nbitq), 
to_sfixed(906.0/65536.0,1,-nbitq), 
to_sfixed(-1376.0/65536.0,1,-nbitq), 
to_sfixed(2905.0/65536.0,1,-nbitq), 
to_sfixed(2003.0/65536.0,1,-nbitq), 
to_sfixed(5098.0/65536.0,1,-nbitq), 
to_sfixed(-2299.0/65536.0,1,-nbitq), 
to_sfixed(-6304.0/65536.0,1,-nbitq), 
to_sfixed(567.0/65536.0,1,-nbitq), 
to_sfixed(9016.0/65536.0,1,-nbitq), 
to_sfixed(372.0/65536.0,1,-nbitq), 
to_sfixed(-354.0/65536.0,1,-nbitq), 
to_sfixed(12059.0/65536.0,1,-nbitq), 
to_sfixed(-2751.0/65536.0,1,-nbitq), 
to_sfixed(890.0/65536.0,1,-nbitq), 
to_sfixed(-7023.0/65536.0,1,-nbitq), 
to_sfixed(8667.0/65536.0,1,-nbitq), 
to_sfixed(2275.0/65536.0,1,-nbitq), 
to_sfixed(-568.0/65536.0,1,-nbitq), 
to_sfixed(-1228.0/65536.0,1,-nbitq), 
to_sfixed(-5314.0/65536.0,1,-nbitq), 
to_sfixed(1636.0/65536.0,1,-nbitq), 
to_sfixed(-1181.0/65536.0,1,-nbitq), 
to_sfixed(-1459.0/65536.0,1,-nbitq), 
to_sfixed(165.0/65536.0,1,-nbitq), 
to_sfixed(777.0/65536.0,1,-nbitq), 
to_sfixed(3623.0/65536.0,1,-nbitq), 
to_sfixed(8062.0/65536.0,1,-nbitq), 
to_sfixed(-1806.0/65536.0,1,-nbitq), 
to_sfixed(3399.0/65536.0,1,-nbitq), 
to_sfixed(-3130.0/65536.0,1,-nbitq), 
to_sfixed(3375.0/65536.0,1,-nbitq), 
to_sfixed(2154.0/65536.0,1,-nbitq), 
to_sfixed(-1156.0/65536.0,1,-nbitq), 
to_sfixed(-1026.0/65536.0,1,-nbitq), 
to_sfixed(777.0/65536.0,1,-nbitq), 
to_sfixed(2299.0/65536.0,1,-nbitq), 
to_sfixed(14840.0/65536.0,1,-nbitq), 
to_sfixed(-295.0/65536.0,1,-nbitq), 
to_sfixed(2526.0/65536.0,1,-nbitq), 
to_sfixed(686.0/65536.0,1,-nbitq), 
to_sfixed(934.0/65536.0,1,-nbitq), 
to_sfixed(1470.0/65536.0,1,-nbitq), 
to_sfixed(-2662.0/65536.0,1,-nbitq), 
to_sfixed(8941.0/65536.0,1,-nbitq), 
to_sfixed(-2053.0/65536.0,1,-nbitq), 
to_sfixed(-1034.0/65536.0,1,-nbitq), 
to_sfixed(-1272.0/65536.0,1,-nbitq), 
to_sfixed(8912.0/65536.0,1,-nbitq), 
to_sfixed(8380.0/65536.0,1,-nbitq), 
to_sfixed(2760.0/65536.0,1,-nbitq), 
to_sfixed(7911.0/65536.0,1,-nbitq), 
to_sfixed(2080.0/65536.0,1,-nbitq), 
to_sfixed(2461.0/65536.0,1,-nbitq), 
to_sfixed(-1070.0/65536.0,1,-nbitq), 
to_sfixed(-3747.0/65536.0,1,-nbitq), 
to_sfixed(3285.0/65536.0,1,-nbitq), 
to_sfixed(2618.0/65536.0,1,-nbitq), 
to_sfixed(1569.0/65536.0,1,-nbitq), 
to_sfixed(1789.0/65536.0,1,-nbitq), 
to_sfixed(-10170.0/65536.0,1,-nbitq), 
to_sfixed(2433.0/65536.0,1,-nbitq), 
to_sfixed(138.0/65536.0,1,-nbitq), 
to_sfixed(-5280.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1570.0/65536.0,1,-nbitq), 
to_sfixed(1169.0/65536.0,1,-nbitq), 
to_sfixed(-598.0/65536.0,1,-nbitq), 
to_sfixed(7802.0/65536.0,1,-nbitq), 
to_sfixed(3527.0/65536.0,1,-nbitq), 
to_sfixed(2918.0/65536.0,1,-nbitq), 
to_sfixed(-433.0/65536.0,1,-nbitq), 
to_sfixed(9307.0/65536.0,1,-nbitq), 
to_sfixed(-232.0/65536.0,1,-nbitq), 
to_sfixed(-1786.0/65536.0,1,-nbitq), 
to_sfixed(6171.0/65536.0,1,-nbitq), 
to_sfixed(-6981.0/65536.0,1,-nbitq), 
to_sfixed(-2373.0/65536.0,1,-nbitq), 
to_sfixed(2569.0/65536.0,1,-nbitq), 
to_sfixed(609.0/65536.0,1,-nbitq), 
to_sfixed(-216.0/65536.0,1,-nbitq), 
to_sfixed(-1778.0/65536.0,1,-nbitq), 
to_sfixed(2848.0/65536.0,1,-nbitq), 
to_sfixed(4219.0/65536.0,1,-nbitq), 
to_sfixed(2470.0/65536.0,1,-nbitq), 
to_sfixed(6511.0/65536.0,1,-nbitq), 
to_sfixed(81.0/65536.0,1,-nbitq), 
to_sfixed(-2734.0/65536.0,1,-nbitq), 
to_sfixed(-1630.0/65536.0,1,-nbitq), 
to_sfixed(-463.0/65536.0,1,-nbitq), 
to_sfixed(10340.0/65536.0,1,-nbitq), 
to_sfixed(-2046.0/65536.0,1,-nbitq), 
to_sfixed(-2695.0/65536.0,1,-nbitq), 
to_sfixed(10555.0/65536.0,1,-nbitq), 
to_sfixed(-384.0/65536.0,1,-nbitq), 
to_sfixed(303.0/65536.0,1,-nbitq), 
to_sfixed(-9292.0/65536.0,1,-nbitq), 
to_sfixed(2801.0/65536.0,1,-nbitq), 
to_sfixed(-1240.0/65536.0,1,-nbitq), 
to_sfixed(-1335.0/65536.0,1,-nbitq), 
to_sfixed(-2567.0/65536.0,1,-nbitq), 
to_sfixed(-3102.0/65536.0,1,-nbitq), 
to_sfixed(2475.0/65536.0,1,-nbitq), 
to_sfixed(-4662.0/65536.0,1,-nbitq), 
to_sfixed(7.0/65536.0,1,-nbitq), 
to_sfixed(1720.0/65536.0,1,-nbitq), 
to_sfixed(-2745.0/65536.0,1,-nbitq), 
to_sfixed(5210.0/65536.0,1,-nbitq), 
to_sfixed(3033.0/65536.0,1,-nbitq), 
to_sfixed(-854.0/65536.0,1,-nbitq), 
to_sfixed(-2529.0/65536.0,1,-nbitq), 
to_sfixed(261.0/65536.0,1,-nbitq), 
to_sfixed(823.0/65536.0,1,-nbitq), 
to_sfixed(534.0/65536.0,1,-nbitq), 
to_sfixed(2195.0/65536.0,1,-nbitq), 
to_sfixed(-1895.0/65536.0,1,-nbitq), 
to_sfixed(5007.0/65536.0,1,-nbitq), 
to_sfixed(-1319.0/65536.0,1,-nbitq), 
to_sfixed(16283.0/65536.0,1,-nbitq), 
to_sfixed(-5819.0/65536.0,1,-nbitq), 
to_sfixed(-3182.0/65536.0,1,-nbitq), 
to_sfixed(2086.0/65536.0,1,-nbitq), 
to_sfixed(3479.0/65536.0,1,-nbitq), 
to_sfixed(-2912.0/65536.0,1,-nbitq), 
to_sfixed(-5982.0/65536.0,1,-nbitq), 
to_sfixed(466.0/65536.0,1,-nbitq), 
to_sfixed(-1853.0/65536.0,1,-nbitq), 
to_sfixed(1255.0/65536.0,1,-nbitq), 
to_sfixed(195.0/65536.0,1,-nbitq), 
to_sfixed(-2718.0/65536.0,1,-nbitq), 
to_sfixed(6638.0/65536.0,1,-nbitq), 
to_sfixed(423.0/65536.0,1,-nbitq), 
to_sfixed(5550.0/65536.0,1,-nbitq), 
to_sfixed(-3086.0/65536.0,1,-nbitq), 
to_sfixed(885.0/65536.0,1,-nbitq), 
to_sfixed(-1579.0/65536.0,1,-nbitq), 
to_sfixed(-6080.0/65536.0,1,-nbitq), 
to_sfixed(4826.0/65536.0,1,-nbitq), 
to_sfixed(2026.0/65536.0,1,-nbitq), 
to_sfixed(931.0/65536.0,1,-nbitq), 
to_sfixed(-245.0/65536.0,1,-nbitq), 
to_sfixed(-4802.0/65536.0,1,-nbitq), 
to_sfixed(1403.0/65536.0,1,-nbitq), 
to_sfixed(-1240.0/65536.0,1,-nbitq), 
to_sfixed(-5052.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2456.0/65536.0,1,-nbitq), 
to_sfixed(-532.0/65536.0,1,-nbitq), 
to_sfixed(-1700.0/65536.0,1,-nbitq), 
to_sfixed(1320.0/65536.0,1,-nbitq), 
to_sfixed(2593.0/65536.0,1,-nbitq), 
to_sfixed(1610.0/65536.0,1,-nbitq), 
to_sfixed(52.0/65536.0,1,-nbitq), 
to_sfixed(6531.0/65536.0,1,-nbitq), 
to_sfixed(-1415.0/65536.0,1,-nbitq), 
to_sfixed(2580.0/65536.0,1,-nbitq), 
to_sfixed(2223.0/65536.0,1,-nbitq), 
to_sfixed(-11839.0/65536.0,1,-nbitq), 
to_sfixed(1431.0/65536.0,1,-nbitq), 
to_sfixed(3671.0/65536.0,1,-nbitq), 
to_sfixed(-1964.0/65536.0,1,-nbitq), 
to_sfixed(1167.0/65536.0,1,-nbitq), 
to_sfixed(-3016.0/65536.0,1,-nbitq), 
to_sfixed(6603.0/65536.0,1,-nbitq), 
to_sfixed(2306.0/65536.0,1,-nbitq), 
to_sfixed(-728.0/65536.0,1,-nbitq), 
to_sfixed(1284.0/65536.0,1,-nbitq), 
to_sfixed(-6566.0/65536.0,1,-nbitq), 
to_sfixed(504.0/65536.0,1,-nbitq), 
to_sfixed(-2207.0/65536.0,1,-nbitq), 
to_sfixed(-1601.0/65536.0,1,-nbitq), 
to_sfixed(4301.0/65536.0,1,-nbitq), 
to_sfixed(-3945.0/65536.0,1,-nbitq), 
to_sfixed(-413.0/65536.0,1,-nbitq), 
to_sfixed(7148.0/65536.0,1,-nbitq), 
to_sfixed(1865.0/65536.0,1,-nbitq), 
to_sfixed(2359.0/65536.0,1,-nbitq), 
to_sfixed(-6516.0/65536.0,1,-nbitq), 
to_sfixed(1623.0/65536.0,1,-nbitq), 
to_sfixed(-5328.0/65536.0,1,-nbitq), 
to_sfixed(-2976.0/65536.0,1,-nbitq), 
to_sfixed(-1965.0/65536.0,1,-nbitq), 
to_sfixed(-933.0/65536.0,1,-nbitq), 
to_sfixed(-1752.0/65536.0,1,-nbitq), 
to_sfixed(-1289.0/65536.0,1,-nbitq), 
to_sfixed(1220.0/65536.0,1,-nbitq), 
to_sfixed(-1631.0/65536.0,1,-nbitq), 
to_sfixed(843.0/65536.0,1,-nbitq), 
to_sfixed(2605.0/65536.0,1,-nbitq), 
to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(-821.0/65536.0,1,-nbitq), 
to_sfixed(-1661.0/65536.0,1,-nbitq), 
to_sfixed(611.0/65536.0,1,-nbitq), 
to_sfixed(-484.0/65536.0,1,-nbitq), 
to_sfixed(1745.0/65536.0,1,-nbitq), 
to_sfixed(1847.0/65536.0,1,-nbitq), 
to_sfixed(-1535.0/65536.0,1,-nbitq), 
to_sfixed(4386.0/65536.0,1,-nbitq), 
to_sfixed(-138.0/65536.0,1,-nbitq), 
to_sfixed(11150.0/65536.0,1,-nbitq), 
to_sfixed(-4490.0/65536.0,1,-nbitq), 
to_sfixed(-1683.0/65536.0,1,-nbitq), 
to_sfixed(667.0/65536.0,1,-nbitq), 
to_sfixed(949.0/65536.0,1,-nbitq), 
to_sfixed(-1675.0/65536.0,1,-nbitq), 
to_sfixed(-4225.0/65536.0,1,-nbitq), 
to_sfixed(-3324.0/65536.0,1,-nbitq), 
to_sfixed(170.0/65536.0,1,-nbitq), 
to_sfixed(-1639.0/65536.0,1,-nbitq), 
to_sfixed(1500.0/65536.0,1,-nbitq), 
to_sfixed(897.0/65536.0,1,-nbitq), 
to_sfixed(-1725.0/65536.0,1,-nbitq), 
to_sfixed(3960.0/65536.0,1,-nbitq), 
to_sfixed(3384.0/65536.0,1,-nbitq), 
to_sfixed(3069.0/65536.0,1,-nbitq), 
to_sfixed(3465.0/65536.0,1,-nbitq), 
to_sfixed(1432.0/65536.0,1,-nbitq), 
to_sfixed(1116.0/65536.0,1,-nbitq), 
to_sfixed(5076.0/65536.0,1,-nbitq), 
to_sfixed(-1633.0/65536.0,1,-nbitq), 
to_sfixed(133.0/65536.0,1,-nbitq), 
to_sfixed(-386.0/65536.0,1,-nbitq), 
to_sfixed(-6138.0/65536.0,1,-nbitq), 
to_sfixed(1336.0/65536.0,1,-nbitq), 
to_sfixed(297.0/65536.0,1,-nbitq), 
to_sfixed(-305.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3670.0/65536.0,1,-nbitq), 
to_sfixed(-838.0/65536.0,1,-nbitq), 
to_sfixed(-5315.0/65536.0,1,-nbitq), 
to_sfixed(531.0/65536.0,1,-nbitq), 
to_sfixed(1335.0/65536.0,1,-nbitq), 
to_sfixed(610.0/65536.0,1,-nbitq), 
to_sfixed(-2818.0/65536.0,1,-nbitq), 
to_sfixed(6393.0/65536.0,1,-nbitq), 
to_sfixed(-3048.0/65536.0,1,-nbitq), 
to_sfixed(-191.0/65536.0,1,-nbitq), 
to_sfixed(1457.0/65536.0,1,-nbitq), 
to_sfixed(-7371.0/65536.0,1,-nbitq), 
to_sfixed(-150.0/65536.0,1,-nbitq), 
to_sfixed(-1411.0/65536.0,1,-nbitq), 
to_sfixed(-2510.0/65536.0,1,-nbitq), 
to_sfixed(883.0/65536.0,1,-nbitq), 
to_sfixed(-937.0/65536.0,1,-nbitq), 
to_sfixed(7118.0/65536.0,1,-nbitq), 
to_sfixed(-1470.0/65536.0,1,-nbitq), 
to_sfixed(2758.0/65536.0,1,-nbitq), 
to_sfixed(-534.0/65536.0,1,-nbitq), 
to_sfixed(2828.0/65536.0,1,-nbitq), 
to_sfixed(-1619.0/65536.0,1,-nbitq), 
to_sfixed(-2625.0/65536.0,1,-nbitq), 
to_sfixed(-873.0/65536.0,1,-nbitq), 
to_sfixed(148.0/65536.0,1,-nbitq), 
to_sfixed(-3356.0/65536.0,1,-nbitq), 
to_sfixed(-1940.0/65536.0,1,-nbitq), 
to_sfixed(5797.0/65536.0,1,-nbitq), 
to_sfixed(-2880.0/65536.0,1,-nbitq), 
to_sfixed(3330.0/65536.0,1,-nbitq), 
to_sfixed(-867.0/65536.0,1,-nbitq), 
to_sfixed(-2119.0/65536.0,1,-nbitq), 
to_sfixed(-8200.0/65536.0,1,-nbitq), 
to_sfixed(-567.0/65536.0,1,-nbitq), 
to_sfixed(-301.0/65536.0,1,-nbitq), 
to_sfixed(-5654.0/65536.0,1,-nbitq), 
to_sfixed(1792.0/65536.0,1,-nbitq), 
to_sfixed(-3332.0/65536.0,1,-nbitq), 
to_sfixed(1508.0/65536.0,1,-nbitq), 
to_sfixed(-381.0/65536.0,1,-nbitq), 
to_sfixed(2384.0/65536.0,1,-nbitq), 
to_sfixed(936.0/65536.0,1,-nbitq), 
to_sfixed(3321.0/65536.0,1,-nbitq), 
to_sfixed(2819.0/65536.0,1,-nbitq), 
to_sfixed(324.0/65536.0,1,-nbitq), 
to_sfixed(794.0/65536.0,1,-nbitq), 
to_sfixed(-2899.0/65536.0,1,-nbitq), 
to_sfixed(2678.0/65536.0,1,-nbitq), 
to_sfixed(3029.0/65536.0,1,-nbitq), 
to_sfixed(-1315.0/65536.0,1,-nbitq), 
to_sfixed(2267.0/65536.0,1,-nbitq), 
to_sfixed(-5178.0/65536.0,1,-nbitq), 
to_sfixed(7291.0/65536.0,1,-nbitq), 
to_sfixed(-3365.0/65536.0,1,-nbitq), 
to_sfixed(-942.0/65536.0,1,-nbitq), 
to_sfixed(-133.0/65536.0,1,-nbitq), 
to_sfixed(860.0/65536.0,1,-nbitq), 
to_sfixed(-121.0/65536.0,1,-nbitq), 
to_sfixed(-1161.0/65536.0,1,-nbitq), 
to_sfixed(-3274.0/65536.0,1,-nbitq), 
to_sfixed(-2154.0/65536.0,1,-nbitq), 
to_sfixed(1241.0/65536.0,1,-nbitq), 
to_sfixed(-1661.0/65536.0,1,-nbitq), 
to_sfixed(-1084.0/65536.0,1,-nbitq), 
to_sfixed(-1708.0/65536.0,1,-nbitq), 
to_sfixed(2773.0/65536.0,1,-nbitq), 
to_sfixed(1738.0/65536.0,1,-nbitq), 
to_sfixed(6040.0/65536.0,1,-nbitq), 
to_sfixed(336.0/65536.0,1,-nbitq), 
to_sfixed(-332.0/65536.0,1,-nbitq), 
to_sfixed(-2532.0/65536.0,1,-nbitq), 
to_sfixed(6374.0/65536.0,1,-nbitq), 
to_sfixed(1780.0/65536.0,1,-nbitq), 
to_sfixed(267.0/65536.0,1,-nbitq), 
to_sfixed(-2764.0/65536.0,1,-nbitq), 
to_sfixed(-5220.0/65536.0,1,-nbitq), 
to_sfixed(4237.0/65536.0,1,-nbitq), 
to_sfixed(942.0/65536.0,1,-nbitq), 
to_sfixed(-1550.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1636.0/65536.0,1,-nbitq), 
to_sfixed(1137.0/65536.0,1,-nbitq), 
to_sfixed(991.0/65536.0,1,-nbitq), 
to_sfixed(-847.0/65536.0,1,-nbitq), 
to_sfixed(-2921.0/65536.0,1,-nbitq), 
to_sfixed(-4020.0/65536.0,1,-nbitq), 
to_sfixed(113.0/65536.0,1,-nbitq), 
to_sfixed(3602.0/65536.0,1,-nbitq), 
to_sfixed(1144.0/65536.0,1,-nbitq), 
to_sfixed(-2357.0/65536.0,1,-nbitq), 
to_sfixed(-1301.0/65536.0,1,-nbitq), 
to_sfixed(-482.0/65536.0,1,-nbitq), 
to_sfixed(-496.0/65536.0,1,-nbitq), 
to_sfixed(-1380.0/65536.0,1,-nbitq), 
to_sfixed(201.0/65536.0,1,-nbitq), 
to_sfixed(-603.0/65536.0,1,-nbitq), 
to_sfixed(233.0/65536.0,1,-nbitq), 
to_sfixed(3675.0/65536.0,1,-nbitq), 
to_sfixed(-612.0/65536.0,1,-nbitq), 
to_sfixed(1523.0/65536.0,1,-nbitq), 
to_sfixed(184.0/65536.0,1,-nbitq), 
to_sfixed(2305.0/65536.0,1,-nbitq), 
to_sfixed(-2400.0/65536.0,1,-nbitq), 
to_sfixed(1232.0/65536.0,1,-nbitq), 
to_sfixed(-1117.0/65536.0,1,-nbitq), 
to_sfixed(2341.0/65536.0,1,-nbitq), 
to_sfixed(177.0/65536.0,1,-nbitq), 
to_sfixed(817.0/65536.0,1,-nbitq), 
to_sfixed(-2044.0/65536.0,1,-nbitq), 
to_sfixed(-1063.0/65536.0,1,-nbitq), 
to_sfixed(1574.0/65536.0,1,-nbitq), 
to_sfixed(-1285.0/65536.0,1,-nbitq), 
to_sfixed(-4183.0/65536.0,1,-nbitq), 
to_sfixed(-3556.0/65536.0,1,-nbitq), 
to_sfixed(-808.0/65536.0,1,-nbitq), 
to_sfixed(-3199.0/65536.0,1,-nbitq), 
to_sfixed(-1416.0/65536.0,1,-nbitq), 
to_sfixed(-765.0/65536.0,1,-nbitq), 
to_sfixed(580.0/65536.0,1,-nbitq), 
to_sfixed(-602.0/65536.0,1,-nbitq), 
to_sfixed(-1732.0/65536.0,1,-nbitq), 
to_sfixed(-2062.0/65536.0,1,-nbitq), 
to_sfixed(-824.0/65536.0,1,-nbitq), 
to_sfixed(136.0/65536.0,1,-nbitq), 
to_sfixed(-1832.0/65536.0,1,-nbitq), 
to_sfixed(1283.0/65536.0,1,-nbitq), 
to_sfixed(668.0/65536.0,1,-nbitq), 
to_sfixed(-453.0/65536.0,1,-nbitq), 
to_sfixed(129.0/65536.0,1,-nbitq), 
to_sfixed(3931.0/65536.0,1,-nbitq), 
to_sfixed(-2488.0/65536.0,1,-nbitq), 
to_sfixed(2320.0/65536.0,1,-nbitq), 
to_sfixed(-3613.0/65536.0,1,-nbitq), 
to_sfixed(344.0/65536.0,1,-nbitq), 
to_sfixed(-100.0/65536.0,1,-nbitq), 
to_sfixed(-2714.0/65536.0,1,-nbitq), 
to_sfixed(-27.0/65536.0,1,-nbitq), 
to_sfixed(1601.0/65536.0,1,-nbitq), 
to_sfixed(1236.0/65536.0,1,-nbitq), 
to_sfixed(3540.0/65536.0,1,-nbitq), 
to_sfixed(-2630.0/65536.0,1,-nbitq), 
to_sfixed(2072.0/65536.0,1,-nbitq), 
to_sfixed(-1704.0/65536.0,1,-nbitq), 
to_sfixed(634.0/65536.0,1,-nbitq), 
to_sfixed(-26.0/65536.0,1,-nbitq), 
to_sfixed(552.0/65536.0,1,-nbitq), 
to_sfixed(1390.0/65536.0,1,-nbitq), 
to_sfixed(-3296.0/65536.0,1,-nbitq), 
to_sfixed(4365.0/65536.0,1,-nbitq), 
to_sfixed(-871.0/65536.0,1,-nbitq), 
to_sfixed(1696.0/65536.0,1,-nbitq), 
to_sfixed(1974.0/65536.0,1,-nbitq), 
to_sfixed(558.0/65536.0,1,-nbitq), 
to_sfixed(-2709.0/65536.0,1,-nbitq), 
to_sfixed(162.0/65536.0,1,-nbitq), 
to_sfixed(2405.0/65536.0,1,-nbitq), 
to_sfixed(-1319.0/65536.0,1,-nbitq), 
to_sfixed(969.0/65536.0,1,-nbitq), 
to_sfixed(-1536.0/65536.0,1,-nbitq), 
to_sfixed(338.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1000.0/65536.0,1,-nbitq), 
to_sfixed(1322.0/65536.0,1,-nbitq), 
to_sfixed(564.0/65536.0,1,-nbitq), 
to_sfixed(2407.0/65536.0,1,-nbitq), 
to_sfixed(1410.0/65536.0,1,-nbitq), 
to_sfixed(-931.0/65536.0,1,-nbitq), 
to_sfixed(812.0/65536.0,1,-nbitq), 
to_sfixed(2757.0/65536.0,1,-nbitq), 
to_sfixed(-2875.0/65536.0,1,-nbitq), 
to_sfixed(-277.0/65536.0,1,-nbitq), 
to_sfixed(1035.0/65536.0,1,-nbitq), 
to_sfixed(-460.0/65536.0,1,-nbitq), 
to_sfixed(1694.0/65536.0,1,-nbitq), 
to_sfixed(-3464.0/65536.0,1,-nbitq), 
to_sfixed(3647.0/65536.0,1,-nbitq), 
to_sfixed(1535.0/65536.0,1,-nbitq), 
to_sfixed(2739.0/65536.0,1,-nbitq), 
to_sfixed(863.0/65536.0,1,-nbitq), 
to_sfixed(1940.0/65536.0,1,-nbitq), 
to_sfixed(376.0/65536.0,1,-nbitq), 
to_sfixed(741.0/65536.0,1,-nbitq), 
to_sfixed(-2298.0/65536.0,1,-nbitq), 
to_sfixed(-348.0/65536.0,1,-nbitq), 
to_sfixed(-149.0/65536.0,1,-nbitq), 
to_sfixed(1210.0/65536.0,1,-nbitq), 
to_sfixed(2697.0/65536.0,1,-nbitq), 
to_sfixed(-3163.0/65536.0,1,-nbitq), 
to_sfixed(-405.0/65536.0,1,-nbitq), 
to_sfixed(2162.0/65536.0,1,-nbitq), 
to_sfixed(-1170.0/65536.0,1,-nbitq), 
to_sfixed(-1747.0/65536.0,1,-nbitq), 
to_sfixed(-1827.0/65536.0,1,-nbitq), 
to_sfixed(-3804.0/65536.0,1,-nbitq), 
to_sfixed(-1234.0/65536.0,1,-nbitq), 
to_sfixed(-438.0/65536.0,1,-nbitq), 
to_sfixed(2114.0/65536.0,1,-nbitq), 
to_sfixed(-1338.0/65536.0,1,-nbitq), 
to_sfixed(-1671.0/65536.0,1,-nbitq), 
to_sfixed(-1034.0/65536.0,1,-nbitq), 
to_sfixed(-237.0/65536.0,1,-nbitq), 
to_sfixed(-3499.0/65536.0,1,-nbitq), 
to_sfixed(-599.0/65536.0,1,-nbitq), 
to_sfixed(454.0/65536.0,1,-nbitq), 
to_sfixed(1185.0/65536.0,1,-nbitq), 
to_sfixed(-1646.0/65536.0,1,-nbitq), 
to_sfixed(1436.0/65536.0,1,-nbitq), 
to_sfixed(304.0/65536.0,1,-nbitq), 
to_sfixed(2929.0/65536.0,1,-nbitq), 
to_sfixed(-2240.0/65536.0,1,-nbitq), 
to_sfixed(-291.0/65536.0,1,-nbitq), 
to_sfixed(-1635.0/65536.0,1,-nbitq), 
to_sfixed(165.0/65536.0,1,-nbitq), 
to_sfixed(-672.0/65536.0,1,-nbitq), 
to_sfixed(1584.0/65536.0,1,-nbitq), 
to_sfixed(-1105.0/65536.0,1,-nbitq), 
to_sfixed(1314.0/65536.0,1,-nbitq), 
to_sfixed(517.0/65536.0,1,-nbitq), 
to_sfixed(2403.0/65536.0,1,-nbitq), 
to_sfixed(559.0/65536.0,1,-nbitq), 
to_sfixed(3583.0/65536.0,1,-nbitq), 
to_sfixed(-34.0/65536.0,1,-nbitq), 
to_sfixed(501.0/65536.0,1,-nbitq), 
to_sfixed(-1358.0/65536.0,1,-nbitq), 
to_sfixed(-2557.0/65536.0,1,-nbitq), 
to_sfixed(502.0/65536.0,1,-nbitq), 
to_sfixed(483.0/65536.0,1,-nbitq), 
to_sfixed(-1966.0/65536.0,1,-nbitq), 
to_sfixed(-3698.0/65536.0,1,-nbitq), 
to_sfixed(1247.0/65536.0,1,-nbitq), 
to_sfixed(-844.0/65536.0,1,-nbitq), 
to_sfixed(-1657.0/65536.0,1,-nbitq), 
to_sfixed(2077.0/65536.0,1,-nbitq), 
to_sfixed(1893.0/65536.0,1,-nbitq), 
to_sfixed(1004.0/65536.0,1,-nbitq), 
to_sfixed(384.0/65536.0,1,-nbitq), 
to_sfixed(2461.0/65536.0,1,-nbitq), 
to_sfixed(1708.0/65536.0,1,-nbitq), 
to_sfixed(193.0/65536.0,1,-nbitq), 
to_sfixed(1382.0/65536.0,1,-nbitq), 
to_sfixed(-466.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(704.0/65536.0,1,-nbitq), 
to_sfixed(2267.0/65536.0,1,-nbitq), 
to_sfixed(-338.0/65536.0,1,-nbitq), 
to_sfixed(2041.0/65536.0,1,-nbitq), 
to_sfixed(1961.0/65536.0,1,-nbitq), 
to_sfixed(-1817.0/65536.0,1,-nbitq), 
to_sfixed(-1589.0/65536.0,1,-nbitq), 
to_sfixed(-2364.0/65536.0,1,-nbitq), 
to_sfixed(963.0/65536.0,1,-nbitq), 
to_sfixed(653.0/65536.0,1,-nbitq), 
to_sfixed(-561.0/65536.0,1,-nbitq), 
to_sfixed(-2900.0/65536.0,1,-nbitq), 
to_sfixed(1925.0/65536.0,1,-nbitq), 
to_sfixed(-4849.0/65536.0,1,-nbitq), 
to_sfixed(48.0/65536.0,1,-nbitq), 
to_sfixed(2689.0/65536.0,1,-nbitq), 
to_sfixed(-2046.0/65536.0,1,-nbitq), 
to_sfixed(-556.0/65536.0,1,-nbitq), 
to_sfixed(3043.0/65536.0,1,-nbitq), 
to_sfixed(1767.0/65536.0,1,-nbitq), 
to_sfixed(-1034.0/65536.0,1,-nbitq), 
to_sfixed(-504.0/65536.0,1,-nbitq), 
to_sfixed(-2289.0/65536.0,1,-nbitq), 
to_sfixed(-427.0/65536.0,1,-nbitq), 
to_sfixed(655.0/65536.0,1,-nbitq), 
to_sfixed(4404.0/65536.0,1,-nbitq), 
to_sfixed(-2188.0/65536.0,1,-nbitq), 
to_sfixed(-2436.0/65536.0,1,-nbitq), 
to_sfixed(1306.0/65536.0,1,-nbitq), 
to_sfixed(-2691.0/65536.0,1,-nbitq), 
to_sfixed(1406.0/65536.0,1,-nbitq), 
to_sfixed(-3217.0/65536.0,1,-nbitq), 
to_sfixed(-4275.0/65536.0,1,-nbitq), 
to_sfixed(-1877.0/65536.0,1,-nbitq), 
to_sfixed(-1905.0/65536.0,1,-nbitq), 
to_sfixed(2590.0/65536.0,1,-nbitq), 
to_sfixed(1018.0/65536.0,1,-nbitq), 
to_sfixed(-2812.0/65536.0,1,-nbitq), 
to_sfixed(-1201.0/65536.0,1,-nbitq), 
to_sfixed(-30.0/65536.0,1,-nbitq), 
to_sfixed(-2572.0/65536.0,1,-nbitq), 
to_sfixed(1504.0/65536.0,1,-nbitq), 
to_sfixed(-1078.0/65536.0,1,-nbitq), 
to_sfixed(862.0/65536.0,1,-nbitq), 
to_sfixed(1790.0/65536.0,1,-nbitq), 
to_sfixed(2153.0/65536.0,1,-nbitq), 
to_sfixed(1227.0/65536.0,1,-nbitq), 
to_sfixed(1907.0/65536.0,1,-nbitq), 
to_sfixed(-284.0/65536.0,1,-nbitq), 
to_sfixed(-141.0/65536.0,1,-nbitq), 
to_sfixed(843.0/65536.0,1,-nbitq), 
to_sfixed(-1937.0/65536.0,1,-nbitq), 
to_sfixed(-309.0/65536.0,1,-nbitq), 
to_sfixed(-1523.0/65536.0,1,-nbitq), 
to_sfixed(-254.0/65536.0,1,-nbitq), 
to_sfixed(-2664.0/65536.0,1,-nbitq), 
to_sfixed(-963.0/65536.0,1,-nbitq), 
to_sfixed(1856.0/65536.0,1,-nbitq), 
to_sfixed(135.0/65536.0,1,-nbitq), 
to_sfixed(4009.0/65536.0,1,-nbitq), 
to_sfixed(-3653.0/65536.0,1,-nbitq), 
to_sfixed(2519.0/65536.0,1,-nbitq), 
to_sfixed(-2054.0/65536.0,1,-nbitq), 
to_sfixed(191.0/65536.0,1,-nbitq), 
to_sfixed(75.0/65536.0,1,-nbitq), 
to_sfixed(1427.0/65536.0,1,-nbitq), 
to_sfixed(2209.0/65536.0,1,-nbitq), 
to_sfixed(-1289.0/65536.0,1,-nbitq), 
to_sfixed(-56.0/65536.0,1,-nbitq), 
to_sfixed(-2892.0/65536.0,1,-nbitq), 
to_sfixed(-839.0/65536.0,1,-nbitq), 
to_sfixed(-860.0/65536.0,1,-nbitq), 
to_sfixed(731.0/65536.0,1,-nbitq), 
to_sfixed(-1910.0/65536.0,1,-nbitq), 
to_sfixed(921.0/65536.0,1,-nbitq), 
to_sfixed(291.0/65536.0,1,-nbitq), 
to_sfixed(-2377.0/65536.0,1,-nbitq), 
to_sfixed(161.0/65536.0,1,-nbitq), 
to_sfixed(732.0/65536.0,1,-nbitq), 
to_sfixed(1077.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3050.0/65536.0,1,-nbitq), 
to_sfixed(647.0/65536.0,1,-nbitq), 
to_sfixed(4597.0/65536.0,1,-nbitq), 
to_sfixed(-2798.0/65536.0,1,-nbitq), 
to_sfixed(-1654.0/65536.0,1,-nbitq), 
to_sfixed(-2955.0/65536.0,1,-nbitq), 
to_sfixed(-2868.0/65536.0,1,-nbitq), 
to_sfixed(-1407.0/65536.0,1,-nbitq), 
to_sfixed(-2513.0/65536.0,1,-nbitq), 
to_sfixed(678.0/65536.0,1,-nbitq), 
to_sfixed(1451.0/65536.0,1,-nbitq), 
to_sfixed(-529.0/65536.0,1,-nbitq), 
to_sfixed(2079.0/65536.0,1,-nbitq), 
to_sfixed(526.0/65536.0,1,-nbitq), 
to_sfixed(-444.0/65536.0,1,-nbitq), 
to_sfixed(-826.0/65536.0,1,-nbitq), 
to_sfixed(-2914.0/65536.0,1,-nbitq), 
to_sfixed(2672.0/65536.0,1,-nbitq), 
to_sfixed(150.0/65536.0,1,-nbitq), 
to_sfixed(258.0/65536.0,1,-nbitq), 
to_sfixed(-3058.0/65536.0,1,-nbitq), 
to_sfixed(2085.0/65536.0,1,-nbitq), 
to_sfixed(673.0/65536.0,1,-nbitq), 
to_sfixed(637.0/65536.0,1,-nbitq), 
to_sfixed(3599.0/65536.0,1,-nbitq), 
to_sfixed(1038.0/65536.0,1,-nbitq), 
to_sfixed(-2603.0/65536.0,1,-nbitq), 
to_sfixed(779.0/65536.0,1,-nbitq), 
to_sfixed(4300.0/65536.0,1,-nbitq), 
to_sfixed(-3638.0/65536.0,1,-nbitq), 
to_sfixed(-902.0/65536.0,1,-nbitq), 
to_sfixed(-1103.0/65536.0,1,-nbitq), 
to_sfixed(-4644.0/65536.0,1,-nbitq), 
to_sfixed(-3988.0/65536.0,1,-nbitq), 
to_sfixed(-1183.0/65536.0,1,-nbitq), 
to_sfixed(1755.0/65536.0,1,-nbitq), 
to_sfixed(947.0/65536.0,1,-nbitq), 
to_sfixed(-1196.0/65536.0,1,-nbitq), 
to_sfixed(-1366.0/65536.0,1,-nbitq), 
to_sfixed(-1740.0/65536.0,1,-nbitq), 
to_sfixed(-2443.0/65536.0,1,-nbitq), 
to_sfixed(-1465.0/65536.0,1,-nbitq), 
to_sfixed(-2928.0/65536.0,1,-nbitq), 
to_sfixed(-2409.0/65536.0,1,-nbitq), 
to_sfixed(2692.0/65536.0,1,-nbitq), 
to_sfixed(6008.0/65536.0,1,-nbitq), 
to_sfixed(2417.0/65536.0,1,-nbitq), 
to_sfixed(2292.0/65536.0,1,-nbitq), 
to_sfixed(-1924.0/65536.0,1,-nbitq), 
to_sfixed(-338.0/65536.0,1,-nbitq), 
to_sfixed(-2411.0/65536.0,1,-nbitq), 
to_sfixed(-1273.0/65536.0,1,-nbitq), 
to_sfixed(-1323.0/65536.0,1,-nbitq), 
to_sfixed(-88.0/65536.0,1,-nbitq), 
to_sfixed(-1853.0/65536.0,1,-nbitq), 
to_sfixed(-1502.0/65536.0,1,-nbitq), 
to_sfixed(767.0/65536.0,1,-nbitq), 
to_sfixed(1267.0/65536.0,1,-nbitq), 
to_sfixed(315.0/65536.0,1,-nbitq), 
to_sfixed(4694.0/65536.0,1,-nbitq), 
to_sfixed(-562.0/65536.0,1,-nbitq), 
to_sfixed(385.0/65536.0,1,-nbitq), 
to_sfixed(-2568.0/65536.0,1,-nbitq), 
to_sfixed(-2068.0/65536.0,1,-nbitq), 
to_sfixed(77.0/65536.0,1,-nbitq), 
to_sfixed(3950.0/65536.0,1,-nbitq), 
to_sfixed(316.0/65536.0,1,-nbitq), 
to_sfixed(211.0/65536.0,1,-nbitq), 
to_sfixed(231.0/65536.0,1,-nbitq), 
to_sfixed(1473.0/65536.0,1,-nbitq), 
to_sfixed(-1551.0/65536.0,1,-nbitq), 
to_sfixed(3061.0/65536.0,1,-nbitq), 
to_sfixed(2290.0/65536.0,1,-nbitq), 
to_sfixed(-1834.0/65536.0,1,-nbitq), 
to_sfixed(-1490.0/65536.0,1,-nbitq), 
to_sfixed(-1325.0/65536.0,1,-nbitq), 
to_sfixed(367.0/65536.0,1,-nbitq), 
to_sfixed(4443.0/65536.0,1,-nbitq), 
to_sfixed(237.0/65536.0,1,-nbitq), 
to_sfixed(4728.0/65536.0,1,-nbitq)  ), 
( to_sfixed(503.0/65536.0,1,-nbitq), 
to_sfixed(2863.0/65536.0,1,-nbitq), 
to_sfixed(3123.0/65536.0,1,-nbitq), 
to_sfixed(2835.0/65536.0,1,-nbitq), 
to_sfixed(1131.0/65536.0,1,-nbitq), 
to_sfixed(3529.0/65536.0,1,-nbitq), 
to_sfixed(-3328.0/65536.0,1,-nbitq), 
to_sfixed(518.0/65536.0,1,-nbitq), 
to_sfixed(-774.0/65536.0,1,-nbitq), 
to_sfixed(-2531.0/65536.0,1,-nbitq), 
to_sfixed(-1203.0/65536.0,1,-nbitq), 
to_sfixed(-698.0/65536.0,1,-nbitq), 
to_sfixed(306.0/65536.0,1,-nbitq), 
to_sfixed(-604.0/65536.0,1,-nbitq), 
to_sfixed(4916.0/65536.0,1,-nbitq), 
to_sfixed(1210.0/65536.0,1,-nbitq), 
to_sfixed(74.0/65536.0,1,-nbitq), 
to_sfixed(3318.0/65536.0,1,-nbitq), 
to_sfixed(224.0/65536.0,1,-nbitq), 
to_sfixed(-2528.0/65536.0,1,-nbitq), 
to_sfixed(759.0/65536.0,1,-nbitq), 
to_sfixed(-1572.0/65536.0,1,-nbitq), 
to_sfixed(718.0/65536.0,1,-nbitq), 
to_sfixed(4383.0/65536.0,1,-nbitq), 
to_sfixed(-344.0/65536.0,1,-nbitq), 
to_sfixed(6865.0/65536.0,1,-nbitq), 
to_sfixed(4459.0/65536.0,1,-nbitq), 
to_sfixed(-1882.0/65536.0,1,-nbitq), 
to_sfixed(3811.0/65536.0,1,-nbitq), 
to_sfixed(2859.0/65536.0,1,-nbitq), 
to_sfixed(-3046.0/65536.0,1,-nbitq), 
to_sfixed(6.0/65536.0,1,-nbitq), 
to_sfixed(312.0/65536.0,1,-nbitq), 
to_sfixed(-5348.0/65536.0,1,-nbitq), 
to_sfixed(645.0/65536.0,1,-nbitq), 
to_sfixed(-528.0/65536.0,1,-nbitq), 
to_sfixed(-1567.0/65536.0,1,-nbitq), 
to_sfixed(-1687.0/65536.0,1,-nbitq), 
to_sfixed(-2136.0/65536.0,1,-nbitq), 
to_sfixed(483.0/65536.0,1,-nbitq), 
to_sfixed(-2918.0/65536.0,1,-nbitq), 
to_sfixed(1573.0/65536.0,1,-nbitq), 
to_sfixed(-3342.0/65536.0,1,-nbitq), 
to_sfixed(588.0/65536.0,1,-nbitq), 
to_sfixed(-345.0/65536.0,1,-nbitq), 
to_sfixed(5609.0/65536.0,1,-nbitq), 
to_sfixed(385.0/65536.0,1,-nbitq), 
to_sfixed(-614.0/65536.0,1,-nbitq), 
to_sfixed(-1495.0/65536.0,1,-nbitq), 
to_sfixed(-619.0/65536.0,1,-nbitq), 
to_sfixed(-730.0/65536.0,1,-nbitq), 
to_sfixed(-3057.0/65536.0,1,-nbitq), 
to_sfixed(-358.0/65536.0,1,-nbitq), 
to_sfixed(1073.0/65536.0,1,-nbitq), 
to_sfixed(-1789.0/65536.0,1,-nbitq), 
to_sfixed(5488.0/65536.0,1,-nbitq), 
to_sfixed(2744.0/65536.0,1,-nbitq), 
to_sfixed(2572.0/65536.0,1,-nbitq), 
to_sfixed(-1324.0/65536.0,1,-nbitq), 
to_sfixed(-115.0/65536.0,1,-nbitq), 
to_sfixed(-2892.0/65536.0,1,-nbitq), 
to_sfixed(2046.0/65536.0,1,-nbitq), 
to_sfixed(-2826.0/65536.0,1,-nbitq), 
to_sfixed(-2560.0/65536.0,1,-nbitq), 
to_sfixed(1019.0/65536.0,1,-nbitq), 
to_sfixed(232.0/65536.0,1,-nbitq), 
to_sfixed(-3354.0/65536.0,1,-nbitq), 
to_sfixed(835.0/65536.0,1,-nbitq), 
to_sfixed(2592.0/65536.0,1,-nbitq), 
to_sfixed(-1977.0/65536.0,1,-nbitq), 
to_sfixed(-2220.0/65536.0,1,-nbitq), 
to_sfixed(2466.0/65536.0,1,-nbitq), 
to_sfixed(2117.0/65536.0,1,-nbitq), 
to_sfixed(782.0/65536.0,1,-nbitq), 
to_sfixed(-743.0/65536.0,1,-nbitq), 
to_sfixed(3727.0/65536.0,1,-nbitq), 
to_sfixed(809.0/65536.0,1,-nbitq), 
to_sfixed(-3303.0/65536.0,1,-nbitq), 
to_sfixed(-673.0/65536.0,1,-nbitq), 
to_sfixed(284.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2494.0/65536.0,1,-nbitq), 
to_sfixed(-581.0/65536.0,1,-nbitq), 
to_sfixed(5521.0/65536.0,1,-nbitq), 
to_sfixed(1247.0/65536.0,1,-nbitq), 
to_sfixed(-357.0/65536.0,1,-nbitq), 
to_sfixed(1442.0/65536.0,1,-nbitq), 
to_sfixed(-5304.0/65536.0,1,-nbitq), 
to_sfixed(-1144.0/65536.0,1,-nbitq), 
to_sfixed(1452.0/65536.0,1,-nbitq), 
to_sfixed(2296.0/65536.0,1,-nbitq), 
to_sfixed(4167.0/65536.0,1,-nbitq), 
to_sfixed(3701.0/65536.0,1,-nbitq), 
to_sfixed(3171.0/65536.0,1,-nbitq), 
to_sfixed(4393.0/65536.0,1,-nbitq), 
to_sfixed(1304.0/65536.0,1,-nbitq), 
to_sfixed(-1955.0/65536.0,1,-nbitq), 
to_sfixed(-2037.0/65536.0,1,-nbitq), 
to_sfixed(-4556.0/65536.0,1,-nbitq), 
to_sfixed(3406.0/65536.0,1,-nbitq), 
to_sfixed(1346.0/65536.0,1,-nbitq), 
to_sfixed(-2979.0/65536.0,1,-nbitq), 
to_sfixed(2164.0/65536.0,1,-nbitq), 
to_sfixed(4697.0/65536.0,1,-nbitq), 
to_sfixed(5478.0/65536.0,1,-nbitq), 
to_sfixed(3343.0/65536.0,1,-nbitq), 
to_sfixed(9316.0/65536.0,1,-nbitq), 
to_sfixed(6873.0/65536.0,1,-nbitq), 
to_sfixed(1979.0/65536.0,1,-nbitq), 
to_sfixed(-894.0/65536.0,1,-nbitq), 
to_sfixed(820.0/65536.0,1,-nbitq), 
to_sfixed(-189.0/65536.0,1,-nbitq), 
to_sfixed(664.0/65536.0,1,-nbitq), 
to_sfixed(2209.0/65536.0,1,-nbitq), 
to_sfixed(-2688.0/65536.0,1,-nbitq), 
to_sfixed(-1161.0/65536.0,1,-nbitq), 
to_sfixed(875.0/65536.0,1,-nbitq), 
to_sfixed(-5361.0/65536.0,1,-nbitq), 
to_sfixed(-2389.0/65536.0,1,-nbitq), 
to_sfixed(-2983.0/65536.0,1,-nbitq), 
to_sfixed(-3110.0/65536.0,1,-nbitq), 
to_sfixed(1298.0/65536.0,1,-nbitq), 
to_sfixed(983.0/65536.0,1,-nbitq), 
to_sfixed(-5218.0/65536.0,1,-nbitq), 
to_sfixed(-714.0/65536.0,1,-nbitq), 
to_sfixed(-1468.0/65536.0,1,-nbitq), 
to_sfixed(3584.0/65536.0,1,-nbitq), 
to_sfixed(1160.0/65536.0,1,-nbitq), 
to_sfixed(2758.0/65536.0,1,-nbitq), 
to_sfixed(1555.0/65536.0,1,-nbitq), 
to_sfixed(-519.0/65536.0,1,-nbitq), 
to_sfixed(808.0/65536.0,1,-nbitq), 
to_sfixed(-749.0/65536.0,1,-nbitq), 
to_sfixed(2966.0/65536.0,1,-nbitq), 
to_sfixed(6834.0/65536.0,1,-nbitq), 
to_sfixed(-1537.0/65536.0,1,-nbitq), 
to_sfixed(9024.0/65536.0,1,-nbitq), 
to_sfixed(1190.0/65536.0,1,-nbitq), 
to_sfixed(-741.0/65536.0,1,-nbitq), 
to_sfixed(-1715.0/65536.0,1,-nbitq), 
to_sfixed(2713.0/65536.0,1,-nbitq), 
to_sfixed(-2726.0/65536.0,1,-nbitq), 
to_sfixed(890.0/65536.0,1,-nbitq), 
to_sfixed(2002.0/65536.0,1,-nbitq), 
to_sfixed(-1180.0/65536.0,1,-nbitq), 
to_sfixed(3105.0/65536.0,1,-nbitq), 
to_sfixed(3719.0/65536.0,1,-nbitq), 
to_sfixed(804.0/65536.0,1,-nbitq), 
to_sfixed(-6170.0/65536.0,1,-nbitq), 
to_sfixed(-3372.0/65536.0,1,-nbitq), 
to_sfixed(-7435.0/65536.0,1,-nbitq), 
to_sfixed(956.0/65536.0,1,-nbitq), 
to_sfixed(-2950.0/65536.0,1,-nbitq), 
to_sfixed(-2888.0/65536.0,1,-nbitq), 
to_sfixed(2622.0/65536.0,1,-nbitq), 
to_sfixed(1034.0/65536.0,1,-nbitq), 
to_sfixed(-1793.0/65536.0,1,-nbitq), 
to_sfixed(-3454.0/65536.0,1,-nbitq), 
to_sfixed(-4545.0/65536.0,1,-nbitq), 
to_sfixed(-89.0/65536.0,1,-nbitq), 
to_sfixed(-1625.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2318.0/65536.0,1,-nbitq), 
to_sfixed(-3300.0/65536.0,1,-nbitq), 
to_sfixed(3229.0/65536.0,1,-nbitq), 
to_sfixed(7758.0/65536.0,1,-nbitq), 
to_sfixed(433.0/65536.0,1,-nbitq), 
to_sfixed(2246.0/65536.0,1,-nbitq), 
to_sfixed(-2144.0/65536.0,1,-nbitq), 
to_sfixed(2725.0/65536.0,1,-nbitq), 
to_sfixed(-4120.0/65536.0,1,-nbitq), 
to_sfixed(-218.0/65536.0,1,-nbitq), 
to_sfixed(3240.0/65536.0,1,-nbitq), 
to_sfixed(6335.0/65536.0,1,-nbitq), 
to_sfixed(648.0/65536.0,1,-nbitq), 
to_sfixed(802.0/65536.0,1,-nbitq), 
to_sfixed(-984.0/65536.0,1,-nbitq), 
to_sfixed(-2569.0/65536.0,1,-nbitq), 
to_sfixed(1742.0/65536.0,1,-nbitq), 
to_sfixed(-2211.0/65536.0,1,-nbitq), 
to_sfixed(310.0/65536.0,1,-nbitq), 
to_sfixed(1646.0/65536.0,1,-nbitq), 
to_sfixed(-915.0/65536.0,1,-nbitq), 
to_sfixed(3242.0/65536.0,1,-nbitq), 
to_sfixed(219.0/65536.0,1,-nbitq), 
to_sfixed(4682.0/65536.0,1,-nbitq), 
to_sfixed(2492.0/65536.0,1,-nbitq), 
to_sfixed(6339.0/65536.0,1,-nbitq), 
to_sfixed(9348.0/65536.0,1,-nbitq), 
to_sfixed(2344.0/65536.0,1,-nbitq), 
to_sfixed(5200.0/65536.0,1,-nbitq), 
to_sfixed(4074.0/65536.0,1,-nbitq), 
to_sfixed(2007.0/65536.0,1,-nbitq), 
to_sfixed(4144.0/65536.0,1,-nbitq), 
to_sfixed(3537.0/65536.0,1,-nbitq), 
to_sfixed(-9149.0/65536.0,1,-nbitq), 
to_sfixed(-1979.0/65536.0,1,-nbitq), 
to_sfixed(-1221.0/65536.0,1,-nbitq), 
to_sfixed(-6800.0/65536.0,1,-nbitq), 
to_sfixed(4433.0/65536.0,1,-nbitq), 
to_sfixed(-8552.0/65536.0,1,-nbitq), 
to_sfixed(-10443.0/65536.0,1,-nbitq), 
to_sfixed(5235.0/65536.0,1,-nbitq), 
to_sfixed(1525.0/65536.0,1,-nbitq), 
to_sfixed(-1885.0/65536.0,1,-nbitq), 
to_sfixed(-693.0/65536.0,1,-nbitq), 
to_sfixed(-96.0/65536.0,1,-nbitq), 
to_sfixed(3322.0/65536.0,1,-nbitq), 
to_sfixed(1299.0/65536.0,1,-nbitq), 
to_sfixed(-2197.0/65536.0,1,-nbitq), 
to_sfixed(-594.0/65536.0,1,-nbitq), 
to_sfixed(643.0/65536.0,1,-nbitq), 
to_sfixed(2036.0/65536.0,1,-nbitq), 
to_sfixed(-825.0/65536.0,1,-nbitq), 
to_sfixed(2102.0/65536.0,1,-nbitq), 
to_sfixed(3546.0/65536.0,1,-nbitq), 
to_sfixed(-5086.0/65536.0,1,-nbitq), 
to_sfixed(9103.0/65536.0,1,-nbitq), 
to_sfixed(-43.0/65536.0,1,-nbitq), 
to_sfixed(-2341.0/65536.0,1,-nbitq), 
to_sfixed(-1060.0/65536.0,1,-nbitq), 
to_sfixed(-4639.0/65536.0,1,-nbitq), 
to_sfixed(-8059.0/65536.0,1,-nbitq), 
to_sfixed(1827.0/65536.0,1,-nbitq), 
to_sfixed(-54.0/65536.0,1,-nbitq), 
to_sfixed(2344.0/65536.0,1,-nbitq), 
to_sfixed(2665.0/65536.0,1,-nbitq), 
to_sfixed(6391.0/65536.0,1,-nbitq), 
to_sfixed(-3948.0/65536.0,1,-nbitq), 
to_sfixed(-5069.0/65536.0,1,-nbitq), 
to_sfixed(-3044.0/65536.0,1,-nbitq), 
to_sfixed(-717.0/65536.0,1,-nbitq), 
to_sfixed(358.0/65536.0,1,-nbitq), 
to_sfixed(420.0/65536.0,1,-nbitq), 
to_sfixed(-508.0/65536.0,1,-nbitq), 
to_sfixed(-3288.0/65536.0,1,-nbitq), 
to_sfixed(-1254.0/65536.0,1,-nbitq), 
to_sfixed(-1653.0/65536.0,1,-nbitq), 
to_sfixed(-291.0/65536.0,1,-nbitq), 
to_sfixed(-1412.0/65536.0,1,-nbitq), 
to_sfixed(1085.0/65536.0,1,-nbitq), 
to_sfixed(-1019.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2112.0/65536.0,1,-nbitq), 
to_sfixed(439.0/65536.0,1,-nbitq), 
to_sfixed(1382.0/65536.0,1,-nbitq), 
to_sfixed(3836.0/65536.0,1,-nbitq), 
to_sfixed(961.0/65536.0,1,-nbitq), 
to_sfixed(3524.0/65536.0,1,-nbitq), 
to_sfixed(-115.0/65536.0,1,-nbitq), 
to_sfixed(-2162.0/65536.0,1,-nbitq), 
to_sfixed(2598.0/65536.0,1,-nbitq), 
to_sfixed(256.0/65536.0,1,-nbitq), 
to_sfixed(2571.0/65536.0,1,-nbitq), 
to_sfixed(18906.0/65536.0,1,-nbitq), 
to_sfixed(-761.0/65536.0,1,-nbitq), 
to_sfixed(6102.0/65536.0,1,-nbitq), 
to_sfixed(-7099.0/65536.0,1,-nbitq), 
to_sfixed(-2559.0/65536.0,1,-nbitq), 
to_sfixed(2583.0/65536.0,1,-nbitq), 
to_sfixed(3390.0/65536.0,1,-nbitq), 
to_sfixed(3670.0/65536.0,1,-nbitq), 
to_sfixed(1624.0/65536.0,1,-nbitq), 
to_sfixed(730.0/65536.0,1,-nbitq), 
to_sfixed(-3741.0/65536.0,1,-nbitq), 
to_sfixed(4423.0/65536.0,1,-nbitq), 
to_sfixed(-6167.0/65536.0,1,-nbitq), 
to_sfixed(139.0/65536.0,1,-nbitq), 
to_sfixed(3741.0/65536.0,1,-nbitq), 
to_sfixed(5923.0/65536.0,1,-nbitq), 
to_sfixed(2799.0/65536.0,1,-nbitq), 
to_sfixed(-3002.0/65536.0,1,-nbitq), 
to_sfixed(606.0/65536.0,1,-nbitq), 
to_sfixed(-1950.0/65536.0,1,-nbitq), 
to_sfixed(-4382.0/65536.0,1,-nbitq), 
to_sfixed(-2004.0/65536.0,1,-nbitq), 
to_sfixed(-6522.0/65536.0,1,-nbitq), 
to_sfixed(-1908.0/65536.0,1,-nbitq), 
to_sfixed(2368.0/65536.0,1,-nbitq), 
to_sfixed(-11597.0/65536.0,1,-nbitq), 
to_sfixed(8496.0/65536.0,1,-nbitq), 
to_sfixed(-11329.0/65536.0,1,-nbitq), 
to_sfixed(-10536.0/65536.0,1,-nbitq), 
to_sfixed(1431.0/65536.0,1,-nbitq), 
to_sfixed(1187.0/65536.0,1,-nbitq), 
to_sfixed(-6368.0/65536.0,1,-nbitq), 
to_sfixed(-2254.0/65536.0,1,-nbitq), 
to_sfixed(-2695.0/65536.0,1,-nbitq), 
to_sfixed(100.0/65536.0,1,-nbitq), 
to_sfixed(-2599.0/65536.0,1,-nbitq), 
to_sfixed(-2185.0/65536.0,1,-nbitq), 
to_sfixed(1850.0/65536.0,1,-nbitq), 
to_sfixed(-571.0/65536.0,1,-nbitq), 
to_sfixed(2066.0/65536.0,1,-nbitq), 
to_sfixed(2958.0/65536.0,1,-nbitq), 
to_sfixed(-1268.0/65536.0,1,-nbitq), 
to_sfixed(9893.0/65536.0,1,-nbitq), 
to_sfixed(-7861.0/65536.0,1,-nbitq), 
to_sfixed(13933.0/65536.0,1,-nbitq), 
to_sfixed(757.0/65536.0,1,-nbitq), 
to_sfixed(879.0/65536.0,1,-nbitq), 
to_sfixed(2552.0/65536.0,1,-nbitq), 
to_sfixed(985.0/65536.0,1,-nbitq), 
to_sfixed(-3997.0/65536.0,1,-nbitq), 
to_sfixed(-8.0/65536.0,1,-nbitq), 
to_sfixed(-1912.0/65536.0,1,-nbitq), 
to_sfixed(-627.0/65536.0,1,-nbitq), 
to_sfixed(-296.0/65536.0,1,-nbitq), 
to_sfixed(3135.0/65536.0,1,-nbitq), 
to_sfixed(-1024.0/65536.0,1,-nbitq), 
to_sfixed(-11450.0/65536.0,1,-nbitq), 
to_sfixed(-8666.0/65536.0,1,-nbitq), 
to_sfixed(6560.0/65536.0,1,-nbitq), 
to_sfixed(666.0/65536.0,1,-nbitq), 
to_sfixed(-196.0/65536.0,1,-nbitq), 
to_sfixed(-494.0/65536.0,1,-nbitq), 
to_sfixed(483.0/65536.0,1,-nbitq), 
to_sfixed(2437.0/65536.0,1,-nbitq), 
to_sfixed(-4102.0/65536.0,1,-nbitq), 
to_sfixed(893.0/65536.0,1,-nbitq), 
to_sfixed(-4500.0/65536.0,1,-nbitq), 
to_sfixed(2614.0/65536.0,1,-nbitq), 
to_sfixed(-4506.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3178.0/65536.0,1,-nbitq), 
to_sfixed(-324.0/65536.0,1,-nbitq), 
to_sfixed(4831.0/65536.0,1,-nbitq), 
to_sfixed(4614.0/65536.0,1,-nbitq), 
to_sfixed(-8734.0/65536.0,1,-nbitq), 
to_sfixed(5611.0/65536.0,1,-nbitq), 
to_sfixed(-955.0/65536.0,1,-nbitq), 
to_sfixed(-9324.0/65536.0,1,-nbitq), 
to_sfixed(2991.0/65536.0,1,-nbitq), 
to_sfixed(-32.0/65536.0,1,-nbitq), 
to_sfixed(3737.0/65536.0,1,-nbitq), 
to_sfixed(15510.0/65536.0,1,-nbitq), 
to_sfixed(2932.0/65536.0,1,-nbitq), 
to_sfixed(4252.0/65536.0,1,-nbitq), 
to_sfixed(-5674.0/65536.0,1,-nbitq), 
to_sfixed(507.0/65536.0,1,-nbitq), 
to_sfixed(637.0/65536.0,1,-nbitq), 
to_sfixed(7348.0/65536.0,1,-nbitq), 
to_sfixed(6805.0/65536.0,1,-nbitq), 
to_sfixed(347.0/65536.0,1,-nbitq), 
to_sfixed(-6012.0/65536.0,1,-nbitq), 
to_sfixed(-9832.0/65536.0,1,-nbitq), 
to_sfixed(-12236.0/65536.0,1,-nbitq), 
to_sfixed(-51.0/65536.0,1,-nbitq), 
to_sfixed(-817.0/65536.0,1,-nbitq), 
to_sfixed(13703.0/65536.0,1,-nbitq), 
to_sfixed(5118.0/65536.0,1,-nbitq), 
to_sfixed(2353.0/65536.0,1,-nbitq), 
to_sfixed(-2834.0/65536.0,1,-nbitq), 
to_sfixed(-7021.0/65536.0,1,-nbitq), 
to_sfixed(-846.0/65536.0,1,-nbitq), 
to_sfixed(-954.0/65536.0,1,-nbitq), 
to_sfixed(-5825.0/65536.0,1,-nbitq), 
to_sfixed(-2223.0/65536.0,1,-nbitq), 
to_sfixed(-4056.0/65536.0,1,-nbitq), 
to_sfixed(3094.0/65536.0,1,-nbitq), 
to_sfixed(-9430.0/65536.0,1,-nbitq), 
to_sfixed(6388.0/65536.0,1,-nbitq), 
to_sfixed(-15705.0/65536.0,1,-nbitq), 
to_sfixed(-8525.0/65536.0,1,-nbitq), 
to_sfixed(8272.0/65536.0,1,-nbitq), 
to_sfixed(1400.0/65536.0,1,-nbitq), 
to_sfixed(-4286.0/65536.0,1,-nbitq), 
to_sfixed(-2962.0/65536.0,1,-nbitq), 
to_sfixed(2328.0/65536.0,1,-nbitq), 
to_sfixed(329.0/65536.0,1,-nbitq), 
to_sfixed(2102.0/65536.0,1,-nbitq), 
to_sfixed(-1886.0/65536.0,1,-nbitq), 
to_sfixed(-518.0/65536.0,1,-nbitq), 
to_sfixed(841.0/65536.0,1,-nbitq), 
to_sfixed(-1848.0/65536.0,1,-nbitq), 
to_sfixed(2436.0/65536.0,1,-nbitq), 
to_sfixed(141.0/65536.0,1,-nbitq), 
to_sfixed(357.0/65536.0,1,-nbitq), 
to_sfixed(-1587.0/65536.0,1,-nbitq), 
to_sfixed(11036.0/65536.0,1,-nbitq), 
to_sfixed(3067.0/65536.0,1,-nbitq), 
to_sfixed(834.0/65536.0,1,-nbitq), 
to_sfixed(-1489.0/65536.0,1,-nbitq), 
to_sfixed(5148.0/65536.0,1,-nbitq), 
to_sfixed(-3014.0/65536.0,1,-nbitq), 
to_sfixed(-2172.0/65536.0,1,-nbitq), 
to_sfixed(413.0/65536.0,1,-nbitq), 
to_sfixed(1005.0/65536.0,1,-nbitq), 
to_sfixed(2438.0/65536.0,1,-nbitq), 
to_sfixed(10377.0/65536.0,1,-nbitq), 
to_sfixed(5866.0/65536.0,1,-nbitq), 
to_sfixed(3612.0/65536.0,1,-nbitq), 
to_sfixed(-9457.0/65536.0,1,-nbitq), 
to_sfixed(-261.0/65536.0,1,-nbitq), 
to_sfixed(-2779.0/65536.0,1,-nbitq), 
to_sfixed(-4692.0/65536.0,1,-nbitq), 
to_sfixed(-1831.0/65536.0,1,-nbitq), 
to_sfixed(1380.0/65536.0,1,-nbitq), 
to_sfixed(-2506.0/65536.0,1,-nbitq), 
to_sfixed(-2498.0/65536.0,1,-nbitq), 
to_sfixed(9189.0/65536.0,1,-nbitq), 
to_sfixed(-3947.0/65536.0,1,-nbitq), 
to_sfixed(-837.0/65536.0,1,-nbitq), 
to_sfixed(-4668.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1369.0/65536.0,1,-nbitq), 
to_sfixed(-775.0/65536.0,1,-nbitq), 
to_sfixed(-984.0/65536.0,1,-nbitq), 
to_sfixed(6314.0/65536.0,1,-nbitq), 
to_sfixed(-7519.0/65536.0,1,-nbitq), 
to_sfixed(2791.0/65536.0,1,-nbitq), 
to_sfixed(-1858.0/65536.0,1,-nbitq), 
to_sfixed(-2187.0/65536.0,1,-nbitq), 
to_sfixed(2245.0/65536.0,1,-nbitq), 
to_sfixed(551.0/65536.0,1,-nbitq), 
to_sfixed(6057.0/65536.0,1,-nbitq), 
to_sfixed(2782.0/65536.0,1,-nbitq), 
to_sfixed(2509.0/65536.0,1,-nbitq), 
to_sfixed(5155.0/65536.0,1,-nbitq), 
to_sfixed(-476.0/65536.0,1,-nbitq), 
to_sfixed(-1152.0/65536.0,1,-nbitq), 
to_sfixed(861.0/65536.0,1,-nbitq), 
to_sfixed(8004.0/65536.0,1,-nbitq), 
to_sfixed(412.0/65536.0,1,-nbitq), 
to_sfixed(234.0/65536.0,1,-nbitq), 
to_sfixed(-7062.0/65536.0,1,-nbitq), 
to_sfixed(-2652.0/65536.0,1,-nbitq), 
to_sfixed(-11875.0/65536.0,1,-nbitq), 
to_sfixed(6430.0/65536.0,1,-nbitq), 
to_sfixed(-765.0/65536.0,1,-nbitq), 
to_sfixed(13491.0/65536.0,1,-nbitq), 
to_sfixed(6342.0/65536.0,1,-nbitq), 
to_sfixed(6255.0/65536.0,1,-nbitq), 
to_sfixed(10183.0/65536.0,1,-nbitq), 
to_sfixed(-11177.0/65536.0,1,-nbitq), 
to_sfixed(-5157.0/65536.0,1,-nbitq), 
to_sfixed(-221.0/65536.0,1,-nbitq), 
to_sfixed(-420.0/65536.0,1,-nbitq), 
to_sfixed(-3217.0/65536.0,1,-nbitq), 
to_sfixed(311.0/65536.0,1,-nbitq), 
to_sfixed(1566.0/65536.0,1,-nbitq), 
to_sfixed(-9414.0/65536.0,1,-nbitq), 
to_sfixed(3958.0/65536.0,1,-nbitq), 
to_sfixed(-12163.0/65536.0,1,-nbitq), 
to_sfixed(-7151.0/65536.0,1,-nbitq), 
to_sfixed(3506.0/65536.0,1,-nbitq), 
to_sfixed(-2252.0/65536.0,1,-nbitq), 
to_sfixed(-2846.0/65536.0,1,-nbitq), 
to_sfixed(-6628.0/65536.0,1,-nbitq), 
to_sfixed(-621.0/65536.0,1,-nbitq), 
to_sfixed(-2721.0/65536.0,1,-nbitq), 
to_sfixed(501.0/65536.0,1,-nbitq), 
to_sfixed(7856.0/65536.0,1,-nbitq), 
to_sfixed(2898.0/65536.0,1,-nbitq), 
to_sfixed(515.0/65536.0,1,-nbitq), 
to_sfixed(1088.0/65536.0,1,-nbitq), 
to_sfixed(2745.0/65536.0,1,-nbitq), 
to_sfixed(-3286.0/65536.0,1,-nbitq), 
to_sfixed(6182.0/65536.0,1,-nbitq), 
to_sfixed(-1790.0/65536.0,1,-nbitq), 
to_sfixed(5851.0/65536.0,1,-nbitq), 
to_sfixed(2420.0/65536.0,1,-nbitq), 
to_sfixed(3007.0/65536.0,1,-nbitq), 
to_sfixed(1822.0/65536.0,1,-nbitq), 
to_sfixed(2522.0/65536.0,1,-nbitq), 
to_sfixed(8656.0/65536.0,1,-nbitq), 
to_sfixed(2820.0/65536.0,1,-nbitq), 
to_sfixed(-2733.0/65536.0,1,-nbitq), 
to_sfixed(-233.0/65536.0,1,-nbitq), 
to_sfixed(-277.0/65536.0,1,-nbitq), 
to_sfixed(1855.0/65536.0,1,-nbitq), 
to_sfixed(591.0/65536.0,1,-nbitq), 
to_sfixed(6203.0/65536.0,1,-nbitq), 
to_sfixed(-2088.0/65536.0,1,-nbitq), 
to_sfixed(3326.0/65536.0,1,-nbitq), 
to_sfixed(-4010.0/65536.0,1,-nbitq), 
to_sfixed(-11170.0/65536.0,1,-nbitq), 
to_sfixed(-877.0/65536.0,1,-nbitq), 
to_sfixed(-2077.0/65536.0,1,-nbitq), 
to_sfixed(-1227.0/65536.0,1,-nbitq), 
to_sfixed(3354.0/65536.0,1,-nbitq), 
to_sfixed(3674.0/65536.0,1,-nbitq), 
to_sfixed(-1877.0/65536.0,1,-nbitq), 
to_sfixed(881.0/65536.0,1,-nbitq), 
to_sfixed(-677.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1242.0/65536.0,1,-nbitq), 
to_sfixed(4620.0/65536.0,1,-nbitq), 
to_sfixed(662.0/65536.0,1,-nbitq), 
to_sfixed(7824.0/65536.0,1,-nbitq), 
to_sfixed(-10591.0/65536.0,1,-nbitq), 
to_sfixed(-809.0/65536.0,1,-nbitq), 
to_sfixed(-2396.0/65536.0,1,-nbitq), 
to_sfixed(2997.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(1932.0/65536.0,1,-nbitq), 
to_sfixed(252.0/65536.0,1,-nbitq), 
to_sfixed(-2724.0/65536.0,1,-nbitq), 
to_sfixed(-2481.0/65536.0,1,-nbitq), 
to_sfixed(9427.0/65536.0,1,-nbitq), 
to_sfixed(4201.0/65536.0,1,-nbitq), 
to_sfixed(-457.0/65536.0,1,-nbitq), 
to_sfixed(1836.0/65536.0,1,-nbitq), 
to_sfixed(7041.0/65536.0,1,-nbitq), 
to_sfixed(2561.0/65536.0,1,-nbitq), 
to_sfixed(1065.0/65536.0,1,-nbitq), 
to_sfixed(-9900.0/65536.0,1,-nbitq), 
to_sfixed(-5506.0/65536.0,1,-nbitq), 
to_sfixed(3421.0/65536.0,1,-nbitq), 
to_sfixed(6738.0/65536.0,1,-nbitq), 
to_sfixed(-3454.0/65536.0,1,-nbitq), 
to_sfixed(9354.0/65536.0,1,-nbitq), 
to_sfixed(2857.0/65536.0,1,-nbitq), 
to_sfixed(2413.0/65536.0,1,-nbitq), 
to_sfixed(2949.0/65536.0,1,-nbitq), 
to_sfixed(-10588.0/65536.0,1,-nbitq), 
to_sfixed(-1818.0/65536.0,1,-nbitq), 
to_sfixed(778.0/65536.0,1,-nbitq), 
to_sfixed(-1368.0/65536.0,1,-nbitq), 
to_sfixed(-8056.0/65536.0,1,-nbitq), 
to_sfixed(319.0/65536.0,1,-nbitq), 
to_sfixed(3476.0/65536.0,1,-nbitq), 
to_sfixed(-6926.0/65536.0,1,-nbitq), 
to_sfixed(-2058.0/65536.0,1,-nbitq), 
to_sfixed(-9326.0/65536.0,1,-nbitq), 
to_sfixed(-2786.0/65536.0,1,-nbitq), 
to_sfixed(1476.0/65536.0,1,-nbitq), 
to_sfixed(2101.0/65536.0,1,-nbitq), 
to_sfixed(-3327.0/65536.0,1,-nbitq), 
to_sfixed(-9509.0/65536.0,1,-nbitq), 
to_sfixed(958.0/65536.0,1,-nbitq), 
to_sfixed(-16096.0/65536.0,1,-nbitq), 
to_sfixed(3517.0/65536.0,1,-nbitq), 
to_sfixed(2859.0/65536.0,1,-nbitq), 
to_sfixed(-1102.0/65536.0,1,-nbitq), 
to_sfixed(2111.0/65536.0,1,-nbitq), 
to_sfixed(249.0/65536.0,1,-nbitq), 
to_sfixed(4815.0/65536.0,1,-nbitq), 
to_sfixed(-3452.0/65536.0,1,-nbitq), 
to_sfixed(8931.0/65536.0,1,-nbitq), 
to_sfixed(-3607.0/65536.0,1,-nbitq), 
to_sfixed(1956.0/65536.0,1,-nbitq), 
to_sfixed(2818.0/65536.0,1,-nbitq), 
to_sfixed(-423.0/65536.0,1,-nbitq), 
to_sfixed(2620.0/65536.0,1,-nbitq), 
to_sfixed(1755.0/65536.0,1,-nbitq), 
to_sfixed(16561.0/65536.0,1,-nbitq), 
to_sfixed(-760.0/65536.0,1,-nbitq), 
to_sfixed(-1829.0/65536.0,1,-nbitq), 
to_sfixed(-3601.0/65536.0,1,-nbitq), 
to_sfixed(3306.0/65536.0,1,-nbitq), 
to_sfixed(2740.0/65536.0,1,-nbitq), 
to_sfixed(-1847.0/65536.0,1,-nbitq), 
to_sfixed(-4579.0/65536.0,1,-nbitq), 
to_sfixed(-3015.0/65536.0,1,-nbitq), 
to_sfixed(2382.0/65536.0,1,-nbitq), 
to_sfixed(-693.0/65536.0,1,-nbitq), 
to_sfixed(-5486.0/65536.0,1,-nbitq), 
to_sfixed(-63.0/65536.0,1,-nbitq), 
to_sfixed(-1422.0/65536.0,1,-nbitq), 
to_sfixed(3070.0/65536.0,1,-nbitq), 
to_sfixed(2634.0/65536.0,1,-nbitq), 
to_sfixed(-6724.0/65536.0,1,-nbitq), 
to_sfixed(-8001.0/65536.0,1,-nbitq), 
to_sfixed(-1965.0/65536.0,1,-nbitq), 
to_sfixed(-929.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2770.0/65536.0,1,-nbitq), 
to_sfixed(5764.0/65536.0,1,-nbitq), 
to_sfixed(-2350.0/65536.0,1,-nbitq), 
to_sfixed(6418.0/65536.0,1,-nbitq), 
to_sfixed(-2093.0/65536.0,1,-nbitq), 
to_sfixed(8039.0/65536.0,1,-nbitq), 
to_sfixed(-1542.0/65536.0,1,-nbitq), 
to_sfixed(291.0/65536.0,1,-nbitq), 
to_sfixed(-3254.0/65536.0,1,-nbitq), 
to_sfixed(-1079.0/65536.0,1,-nbitq), 
to_sfixed(2279.0/65536.0,1,-nbitq), 
to_sfixed(-2729.0/65536.0,1,-nbitq), 
to_sfixed(-1256.0/65536.0,1,-nbitq), 
to_sfixed(-3003.0/65536.0,1,-nbitq), 
to_sfixed(-224.0/65536.0,1,-nbitq), 
to_sfixed(-196.0/65536.0,1,-nbitq), 
to_sfixed(2557.0/65536.0,1,-nbitq), 
to_sfixed(10110.0/65536.0,1,-nbitq), 
to_sfixed(-6480.0/65536.0,1,-nbitq), 
to_sfixed(2650.0/65536.0,1,-nbitq), 
to_sfixed(-6884.0/65536.0,1,-nbitq), 
to_sfixed(-10163.0/65536.0,1,-nbitq), 
to_sfixed(4042.0/65536.0,1,-nbitq), 
to_sfixed(3483.0/65536.0,1,-nbitq), 
to_sfixed(-745.0/65536.0,1,-nbitq), 
to_sfixed(10769.0/65536.0,1,-nbitq), 
to_sfixed(-1333.0/65536.0,1,-nbitq), 
to_sfixed(3646.0/65536.0,1,-nbitq), 
to_sfixed(5667.0/65536.0,1,-nbitq), 
to_sfixed(-3765.0/65536.0,1,-nbitq), 
to_sfixed(1795.0/65536.0,1,-nbitq), 
to_sfixed(2251.0/65536.0,1,-nbitq), 
to_sfixed(6326.0/65536.0,1,-nbitq), 
to_sfixed(10485.0/65536.0,1,-nbitq), 
to_sfixed(-2759.0/65536.0,1,-nbitq), 
to_sfixed(3655.0/65536.0,1,-nbitq), 
to_sfixed(4685.0/65536.0,1,-nbitq), 
to_sfixed(-9042.0/65536.0,1,-nbitq), 
to_sfixed(-13193.0/65536.0,1,-nbitq), 
to_sfixed(-3596.0/65536.0,1,-nbitq), 
to_sfixed(1616.0/65536.0,1,-nbitq), 
to_sfixed(-85.0/65536.0,1,-nbitq), 
to_sfixed(2495.0/65536.0,1,-nbitq), 
to_sfixed(-9034.0/65536.0,1,-nbitq), 
to_sfixed(582.0/65536.0,1,-nbitq), 
to_sfixed(-12747.0/65536.0,1,-nbitq), 
to_sfixed(2829.0/65536.0,1,-nbitq), 
to_sfixed(-2645.0/65536.0,1,-nbitq), 
to_sfixed(3852.0/65536.0,1,-nbitq), 
to_sfixed(1183.0/65536.0,1,-nbitq), 
to_sfixed(2422.0/65536.0,1,-nbitq), 
to_sfixed(5951.0/65536.0,1,-nbitq), 
to_sfixed(1037.0/65536.0,1,-nbitq), 
to_sfixed(-1344.0/65536.0,1,-nbitq), 
to_sfixed(-4648.0/65536.0,1,-nbitq), 
to_sfixed(4145.0/65536.0,1,-nbitq), 
to_sfixed(-695.0/65536.0,1,-nbitq), 
to_sfixed(-7167.0/65536.0,1,-nbitq), 
to_sfixed(-299.0/65536.0,1,-nbitq), 
to_sfixed(331.0/65536.0,1,-nbitq), 
to_sfixed(20128.0/65536.0,1,-nbitq), 
to_sfixed(51.0/65536.0,1,-nbitq), 
to_sfixed(2729.0/65536.0,1,-nbitq), 
to_sfixed(1998.0/65536.0,1,-nbitq), 
to_sfixed(11585.0/65536.0,1,-nbitq), 
to_sfixed(10463.0/65536.0,1,-nbitq), 
to_sfixed(-3691.0/65536.0,1,-nbitq), 
to_sfixed(1264.0/65536.0,1,-nbitq), 
to_sfixed(4075.0/65536.0,1,-nbitq), 
to_sfixed(-3993.0/65536.0,1,-nbitq), 
to_sfixed(-2168.0/65536.0,1,-nbitq), 
to_sfixed(-9550.0/65536.0,1,-nbitq), 
to_sfixed(2159.0/65536.0,1,-nbitq), 
to_sfixed(37.0/65536.0,1,-nbitq), 
to_sfixed(-1965.0/65536.0,1,-nbitq), 
to_sfixed(5366.0/65536.0,1,-nbitq), 
to_sfixed(-10394.0/65536.0,1,-nbitq), 
to_sfixed(-11851.0/65536.0,1,-nbitq), 
to_sfixed(1787.0/65536.0,1,-nbitq), 
to_sfixed(-2752.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4869.0/65536.0,1,-nbitq), 
to_sfixed(9753.0/65536.0,1,-nbitq), 
to_sfixed(3672.0/65536.0,1,-nbitq), 
to_sfixed(11708.0/65536.0,1,-nbitq), 
to_sfixed(975.0/65536.0,1,-nbitq), 
to_sfixed(5653.0/65536.0,1,-nbitq), 
to_sfixed(772.0/65536.0,1,-nbitq), 
to_sfixed(9038.0/65536.0,1,-nbitq), 
to_sfixed(1284.0/65536.0,1,-nbitq), 
to_sfixed(2014.0/65536.0,1,-nbitq), 
to_sfixed(3852.0/65536.0,1,-nbitq), 
to_sfixed(2536.0/65536.0,1,-nbitq), 
to_sfixed(-95.0/65536.0,1,-nbitq), 
to_sfixed(-12718.0/65536.0,1,-nbitq), 
to_sfixed(-1097.0/65536.0,1,-nbitq), 
to_sfixed(1176.0/65536.0,1,-nbitq), 
to_sfixed(239.0/65536.0,1,-nbitq), 
to_sfixed(17526.0/65536.0,1,-nbitq), 
to_sfixed(-12052.0/65536.0,1,-nbitq), 
to_sfixed(1235.0/65536.0,1,-nbitq), 
to_sfixed(-3595.0/65536.0,1,-nbitq), 
to_sfixed(-14990.0/65536.0,1,-nbitq), 
to_sfixed(-1069.0/65536.0,1,-nbitq), 
to_sfixed(5421.0/65536.0,1,-nbitq), 
to_sfixed(-4076.0/65536.0,1,-nbitq), 
to_sfixed(9962.0/65536.0,1,-nbitq), 
to_sfixed(1404.0/65536.0,1,-nbitq), 
to_sfixed(3872.0/65536.0,1,-nbitq), 
to_sfixed(13528.0/65536.0,1,-nbitq), 
to_sfixed(-2537.0/65536.0,1,-nbitq), 
to_sfixed(-148.0/65536.0,1,-nbitq), 
to_sfixed(2728.0/65536.0,1,-nbitq), 
to_sfixed(4066.0/65536.0,1,-nbitq), 
to_sfixed(17894.0/65536.0,1,-nbitq), 
to_sfixed(-2463.0/65536.0,1,-nbitq), 
to_sfixed(2581.0/65536.0,1,-nbitq), 
to_sfixed(6778.0/65536.0,1,-nbitq), 
to_sfixed(-4076.0/65536.0,1,-nbitq), 
to_sfixed(-9023.0/65536.0,1,-nbitq), 
to_sfixed(-2173.0/65536.0,1,-nbitq), 
to_sfixed(3615.0/65536.0,1,-nbitq), 
to_sfixed(635.0/65536.0,1,-nbitq), 
to_sfixed(1164.0/65536.0,1,-nbitq), 
to_sfixed(-13120.0/65536.0,1,-nbitq), 
to_sfixed(1408.0/65536.0,1,-nbitq), 
to_sfixed(-14476.0/65536.0,1,-nbitq), 
to_sfixed(1832.0/65536.0,1,-nbitq), 
to_sfixed(959.0/65536.0,1,-nbitq), 
to_sfixed(1670.0/65536.0,1,-nbitq), 
to_sfixed(311.0/65536.0,1,-nbitq), 
to_sfixed(-1808.0/65536.0,1,-nbitq), 
to_sfixed(3223.0/65536.0,1,-nbitq), 
to_sfixed(989.0/65536.0,1,-nbitq), 
to_sfixed(5754.0/65536.0,1,-nbitq), 
to_sfixed(-5602.0/65536.0,1,-nbitq), 
to_sfixed(7909.0/65536.0,1,-nbitq), 
to_sfixed(2753.0/65536.0,1,-nbitq), 
to_sfixed(-2506.0/65536.0,1,-nbitq), 
to_sfixed(2975.0/65536.0,1,-nbitq), 
to_sfixed(8336.0/65536.0,1,-nbitq), 
to_sfixed(17349.0/65536.0,1,-nbitq), 
to_sfixed(-231.0/65536.0,1,-nbitq), 
to_sfixed(-2679.0/65536.0,1,-nbitq), 
to_sfixed(2120.0/65536.0,1,-nbitq), 
to_sfixed(6841.0/65536.0,1,-nbitq), 
to_sfixed(-1141.0/65536.0,1,-nbitq), 
to_sfixed(-1356.0/65536.0,1,-nbitq), 
to_sfixed(-3868.0/65536.0,1,-nbitq), 
to_sfixed(5407.0/65536.0,1,-nbitq), 
to_sfixed(-15305.0/65536.0,1,-nbitq), 
to_sfixed(636.0/65536.0,1,-nbitq), 
to_sfixed(-6376.0/65536.0,1,-nbitq), 
to_sfixed(2174.0/65536.0,1,-nbitq), 
to_sfixed(1715.0/65536.0,1,-nbitq), 
to_sfixed(-2593.0/65536.0,1,-nbitq), 
to_sfixed(-4306.0/65536.0,1,-nbitq), 
to_sfixed(-5565.0/65536.0,1,-nbitq), 
to_sfixed(-4001.0/65536.0,1,-nbitq), 
to_sfixed(-1587.0/65536.0,1,-nbitq), 
to_sfixed(886.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4687.0/65536.0,1,-nbitq), 
to_sfixed(7302.0/65536.0,1,-nbitq), 
to_sfixed(2716.0/65536.0,1,-nbitq), 
to_sfixed(14397.0/65536.0,1,-nbitq), 
to_sfixed(-433.0/65536.0,1,-nbitq), 
to_sfixed(6762.0/65536.0,1,-nbitq), 
to_sfixed(3009.0/65536.0,1,-nbitq), 
to_sfixed(11936.0/65536.0,1,-nbitq), 
to_sfixed(1845.0/65536.0,1,-nbitq), 
to_sfixed(4203.0/65536.0,1,-nbitq), 
to_sfixed(6278.0/65536.0,1,-nbitq), 
to_sfixed(169.0/65536.0,1,-nbitq), 
to_sfixed(-1085.0/65536.0,1,-nbitq), 
to_sfixed(-12237.0/65536.0,1,-nbitq), 
to_sfixed(-9031.0/65536.0,1,-nbitq), 
to_sfixed(2678.0/65536.0,1,-nbitq), 
to_sfixed(101.0/65536.0,1,-nbitq), 
to_sfixed(-15426.0/65536.0,1,-nbitq), 
to_sfixed(-8245.0/65536.0,1,-nbitq), 
to_sfixed(596.0/65536.0,1,-nbitq), 
to_sfixed(-10380.0/65536.0,1,-nbitq), 
to_sfixed(-16339.0/65536.0,1,-nbitq), 
to_sfixed(-2527.0/65536.0,1,-nbitq), 
to_sfixed(2189.0/65536.0,1,-nbitq), 
to_sfixed(1853.0/65536.0,1,-nbitq), 
to_sfixed(4870.0/65536.0,1,-nbitq), 
to_sfixed(-1449.0/65536.0,1,-nbitq), 
to_sfixed(1239.0/65536.0,1,-nbitq), 
to_sfixed(14537.0/65536.0,1,-nbitq), 
to_sfixed(214.0/65536.0,1,-nbitq), 
to_sfixed(-6049.0/65536.0,1,-nbitq), 
to_sfixed(548.0/65536.0,1,-nbitq), 
to_sfixed(12407.0/65536.0,1,-nbitq), 
to_sfixed(17791.0/65536.0,1,-nbitq), 
to_sfixed(1371.0/65536.0,1,-nbitq), 
to_sfixed(-904.0/65536.0,1,-nbitq), 
to_sfixed(6335.0/65536.0,1,-nbitq), 
to_sfixed(-6526.0/65536.0,1,-nbitq), 
to_sfixed(-11902.0/65536.0,1,-nbitq), 
to_sfixed(958.0/65536.0,1,-nbitq), 
to_sfixed(-1400.0/65536.0,1,-nbitq), 
to_sfixed(-1641.0/65536.0,1,-nbitq), 
to_sfixed(-1898.0/65536.0,1,-nbitq), 
to_sfixed(-16454.0/65536.0,1,-nbitq), 
to_sfixed(653.0/65536.0,1,-nbitq), 
to_sfixed(4264.0/65536.0,1,-nbitq), 
to_sfixed(-1422.0/65536.0,1,-nbitq), 
to_sfixed(-6779.0/65536.0,1,-nbitq), 
to_sfixed(51.0/65536.0,1,-nbitq), 
to_sfixed(-202.0/65536.0,1,-nbitq), 
to_sfixed(1519.0/65536.0,1,-nbitq), 
to_sfixed(5577.0/65536.0,1,-nbitq), 
to_sfixed(-6641.0/65536.0,1,-nbitq), 
to_sfixed(11198.0/65536.0,1,-nbitq), 
to_sfixed(-3083.0/65536.0,1,-nbitq), 
to_sfixed(-1241.0/65536.0,1,-nbitq), 
to_sfixed(-1900.0/65536.0,1,-nbitq), 
to_sfixed(-2358.0/65536.0,1,-nbitq), 
to_sfixed(-445.0/65536.0,1,-nbitq), 
to_sfixed(8046.0/65536.0,1,-nbitq), 
to_sfixed(-1941.0/65536.0,1,-nbitq), 
to_sfixed(-951.0/65536.0,1,-nbitq), 
to_sfixed(-1124.0/65536.0,1,-nbitq), 
to_sfixed(1771.0/65536.0,1,-nbitq), 
to_sfixed(5516.0/65536.0,1,-nbitq), 
to_sfixed(-15290.0/65536.0,1,-nbitq), 
to_sfixed(1721.0/65536.0,1,-nbitq), 
to_sfixed(-520.0/65536.0,1,-nbitq), 
to_sfixed(-1972.0/65536.0,1,-nbitq), 
to_sfixed(-15068.0/65536.0,1,-nbitq), 
to_sfixed(-7584.0/65536.0,1,-nbitq), 
to_sfixed(-5995.0/65536.0,1,-nbitq), 
to_sfixed(989.0/65536.0,1,-nbitq), 
to_sfixed(-1343.0/65536.0,1,-nbitq), 
to_sfixed(1246.0/65536.0,1,-nbitq), 
to_sfixed(-16259.0/65536.0,1,-nbitq), 
to_sfixed(-645.0/65536.0,1,-nbitq), 
to_sfixed(8737.0/65536.0,1,-nbitq), 
to_sfixed(-719.0/65536.0,1,-nbitq), 
to_sfixed(-7079.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2920.0/65536.0,1,-nbitq), 
to_sfixed(1105.0/65536.0,1,-nbitq), 
to_sfixed(-8135.0/65536.0,1,-nbitq), 
to_sfixed(13268.0/65536.0,1,-nbitq), 
to_sfixed(5454.0/65536.0,1,-nbitq), 
to_sfixed(3192.0/65536.0,1,-nbitq), 
to_sfixed(2983.0/65536.0,1,-nbitq), 
to_sfixed(14164.0/65536.0,1,-nbitq), 
to_sfixed(454.0/65536.0,1,-nbitq), 
to_sfixed(1721.0/65536.0,1,-nbitq), 
to_sfixed(5996.0/65536.0,1,-nbitq), 
to_sfixed(11614.0/65536.0,1,-nbitq), 
to_sfixed(429.0/65536.0,1,-nbitq), 
to_sfixed(-4188.0/65536.0,1,-nbitq), 
to_sfixed(-8281.0/65536.0,1,-nbitq), 
to_sfixed(1603.0/65536.0,1,-nbitq), 
to_sfixed(-413.0/65536.0,1,-nbitq), 
to_sfixed(-10444.0/65536.0,1,-nbitq), 
to_sfixed(-7952.0/65536.0,1,-nbitq), 
to_sfixed(539.0/65536.0,1,-nbitq), 
to_sfixed(-6820.0/65536.0,1,-nbitq), 
to_sfixed(-10137.0/65536.0,1,-nbitq), 
to_sfixed(-11164.0/65536.0,1,-nbitq), 
to_sfixed(-8186.0/65536.0,1,-nbitq), 
to_sfixed(-870.0/65536.0,1,-nbitq), 
to_sfixed(251.0/65536.0,1,-nbitq), 
to_sfixed(4477.0/65536.0,1,-nbitq), 
to_sfixed(848.0/65536.0,1,-nbitq), 
to_sfixed(8795.0/65536.0,1,-nbitq), 
to_sfixed(4448.0/65536.0,1,-nbitq), 
to_sfixed(-4992.0/65536.0,1,-nbitq), 
to_sfixed(4767.0/65536.0,1,-nbitq), 
to_sfixed(10917.0/65536.0,1,-nbitq), 
to_sfixed(7438.0/65536.0,1,-nbitq), 
to_sfixed(2485.0/65536.0,1,-nbitq), 
to_sfixed(-1363.0/65536.0,1,-nbitq), 
to_sfixed(-336.0/65536.0,1,-nbitq), 
to_sfixed(99.0/65536.0,1,-nbitq), 
to_sfixed(-8784.0/65536.0,1,-nbitq), 
to_sfixed(465.0/65536.0,1,-nbitq), 
to_sfixed(-9271.0/65536.0,1,-nbitq), 
to_sfixed(-640.0/65536.0,1,-nbitq), 
to_sfixed(8788.0/65536.0,1,-nbitq), 
to_sfixed(-17712.0/65536.0,1,-nbitq), 
to_sfixed(-2113.0/65536.0,1,-nbitq), 
to_sfixed(15093.0/65536.0,1,-nbitq), 
to_sfixed(-3874.0/65536.0,1,-nbitq), 
to_sfixed(-2340.0/65536.0,1,-nbitq), 
to_sfixed(2314.0/65536.0,1,-nbitq), 
to_sfixed(-3032.0/65536.0,1,-nbitq), 
to_sfixed(-437.0/65536.0,1,-nbitq), 
to_sfixed(4008.0/65536.0,1,-nbitq), 
to_sfixed(-4088.0/65536.0,1,-nbitq), 
to_sfixed(13074.0/65536.0,1,-nbitq), 
to_sfixed(-1032.0/65536.0,1,-nbitq), 
to_sfixed(9052.0/65536.0,1,-nbitq), 
to_sfixed(-2425.0/65536.0,1,-nbitq), 
to_sfixed(-1375.0/65536.0,1,-nbitq), 
to_sfixed(2310.0/65536.0,1,-nbitq), 
to_sfixed(16300.0/65536.0,1,-nbitq), 
to_sfixed(-1427.0/65536.0,1,-nbitq), 
to_sfixed(-1097.0/65536.0,1,-nbitq), 
to_sfixed(1731.0/65536.0,1,-nbitq), 
to_sfixed(662.0/65536.0,1,-nbitq), 
to_sfixed(-3430.0/65536.0,1,-nbitq), 
to_sfixed(-18448.0/65536.0,1,-nbitq), 
to_sfixed(-775.0/65536.0,1,-nbitq), 
to_sfixed(-6547.0/65536.0,1,-nbitq), 
to_sfixed(-5890.0/65536.0,1,-nbitq), 
to_sfixed(-106.0/65536.0,1,-nbitq), 
to_sfixed(-5018.0/65536.0,1,-nbitq), 
to_sfixed(2390.0/65536.0,1,-nbitq), 
to_sfixed(-1690.0/65536.0,1,-nbitq), 
to_sfixed(2029.0/65536.0,1,-nbitq), 
to_sfixed(-606.0/65536.0,1,-nbitq), 
to_sfixed(-19688.0/65536.0,1,-nbitq), 
to_sfixed(-9462.0/65536.0,1,-nbitq), 
to_sfixed(3793.0/65536.0,1,-nbitq), 
to_sfixed(1163.0/65536.0,1,-nbitq), 
to_sfixed(-544.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-6012.0/65536.0,1,-nbitq), 
to_sfixed(-4569.0/65536.0,1,-nbitq), 
to_sfixed(-383.0/65536.0,1,-nbitq), 
to_sfixed(9256.0/65536.0,1,-nbitq), 
to_sfixed(12801.0/65536.0,1,-nbitq), 
to_sfixed(-11124.0/65536.0,1,-nbitq), 
to_sfixed(3283.0/65536.0,1,-nbitq), 
to_sfixed(12514.0/65536.0,1,-nbitq), 
to_sfixed(-1991.0/65536.0,1,-nbitq), 
to_sfixed(2087.0/65536.0,1,-nbitq), 
to_sfixed(3964.0/65536.0,1,-nbitq), 
to_sfixed(12642.0/65536.0,1,-nbitq), 
to_sfixed(3684.0/65536.0,1,-nbitq), 
to_sfixed(-1213.0/65536.0,1,-nbitq), 
to_sfixed(1543.0/65536.0,1,-nbitq), 
to_sfixed(1911.0/65536.0,1,-nbitq), 
to_sfixed(-658.0/65536.0,1,-nbitq), 
to_sfixed(1003.0/65536.0,1,-nbitq), 
to_sfixed(-6303.0/65536.0,1,-nbitq), 
to_sfixed(-1057.0/65536.0,1,-nbitq), 
to_sfixed(-454.0/65536.0,1,-nbitq), 
to_sfixed(-13243.0/65536.0,1,-nbitq), 
to_sfixed(-14139.0/65536.0,1,-nbitq), 
to_sfixed(4224.0/65536.0,1,-nbitq), 
to_sfixed(-2753.0/65536.0,1,-nbitq), 
to_sfixed(12651.0/65536.0,1,-nbitq), 
to_sfixed(3586.0/65536.0,1,-nbitq), 
to_sfixed(-2750.0/65536.0,1,-nbitq), 
to_sfixed(7167.0/65536.0,1,-nbitq), 
to_sfixed(3193.0/65536.0,1,-nbitq), 
to_sfixed(-4296.0/65536.0,1,-nbitq), 
to_sfixed(13471.0/65536.0,1,-nbitq), 
to_sfixed(-4805.0/65536.0,1,-nbitq), 
to_sfixed(-8512.0/65536.0,1,-nbitq), 
to_sfixed(1464.0/65536.0,1,-nbitq), 
to_sfixed(-658.0/65536.0,1,-nbitq), 
to_sfixed(-4873.0/65536.0,1,-nbitq), 
to_sfixed(-280.0/65536.0,1,-nbitq), 
to_sfixed(19085.0/65536.0,1,-nbitq), 
to_sfixed(849.0/65536.0,1,-nbitq), 
to_sfixed(-11515.0/65536.0,1,-nbitq), 
to_sfixed(2388.0/65536.0,1,-nbitq), 
to_sfixed(2270.0/65536.0,1,-nbitq), 
to_sfixed(-14446.0/65536.0,1,-nbitq), 
to_sfixed(1288.0/65536.0,1,-nbitq), 
to_sfixed(7108.0/65536.0,1,-nbitq), 
to_sfixed(-1482.0/65536.0,1,-nbitq), 
to_sfixed(-3173.0/65536.0,1,-nbitq), 
to_sfixed(3556.0/65536.0,1,-nbitq), 
to_sfixed(310.0/65536.0,1,-nbitq), 
to_sfixed(235.0/65536.0,1,-nbitq), 
to_sfixed(7386.0/65536.0,1,-nbitq), 
to_sfixed(3670.0/65536.0,1,-nbitq), 
to_sfixed(6133.0/65536.0,1,-nbitq), 
to_sfixed(-353.0/65536.0,1,-nbitq), 
to_sfixed(4017.0/65536.0,1,-nbitq), 
to_sfixed(2270.0/65536.0,1,-nbitq), 
to_sfixed(3580.0/65536.0,1,-nbitq), 
to_sfixed(1480.0/65536.0,1,-nbitq), 
to_sfixed(11638.0/65536.0,1,-nbitq), 
to_sfixed(-5342.0/65536.0,1,-nbitq), 
to_sfixed(-829.0/65536.0,1,-nbitq), 
to_sfixed(1451.0/65536.0,1,-nbitq), 
to_sfixed(525.0/65536.0,1,-nbitq), 
to_sfixed(1223.0/65536.0,1,-nbitq), 
to_sfixed(-8441.0/65536.0,1,-nbitq), 
to_sfixed(-8376.0/65536.0,1,-nbitq), 
to_sfixed(-3048.0/65536.0,1,-nbitq), 
to_sfixed(-9423.0/65536.0,1,-nbitq), 
to_sfixed(-8816.0/65536.0,1,-nbitq), 
to_sfixed(-4491.0/65536.0,1,-nbitq), 
to_sfixed(18489.0/65536.0,1,-nbitq), 
to_sfixed(-11504.0/65536.0,1,-nbitq), 
to_sfixed(2211.0/65536.0,1,-nbitq), 
to_sfixed(826.0/65536.0,1,-nbitq), 
to_sfixed(-18777.0/65536.0,1,-nbitq), 
to_sfixed(-956.0/65536.0,1,-nbitq), 
to_sfixed(2550.0/65536.0,1,-nbitq), 
to_sfixed(2481.0/65536.0,1,-nbitq), 
to_sfixed(4269.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-7945.0/65536.0,1,-nbitq), 
to_sfixed(-4993.0/65536.0,1,-nbitq), 
to_sfixed(4795.0/65536.0,1,-nbitq), 
to_sfixed(8182.0/65536.0,1,-nbitq), 
to_sfixed(1450.0/65536.0,1,-nbitq), 
to_sfixed(2264.0/65536.0,1,-nbitq), 
to_sfixed(3675.0/65536.0,1,-nbitq), 
to_sfixed(16491.0/65536.0,1,-nbitq), 
to_sfixed(-7014.0/65536.0,1,-nbitq), 
to_sfixed(2331.0/65536.0,1,-nbitq), 
to_sfixed(4817.0/65536.0,1,-nbitq), 
to_sfixed(34139.0/65536.0,1,-nbitq), 
to_sfixed(3586.0/65536.0,1,-nbitq), 
to_sfixed(2239.0/65536.0,1,-nbitq), 
to_sfixed(-1300.0/65536.0,1,-nbitq), 
to_sfixed(-2642.0/65536.0,1,-nbitq), 
to_sfixed(-1091.0/65536.0,1,-nbitq), 
to_sfixed(-81.0/65536.0,1,-nbitq), 
to_sfixed(-2228.0/65536.0,1,-nbitq), 
to_sfixed(-485.0/65536.0,1,-nbitq), 
to_sfixed(2068.0/65536.0,1,-nbitq), 
to_sfixed(-1294.0/65536.0,1,-nbitq), 
to_sfixed(-20253.0/65536.0,1,-nbitq), 
to_sfixed(404.0/65536.0,1,-nbitq), 
to_sfixed(1525.0/65536.0,1,-nbitq), 
to_sfixed(584.0/65536.0,1,-nbitq), 
to_sfixed(-3899.0/65536.0,1,-nbitq), 
to_sfixed(509.0/65536.0,1,-nbitq), 
to_sfixed(15969.0/65536.0,1,-nbitq), 
to_sfixed(3699.0/65536.0,1,-nbitq), 
to_sfixed(-1033.0/65536.0,1,-nbitq), 
to_sfixed(9864.0/65536.0,1,-nbitq), 
to_sfixed(-7094.0/65536.0,1,-nbitq), 
to_sfixed(-10536.0/65536.0,1,-nbitq), 
to_sfixed(-2085.0/65536.0,1,-nbitq), 
to_sfixed(-602.0/65536.0,1,-nbitq), 
to_sfixed(-416.0/65536.0,1,-nbitq), 
to_sfixed(10287.0/65536.0,1,-nbitq), 
to_sfixed(-791.0/65536.0,1,-nbitq), 
to_sfixed(940.0/65536.0,1,-nbitq), 
to_sfixed(-12772.0/65536.0,1,-nbitq), 
to_sfixed(-502.0/65536.0,1,-nbitq), 
to_sfixed(-3427.0/65536.0,1,-nbitq), 
to_sfixed(-12115.0/65536.0,1,-nbitq), 
to_sfixed(1070.0/65536.0,1,-nbitq), 
to_sfixed(12028.0/65536.0,1,-nbitq), 
to_sfixed(1643.0/65536.0,1,-nbitq), 
to_sfixed(-2170.0/65536.0,1,-nbitq), 
to_sfixed(1248.0/65536.0,1,-nbitq), 
to_sfixed(-1972.0/65536.0,1,-nbitq), 
to_sfixed(-1044.0/65536.0,1,-nbitq), 
to_sfixed(-4162.0/65536.0,1,-nbitq), 
to_sfixed(6745.0/65536.0,1,-nbitq), 
to_sfixed(5436.0/65536.0,1,-nbitq), 
to_sfixed(7249.0/65536.0,1,-nbitq), 
to_sfixed(-19534.0/65536.0,1,-nbitq), 
to_sfixed(-1731.0/65536.0,1,-nbitq), 
to_sfixed(4096.0/65536.0,1,-nbitq), 
to_sfixed(2946.0/65536.0,1,-nbitq), 
to_sfixed(6399.0/65536.0,1,-nbitq), 
to_sfixed(-7511.0/65536.0,1,-nbitq), 
to_sfixed(1550.0/65536.0,1,-nbitq), 
to_sfixed(728.0/65536.0,1,-nbitq), 
to_sfixed(1346.0/65536.0,1,-nbitq), 
to_sfixed(-5689.0/65536.0,1,-nbitq), 
to_sfixed(-3870.0/65536.0,1,-nbitq), 
to_sfixed(-3292.0/65536.0,1,-nbitq), 
to_sfixed(-8336.0/65536.0,1,-nbitq), 
to_sfixed(-6970.0/65536.0,1,-nbitq), 
to_sfixed(15856.0/65536.0,1,-nbitq), 
to_sfixed(-1819.0/65536.0,1,-nbitq), 
to_sfixed(5790.0/65536.0,1,-nbitq), 
to_sfixed(-12423.0/65536.0,1,-nbitq), 
to_sfixed(65.0/65536.0,1,-nbitq), 
to_sfixed(959.0/65536.0,1,-nbitq), 
to_sfixed(6769.0/65536.0,1,-nbitq), 
to_sfixed(1380.0/65536.0,1,-nbitq), 
to_sfixed(30.0/65536.0,1,-nbitq), 
to_sfixed(-1669.0/65536.0,1,-nbitq), 
to_sfixed(11605.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4721.0/65536.0,1,-nbitq), 
to_sfixed(-4570.0/65536.0,1,-nbitq), 
to_sfixed(465.0/65536.0,1,-nbitq), 
to_sfixed(9428.0/65536.0,1,-nbitq), 
to_sfixed(-2909.0/65536.0,1,-nbitq), 
to_sfixed(16965.0/65536.0,1,-nbitq), 
to_sfixed(2738.0/65536.0,1,-nbitq), 
to_sfixed(7947.0/65536.0,1,-nbitq), 
to_sfixed(-2823.0/65536.0,1,-nbitq), 
to_sfixed(-625.0/65536.0,1,-nbitq), 
to_sfixed(503.0/65536.0,1,-nbitq), 
to_sfixed(8486.0/65536.0,1,-nbitq), 
to_sfixed(2130.0/65536.0,1,-nbitq), 
to_sfixed(8794.0/65536.0,1,-nbitq), 
to_sfixed(-553.0/65536.0,1,-nbitq), 
to_sfixed(2194.0/65536.0,1,-nbitq), 
to_sfixed(1913.0/65536.0,1,-nbitq), 
to_sfixed(5159.0/65536.0,1,-nbitq), 
to_sfixed(-3401.0/65536.0,1,-nbitq), 
to_sfixed(704.0/65536.0,1,-nbitq), 
to_sfixed(-1760.0/65536.0,1,-nbitq), 
to_sfixed(-6282.0/65536.0,1,-nbitq), 
to_sfixed(-27395.0/65536.0,1,-nbitq), 
to_sfixed(-5475.0/65536.0,1,-nbitq), 
to_sfixed(3191.0/65536.0,1,-nbitq), 
to_sfixed(1172.0/65536.0,1,-nbitq), 
to_sfixed(-2650.0/65536.0,1,-nbitq), 
to_sfixed(2661.0/65536.0,1,-nbitq), 
to_sfixed(9364.0/65536.0,1,-nbitq), 
to_sfixed(-99.0/65536.0,1,-nbitq), 
to_sfixed(2340.0/65536.0,1,-nbitq), 
to_sfixed(-1934.0/65536.0,1,-nbitq), 
to_sfixed(-10606.0/65536.0,1,-nbitq), 
to_sfixed(-5197.0/65536.0,1,-nbitq), 
to_sfixed(-2501.0/65536.0,1,-nbitq), 
to_sfixed(1939.0/65536.0,1,-nbitq), 
to_sfixed(-4155.0/65536.0,1,-nbitq), 
to_sfixed(7990.0/65536.0,1,-nbitq), 
to_sfixed(-14592.0/65536.0,1,-nbitq), 
to_sfixed(86.0/65536.0,1,-nbitq), 
to_sfixed(828.0/65536.0,1,-nbitq), 
to_sfixed(483.0/65536.0,1,-nbitq), 
to_sfixed(-4836.0/65536.0,1,-nbitq), 
to_sfixed(-5038.0/65536.0,1,-nbitq), 
to_sfixed(-2450.0/65536.0,1,-nbitq), 
to_sfixed(-1566.0/65536.0,1,-nbitq), 
to_sfixed(-2493.0/65536.0,1,-nbitq), 
to_sfixed(1462.0/65536.0,1,-nbitq), 
to_sfixed(1833.0/65536.0,1,-nbitq), 
to_sfixed(1499.0/65536.0,1,-nbitq), 
to_sfixed(1990.0/65536.0,1,-nbitq), 
to_sfixed(-3866.0/65536.0,1,-nbitq), 
to_sfixed(7074.0/65536.0,1,-nbitq), 
to_sfixed(-6328.0/65536.0,1,-nbitq), 
to_sfixed(9531.0/65536.0,1,-nbitq), 
to_sfixed(-20950.0/65536.0,1,-nbitq), 
to_sfixed(-2171.0/65536.0,1,-nbitq), 
to_sfixed(-1968.0/65536.0,1,-nbitq), 
to_sfixed(2806.0/65536.0,1,-nbitq), 
to_sfixed(5738.0/65536.0,1,-nbitq), 
to_sfixed(-6474.0/65536.0,1,-nbitq), 
to_sfixed(-1927.0/65536.0,1,-nbitq), 
to_sfixed(863.0/65536.0,1,-nbitq), 
to_sfixed(-31.0/65536.0,1,-nbitq), 
to_sfixed(-3628.0/65536.0,1,-nbitq), 
to_sfixed(-3230.0/65536.0,1,-nbitq), 
to_sfixed(5082.0/65536.0,1,-nbitq), 
to_sfixed(230.0/65536.0,1,-nbitq), 
to_sfixed(-5999.0/65536.0,1,-nbitq), 
to_sfixed(16317.0/65536.0,1,-nbitq), 
to_sfixed(2881.0/65536.0,1,-nbitq), 
to_sfixed(3183.0/65536.0,1,-nbitq), 
to_sfixed(7240.0/65536.0,1,-nbitq), 
to_sfixed(2623.0/65536.0,1,-nbitq), 
to_sfixed(-2766.0/65536.0,1,-nbitq), 
to_sfixed(13237.0/65536.0,1,-nbitq), 
to_sfixed(-3551.0/65536.0,1,-nbitq), 
to_sfixed(353.0/65536.0,1,-nbitq), 
to_sfixed(-110.0/65536.0,1,-nbitq), 
to_sfixed(15662.0/65536.0,1,-nbitq)  ), 
( to_sfixed(958.0/65536.0,1,-nbitq), 
to_sfixed(-2065.0/65536.0,1,-nbitq), 
to_sfixed(6032.0/65536.0,1,-nbitq), 
to_sfixed(2934.0/65536.0,1,-nbitq), 
to_sfixed(3919.0/65536.0,1,-nbitq), 
to_sfixed(14568.0/65536.0,1,-nbitq), 
to_sfixed(4527.0/65536.0,1,-nbitq), 
to_sfixed(-5512.0/65536.0,1,-nbitq), 
to_sfixed(606.0/65536.0,1,-nbitq), 
to_sfixed(-2616.0/65536.0,1,-nbitq), 
to_sfixed(-977.0/65536.0,1,-nbitq), 
to_sfixed(7063.0/65536.0,1,-nbitq), 
to_sfixed(-228.0/65536.0,1,-nbitq), 
to_sfixed(2968.0/65536.0,1,-nbitq), 
to_sfixed(-3161.0/65536.0,1,-nbitq), 
to_sfixed(1971.0/65536.0,1,-nbitq), 
to_sfixed(1284.0/65536.0,1,-nbitq), 
to_sfixed(1416.0/65536.0,1,-nbitq), 
to_sfixed(-19.0/65536.0,1,-nbitq), 
to_sfixed(-204.0/65536.0,1,-nbitq), 
to_sfixed(-5072.0/65536.0,1,-nbitq), 
to_sfixed(790.0/65536.0,1,-nbitq), 
to_sfixed(-16434.0/65536.0,1,-nbitq), 
to_sfixed(934.0/65536.0,1,-nbitq), 
to_sfixed(5990.0/65536.0,1,-nbitq), 
to_sfixed(-3376.0/65536.0,1,-nbitq), 
to_sfixed(261.0/65536.0,1,-nbitq), 
to_sfixed(1569.0/65536.0,1,-nbitq), 
to_sfixed(4324.0/65536.0,1,-nbitq), 
to_sfixed(-370.0/65536.0,1,-nbitq), 
to_sfixed(1997.0/65536.0,1,-nbitq), 
to_sfixed(-3918.0/65536.0,1,-nbitq), 
to_sfixed(-7488.0/65536.0,1,-nbitq), 
to_sfixed(-5317.0/65536.0,1,-nbitq), 
to_sfixed(1101.0/65536.0,1,-nbitq), 
to_sfixed(-1386.0/65536.0,1,-nbitq), 
to_sfixed(3251.0/65536.0,1,-nbitq), 
to_sfixed(414.0/65536.0,1,-nbitq), 
to_sfixed(-10791.0/65536.0,1,-nbitq), 
to_sfixed(4185.0/65536.0,1,-nbitq), 
to_sfixed(6626.0/65536.0,1,-nbitq), 
to_sfixed(-2076.0/65536.0,1,-nbitq), 
to_sfixed(1859.0/65536.0,1,-nbitq), 
to_sfixed(-127.0/65536.0,1,-nbitq), 
to_sfixed(1547.0/65536.0,1,-nbitq), 
to_sfixed(-10404.0/65536.0,1,-nbitq), 
to_sfixed(332.0/65536.0,1,-nbitq), 
to_sfixed(1885.0/65536.0,1,-nbitq), 
to_sfixed(-430.0/65536.0,1,-nbitq), 
to_sfixed(2793.0/65536.0,1,-nbitq), 
to_sfixed(-1654.0/65536.0,1,-nbitq), 
to_sfixed(-10471.0/65536.0,1,-nbitq), 
to_sfixed(3798.0/65536.0,1,-nbitq), 
to_sfixed(-3055.0/65536.0,1,-nbitq), 
to_sfixed(4392.0/65536.0,1,-nbitq), 
to_sfixed(-14987.0/65536.0,1,-nbitq), 
to_sfixed(-3289.0/65536.0,1,-nbitq), 
to_sfixed(-3954.0/65536.0,1,-nbitq), 
to_sfixed(-853.0/65536.0,1,-nbitq), 
to_sfixed(4223.0/65536.0,1,-nbitq), 
to_sfixed(-254.0/65536.0,1,-nbitq), 
to_sfixed(632.0/65536.0,1,-nbitq), 
to_sfixed(2195.0/65536.0,1,-nbitq), 
to_sfixed(-864.0/65536.0,1,-nbitq), 
to_sfixed(2266.0/65536.0,1,-nbitq), 
to_sfixed(102.0/65536.0,1,-nbitq), 
to_sfixed(-1362.0/65536.0,1,-nbitq), 
to_sfixed(-4780.0/65536.0,1,-nbitq), 
to_sfixed(-5269.0/65536.0,1,-nbitq), 
to_sfixed(11282.0/65536.0,1,-nbitq), 
to_sfixed(3043.0/65536.0,1,-nbitq), 
to_sfixed(8669.0/65536.0,1,-nbitq), 
to_sfixed(17987.0/65536.0,1,-nbitq), 
to_sfixed(-1182.0/65536.0,1,-nbitq), 
to_sfixed(702.0/65536.0,1,-nbitq), 
to_sfixed(6607.0/65536.0,1,-nbitq), 
to_sfixed(-16351.0/65536.0,1,-nbitq), 
to_sfixed(-11442.0/65536.0,1,-nbitq), 
to_sfixed(-8.0/65536.0,1,-nbitq), 
to_sfixed(14244.0/65536.0,1,-nbitq)  ), 
( to_sfixed(6764.0/65536.0,1,-nbitq), 
to_sfixed(1102.0/65536.0,1,-nbitq), 
to_sfixed(1587.0/65536.0,1,-nbitq), 
to_sfixed(4981.0/65536.0,1,-nbitq), 
to_sfixed(-203.0/65536.0,1,-nbitq), 
to_sfixed(14485.0/65536.0,1,-nbitq), 
to_sfixed(3540.0/65536.0,1,-nbitq), 
to_sfixed(-3019.0/65536.0,1,-nbitq), 
to_sfixed(2389.0/65536.0,1,-nbitq), 
to_sfixed(-960.0/65536.0,1,-nbitq), 
to_sfixed(-3395.0/65536.0,1,-nbitq), 
to_sfixed(421.0/65536.0,1,-nbitq), 
to_sfixed(-381.0/65536.0,1,-nbitq), 
to_sfixed(1603.0/65536.0,1,-nbitq), 
to_sfixed(748.0/65536.0,1,-nbitq), 
to_sfixed(1980.0/65536.0,1,-nbitq), 
to_sfixed(988.0/65536.0,1,-nbitq), 
to_sfixed(2467.0/65536.0,1,-nbitq), 
to_sfixed(-424.0/65536.0,1,-nbitq), 
to_sfixed(-2274.0/65536.0,1,-nbitq), 
to_sfixed(-2357.0/65536.0,1,-nbitq), 
to_sfixed(-1894.0/65536.0,1,-nbitq), 
to_sfixed(-14196.0/65536.0,1,-nbitq), 
to_sfixed(-1855.0/65536.0,1,-nbitq), 
to_sfixed(1208.0/65536.0,1,-nbitq), 
to_sfixed(-1338.0/65536.0,1,-nbitq), 
to_sfixed(-1666.0/65536.0,1,-nbitq), 
to_sfixed(-766.0/65536.0,1,-nbitq), 
to_sfixed(4826.0/65536.0,1,-nbitq), 
to_sfixed(3685.0/65536.0,1,-nbitq), 
to_sfixed(-1799.0/65536.0,1,-nbitq), 
to_sfixed(-4260.0/65536.0,1,-nbitq), 
to_sfixed(-12791.0/65536.0,1,-nbitq), 
to_sfixed(-7604.0/65536.0,1,-nbitq), 
to_sfixed(2168.0/65536.0,1,-nbitq), 
to_sfixed(2179.0/65536.0,1,-nbitq), 
to_sfixed(-720.0/65536.0,1,-nbitq), 
to_sfixed(-1366.0/65536.0,1,-nbitq), 
to_sfixed(-14550.0/65536.0,1,-nbitq), 
to_sfixed(-945.0/65536.0,1,-nbitq), 
to_sfixed(16669.0/65536.0,1,-nbitq), 
to_sfixed(-734.0/65536.0,1,-nbitq), 
to_sfixed(3099.0/65536.0,1,-nbitq), 
to_sfixed(2003.0/65536.0,1,-nbitq), 
to_sfixed(-1271.0/65536.0,1,-nbitq), 
to_sfixed(-18274.0/65536.0,1,-nbitq), 
to_sfixed(-2528.0/65536.0,1,-nbitq), 
to_sfixed(7062.0/65536.0,1,-nbitq), 
to_sfixed(2777.0/65536.0,1,-nbitq), 
to_sfixed(-1699.0/65536.0,1,-nbitq), 
to_sfixed(-1962.0/65536.0,1,-nbitq), 
to_sfixed(-66.0/65536.0,1,-nbitq), 
to_sfixed(15556.0/65536.0,1,-nbitq), 
to_sfixed(5251.0/65536.0,1,-nbitq), 
to_sfixed(6095.0/65536.0,1,-nbitq), 
to_sfixed(-4046.0/65536.0,1,-nbitq), 
to_sfixed(424.0/65536.0,1,-nbitq), 
to_sfixed(-3476.0/65536.0,1,-nbitq), 
to_sfixed(817.0/65536.0,1,-nbitq), 
to_sfixed(332.0/65536.0,1,-nbitq), 
to_sfixed(-1901.0/65536.0,1,-nbitq), 
to_sfixed(875.0/65536.0,1,-nbitq), 
to_sfixed(2291.0/65536.0,1,-nbitq), 
to_sfixed(1271.0/65536.0,1,-nbitq), 
to_sfixed(1488.0/65536.0,1,-nbitq), 
to_sfixed(-478.0/65536.0,1,-nbitq), 
to_sfixed(-5724.0/65536.0,1,-nbitq), 
to_sfixed(-4085.0/65536.0,1,-nbitq), 
to_sfixed(1005.0/65536.0,1,-nbitq), 
to_sfixed(4001.0/65536.0,1,-nbitq), 
to_sfixed(4650.0/65536.0,1,-nbitq), 
to_sfixed(1960.0/65536.0,1,-nbitq), 
to_sfixed(10186.0/65536.0,1,-nbitq), 
to_sfixed(-2951.0/65536.0,1,-nbitq), 
to_sfixed(-680.0/65536.0,1,-nbitq), 
to_sfixed(1622.0/65536.0,1,-nbitq), 
to_sfixed(-7155.0/65536.0,1,-nbitq), 
to_sfixed(-16090.0/65536.0,1,-nbitq), 
to_sfixed(1486.0/65536.0,1,-nbitq), 
to_sfixed(4207.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-395.0/65536.0,1,-nbitq), 
to_sfixed(-1518.0/65536.0,1,-nbitq), 
to_sfixed(-460.0/65536.0,1,-nbitq), 
to_sfixed(4157.0/65536.0,1,-nbitq), 
to_sfixed(-4906.0/65536.0,1,-nbitq), 
to_sfixed(10219.0/65536.0,1,-nbitq), 
to_sfixed(-1937.0/65536.0,1,-nbitq), 
to_sfixed(-1394.0/65536.0,1,-nbitq), 
to_sfixed(6672.0/65536.0,1,-nbitq), 
to_sfixed(-663.0/65536.0,1,-nbitq), 
to_sfixed(694.0/65536.0,1,-nbitq), 
to_sfixed(2490.0/65536.0,1,-nbitq), 
to_sfixed(-140.0/65536.0,1,-nbitq), 
to_sfixed(-1434.0/65536.0,1,-nbitq), 
to_sfixed(-1565.0/65536.0,1,-nbitq), 
to_sfixed(1293.0/65536.0,1,-nbitq), 
to_sfixed(476.0/65536.0,1,-nbitq), 
to_sfixed(-2054.0/65536.0,1,-nbitq), 
to_sfixed(-3903.0/65536.0,1,-nbitq), 
to_sfixed(783.0/65536.0,1,-nbitq), 
to_sfixed(-2928.0/65536.0,1,-nbitq), 
to_sfixed(8571.0/65536.0,1,-nbitq), 
to_sfixed(-7140.0/65536.0,1,-nbitq), 
to_sfixed(-5311.0/65536.0,1,-nbitq), 
to_sfixed(4585.0/65536.0,1,-nbitq), 
to_sfixed(4418.0/65536.0,1,-nbitq), 
to_sfixed(-2958.0/65536.0,1,-nbitq), 
to_sfixed(-1736.0/65536.0,1,-nbitq), 
to_sfixed(8663.0/65536.0,1,-nbitq), 
to_sfixed(-710.0/65536.0,1,-nbitq), 
to_sfixed(1653.0/65536.0,1,-nbitq), 
to_sfixed(-5843.0/65536.0,1,-nbitq), 
to_sfixed(-7650.0/65536.0,1,-nbitq), 
to_sfixed(-1540.0/65536.0,1,-nbitq), 
to_sfixed(830.0/65536.0,1,-nbitq), 
to_sfixed(-1529.0/65536.0,1,-nbitq), 
to_sfixed(-2924.0/65536.0,1,-nbitq), 
to_sfixed(-3025.0/65536.0,1,-nbitq), 
to_sfixed(-4735.0/65536.0,1,-nbitq), 
to_sfixed(-2377.0/65536.0,1,-nbitq), 
to_sfixed(16069.0/65536.0,1,-nbitq), 
to_sfixed(-101.0/65536.0,1,-nbitq), 
to_sfixed(-1367.0/65536.0,1,-nbitq), 
to_sfixed(-4904.0/65536.0,1,-nbitq), 
to_sfixed(1009.0/65536.0,1,-nbitq), 
to_sfixed(-868.0/65536.0,1,-nbitq), 
to_sfixed(-630.0/65536.0,1,-nbitq), 
to_sfixed(8551.0/65536.0,1,-nbitq), 
to_sfixed(1016.0/65536.0,1,-nbitq), 
to_sfixed(1053.0/65536.0,1,-nbitq), 
to_sfixed(-836.0/65536.0,1,-nbitq), 
to_sfixed(-3639.0/65536.0,1,-nbitq), 
to_sfixed(18171.0/65536.0,1,-nbitq), 
to_sfixed(14396.0/65536.0,1,-nbitq), 
to_sfixed(6479.0/65536.0,1,-nbitq), 
to_sfixed(-9582.0/65536.0,1,-nbitq), 
to_sfixed(-2073.0/65536.0,1,-nbitq), 
to_sfixed(-4487.0/65536.0,1,-nbitq), 
to_sfixed(-1371.0/65536.0,1,-nbitq), 
to_sfixed(856.0/65536.0,1,-nbitq), 
to_sfixed(1908.0/65536.0,1,-nbitq), 
to_sfixed(-1999.0/65536.0,1,-nbitq), 
to_sfixed(1260.0/65536.0,1,-nbitq), 
to_sfixed(920.0/65536.0,1,-nbitq), 
to_sfixed(5895.0/65536.0,1,-nbitq), 
to_sfixed(-6116.0/65536.0,1,-nbitq), 
to_sfixed(-2097.0/65536.0,1,-nbitq), 
to_sfixed(-641.0/65536.0,1,-nbitq), 
to_sfixed(3182.0/65536.0,1,-nbitq), 
to_sfixed(530.0/65536.0,1,-nbitq), 
to_sfixed(4440.0/65536.0,1,-nbitq), 
to_sfixed(4338.0/65536.0,1,-nbitq), 
to_sfixed(7935.0/65536.0,1,-nbitq), 
to_sfixed(18.0/65536.0,1,-nbitq), 
to_sfixed(1758.0/65536.0,1,-nbitq), 
to_sfixed(-824.0/65536.0,1,-nbitq), 
to_sfixed(-7911.0/65536.0,1,-nbitq), 
to_sfixed(-11206.0/65536.0,1,-nbitq), 
to_sfixed(-581.0/65536.0,1,-nbitq), 
to_sfixed(-1884.0/65536.0,1,-nbitq)  ), 
( to_sfixed(493.0/65536.0,1,-nbitq), 
to_sfixed(3903.0/65536.0,1,-nbitq), 
to_sfixed(-4628.0/65536.0,1,-nbitq), 
to_sfixed(2037.0/65536.0,1,-nbitq), 
to_sfixed(10171.0/65536.0,1,-nbitq), 
to_sfixed(10701.0/65536.0,1,-nbitq), 
to_sfixed(910.0/65536.0,1,-nbitq), 
to_sfixed(761.0/65536.0,1,-nbitq), 
to_sfixed(4789.0/65536.0,1,-nbitq), 
to_sfixed(-143.0/65536.0,1,-nbitq), 
to_sfixed(3345.0/65536.0,1,-nbitq), 
to_sfixed(-4914.0/65536.0,1,-nbitq), 
to_sfixed(-112.0/65536.0,1,-nbitq), 
to_sfixed(4593.0/65536.0,1,-nbitq), 
to_sfixed(-4308.0/65536.0,1,-nbitq), 
to_sfixed(1324.0/65536.0,1,-nbitq), 
to_sfixed(835.0/65536.0,1,-nbitq), 
to_sfixed(2552.0/65536.0,1,-nbitq), 
to_sfixed(1264.0/65536.0,1,-nbitq), 
to_sfixed(630.0/65536.0,1,-nbitq), 
to_sfixed(2083.0/65536.0,1,-nbitq), 
to_sfixed(6037.0/65536.0,1,-nbitq), 
to_sfixed(-6613.0/65536.0,1,-nbitq), 
to_sfixed(-7188.0/65536.0,1,-nbitq), 
to_sfixed(6022.0/65536.0,1,-nbitq), 
to_sfixed(7869.0/65536.0,1,-nbitq), 
to_sfixed(-9037.0/65536.0,1,-nbitq), 
to_sfixed(1591.0/65536.0,1,-nbitq), 
to_sfixed(11139.0/65536.0,1,-nbitq), 
to_sfixed(-2906.0/65536.0,1,-nbitq), 
to_sfixed(1045.0/65536.0,1,-nbitq), 
to_sfixed(-10142.0/65536.0,1,-nbitq), 
to_sfixed(-1145.0/65536.0,1,-nbitq), 
to_sfixed(12097.0/65536.0,1,-nbitq), 
to_sfixed(-2623.0/65536.0,1,-nbitq), 
to_sfixed(-3522.0/65536.0,1,-nbitq), 
to_sfixed(-5347.0/65536.0,1,-nbitq), 
to_sfixed(-5009.0/65536.0,1,-nbitq), 
to_sfixed(-7518.0/65536.0,1,-nbitq), 
to_sfixed(2553.0/65536.0,1,-nbitq), 
to_sfixed(9201.0/65536.0,1,-nbitq), 
to_sfixed(-1566.0/65536.0,1,-nbitq), 
to_sfixed(1116.0/65536.0,1,-nbitq), 
to_sfixed(6884.0/65536.0,1,-nbitq), 
to_sfixed(-1849.0/65536.0,1,-nbitq), 
to_sfixed(3003.0/65536.0,1,-nbitq), 
to_sfixed(-3369.0/65536.0,1,-nbitq), 
to_sfixed(5527.0/65536.0,1,-nbitq), 
to_sfixed(-745.0/65536.0,1,-nbitq), 
to_sfixed(-464.0/65536.0,1,-nbitq), 
to_sfixed(3120.0/65536.0,1,-nbitq), 
to_sfixed(476.0/65536.0,1,-nbitq), 
to_sfixed(13271.0/65536.0,1,-nbitq), 
to_sfixed(12684.0/65536.0,1,-nbitq), 
to_sfixed(5449.0/65536.0,1,-nbitq), 
to_sfixed(-6817.0/65536.0,1,-nbitq), 
to_sfixed(2118.0/65536.0,1,-nbitq), 
to_sfixed(-4487.0/65536.0,1,-nbitq), 
to_sfixed(1319.0/65536.0,1,-nbitq), 
to_sfixed(5405.0/65536.0,1,-nbitq), 
to_sfixed(1542.0/65536.0,1,-nbitq), 
to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(3024.0/65536.0,1,-nbitq), 
to_sfixed(-80.0/65536.0,1,-nbitq), 
to_sfixed(7281.0/65536.0,1,-nbitq), 
to_sfixed(-7590.0/65536.0,1,-nbitq), 
to_sfixed(-2912.0/65536.0,1,-nbitq), 
to_sfixed(1687.0/65536.0,1,-nbitq), 
to_sfixed(3839.0/65536.0,1,-nbitq), 
to_sfixed(1838.0/65536.0,1,-nbitq), 
to_sfixed(163.0/65536.0,1,-nbitq), 
to_sfixed(-3225.0/65536.0,1,-nbitq), 
to_sfixed(11632.0/65536.0,1,-nbitq), 
to_sfixed(-1959.0/65536.0,1,-nbitq), 
to_sfixed(1808.0/65536.0,1,-nbitq), 
to_sfixed(-2307.0/65536.0,1,-nbitq), 
to_sfixed(-8114.0/65536.0,1,-nbitq), 
to_sfixed(-8298.0/65536.0,1,-nbitq), 
to_sfixed(-523.0/65536.0,1,-nbitq), 
to_sfixed(-6811.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1055.0/65536.0,1,-nbitq), 
to_sfixed(591.0/65536.0,1,-nbitq), 
to_sfixed(-7956.0/65536.0,1,-nbitq), 
to_sfixed(2932.0/65536.0,1,-nbitq), 
to_sfixed(7221.0/65536.0,1,-nbitq), 
to_sfixed(6300.0/65536.0,1,-nbitq), 
to_sfixed(-740.0/65536.0,1,-nbitq), 
to_sfixed(1837.0/65536.0,1,-nbitq), 
to_sfixed(-3627.0/65536.0,1,-nbitq), 
to_sfixed(-765.0/65536.0,1,-nbitq), 
to_sfixed(5054.0/65536.0,1,-nbitq), 
to_sfixed(-6615.0/65536.0,1,-nbitq), 
to_sfixed(357.0/65536.0,1,-nbitq), 
to_sfixed(5888.0/65536.0,1,-nbitq), 
to_sfixed(-1600.0/65536.0,1,-nbitq), 
to_sfixed(-451.0/65536.0,1,-nbitq), 
to_sfixed(-2274.0/65536.0,1,-nbitq), 
to_sfixed(229.0/65536.0,1,-nbitq), 
to_sfixed(1487.0/65536.0,1,-nbitq), 
to_sfixed(2197.0/65536.0,1,-nbitq), 
to_sfixed(2555.0/65536.0,1,-nbitq), 
to_sfixed(-383.0/65536.0,1,-nbitq), 
to_sfixed(-453.0/65536.0,1,-nbitq), 
to_sfixed(-4556.0/65536.0,1,-nbitq), 
to_sfixed(1841.0/65536.0,1,-nbitq), 
to_sfixed(4943.0/65536.0,1,-nbitq), 
to_sfixed(-5410.0/65536.0,1,-nbitq), 
to_sfixed(2441.0/65536.0,1,-nbitq), 
to_sfixed(5727.0/65536.0,1,-nbitq), 
to_sfixed(-5468.0/65536.0,1,-nbitq), 
to_sfixed(1654.0/65536.0,1,-nbitq), 
to_sfixed(-8085.0/65536.0,1,-nbitq), 
to_sfixed(7137.0/65536.0,1,-nbitq), 
to_sfixed(16491.0/65536.0,1,-nbitq), 
to_sfixed(-498.0/65536.0,1,-nbitq), 
to_sfixed(-250.0/65536.0,1,-nbitq), 
to_sfixed(-7846.0/65536.0,1,-nbitq), 
to_sfixed(72.0/65536.0,1,-nbitq), 
to_sfixed(-1190.0/65536.0,1,-nbitq), 
to_sfixed(2253.0/65536.0,1,-nbitq), 
to_sfixed(7436.0/65536.0,1,-nbitq), 
to_sfixed(-2397.0/65536.0,1,-nbitq), 
to_sfixed(8859.0/65536.0,1,-nbitq), 
to_sfixed(5249.0/65536.0,1,-nbitq), 
to_sfixed(2356.0/65536.0,1,-nbitq), 
to_sfixed(7150.0/65536.0,1,-nbitq), 
to_sfixed(-2822.0/65536.0,1,-nbitq), 
to_sfixed(2633.0/65536.0,1,-nbitq), 
to_sfixed(-220.0/65536.0,1,-nbitq), 
to_sfixed(-1867.0/65536.0,1,-nbitq), 
to_sfixed(1077.0/65536.0,1,-nbitq), 
to_sfixed(2412.0/65536.0,1,-nbitq), 
to_sfixed(8033.0/65536.0,1,-nbitq), 
to_sfixed(11269.0/65536.0,1,-nbitq), 
to_sfixed(3839.0/65536.0,1,-nbitq), 
to_sfixed(-6492.0/65536.0,1,-nbitq), 
to_sfixed(-2389.0/65536.0,1,-nbitq), 
to_sfixed(2722.0/65536.0,1,-nbitq), 
to_sfixed(-1066.0/65536.0,1,-nbitq), 
to_sfixed(152.0/65536.0,1,-nbitq), 
to_sfixed(5715.0/65536.0,1,-nbitq), 
to_sfixed(-1591.0/65536.0,1,-nbitq), 
to_sfixed(-791.0/65536.0,1,-nbitq), 
to_sfixed(-225.0/65536.0,1,-nbitq), 
to_sfixed(6171.0/65536.0,1,-nbitq), 
to_sfixed(829.0/65536.0,1,-nbitq), 
to_sfixed(-2297.0/65536.0,1,-nbitq), 
to_sfixed(5629.0/65536.0,1,-nbitq), 
to_sfixed(5409.0/65536.0,1,-nbitq), 
to_sfixed(5675.0/65536.0,1,-nbitq), 
to_sfixed(-679.0/65536.0,1,-nbitq), 
to_sfixed(-3169.0/65536.0,1,-nbitq), 
to_sfixed(9483.0/65536.0,1,-nbitq), 
to_sfixed(505.0/65536.0,1,-nbitq), 
to_sfixed(-2108.0/65536.0,1,-nbitq), 
to_sfixed(-1293.0/65536.0,1,-nbitq), 
to_sfixed(-3530.0/65536.0,1,-nbitq), 
to_sfixed(-421.0/65536.0,1,-nbitq), 
to_sfixed(2008.0/65536.0,1,-nbitq), 
to_sfixed(-12357.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3072.0/65536.0,1,-nbitq), 
to_sfixed(2091.0/65536.0,1,-nbitq), 
to_sfixed(245.0/65536.0,1,-nbitq), 
to_sfixed(6846.0/65536.0,1,-nbitq), 
to_sfixed(-877.0/65536.0,1,-nbitq), 
to_sfixed(8449.0/65536.0,1,-nbitq), 
to_sfixed(-1540.0/65536.0,1,-nbitq), 
to_sfixed(3647.0/65536.0,1,-nbitq), 
to_sfixed(-4065.0/65536.0,1,-nbitq), 
to_sfixed(-405.0/65536.0,1,-nbitq), 
to_sfixed(3020.0/65536.0,1,-nbitq), 
to_sfixed(-7630.0/65536.0,1,-nbitq), 
to_sfixed(-2108.0/65536.0,1,-nbitq), 
to_sfixed(9373.0/65536.0,1,-nbitq), 
to_sfixed(-2230.0/65536.0,1,-nbitq), 
to_sfixed(3143.0/65536.0,1,-nbitq), 
to_sfixed(-2947.0/65536.0,1,-nbitq), 
to_sfixed(6615.0/65536.0,1,-nbitq), 
to_sfixed(1434.0/65536.0,1,-nbitq), 
to_sfixed(1233.0/65536.0,1,-nbitq), 
to_sfixed(2358.0/65536.0,1,-nbitq), 
to_sfixed(-7929.0/65536.0,1,-nbitq), 
to_sfixed(-5684.0/65536.0,1,-nbitq), 
to_sfixed(-2235.0/65536.0,1,-nbitq), 
to_sfixed(-140.0/65536.0,1,-nbitq), 
to_sfixed(11125.0/65536.0,1,-nbitq), 
to_sfixed(-2736.0/65536.0,1,-nbitq), 
to_sfixed(2075.0/65536.0,1,-nbitq), 
to_sfixed(8033.0/65536.0,1,-nbitq), 
to_sfixed(-2415.0/65536.0,1,-nbitq), 
to_sfixed(3221.0/65536.0,1,-nbitq), 
to_sfixed(-10065.0/65536.0,1,-nbitq), 
to_sfixed(7601.0/65536.0,1,-nbitq), 
to_sfixed(7161.0/65536.0,1,-nbitq), 
to_sfixed(-1160.0/65536.0,1,-nbitq), 
to_sfixed(1957.0/65536.0,1,-nbitq), 
to_sfixed(-7630.0/65536.0,1,-nbitq), 
to_sfixed(967.0/65536.0,1,-nbitq), 
to_sfixed(-659.0/65536.0,1,-nbitq), 
to_sfixed(2135.0/65536.0,1,-nbitq), 
to_sfixed(-328.0/65536.0,1,-nbitq), 
to_sfixed(-1196.0/65536.0,1,-nbitq), 
to_sfixed(6162.0/65536.0,1,-nbitq), 
to_sfixed(5457.0/65536.0,1,-nbitq), 
to_sfixed(1980.0/65536.0,1,-nbitq), 
to_sfixed(2999.0/65536.0,1,-nbitq), 
to_sfixed(-3072.0/65536.0,1,-nbitq), 
to_sfixed(4108.0/65536.0,1,-nbitq), 
to_sfixed(-1895.0/65536.0,1,-nbitq), 
to_sfixed(2225.0/65536.0,1,-nbitq), 
to_sfixed(73.0/65536.0,1,-nbitq), 
to_sfixed(2251.0/65536.0,1,-nbitq), 
to_sfixed(4998.0/65536.0,1,-nbitq), 
to_sfixed(12042.0/65536.0,1,-nbitq), 
to_sfixed(-1442.0/65536.0,1,-nbitq), 
to_sfixed(986.0/65536.0,1,-nbitq), 
to_sfixed(2063.0/65536.0,1,-nbitq), 
to_sfixed(914.0/65536.0,1,-nbitq), 
to_sfixed(-2296.0/65536.0,1,-nbitq), 
to_sfixed(-3899.0/65536.0,1,-nbitq), 
to_sfixed(2758.0/65536.0,1,-nbitq), 
to_sfixed(1016.0/65536.0,1,-nbitq), 
to_sfixed(2540.0/65536.0,1,-nbitq), 
to_sfixed(-2547.0/65536.0,1,-nbitq), 
to_sfixed(2672.0/65536.0,1,-nbitq), 
to_sfixed(5233.0/65536.0,1,-nbitq), 
to_sfixed(-1009.0/65536.0,1,-nbitq), 
to_sfixed(2967.0/65536.0,1,-nbitq), 
to_sfixed(-1504.0/65536.0,1,-nbitq), 
to_sfixed(2637.0/65536.0,1,-nbitq), 
to_sfixed(805.0/65536.0,1,-nbitq), 
to_sfixed(-4728.0/65536.0,1,-nbitq), 
to_sfixed(8210.0/65536.0,1,-nbitq), 
to_sfixed(-406.0/65536.0,1,-nbitq), 
to_sfixed(2538.0/65536.0,1,-nbitq), 
to_sfixed(5314.0/65536.0,1,-nbitq), 
to_sfixed(-4366.0/65536.0,1,-nbitq), 
to_sfixed(1295.0/65536.0,1,-nbitq), 
to_sfixed(-1057.0/65536.0,1,-nbitq), 
to_sfixed(-10993.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4250.0/65536.0,1,-nbitq), 
to_sfixed(-3535.0/65536.0,1,-nbitq), 
to_sfixed(-3884.0/65536.0,1,-nbitq), 
to_sfixed(3235.0/65536.0,1,-nbitq), 
to_sfixed(4062.0/65536.0,1,-nbitq), 
to_sfixed(2807.0/65536.0,1,-nbitq), 
to_sfixed(-1265.0/65536.0,1,-nbitq), 
to_sfixed(8347.0/65536.0,1,-nbitq), 
to_sfixed(-247.0/65536.0,1,-nbitq), 
to_sfixed(-2235.0/65536.0,1,-nbitq), 
to_sfixed(3719.0/65536.0,1,-nbitq), 
to_sfixed(-7612.0/65536.0,1,-nbitq), 
to_sfixed(-1662.0/65536.0,1,-nbitq), 
to_sfixed(8139.0/65536.0,1,-nbitq), 
to_sfixed(1260.0/65536.0,1,-nbitq), 
to_sfixed(1894.0/65536.0,1,-nbitq), 
to_sfixed(-1389.0/65536.0,1,-nbitq), 
to_sfixed(10753.0/65536.0,1,-nbitq), 
to_sfixed(617.0/65536.0,1,-nbitq), 
to_sfixed(930.0/65536.0,1,-nbitq), 
to_sfixed(4611.0/65536.0,1,-nbitq), 
to_sfixed(-8153.0/65536.0,1,-nbitq), 
to_sfixed(-3473.0/65536.0,1,-nbitq), 
to_sfixed(7491.0/65536.0,1,-nbitq), 
to_sfixed(678.0/65536.0,1,-nbitq), 
to_sfixed(11912.0/65536.0,1,-nbitq), 
to_sfixed(2332.0/65536.0,1,-nbitq), 
to_sfixed(-28.0/65536.0,1,-nbitq), 
to_sfixed(5638.0/65536.0,1,-nbitq), 
to_sfixed(-315.0/65536.0,1,-nbitq), 
to_sfixed(319.0/65536.0,1,-nbitq), 
to_sfixed(-6099.0/65536.0,1,-nbitq), 
to_sfixed(9209.0/65536.0,1,-nbitq), 
to_sfixed(2129.0/65536.0,1,-nbitq), 
to_sfixed(-6.0/65536.0,1,-nbitq), 
to_sfixed(-859.0/65536.0,1,-nbitq), 
to_sfixed(-5754.0/65536.0,1,-nbitq), 
to_sfixed(-831.0/65536.0,1,-nbitq), 
to_sfixed(-3021.0/65536.0,1,-nbitq), 
to_sfixed(-2705.0/65536.0,1,-nbitq), 
to_sfixed(-320.0/65536.0,1,-nbitq), 
to_sfixed(-2797.0/65536.0,1,-nbitq), 
to_sfixed(8228.0/65536.0,1,-nbitq), 
to_sfixed(5545.0/65536.0,1,-nbitq), 
to_sfixed(-1453.0/65536.0,1,-nbitq), 
to_sfixed(-3639.0/65536.0,1,-nbitq), 
to_sfixed(-152.0/65536.0,1,-nbitq), 
to_sfixed(1210.0/65536.0,1,-nbitq), 
to_sfixed(-2330.0/65536.0,1,-nbitq), 
to_sfixed(2594.0/65536.0,1,-nbitq), 
to_sfixed(1825.0/65536.0,1,-nbitq), 
to_sfixed(3426.0/65536.0,1,-nbitq), 
to_sfixed(6164.0/65536.0,1,-nbitq), 
to_sfixed(10931.0/65536.0,1,-nbitq), 
to_sfixed(-3008.0/65536.0,1,-nbitq), 
to_sfixed(3124.0/65536.0,1,-nbitq), 
to_sfixed(2008.0/65536.0,1,-nbitq), 
to_sfixed(3525.0/65536.0,1,-nbitq), 
to_sfixed(-312.0/65536.0,1,-nbitq), 
to_sfixed(-2326.0/65536.0,1,-nbitq), 
to_sfixed(-2991.0/65536.0,1,-nbitq), 
to_sfixed(-2707.0/65536.0,1,-nbitq), 
to_sfixed(3105.0/65536.0,1,-nbitq), 
to_sfixed(-413.0/65536.0,1,-nbitq), 
to_sfixed(-5440.0/65536.0,1,-nbitq), 
to_sfixed(5308.0/65536.0,1,-nbitq), 
to_sfixed(4084.0/65536.0,1,-nbitq), 
to_sfixed(6091.0/65536.0,1,-nbitq), 
to_sfixed(-4679.0/65536.0,1,-nbitq), 
to_sfixed(-4780.0/65536.0,1,-nbitq), 
to_sfixed(939.0/65536.0,1,-nbitq), 
to_sfixed(-5804.0/65536.0,1,-nbitq), 
to_sfixed(5739.0/65536.0,1,-nbitq), 
to_sfixed(1424.0/65536.0,1,-nbitq), 
to_sfixed(2286.0/65536.0,1,-nbitq), 
to_sfixed(-921.0/65536.0,1,-nbitq), 
to_sfixed(-6493.0/65536.0,1,-nbitq), 
to_sfixed(-620.0/65536.0,1,-nbitq), 
to_sfixed(-16.0/65536.0,1,-nbitq), 
to_sfixed(-7252.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5088.0/65536.0,1,-nbitq), 
to_sfixed(-1579.0/65536.0,1,-nbitq), 
to_sfixed(-888.0/65536.0,1,-nbitq), 
to_sfixed(4049.0/65536.0,1,-nbitq), 
to_sfixed(5044.0/65536.0,1,-nbitq), 
to_sfixed(548.0/65536.0,1,-nbitq), 
to_sfixed(-2696.0/65536.0,1,-nbitq), 
to_sfixed(6303.0/65536.0,1,-nbitq), 
to_sfixed(-6089.0/65536.0,1,-nbitq), 
to_sfixed(272.0/65536.0,1,-nbitq), 
to_sfixed(-9.0/65536.0,1,-nbitq), 
to_sfixed(-7815.0/65536.0,1,-nbitq), 
to_sfixed(1618.0/65536.0,1,-nbitq), 
to_sfixed(1582.0/65536.0,1,-nbitq), 
to_sfixed(-1247.0/65536.0,1,-nbitq), 
to_sfixed(-821.0/65536.0,1,-nbitq), 
to_sfixed(-1741.0/65536.0,1,-nbitq), 
to_sfixed(8131.0/65536.0,1,-nbitq), 
to_sfixed(3572.0/65536.0,1,-nbitq), 
to_sfixed(1214.0/65536.0,1,-nbitq), 
to_sfixed(2063.0/65536.0,1,-nbitq), 
to_sfixed(-4097.0/65536.0,1,-nbitq), 
to_sfixed(-1538.0/65536.0,1,-nbitq), 
to_sfixed(-2168.0/65536.0,1,-nbitq), 
to_sfixed(291.0/65536.0,1,-nbitq), 
to_sfixed(4467.0/65536.0,1,-nbitq), 
to_sfixed(-5988.0/65536.0,1,-nbitq), 
to_sfixed(-3755.0/65536.0,1,-nbitq), 
to_sfixed(7138.0/65536.0,1,-nbitq), 
to_sfixed(-362.0/65536.0,1,-nbitq), 
to_sfixed(4275.0/65536.0,1,-nbitq), 
to_sfixed(-5884.0/65536.0,1,-nbitq), 
to_sfixed(2194.0/65536.0,1,-nbitq), 
to_sfixed(-7272.0/65536.0,1,-nbitq), 
to_sfixed(1210.0/65536.0,1,-nbitq), 
to_sfixed(-1692.0/65536.0,1,-nbitq), 
to_sfixed(-3763.0/65536.0,1,-nbitq), 
to_sfixed(273.0/65536.0,1,-nbitq), 
to_sfixed(242.0/65536.0,1,-nbitq), 
to_sfixed(20.0/65536.0,1,-nbitq), 
to_sfixed(544.0/65536.0,1,-nbitq), 
to_sfixed(1480.0/65536.0,1,-nbitq), 
to_sfixed(2403.0/65536.0,1,-nbitq), 
to_sfixed(3279.0/65536.0,1,-nbitq), 
to_sfixed(150.0/65536.0,1,-nbitq), 
to_sfixed(-4465.0/65536.0,1,-nbitq), 
to_sfixed(-333.0/65536.0,1,-nbitq), 
to_sfixed(-4298.0/65536.0,1,-nbitq), 
to_sfixed(131.0/65536.0,1,-nbitq), 
to_sfixed(4085.0/65536.0,1,-nbitq), 
to_sfixed(-658.0/65536.0,1,-nbitq), 
to_sfixed(2688.0/65536.0,1,-nbitq), 
to_sfixed(1171.0/65536.0,1,-nbitq), 
to_sfixed(11284.0/65536.0,1,-nbitq), 
to_sfixed(-4417.0/65536.0,1,-nbitq), 
to_sfixed(1276.0/65536.0,1,-nbitq), 
to_sfixed(-1244.0/65536.0,1,-nbitq), 
to_sfixed(2694.0/65536.0,1,-nbitq), 
to_sfixed(-1131.0/65536.0,1,-nbitq), 
to_sfixed(-7140.0/65536.0,1,-nbitq), 
to_sfixed(-4941.0/65536.0,1,-nbitq), 
to_sfixed(2507.0/65536.0,1,-nbitq), 
to_sfixed(-1668.0/65536.0,1,-nbitq), 
to_sfixed(427.0/65536.0,1,-nbitq), 
to_sfixed(-2756.0/65536.0,1,-nbitq), 
to_sfixed(69.0/65536.0,1,-nbitq), 
to_sfixed(9063.0/65536.0,1,-nbitq), 
to_sfixed(1738.0/65536.0,1,-nbitq), 
to_sfixed(-792.0/65536.0,1,-nbitq), 
to_sfixed(-1333.0/65536.0,1,-nbitq), 
to_sfixed(4191.0/65536.0,1,-nbitq), 
to_sfixed(-3942.0/65536.0,1,-nbitq), 
to_sfixed(6814.0/65536.0,1,-nbitq), 
to_sfixed(-1920.0/65536.0,1,-nbitq), 
to_sfixed(1107.0/65536.0,1,-nbitq), 
to_sfixed(-4295.0/65536.0,1,-nbitq), 
to_sfixed(-906.0/65536.0,1,-nbitq), 
to_sfixed(1216.0/65536.0,1,-nbitq), 
to_sfixed(1971.0/65536.0,1,-nbitq), 
to_sfixed(-2896.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1864.0/65536.0,1,-nbitq), 
to_sfixed(703.0/65536.0,1,-nbitq), 
to_sfixed(-6871.0/65536.0,1,-nbitq), 
to_sfixed(2349.0/65536.0,1,-nbitq), 
to_sfixed(4122.0/65536.0,1,-nbitq), 
to_sfixed(1598.0/65536.0,1,-nbitq), 
to_sfixed(150.0/65536.0,1,-nbitq), 
to_sfixed(2553.0/65536.0,1,-nbitq), 
to_sfixed(-3502.0/65536.0,1,-nbitq), 
to_sfixed(-1082.0/65536.0,1,-nbitq), 
to_sfixed(2029.0/65536.0,1,-nbitq), 
to_sfixed(-5457.0/65536.0,1,-nbitq), 
to_sfixed(-3333.0/65536.0,1,-nbitq), 
to_sfixed(562.0/65536.0,1,-nbitq), 
to_sfixed(1795.0/65536.0,1,-nbitq), 
to_sfixed(-740.0/65536.0,1,-nbitq), 
to_sfixed(956.0/65536.0,1,-nbitq), 
to_sfixed(4503.0/65536.0,1,-nbitq), 
to_sfixed(2847.0/65536.0,1,-nbitq), 
to_sfixed(1410.0/65536.0,1,-nbitq), 
to_sfixed(1031.0/65536.0,1,-nbitq), 
to_sfixed(-3325.0/65536.0,1,-nbitq), 
to_sfixed(-2932.0/65536.0,1,-nbitq), 
to_sfixed(-523.0/65536.0,1,-nbitq), 
to_sfixed(2386.0/65536.0,1,-nbitq), 
to_sfixed(1680.0/65536.0,1,-nbitq), 
to_sfixed(-2538.0/65536.0,1,-nbitq), 
to_sfixed(-1473.0/65536.0,1,-nbitq), 
to_sfixed(5854.0/65536.0,1,-nbitq), 
to_sfixed(-3745.0/65536.0,1,-nbitq), 
to_sfixed(1511.0/65536.0,1,-nbitq), 
to_sfixed(-2598.0/65536.0,1,-nbitq), 
to_sfixed(975.0/65536.0,1,-nbitq), 
to_sfixed(-3706.0/65536.0,1,-nbitq), 
to_sfixed(1659.0/65536.0,1,-nbitq), 
to_sfixed(2871.0/65536.0,1,-nbitq), 
to_sfixed(-1722.0/65536.0,1,-nbitq), 
to_sfixed(-2368.0/65536.0,1,-nbitq), 
to_sfixed(-5907.0/65536.0,1,-nbitq), 
to_sfixed(3216.0/65536.0,1,-nbitq), 
to_sfixed(-2498.0/65536.0,1,-nbitq), 
to_sfixed(110.0/65536.0,1,-nbitq), 
to_sfixed(1850.0/65536.0,1,-nbitq), 
to_sfixed(2477.0/65536.0,1,-nbitq), 
to_sfixed(171.0/65536.0,1,-nbitq), 
to_sfixed(2046.0/65536.0,1,-nbitq), 
to_sfixed(-1642.0/65536.0,1,-nbitq), 
to_sfixed(-1546.0/65536.0,1,-nbitq), 
to_sfixed(1793.0/65536.0,1,-nbitq), 
to_sfixed(2009.0/65536.0,1,-nbitq), 
to_sfixed(3263.0/65536.0,1,-nbitq), 
to_sfixed(5873.0/65536.0,1,-nbitq), 
to_sfixed(526.0/65536.0,1,-nbitq), 
to_sfixed(6885.0/65536.0,1,-nbitq), 
to_sfixed(-6499.0/65536.0,1,-nbitq), 
to_sfixed(-2535.0/65536.0,1,-nbitq), 
to_sfixed(2018.0/65536.0,1,-nbitq), 
to_sfixed(564.0/65536.0,1,-nbitq), 
to_sfixed(2033.0/65536.0,1,-nbitq), 
to_sfixed(-1862.0/65536.0,1,-nbitq), 
to_sfixed(-5690.0/65536.0,1,-nbitq), 
to_sfixed(2636.0/65536.0,1,-nbitq), 
to_sfixed(-1608.0/65536.0,1,-nbitq), 
to_sfixed(-40.0/65536.0,1,-nbitq), 
to_sfixed(-3613.0/65536.0,1,-nbitq), 
to_sfixed(-403.0/65536.0,1,-nbitq), 
to_sfixed(4609.0/65536.0,1,-nbitq), 
to_sfixed(-1599.0/65536.0,1,-nbitq), 
to_sfixed(5636.0/65536.0,1,-nbitq), 
to_sfixed(3730.0/65536.0,1,-nbitq), 
to_sfixed(1443.0/65536.0,1,-nbitq), 
to_sfixed(-1407.0/65536.0,1,-nbitq), 
to_sfixed(1311.0/65536.0,1,-nbitq), 
to_sfixed(-2876.0/65536.0,1,-nbitq), 
to_sfixed(851.0/65536.0,1,-nbitq), 
to_sfixed(-1361.0/65536.0,1,-nbitq), 
to_sfixed(-4214.0/65536.0,1,-nbitq), 
to_sfixed(2887.0/65536.0,1,-nbitq), 
to_sfixed(1771.0/65536.0,1,-nbitq), 
to_sfixed(2577.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1726.0/65536.0,1,-nbitq), 
to_sfixed(-15.0/65536.0,1,-nbitq), 
to_sfixed(-3205.0/65536.0,1,-nbitq), 
to_sfixed(2826.0/65536.0,1,-nbitq), 
to_sfixed(922.0/65536.0,1,-nbitq), 
to_sfixed(1241.0/65536.0,1,-nbitq), 
to_sfixed(411.0/65536.0,1,-nbitq), 
to_sfixed(3262.0/65536.0,1,-nbitq), 
to_sfixed(-1574.0/65536.0,1,-nbitq), 
to_sfixed(1774.0/65536.0,1,-nbitq), 
to_sfixed(-2273.0/65536.0,1,-nbitq), 
to_sfixed(-4818.0/65536.0,1,-nbitq), 
to_sfixed(1530.0/65536.0,1,-nbitq), 
to_sfixed(2155.0/65536.0,1,-nbitq), 
to_sfixed(1554.0/65536.0,1,-nbitq), 
to_sfixed(-2561.0/65536.0,1,-nbitq), 
to_sfixed(1875.0/65536.0,1,-nbitq), 
to_sfixed(5862.0/65536.0,1,-nbitq), 
to_sfixed(-1233.0/65536.0,1,-nbitq), 
to_sfixed(3060.0/65536.0,1,-nbitq), 
to_sfixed(1687.0/65536.0,1,-nbitq), 
to_sfixed(-997.0/65536.0,1,-nbitq), 
to_sfixed(-1371.0/65536.0,1,-nbitq), 
to_sfixed(-2077.0/65536.0,1,-nbitq), 
to_sfixed(2857.0/65536.0,1,-nbitq), 
to_sfixed(-457.0/65536.0,1,-nbitq), 
to_sfixed(-2079.0/65536.0,1,-nbitq), 
to_sfixed(-850.0/65536.0,1,-nbitq), 
to_sfixed(1164.0/65536.0,1,-nbitq), 
to_sfixed(-831.0/65536.0,1,-nbitq), 
to_sfixed(-2113.0/65536.0,1,-nbitq), 
to_sfixed(-1211.0/65536.0,1,-nbitq), 
to_sfixed(-1529.0/65536.0,1,-nbitq), 
to_sfixed(-5134.0/65536.0,1,-nbitq), 
to_sfixed(373.0/65536.0,1,-nbitq), 
to_sfixed(-2597.0/65536.0,1,-nbitq), 
to_sfixed(-4108.0/65536.0,1,-nbitq), 
to_sfixed(-1462.0/65536.0,1,-nbitq), 
to_sfixed(-3771.0/65536.0,1,-nbitq), 
to_sfixed(-2137.0/65536.0,1,-nbitq), 
to_sfixed(962.0/65536.0,1,-nbitq), 
to_sfixed(-1599.0/65536.0,1,-nbitq), 
to_sfixed(-1152.0/65536.0,1,-nbitq), 
to_sfixed(-1187.0/65536.0,1,-nbitq), 
to_sfixed(3025.0/65536.0,1,-nbitq), 
to_sfixed(2058.0/65536.0,1,-nbitq), 
to_sfixed(861.0/65536.0,1,-nbitq), 
to_sfixed(2607.0/65536.0,1,-nbitq), 
to_sfixed(438.0/65536.0,1,-nbitq), 
to_sfixed(-1135.0/65536.0,1,-nbitq), 
to_sfixed(-584.0/65536.0,1,-nbitq), 
to_sfixed(-805.0/65536.0,1,-nbitq), 
to_sfixed(1132.0/65536.0,1,-nbitq), 
to_sfixed(1053.0/65536.0,1,-nbitq), 
to_sfixed(-2089.0/65536.0,1,-nbitq), 
to_sfixed(652.0/65536.0,1,-nbitq), 
to_sfixed(952.0/65536.0,1,-nbitq), 
to_sfixed(-680.0/65536.0,1,-nbitq), 
to_sfixed(-212.0/65536.0,1,-nbitq), 
to_sfixed(2061.0/65536.0,1,-nbitq), 
to_sfixed(-2371.0/65536.0,1,-nbitq), 
to_sfixed(2087.0/65536.0,1,-nbitq), 
to_sfixed(-680.0/65536.0,1,-nbitq), 
to_sfixed(1200.0/65536.0,1,-nbitq), 
to_sfixed(-2344.0/65536.0,1,-nbitq), 
to_sfixed(-2193.0/65536.0,1,-nbitq), 
to_sfixed(2590.0/65536.0,1,-nbitq), 
to_sfixed(1077.0/65536.0,1,-nbitq), 
to_sfixed(2477.0/65536.0,1,-nbitq), 
to_sfixed(3996.0/65536.0,1,-nbitq), 
to_sfixed(-1209.0/65536.0,1,-nbitq), 
to_sfixed(-670.0/65536.0,1,-nbitq), 
to_sfixed(3238.0/65536.0,1,-nbitq), 
to_sfixed(-2399.0/65536.0,1,-nbitq), 
to_sfixed(2787.0/65536.0,1,-nbitq), 
to_sfixed(-1681.0/65536.0,1,-nbitq), 
to_sfixed(-4248.0/65536.0,1,-nbitq), 
to_sfixed(3960.0/65536.0,1,-nbitq), 
to_sfixed(-2163.0/65536.0,1,-nbitq), 
to_sfixed(3324.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1227.0/65536.0,1,-nbitq), 
to_sfixed(-2696.0/65536.0,1,-nbitq), 
to_sfixed(4398.0/65536.0,1,-nbitq), 
to_sfixed(741.0/65536.0,1,-nbitq), 
to_sfixed(-2608.0/65536.0,1,-nbitq), 
to_sfixed(-2892.0/65536.0,1,-nbitq), 
to_sfixed(-433.0/65536.0,1,-nbitq), 
to_sfixed(816.0/65536.0,1,-nbitq), 
to_sfixed(-2412.0/65536.0,1,-nbitq), 
to_sfixed(652.0/65536.0,1,-nbitq), 
to_sfixed(-1413.0/65536.0,1,-nbitq), 
to_sfixed(-3658.0/65536.0,1,-nbitq), 
to_sfixed(-2197.0/65536.0,1,-nbitq), 
to_sfixed(-2612.0/65536.0,1,-nbitq), 
to_sfixed(-578.0/65536.0,1,-nbitq), 
to_sfixed(1907.0/65536.0,1,-nbitq), 
to_sfixed(-1229.0/65536.0,1,-nbitq), 
to_sfixed(2196.0/65536.0,1,-nbitq), 
to_sfixed(2102.0/65536.0,1,-nbitq), 
to_sfixed(-507.0/65536.0,1,-nbitq), 
to_sfixed(1742.0/65536.0,1,-nbitq), 
to_sfixed(1530.0/65536.0,1,-nbitq), 
to_sfixed(504.0/65536.0,1,-nbitq), 
to_sfixed(734.0/65536.0,1,-nbitq), 
to_sfixed(-1836.0/65536.0,1,-nbitq), 
to_sfixed(-396.0/65536.0,1,-nbitq), 
to_sfixed(-3265.0/65536.0,1,-nbitq), 
to_sfixed(1858.0/65536.0,1,-nbitq), 
to_sfixed(-2330.0/65536.0,1,-nbitq), 
to_sfixed(-2528.0/65536.0,1,-nbitq), 
to_sfixed(-2774.0/65536.0,1,-nbitq), 
to_sfixed(1603.0/65536.0,1,-nbitq), 
to_sfixed(-4128.0/65536.0,1,-nbitq), 
to_sfixed(-4654.0/65536.0,1,-nbitq), 
to_sfixed(1286.0/65536.0,1,-nbitq), 
to_sfixed(960.0/65536.0,1,-nbitq), 
to_sfixed(-2671.0/65536.0,1,-nbitq), 
to_sfixed(-1761.0/65536.0,1,-nbitq), 
to_sfixed(-1052.0/65536.0,1,-nbitq), 
to_sfixed(81.0/65536.0,1,-nbitq), 
to_sfixed(1899.0/65536.0,1,-nbitq), 
to_sfixed(2100.0/65536.0,1,-nbitq), 
to_sfixed(-659.0/65536.0,1,-nbitq), 
to_sfixed(-1289.0/65536.0,1,-nbitq), 
to_sfixed(-750.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(-2238.0/65536.0,1,-nbitq), 
to_sfixed(-984.0/65536.0,1,-nbitq), 
to_sfixed(3445.0/65536.0,1,-nbitq), 
to_sfixed(1351.0/65536.0,1,-nbitq), 
to_sfixed(-1356.0/65536.0,1,-nbitq), 
to_sfixed(1705.0/65536.0,1,-nbitq), 
to_sfixed(2879.0/65536.0,1,-nbitq), 
to_sfixed(-1.0/65536.0,1,-nbitq), 
to_sfixed(3814.0/65536.0,1,-nbitq), 
to_sfixed(2811.0/65536.0,1,-nbitq), 
to_sfixed(154.0/65536.0,1,-nbitq), 
to_sfixed(-515.0/65536.0,1,-nbitq), 
to_sfixed(732.0/65536.0,1,-nbitq), 
to_sfixed(866.0/65536.0,1,-nbitq), 
to_sfixed(-2438.0/65536.0,1,-nbitq), 
to_sfixed(1554.0/65536.0,1,-nbitq), 
to_sfixed(-1419.0/65536.0,1,-nbitq), 
to_sfixed(-2282.0/65536.0,1,-nbitq), 
to_sfixed(2820.0/65536.0,1,-nbitq), 
to_sfixed(-1798.0/65536.0,1,-nbitq), 
to_sfixed(2488.0/65536.0,1,-nbitq), 
to_sfixed(-1131.0/65536.0,1,-nbitq), 
to_sfixed(-168.0/65536.0,1,-nbitq), 
to_sfixed(-219.0/65536.0,1,-nbitq), 
to_sfixed(-950.0/65536.0,1,-nbitq), 
to_sfixed(385.0/65536.0,1,-nbitq), 
to_sfixed(-2.0/65536.0,1,-nbitq), 
to_sfixed(-1479.0/65536.0,1,-nbitq), 
to_sfixed(1797.0/65536.0,1,-nbitq), 
to_sfixed(1068.0/65536.0,1,-nbitq), 
to_sfixed(-80.0/65536.0,1,-nbitq), 
to_sfixed(3475.0/65536.0,1,-nbitq), 
to_sfixed(-2001.0/65536.0,1,-nbitq), 
to_sfixed(1561.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(163.0/65536.0,1,-nbitq), 
to_sfixed(-926.0/65536.0,1,-nbitq), 
to_sfixed(2419.0/65536.0,1,-nbitq), 
to_sfixed(-3496.0/65536.0,1,-nbitq), 
to_sfixed(-535.0/65536.0,1,-nbitq), 
to_sfixed(-1231.0/65536.0,1,-nbitq), 
to_sfixed(2470.0/65536.0,1,-nbitq), 
to_sfixed(2842.0/65536.0,1,-nbitq), 
to_sfixed(-1574.0/65536.0,1,-nbitq), 
to_sfixed(-1125.0/65536.0,1,-nbitq), 
to_sfixed(-3951.0/65536.0,1,-nbitq), 
to_sfixed(-2915.0/65536.0,1,-nbitq), 
to_sfixed(-213.0/65536.0,1,-nbitq), 
to_sfixed(-4749.0/65536.0,1,-nbitq), 
to_sfixed(-114.0/65536.0,1,-nbitq), 
to_sfixed(1065.0/65536.0,1,-nbitq), 
to_sfixed(2501.0/65536.0,1,-nbitq), 
to_sfixed(3588.0/65536.0,1,-nbitq), 
to_sfixed(376.0/65536.0,1,-nbitq), 
to_sfixed(-2385.0/65536.0,1,-nbitq), 
to_sfixed(-2474.0/65536.0,1,-nbitq), 
to_sfixed(1194.0/65536.0,1,-nbitq), 
to_sfixed(169.0/65536.0,1,-nbitq), 
to_sfixed(589.0/65536.0,1,-nbitq), 
to_sfixed(-82.0/65536.0,1,-nbitq), 
to_sfixed(2332.0/65536.0,1,-nbitq), 
to_sfixed(1445.0/65536.0,1,-nbitq), 
to_sfixed(1266.0/65536.0,1,-nbitq), 
to_sfixed(-1003.0/65536.0,1,-nbitq), 
to_sfixed(-3162.0/65536.0,1,-nbitq), 
to_sfixed(-1950.0/65536.0,1,-nbitq), 
to_sfixed(-1658.0/65536.0,1,-nbitq), 
to_sfixed(-511.0/65536.0,1,-nbitq), 
to_sfixed(-1314.0/65536.0,1,-nbitq), 
to_sfixed(-4.0/65536.0,1,-nbitq), 
to_sfixed(-511.0/65536.0,1,-nbitq), 
to_sfixed(-3414.0/65536.0,1,-nbitq), 
to_sfixed(-2224.0/65536.0,1,-nbitq), 
to_sfixed(-2941.0/65536.0,1,-nbitq), 
to_sfixed(-670.0/65536.0,1,-nbitq), 
to_sfixed(-2882.0/65536.0,1,-nbitq), 
to_sfixed(1135.0/65536.0,1,-nbitq), 
to_sfixed(-3070.0/65536.0,1,-nbitq), 
to_sfixed(226.0/65536.0,1,-nbitq), 
to_sfixed(1328.0/65536.0,1,-nbitq), 
to_sfixed(4527.0/65536.0,1,-nbitq), 
to_sfixed(547.0/65536.0,1,-nbitq), 
to_sfixed(2143.0/65536.0,1,-nbitq), 
to_sfixed(3162.0/65536.0,1,-nbitq), 
to_sfixed(4462.0/65536.0,1,-nbitq), 
to_sfixed(-2476.0/65536.0,1,-nbitq), 
to_sfixed(-3318.0/65536.0,1,-nbitq), 
to_sfixed(3047.0/65536.0,1,-nbitq), 
to_sfixed(-1226.0/65536.0,1,-nbitq), 
to_sfixed(1640.0/65536.0,1,-nbitq), 
to_sfixed(695.0/65536.0,1,-nbitq), 
to_sfixed(-370.0/65536.0,1,-nbitq), 
to_sfixed(1046.0/65536.0,1,-nbitq), 
to_sfixed(-699.0/65536.0,1,-nbitq), 
to_sfixed(3780.0/65536.0,1,-nbitq), 
to_sfixed(-720.0/65536.0,1,-nbitq), 
to_sfixed(-2432.0/65536.0,1,-nbitq), 
to_sfixed(1486.0/65536.0,1,-nbitq), 
to_sfixed(-2905.0/65536.0,1,-nbitq), 
to_sfixed(-647.0/65536.0,1,-nbitq), 
to_sfixed(-395.0/65536.0,1,-nbitq), 
to_sfixed(-63.0/65536.0,1,-nbitq), 
to_sfixed(-577.0/65536.0,1,-nbitq), 
to_sfixed(2905.0/65536.0,1,-nbitq), 
to_sfixed(-1489.0/65536.0,1,-nbitq), 
to_sfixed(-880.0/65536.0,1,-nbitq), 
to_sfixed(1149.0/65536.0,1,-nbitq), 
to_sfixed(2587.0/65536.0,1,-nbitq), 
to_sfixed(-1568.0/65536.0,1,-nbitq), 
to_sfixed(-2048.0/65536.0,1,-nbitq), 
to_sfixed(1369.0/65536.0,1,-nbitq), 
to_sfixed(-1806.0/65536.0,1,-nbitq), 
to_sfixed(2142.0/65536.0,1,-nbitq), 
to_sfixed(-2953.0/65536.0,1,-nbitq), 
to_sfixed(4990.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2791.0/65536.0,1,-nbitq), 
to_sfixed(-482.0/65536.0,1,-nbitq), 
to_sfixed(3786.0/65536.0,1,-nbitq), 
to_sfixed(-1501.0/65536.0,1,-nbitq), 
to_sfixed(809.0/65536.0,1,-nbitq), 
to_sfixed(-4107.0/65536.0,1,-nbitq), 
to_sfixed(-3848.0/65536.0,1,-nbitq), 
to_sfixed(-2480.0/65536.0,1,-nbitq), 
to_sfixed(2417.0/65536.0,1,-nbitq), 
to_sfixed(1875.0/65536.0,1,-nbitq), 
to_sfixed(-1785.0/65536.0,1,-nbitq), 
to_sfixed(-189.0/65536.0,1,-nbitq), 
to_sfixed(1988.0/65536.0,1,-nbitq), 
to_sfixed(-3706.0/65536.0,1,-nbitq), 
to_sfixed(3313.0/65536.0,1,-nbitq), 
to_sfixed(2176.0/65536.0,1,-nbitq), 
to_sfixed(-2618.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(2219.0/65536.0,1,-nbitq), 
to_sfixed(1279.0/65536.0,1,-nbitq), 
to_sfixed(-3181.0/65536.0,1,-nbitq), 
to_sfixed(2605.0/65536.0,1,-nbitq), 
to_sfixed(-2438.0/65536.0,1,-nbitq), 
to_sfixed(-872.0/65536.0,1,-nbitq), 
to_sfixed(1280.0/65536.0,1,-nbitq), 
to_sfixed(5080.0/65536.0,1,-nbitq), 
to_sfixed(-298.0/65536.0,1,-nbitq), 
to_sfixed(2340.0/65536.0,1,-nbitq), 
to_sfixed(2484.0/65536.0,1,-nbitq), 
to_sfixed(-3576.0/65536.0,1,-nbitq), 
to_sfixed(-2497.0/65536.0,1,-nbitq), 
to_sfixed(432.0/65536.0,1,-nbitq), 
to_sfixed(195.0/65536.0,1,-nbitq), 
to_sfixed(-103.0/65536.0,1,-nbitq), 
to_sfixed(-2902.0/65536.0,1,-nbitq), 
to_sfixed(2534.0/65536.0,1,-nbitq), 
to_sfixed(-44.0/65536.0,1,-nbitq), 
to_sfixed(-29.0/65536.0,1,-nbitq), 
to_sfixed(-3588.0/65536.0,1,-nbitq), 
to_sfixed(-2043.0/65536.0,1,-nbitq), 
to_sfixed(-3674.0/65536.0,1,-nbitq), 
to_sfixed(2019.0/65536.0,1,-nbitq), 
to_sfixed(-4502.0/65536.0,1,-nbitq), 
to_sfixed(-323.0/65536.0,1,-nbitq), 
to_sfixed(-1619.0/65536.0,1,-nbitq), 
to_sfixed(1590.0/65536.0,1,-nbitq), 
to_sfixed(-2376.0/65536.0,1,-nbitq), 
to_sfixed(-162.0/65536.0,1,-nbitq), 
to_sfixed(1105.0/65536.0,1,-nbitq), 
to_sfixed(353.0/65536.0,1,-nbitq), 
to_sfixed(-1187.0/65536.0,1,-nbitq), 
to_sfixed(-1933.0/65536.0,1,-nbitq), 
to_sfixed(-660.0/65536.0,1,-nbitq), 
to_sfixed(2143.0/65536.0,1,-nbitq), 
to_sfixed(125.0/65536.0,1,-nbitq), 
to_sfixed(-2304.0/65536.0,1,-nbitq), 
to_sfixed(-1088.0/65536.0,1,-nbitq), 
to_sfixed(2869.0/65536.0,1,-nbitq), 
to_sfixed(-153.0/65536.0,1,-nbitq), 
to_sfixed(2449.0/65536.0,1,-nbitq), 
to_sfixed(-3562.0/65536.0,1,-nbitq), 
to_sfixed(2281.0/65536.0,1,-nbitq), 
to_sfixed(-1858.0/65536.0,1,-nbitq), 
to_sfixed(-1702.0/65536.0,1,-nbitq), 
to_sfixed(-2943.0/65536.0,1,-nbitq), 
to_sfixed(2112.0/65536.0,1,-nbitq), 
to_sfixed(-766.0/65536.0,1,-nbitq), 
to_sfixed(2321.0/65536.0,1,-nbitq), 
to_sfixed(-787.0/65536.0,1,-nbitq), 
to_sfixed(-1992.0/65536.0,1,-nbitq), 
to_sfixed(-2154.0/65536.0,1,-nbitq), 
to_sfixed(-1832.0/65536.0,1,-nbitq), 
to_sfixed(4041.0/65536.0,1,-nbitq), 
to_sfixed(1534.0/65536.0,1,-nbitq), 
to_sfixed(2049.0/65536.0,1,-nbitq), 
to_sfixed(4326.0/65536.0,1,-nbitq), 
to_sfixed(-2235.0/65536.0,1,-nbitq), 
to_sfixed(2799.0/65536.0,1,-nbitq), 
to_sfixed(-1402.0/65536.0,1,-nbitq), 
to_sfixed(3495.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1596.0/65536.0,1,-nbitq), 
to_sfixed(738.0/65536.0,1,-nbitq), 
to_sfixed(2701.0/65536.0,1,-nbitq), 
to_sfixed(-1036.0/65536.0,1,-nbitq), 
to_sfixed(3708.0/65536.0,1,-nbitq), 
to_sfixed(-1024.0/65536.0,1,-nbitq), 
to_sfixed(-5183.0/65536.0,1,-nbitq), 
to_sfixed(-2594.0/65536.0,1,-nbitq), 
to_sfixed(-84.0/65536.0,1,-nbitq), 
to_sfixed(-2029.0/65536.0,1,-nbitq), 
to_sfixed(-1409.0/65536.0,1,-nbitq), 
to_sfixed(399.0/65536.0,1,-nbitq), 
to_sfixed(2889.0/65536.0,1,-nbitq), 
to_sfixed(1007.0/65536.0,1,-nbitq), 
to_sfixed(5685.0/65536.0,1,-nbitq), 
to_sfixed(19.0/65536.0,1,-nbitq), 
to_sfixed(-1651.0/65536.0,1,-nbitq), 
to_sfixed(-2118.0/65536.0,1,-nbitq), 
to_sfixed(942.0/65536.0,1,-nbitq), 
to_sfixed(698.0/65536.0,1,-nbitq), 
to_sfixed(-3613.0/65536.0,1,-nbitq), 
to_sfixed(-1538.0/65536.0,1,-nbitq), 
to_sfixed(-773.0/65536.0,1,-nbitq), 
to_sfixed(3763.0/65536.0,1,-nbitq), 
to_sfixed(446.0/65536.0,1,-nbitq), 
to_sfixed(7993.0/65536.0,1,-nbitq), 
to_sfixed(4153.0/65536.0,1,-nbitq), 
to_sfixed(-137.0/65536.0,1,-nbitq), 
to_sfixed(56.0/65536.0,1,-nbitq), 
to_sfixed(-1805.0/65536.0,1,-nbitq), 
to_sfixed(-3928.0/65536.0,1,-nbitq), 
to_sfixed(493.0/65536.0,1,-nbitq), 
to_sfixed(-3032.0/65536.0,1,-nbitq), 
to_sfixed(1310.0/65536.0,1,-nbitq), 
to_sfixed(-502.0/65536.0,1,-nbitq), 
to_sfixed(1355.0/65536.0,1,-nbitq), 
to_sfixed(-1378.0/65536.0,1,-nbitq), 
to_sfixed(-6272.0/65536.0,1,-nbitq), 
to_sfixed(-1132.0/65536.0,1,-nbitq), 
to_sfixed(1574.0/65536.0,1,-nbitq), 
to_sfixed(259.0/65536.0,1,-nbitq), 
to_sfixed(-998.0/65536.0,1,-nbitq), 
to_sfixed(-1267.0/65536.0,1,-nbitq), 
to_sfixed(-571.0/65536.0,1,-nbitq), 
to_sfixed(2429.0/65536.0,1,-nbitq), 
to_sfixed(2708.0/65536.0,1,-nbitq), 
to_sfixed(2639.0/65536.0,1,-nbitq), 
to_sfixed(-63.0/65536.0,1,-nbitq), 
to_sfixed(-1443.0/65536.0,1,-nbitq), 
to_sfixed(81.0/65536.0,1,-nbitq), 
to_sfixed(-543.0/65536.0,1,-nbitq), 
to_sfixed(-3660.0/65536.0,1,-nbitq), 
to_sfixed(-1301.0/65536.0,1,-nbitq), 
to_sfixed(1282.0/65536.0,1,-nbitq), 
to_sfixed(1044.0/65536.0,1,-nbitq), 
to_sfixed(5146.0/65536.0,1,-nbitq), 
to_sfixed(-1016.0/65536.0,1,-nbitq), 
to_sfixed(-1101.0/65536.0,1,-nbitq), 
to_sfixed(-1923.0/65536.0,1,-nbitq), 
to_sfixed(6430.0/65536.0,1,-nbitq), 
to_sfixed(-4256.0/65536.0,1,-nbitq), 
to_sfixed(-3161.0/65536.0,1,-nbitq), 
to_sfixed(2947.0/65536.0,1,-nbitq), 
to_sfixed(2473.0/65536.0,1,-nbitq), 
to_sfixed(2700.0/65536.0,1,-nbitq), 
to_sfixed(203.0/65536.0,1,-nbitq), 
to_sfixed(-3288.0/65536.0,1,-nbitq), 
to_sfixed(-4153.0/65536.0,1,-nbitq), 
to_sfixed(732.0/65536.0,1,-nbitq), 
to_sfixed(899.0/65536.0,1,-nbitq), 
to_sfixed(-394.0/65536.0,1,-nbitq), 
to_sfixed(-842.0/65536.0,1,-nbitq), 
to_sfixed(-2079.0/65536.0,1,-nbitq), 
to_sfixed(-2668.0/65536.0,1,-nbitq), 
to_sfixed(2075.0/65536.0,1,-nbitq), 
to_sfixed(-235.0/65536.0,1,-nbitq), 
to_sfixed(1311.0/65536.0,1,-nbitq), 
to_sfixed(-185.0/65536.0,1,-nbitq), 
to_sfixed(-1999.0/65536.0,1,-nbitq), 
to_sfixed(-731.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1455.0/65536.0,1,-nbitq), 
to_sfixed(344.0/65536.0,1,-nbitq), 
to_sfixed(6723.0/65536.0,1,-nbitq), 
to_sfixed(4880.0/65536.0,1,-nbitq), 
to_sfixed(-232.0/65536.0,1,-nbitq), 
to_sfixed(523.0/65536.0,1,-nbitq), 
to_sfixed(-4897.0/65536.0,1,-nbitq), 
to_sfixed(-615.0/65536.0,1,-nbitq), 
to_sfixed(-1510.0/65536.0,1,-nbitq), 
to_sfixed(179.0/65536.0,1,-nbitq), 
to_sfixed(-490.0/65536.0,1,-nbitq), 
to_sfixed(9040.0/65536.0,1,-nbitq), 
to_sfixed(1476.0/65536.0,1,-nbitq), 
to_sfixed(5622.0/65536.0,1,-nbitq), 
to_sfixed(3284.0/65536.0,1,-nbitq), 
to_sfixed(-1160.0/65536.0,1,-nbitq), 
to_sfixed(-1895.0/65536.0,1,-nbitq), 
to_sfixed(-5686.0/65536.0,1,-nbitq), 
to_sfixed(2732.0/65536.0,1,-nbitq), 
to_sfixed(3237.0/65536.0,1,-nbitq), 
to_sfixed(-4515.0/65536.0,1,-nbitq), 
to_sfixed(4054.0/65536.0,1,-nbitq), 
to_sfixed(983.0/65536.0,1,-nbitq), 
to_sfixed(12091.0/65536.0,1,-nbitq), 
to_sfixed(-885.0/65536.0,1,-nbitq), 
to_sfixed(17204.0/65536.0,1,-nbitq), 
to_sfixed(3577.0/65536.0,1,-nbitq), 
to_sfixed(1632.0/65536.0,1,-nbitq), 
to_sfixed(-2998.0/65536.0,1,-nbitq), 
to_sfixed(1088.0/65536.0,1,-nbitq), 
to_sfixed(-2314.0/65536.0,1,-nbitq), 
to_sfixed(1733.0/65536.0,1,-nbitq), 
to_sfixed(2615.0/65536.0,1,-nbitq), 
to_sfixed(-125.0/65536.0,1,-nbitq), 
to_sfixed(2191.0/65536.0,1,-nbitq), 
to_sfixed(-2682.0/65536.0,1,-nbitq), 
to_sfixed(-4781.0/65536.0,1,-nbitq), 
to_sfixed(-6593.0/65536.0,1,-nbitq), 
to_sfixed(-3292.0/65536.0,1,-nbitq), 
to_sfixed(-3401.0/65536.0,1,-nbitq), 
to_sfixed(3453.0/65536.0,1,-nbitq), 
to_sfixed(-133.0/65536.0,1,-nbitq), 
to_sfixed(-1861.0/65536.0,1,-nbitq), 
to_sfixed(1513.0/65536.0,1,-nbitq), 
to_sfixed(-2417.0/65536.0,1,-nbitq), 
to_sfixed(2875.0/65536.0,1,-nbitq), 
to_sfixed(-1422.0/65536.0,1,-nbitq), 
to_sfixed(2327.0/65536.0,1,-nbitq), 
to_sfixed(-1096.0/65536.0,1,-nbitq), 
to_sfixed(2168.0/65536.0,1,-nbitq), 
to_sfixed(1264.0/65536.0,1,-nbitq), 
to_sfixed(-1768.0/65536.0,1,-nbitq), 
to_sfixed(-403.0/65536.0,1,-nbitq), 
to_sfixed(9432.0/65536.0,1,-nbitq), 
to_sfixed(-2904.0/65536.0,1,-nbitq), 
to_sfixed(7445.0/65536.0,1,-nbitq), 
to_sfixed(-1905.0/65536.0,1,-nbitq), 
to_sfixed(19.0/65536.0,1,-nbitq), 
to_sfixed(-2650.0/65536.0,1,-nbitq), 
to_sfixed(1954.0/65536.0,1,-nbitq), 
to_sfixed(-3620.0/65536.0,1,-nbitq), 
to_sfixed(-2393.0/65536.0,1,-nbitq), 
to_sfixed(2984.0/65536.0,1,-nbitq), 
to_sfixed(-1016.0/65536.0,1,-nbitq), 
to_sfixed(4847.0/65536.0,1,-nbitq), 
to_sfixed(4757.0/65536.0,1,-nbitq), 
to_sfixed(-2697.0/65536.0,1,-nbitq), 
to_sfixed(-9510.0/65536.0,1,-nbitq), 
to_sfixed(-3560.0/65536.0,1,-nbitq), 
to_sfixed(-3811.0/65536.0,1,-nbitq), 
to_sfixed(-2102.0/65536.0,1,-nbitq), 
to_sfixed(-3458.0/65536.0,1,-nbitq), 
to_sfixed(304.0/65536.0,1,-nbitq), 
to_sfixed(864.0/65536.0,1,-nbitq), 
to_sfixed(-338.0/65536.0,1,-nbitq), 
to_sfixed(25.0/65536.0,1,-nbitq), 
to_sfixed(-3243.0/65536.0,1,-nbitq), 
to_sfixed(-2834.0/65536.0,1,-nbitq), 
to_sfixed(82.0/65536.0,1,-nbitq), 
to_sfixed(583.0/65536.0,1,-nbitq)  ), 
( to_sfixed(781.0/65536.0,1,-nbitq), 
to_sfixed(-540.0/65536.0,1,-nbitq), 
to_sfixed(2446.0/65536.0,1,-nbitq), 
to_sfixed(6428.0/65536.0,1,-nbitq), 
to_sfixed(3044.0/65536.0,1,-nbitq), 
to_sfixed(3750.0/65536.0,1,-nbitq), 
to_sfixed(-4647.0/65536.0,1,-nbitq), 
to_sfixed(3790.0/65536.0,1,-nbitq), 
to_sfixed(1298.0/65536.0,1,-nbitq), 
to_sfixed(-2046.0/65536.0,1,-nbitq), 
to_sfixed(1535.0/65536.0,1,-nbitq), 
to_sfixed(13110.0/65536.0,1,-nbitq), 
to_sfixed(-2264.0/65536.0,1,-nbitq), 
to_sfixed(3711.0/65536.0,1,-nbitq), 
to_sfixed(3584.0/65536.0,1,-nbitq), 
to_sfixed(3109.0/65536.0,1,-nbitq), 
to_sfixed(-2729.0/65536.0,1,-nbitq), 
to_sfixed(-6349.0/65536.0,1,-nbitq), 
to_sfixed(-820.0/65536.0,1,-nbitq), 
to_sfixed(-803.0/65536.0,1,-nbitq), 
to_sfixed(-1436.0/65536.0,1,-nbitq), 
to_sfixed(146.0/65536.0,1,-nbitq), 
to_sfixed(4776.0/65536.0,1,-nbitq), 
to_sfixed(6742.0/65536.0,1,-nbitq), 
to_sfixed(-310.0/65536.0,1,-nbitq), 
to_sfixed(13373.0/65536.0,1,-nbitq), 
to_sfixed(11103.0/65536.0,1,-nbitq), 
to_sfixed(-274.0/65536.0,1,-nbitq), 
to_sfixed(4305.0/65536.0,1,-nbitq), 
to_sfixed(5183.0/65536.0,1,-nbitq), 
to_sfixed(-2111.0/65536.0,1,-nbitq), 
to_sfixed(1422.0/65536.0,1,-nbitq), 
to_sfixed(5076.0/65536.0,1,-nbitq), 
to_sfixed(-2060.0/65536.0,1,-nbitq), 
to_sfixed(-777.0/65536.0,1,-nbitq), 
to_sfixed(1592.0/65536.0,1,-nbitq), 
to_sfixed(-4604.0/65536.0,1,-nbitq), 
to_sfixed(1721.0/65536.0,1,-nbitq), 
to_sfixed(-5285.0/65536.0,1,-nbitq), 
to_sfixed(-7962.0/65536.0,1,-nbitq), 
to_sfixed(2154.0/65536.0,1,-nbitq), 
to_sfixed(2554.0/65536.0,1,-nbitq), 
to_sfixed(-1962.0/65536.0,1,-nbitq), 
to_sfixed(-3143.0/65536.0,1,-nbitq), 
to_sfixed(-1465.0/65536.0,1,-nbitq), 
to_sfixed(2135.0/65536.0,1,-nbitq), 
to_sfixed(-1791.0/65536.0,1,-nbitq), 
to_sfixed(3011.0/65536.0,1,-nbitq), 
to_sfixed(-775.0/65536.0,1,-nbitq), 
to_sfixed(4548.0/65536.0,1,-nbitq), 
to_sfixed(-1319.0/65536.0,1,-nbitq), 
to_sfixed(-2312.0/65536.0,1,-nbitq), 
to_sfixed(1146.0/65536.0,1,-nbitq), 
to_sfixed(7108.0/65536.0,1,-nbitq), 
to_sfixed(-2951.0/65536.0,1,-nbitq), 
to_sfixed(12754.0/65536.0,1,-nbitq), 
to_sfixed(-1647.0/65536.0,1,-nbitq), 
to_sfixed(-1973.0/65536.0,1,-nbitq), 
to_sfixed(1199.0/65536.0,1,-nbitq), 
to_sfixed(-2362.0/65536.0,1,-nbitq), 
to_sfixed(-3688.0/65536.0,1,-nbitq), 
to_sfixed(-597.0/65536.0,1,-nbitq), 
to_sfixed(2096.0/65536.0,1,-nbitq), 
to_sfixed(-2372.0/65536.0,1,-nbitq), 
to_sfixed(5851.0/65536.0,1,-nbitq), 
to_sfixed(10477.0/65536.0,1,-nbitq), 
to_sfixed(-1111.0/65536.0,1,-nbitq), 
to_sfixed(-15304.0/65536.0,1,-nbitq), 
to_sfixed(-7430.0/65536.0,1,-nbitq), 
to_sfixed(-2245.0/65536.0,1,-nbitq), 
to_sfixed(2073.0/65536.0,1,-nbitq), 
to_sfixed(-4074.0/65536.0,1,-nbitq), 
to_sfixed(-2865.0/65536.0,1,-nbitq), 
to_sfixed(1947.0/65536.0,1,-nbitq), 
to_sfixed(-1997.0/65536.0,1,-nbitq), 
to_sfixed(-1574.0/65536.0,1,-nbitq), 
to_sfixed(1972.0/65536.0,1,-nbitq), 
to_sfixed(-294.0/65536.0,1,-nbitq), 
to_sfixed(1162.0/65536.0,1,-nbitq), 
to_sfixed(-1259.0/65536.0,1,-nbitq)  ), 
( to_sfixed(716.0/65536.0,1,-nbitq), 
to_sfixed(159.0/65536.0,1,-nbitq), 
to_sfixed(4559.0/65536.0,1,-nbitq), 
to_sfixed(8162.0/65536.0,1,-nbitq), 
to_sfixed(3357.0/65536.0,1,-nbitq), 
to_sfixed(8069.0/65536.0,1,-nbitq), 
to_sfixed(-3926.0/65536.0,1,-nbitq), 
to_sfixed(4117.0/65536.0,1,-nbitq), 
to_sfixed(4787.0/65536.0,1,-nbitq), 
to_sfixed(-869.0/65536.0,1,-nbitq), 
to_sfixed(5359.0/65536.0,1,-nbitq), 
to_sfixed(21305.0/65536.0,1,-nbitq), 
to_sfixed(2044.0/65536.0,1,-nbitq), 
to_sfixed(-1167.0/65536.0,1,-nbitq), 
to_sfixed(-1896.0/65536.0,1,-nbitq), 
to_sfixed(2888.0/65536.0,1,-nbitq), 
to_sfixed(817.0/65536.0,1,-nbitq), 
to_sfixed(988.0/65536.0,1,-nbitq), 
to_sfixed(5321.0/65536.0,1,-nbitq), 
to_sfixed(1121.0/65536.0,1,-nbitq), 
to_sfixed(-3111.0/65536.0,1,-nbitq), 
to_sfixed(207.0/65536.0,1,-nbitq), 
to_sfixed(-3386.0/65536.0,1,-nbitq), 
to_sfixed(-5717.0/65536.0,1,-nbitq), 
to_sfixed(852.0/65536.0,1,-nbitq), 
to_sfixed(14450.0/65536.0,1,-nbitq), 
to_sfixed(17793.0/65536.0,1,-nbitq), 
to_sfixed(2674.0/65536.0,1,-nbitq), 
to_sfixed(2419.0/65536.0,1,-nbitq), 
to_sfixed(5758.0/65536.0,1,-nbitq), 
to_sfixed(-4960.0/65536.0,1,-nbitq), 
to_sfixed(-618.0/65536.0,1,-nbitq), 
to_sfixed(1163.0/65536.0,1,-nbitq), 
to_sfixed(-10764.0/65536.0,1,-nbitq), 
to_sfixed(-2619.0/65536.0,1,-nbitq), 
to_sfixed(2230.0/65536.0,1,-nbitq), 
to_sfixed(-8718.0/65536.0,1,-nbitq), 
to_sfixed(6487.0/65536.0,1,-nbitq), 
to_sfixed(-15231.0/65536.0,1,-nbitq), 
to_sfixed(-6889.0/65536.0,1,-nbitq), 
to_sfixed(446.0/65536.0,1,-nbitq), 
to_sfixed(1417.0/65536.0,1,-nbitq), 
to_sfixed(-591.0/65536.0,1,-nbitq), 
to_sfixed(1015.0/65536.0,1,-nbitq), 
to_sfixed(-1951.0/65536.0,1,-nbitq), 
to_sfixed(-733.0/65536.0,1,-nbitq), 
to_sfixed(-2446.0/65536.0,1,-nbitq), 
to_sfixed(-344.0/65536.0,1,-nbitq), 
to_sfixed(4113.0/65536.0,1,-nbitq), 
to_sfixed(1219.0/65536.0,1,-nbitq), 
to_sfixed(-812.0/65536.0,1,-nbitq), 
to_sfixed(4253.0/65536.0,1,-nbitq), 
to_sfixed(-2333.0/65536.0,1,-nbitq), 
to_sfixed(5426.0/65536.0,1,-nbitq), 
to_sfixed(-4033.0/65536.0,1,-nbitq), 
to_sfixed(10646.0/65536.0,1,-nbitq), 
to_sfixed(-1851.0/65536.0,1,-nbitq), 
to_sfixed(1336.0/65536.0,1,-nbitq), 
to_sfixed(4049.0/65536.0,1,-nbitq), 
to_sfixed(-1770.0/65536.0,1,-nbitq), 
to_sfixed(-6818.0/65536.0,1,-nbitq), 
to_sfixed(-823.0/65536.0,1,-nbitq), 
to_sfixed(-1627.0/65536.0,1,-nbitq), 
to_sfixed(-2379.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(6847.0/65536.0,1,-nbitq), 
to_sfixed(-1883.0/65536.0,1,-nbitq), 
to_sfixed(-14923.0/65536.0,1,-nbitq), 
to_sfixed(-6997.0/65536.0,1,-nbitq), 
to_sfixed(-412.0/65536.0,1,-nbitq), 
to_sfixed(899.0/65536.0,1,-nbitq), 
to_sfixed(-6705.0/65536.0,1,-nbitq), 
to_sfixed(-1319.0/65536.0,1,-nbitq), 
to_sfixed(2299.0/65536.0,1,-nbitq), 
to_sfixed(-2277.0/65536.0,1,-nbitq), 
to_sfixed(2244.0/65536.0,1,-nbitq), 
to_sfixed(-2236.0/65536.0,1,-nbitq), 
to_sfixed(-2288.0/65536.0,1,-nbitq), 
to_sfixed(1030.0/65536.0,1,-nbitq), 
to_sfixed(-6024.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1980.0/65536.0,1,-nbitq), 
to_sfixed(1104.0/65536.0,1,-nbitq), 
to_sfixed(5563.0/65536.0,1,-nbitq), 
to_sfixed(3641.0/65536.0,1,-nbitq), 
to_sfixed(-3123.0/65536.0,1,-nbitq), 
to_sfixed(2117.0/65536.0,1,-nbitq), 
to_sfixed(1296.0/65536.0,1,-nbitq), 
to_sfixed(2656.0/65536.0,1,-nbitq), 
to_sfixed(8239.0/65536.0,1,-nbitq), 
to_sfixed(-2193.0/65536.0,1,-nbitq), 
to_sfixed(2980.0/65536.0,1,-nbitq), 
to_sfixed(17248.0/65536.0,1,-nbitq), 
to_sfixed(598.0/65536.0,1,-nbitq), 
to_sfixed(4984.0/65536.0,1,-nbitq), 
to_sfixed(-2905.0/65536.0,1,-nbitq), 
to_sfixed(-168.0/65536.0,1,-nbitq), 
to_sfixed(-829.0/65536.0,1,-nbitq), 
to_sfixed(11582.0/65536.0,1,-nbitq), 
to_sfixed(3932.0/65536.0,1,-nbitq), 
to_sfixed(-2518.0/65536.0,1,-nbitq), 
to_sfixed(-838.0/65536.0,1,-nbitq), 
to_sfixed(-4424.0/65536.0,1,-nbitq), 
to_sfixed(-3974.0/65536.0,1,-nbitq), 
to_sfixed(-9417.0/65536.0,1,-nbitq), 
to_sfixed(994.0/65536.0,1,-nbitq), 
to_sfixed(15245.0/65536.0,1,-nbitq), 
to_sfixed(7547.0/65536.0,1,-nbitq), 
to_sfixed(3487.0/65536.0,1,-nbitq), 
to_sfixed(-3929.0/65536.0,1,-nbitq), 
to_sfixed(-1028.0/65536.0,1,-nbitq), 
to_sfixed(-3078.0/65536.0,1,-nbitq), 
to_sfixed(-4201.0/65536.0,1,-nbitq), 
to_sfixed(-4314.0/65536.0,1,-nbitq), 
to_sfixed(-1732.0/65536.0,1,-nbitq), 
to_sfixed(165.0/65536.0,1,-nbitq), 
to_sfixed(561.0/65536.0,1,-nbitq), 
to_sfixed(-4861.0/65536.0,1,-nbitq), 
to_sfixed(7913.0/65536.0,1,-nbitq), 
to_sfixed(-13599.0/65536.0,1,-nbitq), 
to_sfixed(-3377.0/65536.0,1,-nbitq), 
to_sfixed(3601.0/65536.0,1,-nbitq), 
to_sfixed(-2436.0/65536.0,1,-nbitq), 
to_sfixed(-3484.0/65536.0,1,-nbitq), 
to_sfixed(4022.0/65536.0,1,-nbitq), 
to_sfixed(-428.0/65536.0,1,-nbitq), 
to_sfixed(3895.0/65536.0,1,-nbitq), 
to_sfixed(1420.0/65536.0,1,-nbitq), 
to_sfixed(1830.0/65536.0,1,-nbitq), 
to_sfixed(-302.0/65536.0,1,-nbitq), 
to_sfixed(-2308.0/65536.0,1,-nbitq), 
to_sfixed(-1621.0/65536.0,1,-nbitq), 
to_sfixed(7525.0/65536.0,1,-nbitq), 
to_sfixed(-1836.0/65536.0,1,-nbitq), 
to_sfixed(6473.0/65536.0,1,-nbitq), 
to_sfixed(-2849.0/65536.0,1,-nbitq), 
to_sfixed(12433.0/65536.0,1,-nbitq), 
to_sfixed(2846.0/65536.0,1,-nbitq), 
to_sfixed(945.0/65536.0,1,-nbitq), 
to_sfixed(1111.0/65536.0,1,-nbitq), 
to_sfixed(-329.0/65536.0,1,-nbitq), 
to_sfixed(-4889.0/65536.0,1,-nbitq), 
to_sfixed(-382.0/65536.0,1,-nbitq), 
to_sfixed(-1743.0/65536.0,1,-nbitq), 
to_sfixed(-600.0/65536.0,1,-nbitq), 
to_sfixed(-3610.0/65536.0,1,-nbitq), 
to_sfixed(2491.0/65536.0,1,-nbitq), 
to_sfixed(-824.0/65536.0,1,-nbitq), 
to_sfixed(-12130.0/65536.0,1,-nbitq), 
to_sfixed(-5753.0/65536.0,1,-nbitq), 
to_sfixed(-618.0/65536.0,1,-nbitq), 
to_sfixed(-3613.0/65536.0,1,-nbitq), 
to_sfixed(-5193.0/65536.0,1,-nbitq), 
to_sfixed(-1555.0/65536.0,1,-nbitq), 
to_sfixed(-1476.0/65536.0,1,-nbitq), 
to_sfixed(1315.0/65536.0,1,-nbitq), 
to_sfixed(-3090.0/65536.0,1,-nbitq), 
to_sfixed(5558.0/65536.0,1,-nbitq), 
to_sfixed(-4084.0/65536.0,1,-nbitq), 
to_sfixed(-1451.0/65536.0,1,-nbitq), 
to_sfixed(-4999.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-430.0/65536.0,1,-nbitq), 
to_sfixed(1984.0/65536.0,1,-nbitq), 
to_sfixed(2607.0/65536.0,1,-nbitq), 
to_sfixed(9340.0/65536.0,1,-nbitq), 
to_sfixed(-2952.0/65536.0,1,-nbitq), 
to_sfixed(751.0/65536.0,1,-nbitq), 
to_sfixed(-1015.0/65536.0,1,-nbitq), 
to_sfixed(-2432.0/65536.0,1,-nbitq), 
to_sfixed(3572.0/65536.0,1,-nbitq), 
to_sfixed(3089.0/65536.0,1,-nbitq), 
to_sfixed(2513.0/65536.0,1,-nbitq), 
to_sfixed(8160.0/65536.0,1,-nbitq), 
to_sfixed(-255.0/65536.0,1,-nbitq), 
to_sfixed(9638.0/65536.0,1,-nbitq), 
to_sfixed(2542.0/65536.0,1,-nbitq), 
to_sfixed(-2926.0/65536.0,1,-nbitq), 
to_sfixed(-2563.0/65536.0,1,-nbitq), 
to_sfixed(10524.0/65536.0,1,-nbitq), 
to_sfixed(2740.0/65536.0,1,-nbitq), 
to_sfixed(-2395.0/65536.0,1,-nbitq), 
to_sfixed(-3558.0/65536.0,1,-nbitq), 
to_sfixed(-549.0/65536.0,1,-nbitq), 
to_sfixed(-1554.0/65536.0,1,-nbitq), 
to_sfixed(-2093.0/65536.0,1,-nbitq), 
to_sfixed(-4120.0/65536.0,1,-nbitq), 
to_sfixed(9567.0/65536.0,1,-nbitq), 
to_sfixed(15077.0/65536.0,1,-nbitq), 
to_sfixed(1047.0/65536.0,1,-nbitq), 
to_sfixed(7695.0/65536.0,1,-nbitq), 
to_sfixed(-6497.0/65536.0,1,-nbitq), 
to_sfixed(-6461.0/65536.0,1,-nbitq), 
to_sfixed(-1604.0/65536.0,1,-nbitq), 
to_sfixed(-4327.0/65536.0,1,-nbitq), 
to_sfixed(1148.0/65536.0,1,-nbitq), 
to_sfixed(2055.0/65536.0,1,-nbitq), 
to_sfixed(109.0/65536.0,1,-nbitq), 
to_sfixed(-5176.0/65536.0,1,-nbitq), 
to_sfixed(3614.0/65536.0,1,-nbitq), 
to_sfixed(-10936.0/65536.0,1,-nbitq), 
to_sfixed(-1778.0/65536.0,1,-nbitq), 
to_sfixed(-389.0/65536.0,1,-nbitq), 
to_sfixed(1098.0/65536.0,1,-nbitq), 
to_sfixed(-6644.0/65536.0,1,-nbitq), 
to_sfixed(-149.0/65536.0,1,-nbitq), 
to_sfixed(2889.0/65536.0,1,-nbitq), 
to_sfixed(686.0/65536.0,1,-nbitq), 
to_sfixed(257.0/65536.0,1,-nbitq), 
to_sfixed(4279.0/65536.0,1,-nbitq), 
to_sfixed(1014.0/65536.0,1,-nbitq), 
to_sfixed(1805.0/65536.0,1,-nbitq), 
to_sfixed(1512.0/65536.0,1,-nbitq), 
to_sfixed(7748.0/65536.0,1,-nbitq), 
to_sfixed(45.0/65536.0,1,-nbitq), 
to_sfixed(8164.0/65536.0,1,-nbitq), 
to_sfixed(1097.0/65536.0,1,-nbitq), 
to_sfixed(15612.0/65536.0,1,-nbitq), 
to_sfixed(1101.0/65536.0,1,-nbitq), 
to_sfixed(520.0/65536.0,1,-nbitq), 
to_sfixed(-852.0/65536.0,1,-nbitq), 
to_sfixed(4400.0/65536.0,1,-nbitq), 
to_sfixed(475.0/65536.0,1,-nbitq), 
to_sfixed(665.0/65536.0,1,-nbitq), 
to_sfixed(1785.0/65536.0,1,-nbitq), 
to_sfixed(-660.0/65536.0,1,-nbitq), 
to_sfixed(-7228.0/65536.0,1,-nbitq), 
to_sfixed(4260.0/65536.0,1,-nbitq), 
to_sfixed(2935.0/65536.0,1,-nbitq), 
to_sfixed(-8517.0/65536.0,1,-nbitq), 
to_sfixed(-2515.0/65536.0,1,-nbitq), 
to_sfixed(-611.0/65536.0,1,-nbitq), 
to_sfixed(-239.0/65536.0,1,-nbitq), 
to_sfixed(-8900.0/65536.0,1,-nbitq), 
to_sfixed(-939.0/65536.0,1,-nbitq), 
to_sfixed(-786.0/65536.0,1,-nbitq), 
to_sfixed(2336.0/65536.0,1,-nbitq), 
to_sfixed(2244.0/65536.0,1,-nbitq), 
to_sfixed(12114.0/65536.0,1,-nbitq), 
to_sfixed(-2056.0/65536.0,1,-nbitq), 
to_sfixed(-1401.0/65536.0,1,-nbitq), 
to_sfixed(-1001.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2174.0/65536.0,1,-nbitq), 
to_sfixed(-3872.0/65536.0,1,-nbitq), 
to_sfixed(-4952.0/65536.0,1,-nbitq), 
to_sfixed(9431.0/65536.0,1,-nbitq), 
to_sfixed(-7360.0/65536.0,1,-nbitq), 
to_sfixed(6632.0/65536.0,1,-nbitq), 
to_sfixed(-4613.0/65536.0,1,-nbitq), 
to_sfixed(-8083.0/65536.0,1,-nbitq), 
to_sfixed(2739.0/65536.0,1,-nbitq), 
to_sfixed(-472.0/65536.0,1,-nbitq), 
to_sfixed(408.0/65536.0,1,-nbitq), 
to_sfixed(1168.0/65536.0,1,-nbitq), 
to_sfixed(600.0/65536.0,1,-nbitq), 
to_sfixed(6275.0/65536.0,1,-nbitq), 
to_sfixed(4669.0/65536.0,1,-nbitq), 
to_sfixed(-2089.0/65536.0,1,-nbitq), 
to_sfixed(677.0/65536.0,1,-nbitq), 
to_sfixed(2207.0/65536.0,1,-nbitq), 
to_sfixed(5806.0/65536.0,1,-nbitq), 
to_sfixed(-89.0/65536.0,1,-nbitq), 
to_sfixed(-4832.0/65536.0,1,-nbitq), 
to_sfixed(-4413.0/65536.0,1,-nbitq), 
to_sfixed(5536.0/65536.0,1,-nbitq), 
to_sfixed(-2900.0/65536.0,1,-nbitq), 
to_sfixed(-2699.0/65536.0,1,-nbitq), 
to_sfixed(8195.0/65536.0,1,-nbitq), 
to_sfixed(16015.0/65536.0,1,-nbitq), 
to_sfixed(2914.0/65536.0,1,-nbitq), 
to_sfixed(6607.0/65536.0,1,-nbitq), 
to_sfixed(-9730.0/65536.0,1,-nbitq), 
to_sfixed(-6603.0/65536.0,1,-nbitq), 
to_sfixed(1138.0/65536.0,1,-nbitq), 
to_sfixed(-145.0/65536.0,1,-nbitq), 
to_sfixed(1585.0/65536.0,1,-nbitq), 
to_sfixed(2340.0/65536.0,1,-nbitq), 
to_sfixed(-1427.0/65536.0,1,-nbitq), 
to_sfixed(2052.0/65536.0,1,-nbitq), 
to_sfixed(-2510.0/65536.0,1,-nbitq), 
to_sfixed(-5344.0/65536.0,1,-nbitq), 
to_sfixed(-2243.0/65536.0,1,-nbitq), 
to_sfixed(5949.0/65536.0,1,-nbitq), 
to_sfixed(425.0/65536.0,1,-nbitq), 
to_sfixed(-3986.0/65536.0,1,-nbitq), 
to_sfixed(-2557.0/65536.0,1,-nbitq), 
to_sfixed(1397.0/65536.0,1,-nbitq), 
to_sfixed(-9209.0/65536.0,1,-nbitq), 
to_sfixed(-871.0/65536.0,1,-nbitq), 
to_sfixed(1642.0/65536.0,1,-nbitq), 
to_sfixed(-263.0/65536.0,1,-nbitq), 
to_sfixed(1702.0/65536.0,1,-nbitq), 
to_sfixed(-932.0/65536.0,1,-nbitq), 
to_sfixed(11435.0/65536.0,1,-nbitq), 
to_sfixed(702.0/65536.0,1,-nbitq), 
to_sfixed(2476.0/65536.0,1,-nbitq), 
to_sfixed(-2021.0/65536.0,1,-nbitq), 
to_sfixed(11341.0/65536.0,1,-nbitq), 
to_sfixed(-1831.0/65536.0,1,-nbitq), 
to_sfixed(-1070.0/65536.0,1,-nbitq), 
to_sfixed(2403.0/65536.0,1,-nbitq), 
to_sfixed(6979.0/65536.0,1,-nbitq), 
to_sfixed(4185.0/65536.0,1,-nbitq), 
to_sfixed(443.0/65536.0,1,-nbitq), 
to_sfixed(-1682.0/65536.0,1,-nbitq), 
to_sfixed(-1925.0/65536.0,1,-nbitq), 
to_sfixed(-838.0/65536.0,1,-nbitq), 
to_sfixed(4523.0/65536.0,1,-nbitq), 
to_sfixed(-3205.0/65536.0,1,-nbitq), 
to_sfixed(-9988.0/65536.0,1,-nbitq), 
to_sfixed(-3466.0/65536.0,1,-nbitq), 
to_sfixed(-5435.0/65536.0,1,-nbitq), 
to_sfixed(-2203.0/65536.0,1,-nbitq), 
to_sfixed(-7935.0/65536.0,1,-nbitq), 
to_sfixed(-548.0/65536.0,1,-nbitq), 
to_sfixed(1343.0/65536.0,1,-nbitq), 
to_sfixed(-2258.0/65536.0,1,-nbitq), 
to_sfixed(4899.0/65536.0,1,-nbitq), 
to_sfixed(4536.0/65536.0,1,-nbitq), 
to_sfixed(-12261.0/65536.0,1,-nbitq), 
to_sfixed(-195.0/65536.0,1,-nbitq), 
to_sfixed(-185.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4590.0/65536.0,1,-nbitq), 
to_sfixed(-1300.0/65536.0,1,-nbitq), 
to_sfixed(1572.0/65536.0,1,-nbitq), 
to_sfixed(13636.0/65536.0,1,-nbitq), 
to_sfixed(-7983.0/65536.0,1,-nbitq), 
to_sfixed(1010.0/65536.0,1,-nbitq), 
to_sfixed(-3819.0/65536.0,1,-nbitq), 
to_sfixed(-8762.0/65536.0,1,-nbitq), 
to_sfixed(1986.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(3890.0/65536.0,1,-nbitq), 
to_sfixed(6349.0/65536.0,1,-nbitq), 
to_sfixed(1976.0/65536.0,1,-nbitq), 
to_sfixed(2358.0/65536.0,1,-nbitq), 
to_sfixed(978.0/65536.0,1,-nbitq), 
to_sfixed(1080.0/65536.0,1,-nbitq), 
to_sfixed(659.0/65536.0,1,-nbitq), 
to_sfixed(8073.0/65536.0,1,-nbitq), 
to_sfixed(-8421.0/65536.0,1,-nbitq), 
to_sfixed(-6.0/65536.0,1,-nbitq), 
to_sfixed(477.0/65536.0,1,-nbitq), 
to_sfixed(-11743.0/65536.0,1,-nbitq), 
to_sfixed(4468.0/65536.0,1,-nbitq), 
to_sfixed(-4291.0/65536.0,1,-nbitq), 
to_sfixed(-2280.0/65536.0,1,-nbitq), 
to_sfixed(2466.0/65536.0,1,-nbitq), 
to_sfixed(12154.0/65536.0,1,-nbitq), 
to_sfixed(-522.0/65536.0,1,-nbitq), 
to_sfixed(9768.0/65536.0,1,-nbitq), 
to_sfixed(-10580.0/65536.0,1,-nbitq), 
to_sfixed(-3845.0/65536.0,1,-nbitq), 
to_sfixed(5765.0/65536.0,1,-nbitq), 
to_sfixed(3096.0/65536.0,1,-nbitq), 
to_sfixed(9718.0/65536.0,1,-nbitq), 
to_sfixed(1118.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(7852.0/65536.0,1,-nbitq), 
to_sfixed(-5877.0/65536.0,1,-nbitq), 
to_sfixed(-12294.0/65536.0,1,-nbitq), 
to_sfixed(-4765.0/65536.0,1,-nbitq), 
to_sfixed(11485.0/65536.0,1,-nbitq), 
to_sfixed(514.0/65536.0,1,-nbitq), 
to_sfixed(-1349.0/65536.0,1,-nbitq), 
to_sfixed(-7198.0/65536.0,1,-nbitq), 
to_sfixed(-1186.0/65536.0,1,-nbitq), 
to_sfixed(-16718.0/65536.0,1,-nbitq), 
to_sfixed(3849.0/65536.0,1,-nbitq), 
to_sfixed(1766.0/65536.0,1,-nbitq), 
to_sfixed(480.0/65536.0,1,-nbitq), 
to_sfixed(2307.0/65536.0,1,-nbitq), 
to_sfixed(-1687.0/65536.0,1,-nbitq), 
to_sfixed(11325.0/65536.0,1,-nbitq), 
to_sfixed(687.0/65536.0,1,-nbitq), 
to_sfixed(5007.0/65536.0,1,-nbitq), 
to_sfixed(-972.0/65536.0,1,-nbitq), 
to_sfixed(-2099.0/65536.0,1,-nbitq), 
to_sfixed(653.0/65536.0,1,-nbitq), 
to_sfixed(-545.0/65536.0,1,-nbitq), 
to_sfixed(503.0/65536.0,1,-nbitq), 
to_sfixed(8932.0/65536.0,1,-nbitq), 
to_sfixed(13253.0/65536.0,1,-nbitq), 
to_sfixed(-247.0/65536.0,1,-nbitq), 
to_sfixed(-2485.0/65536.0,1,-nbitq), 
to_sfixed(-1241.0/65536.0,1,-nbitq), 
to_sfixed(698.0/65536.0,1,-nbitq), 
to_sfixed(2276.0/65536.0,1,-nbitq), 
to_sfixed(-3938.0/65536.0,1,-nbitq), 
to_sfixed(-7568.0/65536.0,1,-nbitq), 
to_sfixed(-3642.0/65536.0,1,-nbitq), 
to_sfixed(-7609.0/65536.0,1,-nbitq), 
to_sfixed(3080.0/65536.0,1,-nbitq), 
to_sfixed(-4802.0/65536.0,1,-nbitq), 
to_sfixed(550.0/65536.0,1,-nbitq), 
to_sfixed(1099.0/65536.0,1,-nbitq), 
to_sfixed(-2743.0/65536.0,1,-nbitq), 
to_sfixed(3084.0/65536.0,1,-nbitq), 
to_sfixed(-15669.0/65536.0,1,-nbitq), 
to_sfixed(-17914.0/65536.0,1,-nbitq), 
to_sfixed(912.0/65536.0,1,-nbitq), 
to_sfixed(-1978.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1713.0/65536.0,1,-nbitq), 
to_sfixed(-3869.0/65536.0,1,-nbitq), 
to_sfixed(8347.0/65536.0,1,-nbitq), 
to_sfixed(9231.0/65536.0,1,-nbitq), 
to_sfixed(194.0/65536.0,1,-nbitq), 
to_sfixed(1096.0/65536.0,1,-nbitq), 
to_sfixed(308.0/65536.0,1,-nbitq), 
to_sfixed(-2039.0/65536.0,1,-nbitq), 
to_sfixed(4158.0/65536.0,1,-nbitq), 
to_sfixed(-1489.0/65536.0,1,-nbitq), 
to_sfixed(1472.0/65536.0,1,-nbitq), 
to_sfixed(7287.0/65536.0,1,-nbitq), 
to_sfixed(-187.0/65536.0,1,-nbitq), 
to_sfixed(-12686.0/65536.0,1,-nbitq), 
to_sfixed(2205.0/65536.0,1,-nbitq), 
to_sfixed(1599.0/65536.0,1,-nbitq), 
to_sfixed(1596.0/65536.0,1,-nbitq), 
to_sfixed(13685.0/65536.0,1,-nbitq), 
to_sfixed(-10091.0/65536.0,1,-nbitq), 
to_sfixed(-154.0/65536.0,1,-nbitq), 
to_sfixed(3033.0/65536.0,1,-nbitq), 
to_sfixed(-11947.0/65536.0,1,-nbitq), 
to_sfixed(5474.0/65536.0,1,-nbitq), 
to_sfixed(-5068.0/65536.0,1,-nbitq), 
to_sfixed(-2278.0/65536.0,1,-nbitq), 
to_sfixed(-684.0/65536.0,1,-nbitq), 
to_sfixed(9452.0/65536.0,1,-nbitq), 
to_sfixed(-751.0/65536.0,1,-nbitq), 
to_sfixed(11316.0/65536.0,1,-nbitq), 
to_sfixed(-7250.0/65536.0,1,-nbitq), 
to_sfixed(-962.0/65536.0,1,-nbitq), 
to_sfixed(11475.0/65536.0,1,-nbitq), 
to_sfixed(7461.0/65536.0,1,-nbitq), 
to_sfixed(20374.0/65536.0,1,-nbitq), 
to_sfixed(-2842.0/65536.0,1,-nbitq), 
to_sfixed(1814.0/65536.0,1,-nbitq), 
to_sfixed(11125.0/65536.0,1,-nbitq), 
to_sfixed(-4664.0/65536.0,1,-nbitq), 
to_sfixed(-9528.0/65536.0,1,-nbitq), 
to_sfixed(-4881.0/65536.0,1,-nbitq), 
to_sfixed(6977.0/65536.0,1,-nbitq), 
to_sfixed(-1501.0/65536.0,1,-nbitq), 
to_sfixed(-725.0/65536.0,1,-nbitq), 
to_sfixed(-2791.0/65536.0,1,-nbitq), 
to_sfixed(2017.0/65536.0,1,-nbitq), 
to_sfixed(-14395.0/65536.0,1,-nbitq), 
to_sfixed(1531.0/65536.0,1,-nbitq), 
to_sfixed(-3909.0/65536.0,1,-nbitq), 
to_sfixed(-1778.0/65536.0,1,-nbitq), 
to_sfixed(2.0/65536.0,1,-nbitq), 
to_sfixed(716.0/65536.0,1,-nbitq), 
to_sfixed(3680.0/65536.0,1,-nbitq), 
to_sfixed(-4495.0/65536.0,1,-nbitq), 
to_sfixed(6367.0/65536.0,1,-nbitq), 
to_sfixed(3678.0/65536.0,1,-nbitq), 
to_sfixed(2197.0/65536.0,1,-nbitq), 
to_sfixed(1178.0/65536.0,1,-nbitq), 
to_sfixed(-916.0/65536.0,1,-nbitq), 
to_sfixed(-2063.0/65536.0,1,-nbitq), 
to_sfixed(6560.0/65536.0,1,-nbitq), 
to_sfixed(13094.0/65536.0,1,-nbitq), 
to_sfixed(1962.0/65536.0,1,-nbitq), 
to_sfixed(-2077.0/65536.0,1,-nbitq), 
to_sfixed(-1137.0/65536.0,1,-nbitq), 
to_sfixed(-12434.0/65536.0,1,-nbitq), 
to_sfixed(-6454.0/65536.0,1,-nbitq), 
to_sfixed(4265.0/65536.0,1,-nbitq), 
to_sfixed(-3234.0/65536.0,1,-nbitq), 
to_sfixed(-6326.0/65536.0,1,-nbitq), 
to_sfixed(-3204.0/65536.0,1,-nbitq), 
to_sfixed(-355.0/65536.0,1,-nbitq), 
to_sfixed(6420.0/65536.0,1,-nbitq), 
to_sfixed(-1123.0/65536.0,1,-nbitq), 
to_sfixed(-1089.0/65536.0,1,-nbitq), 
to_sfixed(-2761.0/65536.0,1,-nbitq), 
to_sfixed(-5223.0/65536.0,1,-nbitq), 
to_sfixed(-8968.0/65536.0,1,-nbitq), 
to_sfixed(-12180.0/65536.0,1,-nbitq), 
to_sfixed(-2110.0/65536.0,1,-nbitq), 
to_sfixed(-636.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-7054.0/65536.0,1,-nbitq), 
to_sfixed(1288.0/65536.0,1,-nbitq), 
to_sfixed(-5709.0/65536.0,1,-nbitq), 
to_sfixed(13540.0/65536.0,1,-nbitq), 
to_sfixed(10422.0/65536.0,1,-nbitq), 
to_sfixed(7198.0/65536.0,1,-nbitq), 
to_sfixed(1762.0/65536.0,1,-nbitq), 
to_sfixed(5661.0/65536.0,1,-nbitq), 
to_sfixed(-4324.0/65536.0,1,-nbitq), 
to_sfixed(1045.0/65536.0,1,-nbitq), 
to_sfixed(4896.0/65536.0,1,-nbitq), 
to_sfixed(9276.0/65536.0,1,-nbitq), 
to_sfixed(-666.0/65536.0,1,-nbitq), 
to_sfixed(-9368.0/65536.0,1,-nbitq), 
to_sfixed(-3377.0/65536.0,1,-nbitq), 
to_sfixed(408.0/65536.0,1,-nbitq), 
to_sfixed(514.0/65536.0,1,-nbitq), 
to_sfixed(-9666.0/65536.0,1,-nbitq), 
to_sfixed(-6081.0/65536.0,1,-nbitq), 
to_sfixed(1220.0/65536.0,1,-nbitq), 
to_sfixed(-5910.0/65536.0,1,-nbitq), 
to_sfixed(-21993.0/65536.0,1,-nbitq), 
to_sfixed(-3310.0/65536.0,1,-nbitq), 
to_sfixed(28.0/65536.0,1,-nbitq), 
to_sfixed(-846.0/65536.0,1,-nbitq), 
to_sfixed(8769.0/65536.0,1,-nbitq), 
to_sfixed(6476.0/65536.0,1,-nbitq), 
to_sfixed(5779.0/65536.0,1,-nbitq), 
to_sfixed(6412.0/65536.0,1,-nbitq), 
to_sfixed(1683.0/65536.0,1,-nbitq), 
to_sfixed(1651.0/65536.0,1,-nbitq), 
to_sfixed(6953.0/65536.0,1,-nbitq), 
to_sfixed(9266.0/65536.0,1,-nbitq), 
to_sfixed(14626.0/65536.0,1,-nbitq), 
to_sfixed(-458.0/65536.0,1,-nbitq), 
to_sfixed(1657.0/65536.0,1,-nbitq), 
to_sfixed(12216.0/65536.0,1,-nbitq), 
to_sfixed(-3031.0/65536.0,1,-nbitq), 
to_sfixed(-22677.0/65536.0,1,-nbitq), 
to_sfixed(-3980.0/65536.0,1,-nbitq), 
to_sfixed(-2238.0/65536.0,1,-nbitq), 
to_sfixed(1265.0/65536.0,1,-nbitq), 
to_sfixed(1247.0/65536.0,1,-nbitq), 
to_sfixed(1.0/65536.0,1,-nbitq), 
to_sfixed(-1388.0/65536.0,1,-nbitq), 
to_sfixed(11878.0/65536.0,1,-nbitq), 
to_sfixed(857.0/65536.0,1,-nbitq), 
to_sfixed(-2365.0/65536.0,1,-nbitq), 
to_sfixed(-1269.0/65536.0,1,-nbitq), 
to_sfixed(295.0/65536.0,1,-nbitq), 
to_sfixed(-380.0/65536.0,1,-nbitq), 
to_sfixed(3737.0/65536.0,1,-nbitq), 
to_sfixed(-8943.0/65536.0,1,-nbitq), 
to_sfixed(4677.0/65536.0,1,-nbitq), 
to_sfixed(726.0/65536.0,1,-nbitq), 
to_sfixed(1791.0/65536.0,1,-nbitq), 
to_sfixed(3642.0/65536.0,1,-nbitq), 
to_sfixed(-2044.0/65536.0,1,-nbitq), 
to_sfixed(2742.0/65536.0,1,-nbitq), 
to_sfixed(6832.0/65536.0,1,-nbitq), 
to_sfixed(5414.0/65536.0,1,-nbitq), 
to_sfixed(-958.0/65536.0,1,-nbitq), 
to_sfixed(-1050.0/65536.0,1,-nbitq), 
to_sfixed(1238.0/65536.0,1,-nbitq), 
to_sfixed(-7432.0/65536.0,1,-nbitq), 
to_sfixed(-17465.0/65536.0,1,-nbitq), 
to_sfixed(1295.0/65536.0,1,-nbitq), 
to_sfixed(-6573.0/65536.0,1,-nbitq), 
to_sfixed(-12225.0/65536.0,1,-nbitq), 
to_sfixed(-10506.0/65536.0,1,-nbitq), 
to_sfixed(-4598.0/65536.0,1,-nbitq), 
to_sfixed(5203.0/65536.0,1,-nbitq), 
to_sfixed(-4701.0/65536.0,1,-nbitq), 
to_sfixed(-681.0/65536.0,1,-nbitq), 
to_sfixed(476.0/65536.0,1,-nbitq), 
to_sfixed(-17667.0/65536.0,1,-nbitq), 
to_sfixed(-6645.0/65536.0,1,-nbitq), 
to_sfixed(4648.0/65536.0,1,-nbitq), 
to_sfixed(3452.0/65536.0,1,-nbitq), 
to_sfixed(-6678.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-6424.0/65536.0,1,-nbitq), 
to_sfixed(1317.0/65536.0,1,-nbitq), 
to_sfixed(-14685.0/65536.0,1,-nbitq), 
to_sfixed(13216.0/65536.0,1,-nbitq), 
to_sfixed(23895.0/65536.0,1,-nbitq), 
to_sfixed(6296.0/65536.0,1,-nbitq), 
to_sfixed(1614.0/65536.0,1,-nbitq), 
to_sfixed(16068.0/65536.0,1,-nbitq), 
to_sfixed(-1185.0/65536.0,1,-nbitq), 
to_sfixed(3162.0/65536.0,1,-nbitq), 
to_sfixed(5985.0/65536.0,1,-nbitq), 
to_sfixed(15462.0/65536.0,1,-nbitq), 
to_sfixed(560.0/65536.0,1,-nbitq), 
to_sfixed(1039.0/65536.0,1,-nbitq), 
to_sfixed(-6924.0/65536.0,1,-nbitq), 
to_sfixed(1953.0/65536.0,1,-nbitq), 
to_sfixed(-2355.0/65536.0,1,-nbitq), 
to_sfixed(-8030.0/65536.0,1,-nbitq), 
to_sfixed(-6718.0/65536.0,1,-nbitq), 
to_sfixed(-2037.0/65536.0,1,-nbitq), 
to_sfixed(-4723.0/65536.0,1,-nbitq), 
to_sfixed(-21761.0/65536.0,1,-nbitq), 
to_sfixed(-8537.0/65536.0,1,-nbitq), 
to_sfixed(-5115.0/65536.0,1,-nbitq), 
to_sfixed(-1903.0/65536.0,1,-nbitq), 
to_sfixed(773.0/65536.0,1,-nbitq), 
to_sfixed(5917.0/65536.0,1,-nbitq), 
to_sfixed(3487.0/65536.0,1,-nbitq), 
to_sfixed(5212.0/65536.0,1,-nbitq), 
to_sfixed(3116.0/65536.0,1,-nbitq), 
to_sfixed(-9130.0/65536.0,1,-nbitq), 
to_sfixed(6088.0/65536.0,1,-nbitq), 
to_sfixed(10203.0/65536.0,1,-nbitq), 
to_sfixed(-3965.0/65536.0,1,-nbitq), 
to_sfixed(1825.0/65536.0,1,-nbitq), 
to_sfixed(586.0/65536.0,1,-nbitq), 
to_sfixed(6834.0/65536.0,1,-nbitq), 
to_sfixed(-5741.0/65536.0,1,-nbitq), 
to_sfixed(-3571.0/65536.0,1,-nbitq), 
to_sfixed(329.0/65536.0,1,-nbitq), 
to_sfixed(1029.0/65536.0,1,-nbitq), 
to_sfixed(-2215.0/65536.0,1,-nbitq), 
to_sfixed(112.0/65536.0,1,-nbitq), 
to_sfixed(-11178.0/65536.0,1,-nbitq), 
to_sfixed(-1881.0/65536.0,1,-nbitq), 
to_sfixed(17990.0/65536.0,1,-nbitq), 
to_sfixed(1372.0/65536.0,1,-nbitq), 
to_sfixed(-8515.0/65536.0,1,-nbitq), 
to_sfixed(-322.0/65536.0,1,-nbitq), 
to_sfixed(824.0/65536.0,1,-nbitq), 
to_sfixed(-1557.0/65536.0,1,-nbitq), 
to_sfixed(3903.0/65536.0,1,-nbitq), 
to_sfixed(-7140.0/65536.0,1,-nbitq), 
to_sfixed(3485.0/65536.0,1,-nbitq), 
to_sfixed(2574.0/65536.0,1,-nbitq), 
to_sfixed(7633.0/65536.0,1,-nbitq), 
to_sfixed(3721.0/65536.0,1,-nbitq), 
to_sfixed(3460.0/65536.0,1,-nbitq), 
to_sfixed(2185.0/65536.0,1,-nbitq), 
to_sfixed(3719.0/65536.0,1,-nbitq), 
to_sfixed(-7354.0/65536.0,1,-nbitq), 
to_sfixed(1928.0/65536.0,1,-nbitq), 
to_sfixed(-516.0/65536.0,1,-nbitq), 
to_sfixed(-90.0/65536.0,1,-nbitq), 
to_sfixed(-10557.0/65536.0,1,-nbitq), 
to_sfixed(-10896.0/65536.0,1,-nbitq), 
to_sfixed(-3902.0/65536.0,1,-nbitq), 
to_sfixed(-10588.0/65536.0,1,-nbitq), 
to_sfixed(-21740.0/65536.0,1,-nbitq), 
to_sfixed(369.0/65536.0,1,-nbitq), 
to_sfixed(-4771.0/65536.0,1,-nbitq), 
to_sfixed(10970.0/65536.0,1,-nbitq), 
to_sfixed(-2056.0/65536.0,1,-nbitq), 
to_sfixed(428.0/65536.0,1,-nbitq), 
to_sfixed(-607.0/65536.0,1,-nbitq), 
to_sfixed(-17514.0/65536.0,1,-nbitq), 
to_sfixed(-9365.0/65536.0,1,-nbitq), 
to_sfixed(7488.0/65536.0,1,-nbitq), 
to_sfixed(2545.0/65536.0,1,-nbitq), 
to_sfixed(-1581.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-6566.0/65536.0,1,-nbitq), 
to_sfixed(-2508.0/65536.0,1,-nbitq), 
to_sfixed(-772.0/65536.0,1,-nbitq), 
to_sfixed(8060.0/65536.0,1,-nbitq), 
to_sfixed(11515.0/65536.0,1,-nbitq), 
to_sfixed(-13836.0/65536.0,1,-nbitq), 
to_sfixed(-807.0/65536.0,1,-nbitq), 
to_sfixed(7740.0/65536.0,1,-nbitq), 
to_sfixed(-127.0/65536.0,1,-nbitq), 
to_sfixed(-1057.0/65536.0,1,-nbitq), 
to_sfixed(5236.0/65536.0,1,-nbitq), 
to_sfixed(22150.0/65536.0,1,-nbitq), 
to_sfixed(-867.0/65536.0,1,-nbitq), 
to_sfixed(-8747.0/65536.0,1,-nbitq), 
to_sfixed(-5368.0/65536.0,1,-nbitq), 
to_sfixed(1670.0/65536.0,1,-nbitq), 
to_sfixed(1379.0/65536.0,1,-nbitq), 
to_sfixed(-1528.0/65536.0,1,-nbitq), 
to_sfixed(-9870.0/65536.0,1,-nbitq), 
to_sfixed(-1212.0/65536.0,1,-nbitq), 
to_sfixed(-4884.0/65536.0,1,-nbitq), 
to_sfixed(-10711.0/65536.0,1,-nbitq), 
to_sfixed(-9555.0/65536.0,1,-nbitq), 
to_sfixed(-4882.0/65536.0,1,-nbitq), 
to_sfixed(-1914.0/65536.0,1,-nbitq), 
to_sfixed(3899.0/65536.0,1,-nbitq), 
to_sfixed(9513.0/65536.0,1,-nbitq), 
to_sfixed(3376.0/65536.0,1,-nbitq), 
to_sfixed(6939.0/65536.0,1,-nbitq), 
to_sfixed(2885.0/65536.0,1,-nbitq), 
to_sfixed(-7526.0/65536.0,1,-nbitq), 
to_sfixed(14671.0/65536.0,1,-nbitq), 
to_sfixed(1645.0/65536.0,1,-nbitq), 
to_sfixed(-5637.0/65536.0,1,-nbitq), 
to_sfixed(-1144.0/65536.0,1,-nbitq), 
to_sfixed(1139.0/65536.0,1,-nbitq), 
to_sfixed(-6878.0/65536.0,1,-nbitq), 
to_sfixed(-3012.0/65536.0,1,-nbitq), 
to_sfixed(23151.0/65536.0,1,-nbitq), 
to_sfixed(-233.0/65536.0,1,-nbitq), 
to_sfixed(-3066.0/65536.0,1,-nbitq), 
to_sfixed(-3027.0/65536.0,1,-nbitq), 
to_sfixed(1626.0/65536.0,1,-nbitq), 
to_sfixed(-13182.0/65536.0,1,-nbitq), 
to_sfixed(3096.0/65536.0,1,-nbitq), 
to_sfixed(13189.0/65536.0,1,-nbitq), 
to_sfixed(556.0/65536.0,1,-nbitq), 
to_sfixed(-4899.0/65536.0,1,-nbitq), 
to_sfixed(1479.0/65536.0,1,-nbitq), 
to_sfixed(571.0/65536.0,1,-nbitq), 
to_sfixed(-1518.0/65536.0,1,-nbitq), 
to_sfixed(5433.0/65536.0,1,-nbitq), 
to_sfixed(-3626.0/65536.0,1,-nbitq), 
to_sfixed(-6503.0/65536.0,1,-nbitq), 
to_sfixed(659.0/65536.0,1,-nbitq), 
to_sfixed(3543.0/65536.0,1,-nbitq), 
to_sfixed(3437.0/65536.0,1,-nbitq), 
to_sfixed(801.0/65536.0,1,-nbitq), 
to_sfixed(-1899.0/65536.0,1,-nbitq), 
to_sfixed(10876.0/65536.0,1,-nbitq), 
to_sfixed(-4514.0/65536.0,1,-nbitq), 
to_sfixed(-2586.0/65536.0,1,-nbitq), 
to_sfixed(36.0/65536.0,1,-nbitq), 
to_sfixed(329.0/65536.0,1,-nbitq), 
to_sfixed(-12894.0/65536.0,1,-nbitq), 
to_sfixed(-7190.0/65536.0,1,-nbitq), 
to_sfixed(-5985.0/65536.0,1,-nbitq), 
to_sfixed(-8874.0/65536.0,1,-nbitq), 
to_sfixed(-15569.0/65536.0,1,-nbitq), 
to_sfixed(5029.0/65536.0,1,-nbitq), 
to_sfixed(-4903.0/65536.0,1,-nbitq), 
to_sfixed(10980.0/65536.0,1,-nbitq), 
to_sfixed(-12750.0/65536.0,1,-nbitq), 
to_sfixed(554.0/65536.0,1,-nbitq), 
to_sfixed(75.0/65536.0,1,-nbitq), 
to_sfixed(-13896.0/65536.0,1,-nbitq), 
to_sfixed(-4249.0/65536.0,1,-nbitq), 
to_sfixed(2421.0/65536.0,1,-nbitq), 
to_sfixed(2071.0/65536.0,1,-nbitq), 
to_sfixed(3283.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-7992.0/65536.0,1,-nbitq), 
to_sfixed(-6779.0/65536.0,1,-nbitq), 
to_sfixed(6353.0/65536.0,1,-nbitq), 
to_sfixed(6278.0/65536.0,1,-nbitq), 
to_sfixed(-2366.0/65536.0,1,-nbitq), 
to_sfixed(-2667.0/65536.0,1,-nbitq), 
to_sfixed(4680.0/65536.0,1,-nbitq), 
to_sfixed(9494.0/65536.0,1,-nbitq), 
to_sfixed(-2245.0/65536.0,1,-nbitq), 
to_sfixed(-2047.0/65536.0,1,-nbitq), 
to_sfixed(925.0/65536.0,1,-nbitq), 
to_sfixed(22618.0/65536.0,1,-nbitq), 
to_sfixed(-1465.0/65536.0,1,-nbitq), 
to_sfixed(-6291.0/65536.0,1,-nbitq), 
to_sfixed(1874.0/65536.0,1,-nbitq), 
to_sfixed(-407.0/65536.0,1,-nbitq), 
to_sfixed(-350.0/65536.0,1,-nbitq), 
to_sfixed(1705.0/65536.0,1,-nbitq), 
to_sfixed(-4955.0/65536.0,1,-nbitq), 
to_sfixed(414.0/65536.0,1,-nbitq), 
to_sfixed(-3064.0/65536.0,1,-nbitq), 
to_sfixed(-15597.0/65536.0,1,-nbitq), 
to_sfixed(-14635.0/65536.0,1,-nbitq), 
to_sfixed(-6974.0/65536.0,1,-nbitq), 
to_sfixed(-1331.0/65536.0,1,-nbitq), 
to_sfixed(1519.0/65536.0,1,-nbitq), 
to_sfixed(3084.0/65536.0,1,-nbitq), 
to_sfixed(4078.0/65536.0,1,-nbitq), 
to_sfixed(8455.0/65536.0,1,-nbitq), 
to_sfixed(8338.0/65536.0,1,-nbitq), 
to_sfixed(-1173.0/65536.0,1,-nbitq), 
to_sfixed(-150.0/65536.0,1,-nbitq), 
to_sfixed(-7319.0/65536.0,1,-nbitq), 
to_sfixed(-4424.0/65536.0,1,-nbitq), 
to_sfixed(-2953.0/65536.0,1,-nbitq), 
to_sfixed(904.0/65536.0,1,-nbitq), 
to_sfixed(-3956.0/65536.0,1,-nbitq), 
to_sfixed(9289.0/65536.0,1,-nbitq), 
to_sfixed(-1889.0/65536.0,1,-nbitq), 
to_sfixed(1146.0/65536.0,1,-nbitq), 
to_sfixed(-5260.0/65536.0,1,-nbitq), 
to_sfixed(1861.0/65536.0,1,-nbitq), 
to_sfixed(-4621.0/65536.0,1,-nbitq), 
to_sfixed(-13113.0/65536.0,1,-nbitq), 
to_sfixed(2778.0/65536.0,1,-nbitq), 
to_sfixed(18267.0/65536.0,1,-nbitq), 
to_sfixed(10.0/65536.0,1,-nbitq), 
to_sfixed(-6140.0/65536.0,1,-nbitq), 
to_sfixed(-180.0/65536.0,1,-nbitq), 
to_sfixed(-1771.0/65536.0,1,-nbitq), 
to_sfixed(-2786.0/65536.0,1,-nbitq), 
to_sfixed(5032.0/65536.0,1,-nbitq), 
to_sfixed(-969.0/65536.0,1,-nbitq), 
to_sfixed(-3261.0/65536.0,1,-nbitq), 
to_sfixed(-659.0/65536.0,1,-nbitq), 
to_sfixed(-16572.0/65536.0,1,-nbitq), 
to_sfixed(1619.0/65536.0,1,-nbitq), 
to_sfixed(3184.0/65536.0,1,-nbitq), 
to_sfixed(256.0/65536.0,1,-nbitq), 
to_sfixed(15136.0/65536.0,1,-nbitq), 
to_sfixed(-2459.0/65536.0,1,-nbitq), 
to_sfixed(-2348.0/65536.0,1,-nbitq), 
to_sfixed(2208.0/65536.0,1,-nbitq), 
to_sfixed(1772.0/65536.0,1,-nbitq), 
to_sfixed(-6580.0/65536.0,1,-nbitq), 
to_sfixed(4326.0/65536.0,1,-nbitq), 
to_sfixed(-535.0/65536.0,1,-nbitq), 
to_sfixed(-5331.0/65536.0,1,-nbitq), 
to_sfixed(-2870.0/65536.0,1,-nbitq), 
to_sfixed(13353.0/65536.0,1,-nbitq), 
to_sfixed(-709.0/65536.0,1,-nbitq), 
to_sfixed(14912.0/65536.0,1,-nbitq), 
to_sfixed(-12092.0/65536.0,1,-nbitq), 
to_sfixed(2184.0/65536.0,1,-nbitq), 
to_sfixed(-229.0/65536.0,1,-nbitq), 
to_sfixed(-3713.0/65536.0,1,-nbitq), 
to_sfixed(7218.0/65536.0,1,-nbitq), 
to_sfixed(7226.0/65536.0,1,-nbitq), 
to_sfixed(-1327.0/65536.0,1,-nbitq), 
to_sfixed(12133.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-7095.0/65536.0,1,-nbitq), 
to_sfixed(-2495.0/65536.0,1,-nbitq), 
to_sfixed(-2558.0/65536.0,1,-nbitq), 
to_sfixed(1200.0/65536.0,1,-nbitq), 
to_sfixed(-9309.0/65536.0,1,-nbitq), 
to_sfixed(15183.0/65536.0,1,-nbitq), 
to_sfixed(1743.0/65536.0,1,-nbitq), 
to_sfixed(14021.0/65536.0,1,-nbitq), 
to_sfixed(885.0/65536.0,1,-nbitq), 
to_sfixed(2915.0/65536.0,1,-nbitq), 
to_sfixed(735.0/65536.0,1,-nbitq), 
to_sfixed(10944.0/65536.0,1,-nbitq), 
to_sfixed(983.0/65536.0,1,-nbitq), 
to_sfixed(-1075.0/65536.0,1,-nbitq), 
to_sfixed(868.0/65536.0,1,-nbitq), 
to_sfixed(470.0/65536.0,1,-nbitq), 
to_sfixed(-2898.0/65536.0,1,-nbitq), 
to_sfixed(-877.0/65536.0,1,-nbitq), 
to_sfixed(589.0/65536.0,1,-nbitq), 
to_sfixed(-2264.0/65536.0,1,-nbitq), 
to_sfixed(-1744.0/65536.0,1,-nbitq), 
to_sfixed(-7443.0/65536.0,1,-nbitq), 
to_sfixed(-20705.0/65536.0,1,-nbitq), 
to_sfixed(-6013.0/65536.0,1,-nbitq), 
to_sfixed(440.0/65536.0,1,-nbitq), 
to_sfixed(-5775.0/65536.0,1,-nbitq), 
to_sfixed(-4556.0/65536.0,1,-nbitq), 
to_sfixed(4300.0/65536.0,1,-nbitq), 
to_sfixed(5060.0/65536.0,1,-nbitq), 
to_sfixed(3076.0/65536.0,1,-nbitq), 
to_sfixed(1695.0/65536.0,1,-nbitq), 
to_sfixed(-5861.0/65536.0,1,-nbitq), 
to_sfixed(-10727.0/65536.0,1,-nbitq), 
to_sfixed(-4717.0/65536.0,1,-nbitq), 
to_sfixed(-133.0/65536.0,1,-nbitq), 
to_sfixed(133.0/65536.0,1,-nbitq), 
to_sfixed(-714.0/65536.0,1,-nbitq), 
to_sfixed(7796.0/65536.0,1,-nbitq), 
to_sfixed(-8058.0/65536.0,1,-nbitq), 
to_sfixed(1982.0/65536.0,1,-nbitq), 
to_sfixed(2134.0/65536.0,1,-nbitq), 
to_sfixed(1946.0/65536.0,1,-nbitq), 
to_sfixed(-744.0/65536.0,1,-nbitq), 
to_sfixed(-9577.0/65536.0,1,-nbitq), 
to_sfixed(-1711.0/65536.0,1,-nbitq), 
to_sfixed(-731.0/65536.0,1,-nbitq), 
to_sfixed(-4780.0/65536.0,1,-nbitq), 
to_sfixed(2296.0/65536.0,1,-nbitq), 
to_sfixed(458.0/65536.0,1,-nbitq), 
to_sfixed(101.0/65536.0,1,-nbitq), 
to_sfixed(3042.0/65536.0,1,-nbitq), 
to_sfixed(-3674.0/65536.0,1,-nbitq), 
to_sfixed(479.0/65536.0,1,-nbitq), 
to_sfixed(-9921.0/65536.0,1,-nbitq), 
to_sfixed(5895.0/65536.0,1,-nbitq), 
to_sfixed(-22380.0/65536.0,1,-nbitq), 
to_sfixed(335.0/65536.0,1,-nbitq), 
to_sfixed(-4560.0/65536.0,1,-nbitq), 
to_sfixed(1252.0/65536.0,1,-nbitq), 
to_sfixed(5557.0/65536.0,1,-nbitq), 
to_sfixed(120.0/65536.0,1,-nbitq), 
to_sfixed(-920.0/65536.0,1,-nbitq), 
to_sfixed(337.0/65536.0,1,-nbitq), 
to_sfixed(652.0/65536.0,1,-nbitq), 
to_sfixed(-9402.0/65536.0,1,-nbitq), 
to_sfixed(2037.0/65536.0,1,-nbitq), 
to_sfixed(1855.0/65536.0,1,-nbitq), 
to_sfixed(-2485.0/65536.0,1,-nbitq), 
to_sfixed(-2314.0/65536.0,1,-nbitq), 
to_sfixed(16150.0/65536.0,1,-nbitq), 
to_sfixed(1266.0/65536.0,1,-nbitq), 
to_sfixed(9669.0/65536.0,1,-nbitq), 
to_sfixed(8720.0/65536.0,1,-nbitq), 
to_sfixed(-2904.0/65536.0,1,-nbitq), 
to_sfixed(1200.0/65536.0,1,-nbitq), 
to_sfixed(1293.0/65536.0,1,-nbitq), 
to_sfixed(-5344.0/65536.0,1,-nbitq), 
to_sfixed(7898.0/65536.0,1,-nbitq), 
to_sfixed(-2102.0/65536.0,1,-nbitq), 
to_sfixed(12635.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-7731.0/65536.0,1,-nbitq), 
to_sfixed(-1887.0/65536.0,1,-nbitq), 
to_sfixed(1975.0/65536.0,1,-nbitq), 
to_sfixed(9340.0/65536.0,1,-nbitq), 
to_sfixed(-8599.0/65536.0,1,-nbitq), 
to_sfixed(18420.0/65536.0,1,-nbitq), 
to_sfixed(266.0/65536.0,1,-nbitq), 
to_sfixed(12207.0/65536.0,1,-nbitq), 
to_sfixed(1879.0/65536.0,1,-nbitq), 
to_sfixed(1175.0/65536.0,1,-nbitq), 
to_sfixed(2149.0/65536.0,1,-nbitq), 
to_sfixed(-1612.0/65536.0,1,-nbitq), 
to_sfixed(1810.0/65536.0,1,-nbitq), 
to_sfixed(3967.0/65536.0,1,-nbitq), 
to_sfixed(-2954.0/65536.0,1,-nbitq), 
to_sfixed(-2928.0/65536.0,1,-nbitq), 
to_sfixed(-2072.0/65536.0,1,-nbitq), 
to_sfixed(-2444.0/65536.0,1,-nbitq), 
to_sfixed(2079.0/65536.0,1,-nbitq), 
to_sfixed(-577.0/65536.0,1,-nbitq), 
to_sfixed(301.0/65536.0,1,-nbitq), 
to_sfixed(-240.0/65536.0,1,-nbitq), 
to_sfixed(-21682.0/65536.0,1,-nbitq), 
to_sfixed(-1266.0/65536.0,1,-nbitq), 
to_sfixed(770.0/65536.0,1,-nbitq), 
to_sfixed(1287.0/65536.0,1,-nbitq), 
to_sfixed(150.0/65536.0,1,-nbitq), 
to_sfixed(689.0/65536.0,1,-nbitq), 
to_sfixed(11163.0/65536.0,1,-nbitq), 
to_sfixed(925.0/65536.0,1,-nbitq), 
to_sfixed(2040.0/65536.0,1,-nbitq), 
to_sfixed(1947.0/65536.0,1,-nbitq), 
to_sfixed(-8333.0/65536.0,1,-nbitq), 
to_sfixed(200.0/65536.0,1,-nbitq), 
to_sfixed(1022.0/65536.0,1,-nbitq), 
to_sfixed(-595.0/65536.0,1,-nbitq), 
to_sfixed(-6584.0/65536.0,1,-nbitq), 
to_sfixed(-4192.0/65536.0,1,-nbitq), 
to_sfixed(-8488.0/65536.0,1,-nbitq), 
to_sfixed(-2489.0/65536.0,1,-nbitq), 
to_sfixed(10954.0/65536.0,1,-nbitq), 
to_sfixed(1216.0/65536.0,1,-nbitq), 
to_sfixed(7836.0/65536.0,1,-nbitq), 
to_sfixed(-5172.0/65536.0,1,-nbitq), 
to_sfixed(-1933.0/65536.0,1,-nbitq), 
to_sfixed(-13742.0/65536.0,1,-nbitq), 
to_sfixed(-1947.0/65536.0,1,-nbitq), 
to_sfixed(11545.0/65536.0,1,-nbitq), 
to_sfixed(-1383.0/65536.0,1,-nbitq), 
to_sfixed(2005.0/65536.0,1,-nbitq), 
to_sfixed(832.0/65536.0,1,-nbitq), 
to_sfixed(-6154.0/65536.0,1,-nbitq), 
to_sfixed(-220.0/65536.0,1,-nbitq), 
to_sfixed(-1731.0/65536.0,1,-nbitq), 
to_sfixed(13851.0/65536.0,1,-nbitq), 
to_sfixed(-13901.0/65536.0,1,-nbitq), 
to_sfixed(-3397.0/65536.0,1,-nbitq), 
to_sfixed(-4984.0/65536.0,1,-nbitq), 
to_sfixed(-778.0/65536.0,1,-nbitq), 
to_sfixed(4645.0/65536.0,1,-nbitq), 
to_sfixed(-292.0/65536.0,1,-nbitq), 
to_sfixed(-1196.0/65536.0,1,-nbitq), 
to_sfixed(3085.0/65536.0,1,-nbitq), 
to_sfixed(823.0/65536.0,1,-nbitq), 
to_sfixed(-5036.0/65536.0,1,-nbitq), 
to_sfixed(6319.0/65536.0,1,-nbitq), 
to_sfixed(-2111.0/65536.0,1,-nbitq), 
to_sfixed(-4905.0/65536.0,1,-nbitq), 
to_sfixed(-10295.0/65536.0,1,-nbitq), 
to_sfixed(13989.0/65536.0,1,-nbitq), 
to_sfixed(6095.0/65536.0,1,-nbitq), 
to_sfixed(688.0/65536.0,1,-nbitq), 
to_sfixed(18192.0/65536.0,1,-nbitq), 
to_sfixed(2108.0/65536.0,1,-nbitq), 
to_sfixed(1789.0/65536.0,1,-nbitq), 
to_sfixed(2617.0/65536.0,1,-nbitq), 
to_sfixed(-15465.0/65536.0,1,-nbitq), 
to_sfixed(-4577.0/65536.0,1,-nbitq), 
to_sfixed(-671.0/65536.0,1,-nbitq), 
to_sfixed(8132.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-166.0/65536.0,1,-nbitq), 
to_sfixed(1387.0/65536.0,1,-nbitq), 
to_sfixed(-534.0/65536.0,1,-nbitq), 
to_sfixed(7275.0/65536.0,1,-nbitq), 
to_sfixed(-6268.0/65536.0,1,-nbitq), 
to_sfixed(20276.0/65536.0,1,-nbitq), 
to_sfixed(-941.0/65536.0,1,-nbitq), 
to_sfixed(1839.0/65536.0,1,-nbitq), 
to_sfixed(3455.0/65536.0,1,-nbitq), 
to_sfixed(-1132.0/65536.0,1,-nbitq), 
to_sfixed(1003.0/65536.0,1,-nbitq), 
to_sfixed(8257.0/65536.0,1,-nbitq), 
to_sfixed(2754.0/65536.0,1,-nbitq), 
to_sfixed(1554.0/65536.0,1,-nbitq), 
to_sfixed(2112.0/65536.0,1,-nbitq), 
to_sfixed(732.0/65536.0,1,-nbitq), 
to_sfixed(-1571.0/65536.0,1,-nbitq), 
to_sfixed(1387.0/65536.0,1,-nbitq), 
to_sfixed(-1275.0/65536.0,1,-nbitq), 
to_sfixed(-2406.0/65536.0,1,-nbitq), 
to_sfixed(3774.0/65536.0,1,-nbitq), 
to_sfixed(-3131.0/65536.0,1,-nbitq), 
to_sfixed(-20866.0/65536.0,1,-nbitq), 
to_sfixed(-7183.0/65536.0,1,-nbitq), 
to_sfixed(-3121.0/65536.0,1,-nbitq), 
to_sfixed(8423.0/65536.0,1,-nbitq), 
to_sfixed(-2527.0/65536.0,1,-nbitq), 
to_sfixed(550.0/65536.0,1,-nbitq), 
to_sfixed(10800.0/65536.0,1,-nbitq), 
to_sfixed(2438.0/65536.0,1,-nbitq), 
to_sfixed(-639.0/65536.0,1,-nbitq), 
to_sfixed(-3536.0/65536.0,1,-nbitq), 
to_sfixed(-12744.0/65536.0,1,-nbitq), 
to_sfixed(-4889.0/65536.0,1,-nbitq), 
to_sfixed(403.0/65536.0,1,-nbitq), 
to_sfixed(-3232.0/65536.0,1,-nbitq), 
to_sfixed(-3487.0/65536.0,1,-nbitq), 
to_sfixed(-6528.0/65536.0,1,-nbitq), 
to_sfixed(-2939.0/65536.0,1,-nbitq), 
to_sfixed(-1937.0/65536.0,1,-nbitq), 
to_sfixed(11218.0/65536.0,1,-nbitq), 
to_sfixed(-964.0/65536.0,1,-nbitq), 
to_sfixed(8898.0/65536.0,1,-nbitq), 
to_sfixed(-4233.0/65536.0,1,-nbitq), 
to_sfixed(3038.0/65536.0,1,-nbitq), 
to_sfixed(-15094.0/65536.0,1,-nbitq), 
to_sfixed(-162.0/65536.0,1,-nbitq), 
to_sfixed(8223.0/65536.0,1,-nbitq), 
to_sfixed(2944.0/65536.0,1,-nbitq), 
to_sfixed(-510.0/65536.0,1,-nbitq), 
to_sfixed(-1351.0/65536.0,1,-nbitq), 
to_sfixed(-5713.0/65536.0,1,-nbitq), 
to_sfixed(4974.0/65536.0,1,-nbitq), 
to_sfixed(3674.0/65536.0,1,-nbitq), 
to_sfixed(10986.0/65536.0,1,-nbitq), 
to_sfixed(-7673.0/65536.0,1,-nbitq), 
to_sfixed(-3713.0/65536.0,1,-nbitq), 
to_sfixed(-1072.0/65536.0,1,-nbitq), 
to_sfixed(-1589.0/65536.0,1,-nbitq), 
to_sfixed(4951.0/65536.0,1,-nbitq), 
to_sfixed(-2142.0/65536.0,1,-nbitq), 
to_sfixed(114.0/65536.0,1,-nbitq), 
to_sfixed(2371.0/65536.0,1,-nbitq), 
to_sfixed(-602.0/65536.0,1,-nbitq), 
to_sfixed(-2007.0/65536.0,1,-nbitq), 
to_sfixed(1841.0/65536.0,1,-nbitq), 
to_sfixed(-4242.0/65536.0,1,-nbitq), 
to_sfixed(-1623.0/65536.0,1,-nbitq), 
to_sfixed(516.0/65536.0,1,-nbitq), 
to_sfixed(11646.0/65536.0,1,-nbitq), 
to_sfixed(9956.0/65536.0,1,-nbitq), 
to_sfixed(-3784.0/65536.0,1,-nbitq), 
to_sfixed(13871.0/65536.0,1,-nbitq), 
to_sfixed(1403.0/65536.0,1,-nbitq), 
to_sfixed(2649.0/65536.0,1,-nbitq), 
to_sfixed(4342.0/65536.0,1,-nbitq), 
to_sfixed(-10271.0/65536.0,1,-nbitq), 
to_sfixed(-15575.0/65536.0,1,-nbitq), 
to_sfixed(808.0/65536.0,1,-nbitq), 
to_sfixed(4154.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5057.0/65536.0,1,-nbitq), 
to_sfixed(2970.0/65536.0,1,-nbitq), 
to_sfixed(-6909.0/65536.0,1,-nbitq), 
to_sfixed(5613.0/65536.0,1,-nbitq), 
to_sfixed(1441.0/65536.0,1,-nbitq), 
to_sfixed(13429.0/65536.0,1,-nbitq), 
to_sfixed(1695.0/65536.0,1,-nbitq), 
to_sfixed(6822.0/65536.0,1,-nbitq), 
to_sfixed(4741.0/65536.0,1,-nbitq), 
to_sfixed(2326.0/65536.0,1,-nbitq), 
to_sfixed(1329.0/65536.0,1,-nbitq), 
to_sfixed(9138.0/65536.0,1,-nbitq), 
to_sfixed(-15.0/65536.0,1,-nbitq), 
to_sfixed(3102.0/65536.0,1,-nbitq), 
to_sfixed(-276.0/65536.0,1,-nbitq), 
to_sfixed(457.0/65536.0,1,-nbitq), 
to_sfixed(-311.0/65536.0,1,-nbitq), 
to_sfixed(-591.0/65536.0,1,-nbitq), 
to_sfixed(-3013.0/65536.0,1,-nbitq), 
to_sfixed(-2444.0/65536.0,1,-nbitq), 
to_sfixed(2532.0/65536.0,1,-nbitq), 
to_sfixed(2721.0/65536.0,1,-nbitq), 
to_sfixed(-9746.0/65536.0,1,-nbitq), 
to_sfixed(-3162.0/65536.0,1,-nbitq), 
to_sfixed(-1775.0/65536.0,1,-nbitq), 
to_sfixed(8095.0/65536.0,1,-nbitq), 
to_sfixed(-3085.0/65536.0,1,-nbitq), 
to_sfixed(2117.0/65536.0,1,-nbitq), 
to_sfixed(11893.0/65536.0,1,-nbitq), 
to_sfixed(-1060.0/65536.0,1,-nbitq), 
to_sfixed(1727.0/65536.0,1,-nbitq), 
to_sfixed(-10493.0/65536.0,1,-nbitq), 
to_sfixed(-8425.0/65536.0,1,-nbitq), 
to_sfixed(2668.0/65536.0,1,-nbitq), 
to_sfixed(-1100.0/65536.0,1,-nbitq), 
to_sfixed(1824.0/65536.0,1,-nbitq), 
to_sfixed(-5218.0/65536.0,1,-nbitq), 
to_sfixed(-6132.0/65536.0,1,-nbitq), 
to_sfixed(-4227.0/65536.0,1,-nbitq), 
to_sfixed(2684.0/65536.0,1,-nbitq), 
to_sfixed(11878.0/65536.0,1,-nbitq), 
to_sfixed(-309.0/65536.0,1,-nbitq), 
to_sfixed(3076.0/65536.0,1,-nbitq), 
to_sfixed(-1617.0/65536.0,1,-nbitq), 
to_sfixed(-1331.0/65536.0,1,-nbitq), 
to_sfixed(-4654.0/65536.0,1,-nbitq), 
to_sfixed(-1471.0/65536.0,1,-nbitq), 
to_sfixed(5759.0/65536.0,1,-nbitq), 
to_sfixed(-1199.0/65536.0,1,-nbitq), 
to_sfixed(523.0/65536.0,1,-nbitq), 
to_sfixed(2693.0/65536.0,1,-nbitq), 
to_sfixed(-151.0/65536.0,1,-nbitq), 
to_sfixed(9217.0/65536.0,1,-nbitq), 
to_sfixed(6493.0/65536.0,1,-nbitq), 
to_sfixed(3785.0/65536.0,1,-nbitq), 
to_sfixed(-10288.0/65536.0,1,-nbitq), 
to_sfixed(-370.0/65536.0,1,-nbitq), 
to_sfixed(1490.0/65536.0,1,-nbitq), 
to_sfixed(1130.0/65536.0,1,-nbitq), 
to_sfixed(4954.0/65536.0,1,-nbitq), 
to_sfixed(-650.0/65536.0,1,-nbitq), 
to_sfixed(867.0/65536.0,1,-nbitq), 
to_sfixed(1079.0/65536.0,1,-nbitq), 
to_sfixed(-748.0/65536.0,1,-nbitq), 
to_sfixed(-5056.0/65536.0,1,-nbitq), 
to_sfixed(-6354.0/65536.0,1,-nbitq), 
to_sfixed(-729.0/65536.0,1,-nbitq), 
to_sfixed(7179.0/65536.0,1,-nbitq), 
to_sfixed(-1104.0/65536.0,1,-nbitq), 
to_sfixed(5103.0/65536.0,1,-nbitq), 
to_sfixed(7504.0/65536.0,1,-nbitq), 
to_sfixed(-3944.0/65536.0,1,-nbitq), 
to_sfixed(11543.0/65536.0,1,-nbitq), 
to_sfixed(662.0/65536.0,1,-nbitq), 
to_sfixed(-551.0/65536.0,1,-nbitq), 
to_sfixed(348.0/65536.0,1,-nbitq), 
to_sfixed(-12540.0/65536.0,1,-nbitq), 
to_sfixed(-11829.0/65536.0,1,-nbitq), 
to_sfixed(-211.0/65536.0,1,-nbitq), 
to_sfixed(-5017.0/65536.0,1,-nbitq)  ), 
( to_sfixed(6958.0/65536.0,1,-nbitq), 
to_sfixed(33.0/65536.0,1,-nbitq), 
to_sfixed(-5216.0/65536.0,1,-nbitq), 
to_sfixed(109.0/65536.0,1,-nbitq), 
to_sfixed(1667.0/65536.0,1,-nbitq), 
to_sfixed(10956.0/65536.0,1,-nbitq), 
to_sfixed(-926.0/65536.0,1,-nbitq), 
to_sfixed(3571.0/65536.0,1,-nbitq), 
to_sfixed(-504.0/65536.0,1,-nbitq), 
to_sfixed(1016.0/65536.0,1,-nbitq), 
to_sfixed(3518.0/65536.0,1,-nbitq), 
to_sfixed(-718.0/65536.0,1,-nbitq), 
to_sfixed(681.0/65536.0,1,-nbitq), 
to_sfixed(4004.0/65536.0,1,-nbitq), 
to_sfixed(-401.0/65536.0,1,-nbitq), 
to_sfixed(3311.0/65536.0,1,-nbitq), 
to_sfixed(-25.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(3893.0/65536.0,1,-nbitq), 
to_sfixed(683.0/65536.0,1,-nbitq), 
to_sfixed(3365.0/65536.0,1,-nbitq), 
to_sfixed(-2458.0/65536.0,1,-nbitq), 
to_sfixed(-10355.0/65536.0,1,-nbitq), 
to_sfixed(-2369.0/65536.0,1,-nbitq), 
to_sfixed(2982.0/65536.0,1,-nbitq), 
to_sfixed(12332.0/65536.0,1,-nbitq), 
to_sfixed(-628.0/65536.0,1,-nbitq), 
to_sfixed(-1703.0/65536.0,1,-nbitq), 
to_sfixed(9346.0/65536.0,1,-nbitq), 
to_sfixed(-858.0/65536.0,1,-nbitq), 
to_sfixed(6108.0/65536.0,1,-nbitq), 
to_sfixed(-9072.0/65536.0,1,-nbitq), 
to_sfixed(159.0/65536.0,1,-nbitq), 
to_sfixed(12069.0/65536.0,1,-nbitq), 
to_sfixed(-2103.0/65536.0,1,-nbitq), 
to_sfixed(262.0/65536.0,1,-nbitq), 
to_sfixed(36.0/65536.0,1,-nbitq), 
to_sfixed(-5213.0/65536.0,1,-nbitq), 
to_sfixed(-3649.0/65536.0,1,-nbitq), 
to_sfixed(-92.0/65536.0,1,-nbitq), 
to_sfixed(6713.0/65536.0,1,-nbitq), 
to_sfixed(-2160.0/65536.0,1,-nbitq), 
to_sfixed(7498.0/65536.0,1,-nbitq), 
to_sfixed(1217.0/65536.0,1,-nbitq), 
to_sfixed(1931.0/65536.0,1,-nbitq), 
to_sfixed(361.0/65536.0,1,-nbitq), 
to_sfixed(2076.0/65536.0,1,-nbitq), 
to_sfixed(-1421.0/65536.0,1,-nbitq), 
to_sfixed(666.0/65536.0,1,-nbitq), 
to_sfixed(1622.0/65536.0,1,-nbitq), 
to_sfixed(-2200.0/65536.0,1,-nbitq), 
to_sfixed(8501.0/65536.0,1,-nbitq), 
to_sfixed(9192.0/65536.0,1,-nbitq), 
to_sfixed(4298.0/65536.0,1,-nbitq), 
to_sfixed(3291.0/65536.0,1,-nbitq), 
to_sfixed(2116.0/65536.0,1,-nbitq), 
to_sfixed(-972.0/65536.0,1,-nbitq), 
to_sfixed(1416.0/65536.0,1,-nbitq), 
to_sfixed(1855.0/65536.0,1,-nbitq), 
to_sfixed(-951.0/65536.0,1,-nbitq), 
to_sfixed(1164.0/65536.0,1,-nbitq), 
to_sfixed(-1841.0/65536.0,1,-nbitq), 
to_sfixed(2144.0/65536.0,1,-nbitq), 
to_sfixed(2022.0/65536.0,1,-nbitq), 
to_sfixed(6281.0/65536.0,1,-nbitq), 
to_sfixed(-1129.0/65536.0,1,-nbitq), 
to_sfixed(2635.0/65536.0,1,-nbitq), 
to_sfixed(7336.0/65536.0,1,-nbitq), 
to_sfixed(1705.0/65536.0,1,-nbitq), 
to_sfixed(-2870.0/65536.0,1,-nbitq), 
to_sfixed(7100.0/65536.0,1,-nbitq), 
to_sfixed(-2819.0/65536.0,1,-nbitq), 
to_sfixed(11348.0/65536.0,1,-nbitq), 
to_sfixed(-94.0/65536.0,1,-nbitq), 
to_sfixed(-2528.0/65536.0,1,-nbitq), 
to_sfixed(4208.0/65536.0,1,-nbitq), 
to_sfixed(-9174.0/65536.0,1,-nbitq), 
to_sfixed(-10750.0/65536.0,1,-nbitq), 
to_sfixed(2208.0/65536.0,1,-nbitq), 
to_sfixed(-11469.0/65536.0,1,-nbitq)  ), 
( to_sfixed(807.0/65536.0,1,-nbitq), 
to_sfixed(5663.0/65536.0,1,-nbitq), 
to_sfixed(-4218.0/65536.0,1,-nbitq), 
to_sfixed(-191.0/65536.0,1,-nbitq), 
to_sfixed(1215.0/65536.0,1,-nbitq), 
to_sfixed(10205.0/65536.0,1,-nbitq), 
to_sfixed(-5149.0/65536.0,1,-nbitq), 
to_sfixed(1055.0/65536.0,1,-nbitq), 
to_sfixed(-4594.0/65536.0,1,-nbitq), 
to_sfixed(681.0/65536.0,1,-nbitq), 
to_sfixed(6023.0/65536.0,1,-nbitq), 
to_sfixed(-10290.0/65536.0,1,-nbitq), 
to_sfixed(-756.0/65536.0,1,-nbitq), 
to_sfixed(13046.0/65536.0,1,-nbitq), 
to_sfixed(-2303.0/65536.0,1,-nbitq), 
to_sfixed(-685.0/65536.0,1,-nbitq), 
to_sfixed(2475.0/65536.0,1,-nbitq), 
to_sfixed(5577.0/65536.0,1,-nbitq), 
to_sfixed(1854.0/65536.0,1,-nbitq), 
to_sfixed(-2827.0/65536.0,1,-nbitq), 
to_sfixed(5639.0/65536.0,1,-nbitq), 
to_sfixed(-14637.0/65536.0,1,-nbitq), 
to_sfixed(-749.0/65536.0,1,-nbitq), 
to_sfixed(-2743.0/65536.0,1,-nbitq), 
to_sfixed(-542.0/65536.0,1,-nbitq), 
to_sfixed(8298.0/65536.0,1,-nbitq), 
to_sfixed(-2204.0/65536.0,1,-nbitq), 
to_sfixed(997.0/65536.0,1,-nbitq), 
to_sfixed(4649.0/65536.0,1,-nbitq), 
to_sfixed(-660.0/65536.0,1,-nbitq), 
to_sfixed(6352.0/65536.0,1,-nbitq), 
to_sfixed(-8905.0/65536.0,1,-nbitq), 
to_sfixed(7650.0/65536.0,1,-nbitq), 
to_sfixed(17900.0/65536.0,1,-nbitq), 
to_sfixed(-13.0/65536.0,1,-nbitq), 
to_sfixed(-26.0/65536.0,1,-nbitq), 
to_sfixed(-7367.0/65536.0,1,-nbitq), 
to_sfixed(-3473.0/65536.0,1,-nbitq), 
to_sfixed(3253.0/65536.0,1,-nbitq), 
to_sfixed(-2144.0/65536.0,1,-nbitq), 
to_sfixed(5013.0/65536.0,1,-nbitq), 
to_sfixed(1693.0/65536.0,1,-nbitq), 
to_sfixed(10653.0/65536.0,1,-nbitq), 
to_sfixed(5336.0/65536.0,1,-nbitq), 
to_sfixed(2464.0/65536.0,1,-nbitq), 
to_sfixed(3504.0/65536.0,1,-nbitq), 
to_sfixed(1687.0/65536.0,1,-nbitq), 
to_sfixed(-2082.0/65536.0,1,-nbitq), 
to_sfixed(-1495.0/65536.0,1,-nbitq), 
to_sfixed(667.0/65536.0,1,-nbitq), 
to_sfixed(1613.0/65536.0,1,-nbitq), 
to_sfixed(4972.0/65536.0,1,-nbitq), 
to_sfixed(7512.0/65536.0,1,-nbitq), 
to_sfixed(2175.0/65536.0,1,-nbitq), 
to_sfixed(739.0/65536.0,1,-nbitq), 
to_sfixed(2348.0/65536.0,1,-nbitq), 
to_sfixed(-2341.0/65536.0,1,-nbitq), 
to_sfixed(4270.0/65536.0,1,-nbitq), 
to_sfixed(-2291.0/65536.0,1,-nbitq), 
to_sfixed(-1033.0/65536.0,1,-nbitq), 
to_sfixed(-848.0/65536.0,1,-nbitq), 
to_sfixed(1693.0/65536.0,1,-nbitq), 
to_sfixed(689.0/65536.0,1,-nbitq), 
to_sfixed(-703.0/65536.0,1,-nbitq), 
to_sfixed(4558.0/65536.0,1,-nbitq), 
to_sfixed(-1530.0/65536.0,1,-nbitq), 
to_sfixed(5132.0/65536.0,1,-nbitq), 
to_sfixed(7844.0/65536.0,1,-nbitq), 
to_sfixed(-2751.0/65536.0,1,-nbitq), 
to_sfixed(-1470.0/65536.0,1,-nbitq), 
to_sfixed(133.0/65536.0,1,-nbitq), 
to_sfixed(-4373.0/65536.0,1,-nbitq), 
to_sfixed(12233.0/65536.0,1,-nbitq), 
to_sfixed(-3211.0/65536.0,1,-nbitq), 
to_sfixed(1603.0/65536.0,1,-nbitq), 
to_sfixed(629.0/65536.0,1,-nbitq), 
to_sfixed(-5299.0/65536.0,1,-nbitq), 
to_sfixed(-1432.0/65536.0,1,-nbitq), 
to_sfixed(-1872.0/65536.0,1,-nbitq), 
to_sfixed(-10285.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5903.0/65536.0,1,-nbitq), 
to_sfixed(1336.0/65536.0,1,-nbitq), 
to_sfixed(-2226.0/65536.0,1,-nbitq), 
to_sfixed(4524.0/65536.0,1,-nbitq), 
to_sfixed(-3445.0/65536.0,1,-nbitq), 
to_sfixed(6150.0/65536.0,1,-nbitq), 
to_sfixed(-4118.0/65536.0,1,-nbitq), 
to_sfixed(10074.0/65536.0,1,-nbitq), 
to_sfixed(-6053.0/65536.0,1,-nbitq), 
to_sfixed(-2579.0/65536.0,1,-nbitq), 
to_sfixed(4368.0/65536.0,1,-nbitq), 
to_sfixed(-6327.0/65536.0,1,-nbitq), 
to_sfixed(2250.0/65536.0,1,-nbitq), 
to_sfixed(11334.0/65536.0,1,-nbitq), 
to_sfixed(-3794.0/65536.0,1,-nbitq), 
to_sfixed(1821.0/65536.0,1,-nbitq), 
to_sfixed(2332.0/65536.0,1,-nbitq), 
to_sfixed(13527.0/65536.0,1,-nbitq), 
to_sfixed(1302.0/65536.0,1,-nbitq), 
to_sfixed(-2288.0/65536.0,1,-nbitq), 
to_sfixed(3075.0/65536.0,1,-nbitq), 
to_sfixed(-12813.0/65536.0,1,-nbitq), 
to_sfixed(-8035.0/65536.0,1,-nbitq), 
to_sfixed(-1141.0/65536.0,1,-nbitq), 
to_sfixed(1484.0/65536.0,1,-nbitq), 
to_sfixed(11356.0/65536.0,1,-nbitq), 
to_sfixed(-1436.0/65536.0,1,-nbitq), 
to_sfixed(2246.0/65536.0,1,-nbitq), 
to_sfixed(4430.0/65536.0,1,-nbitq), 
to_sfixed(-2801.0/65536.0,1,-nbitq), 
to_sfixed(2092.0/65536.0,1,-nbitq), 
to_sfixed(-7811.0/65536.0,1,-nbitq), 
to_sfixed(9669.0/65536.0,1,-nbitq), 
to_sfixed(6826.0/65536.0,1,-nbitq), 
to_sfixed(-3012.0/65536.0,1,-nbitq), 
to_sfixed(-2160.0/65536.0,1,-nbitq), 
to_sfixed(-3765.0/65536.0,1,-nbitq), 
to_sfixed(2407.0/65536.0,1,-nbitq), 
to_sfixed(137.0/65536.0,1,-nbitq), 
to_sfixed(1985.0/65536.0,1,-nbitq), 
to_sfixed(4103.0/65536.0,1,-nbitq), 
to_sfixed(2417.0/65536.0,1,-nbitq), 
to_sfixed(11674.0/65536.0,1,-nbitq), 
to_sfixed(1845.0/65536.0,1,-nbitq), 
to_sfixed(1698.0/65536.0,1,-nbitq), 
to_sfixed(3283.0/65536.0,1,-nbitq), 
to_sfixed(-2374.0/65536.0,1,-nbitq), 
to_sfixed(-557.0/65536.0,1,-nbitq), 
to_sfixed(-1333.0/65536.0,1,-nbitq), 
to_sfixed(713.0/65536.0,1,-nbitq), 
to_sfixed(2800.0/65536.0,1,-nbitq), 
to_sfixed(632.0/65536.0,1,-nbitq), 
to_sfixed(6061.0/65536.0,1,-nbitq), 
to_sfixed(4753.0/65536.0,1,-nbitq), 
to_sfixed(-5052.0/65536.0,1,-nbitq), 
to_sfixed(-1754.0/65536.0,1,-nbitq), 
to_sfixed(-1239.0/65536.0,1,-nbitq), 
to_sfixed(2023.0/65536.0,1,-nbitq), 
to_sfixed(-2007.0/65536.0,1,-nbitq), 
to_sfixed(-2436.0/65536.0,1,-nbitq), 
to_sfixed(1548.0/65536.0,1,-nbitq), 
to_sfixed(2234.0/65536.0,1,-nbitq), 
to_sfixed(1351.0/65536.0,1,-nbitq), 
to_sfixed(2139.0/65536.0,1,-nbitq), 
to_sfixed(-3902.0/65536.0,1,-nbitq), 
to_sfixed(2804.0/65536.0,1,-nbitq), 
to_sfixed(-1471.0/65536.0,1,-nbitq), 
to_sfixed(5262.0/65536.0,1,-nbitq), 
to_sfixed(-3376.0/65536.0,1,-nbitq), 
to_sfixed(179.0/65536.0,1,-nbitq), 
to_sfixed(-1166.0/65536.0,1,-nbitq), 
to_sfixed(-4563.0/65536.0,1,-nbitq), 
to_sfixed(11786.0/65536.0,1,-nbitq), 
to_sfixed(2322.0/65536.0,1,-nbitq), 
to_sfixed(2008.0/65536.0,1,-nbitq), 
to_sfixed(2851.0/65536.0,1,-nbitq), 
to_sfixed(-2370.0/65536.0,1,-nbitq), 
to_sfixed(416.0/65536.0,1,-nbitq), 
to_sfixed(433.0/65536.0,1,-nbitq), 
to_sfixed(-11175.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3837.0/65536.0,1,-nbitq), 
to_sfixed(-2592.0/65536.0,1,-nbitq), 
to_sfixed(-2133.0/65536.0,1,-nbitq), 
to_sfixed(2467.0/65536.0,1,-nbitq), 
to_sfixed(2995.0/65536.0,1,-nbitq), 
to_sfixed(7436.0/65536.0,1,-nbitq), 
to_sfixed(-967.0/65536.0,1,-nbitq), 
to_sfixed(8574.0/65536.0,1,-nbitq), 
to_sfixed(-2961.0/65536.0,1,-nbitq), 
to_sfixed(548.0/65536.0,1,-nbitq), 
to_sfixed(5257.0/65536.0,1,-nbitq), 
to_sfixed(-6560.0/65536.0,1,-nbitq), 
to_sfixed(-260.0/65536.0,1,-nbitq), 
to_sfixed(7029.0/65536.0,1,-nbitq), 
to_sfixed(891.0/65536.0,1,-nbitq), 
to_sfixed(939.0/65536.0,1,-nbitq), 
to_sfixed(2095.0/65536.0,1,-nbitq), 
to_sfixed(7605.0/65536.0,1,-nbitq), 
to_sfixed(1457.0/65536.0,1,-nbitq), 
to_sfixed(1065.0/65536.0,1,-nbitq), 
to_sfixed(1520.0/65536.0,1,-nbitq), 
to_sfixed(-7504.0/65536.0,1,-nbitq), 
to_sfixed(-1869.0/65536.0,1,-nbitq), 
to_sfixed(2296.0/65536.0,1,-nbitq), 
to_sfixed(1414.0/65536.0,1,-nbitq), 
to_sfixed(8983.0/65536.0,1,-nbitq), 
to_sfixed(-1095.0/65536.0,1,-nbitq), 
to_sfixed(1012.0/65536.0,1,-nbitq), 
to_sfixed(4533.0/65536.0,1,-nbitq), 
to_sfixed(1909.0/65536.0,1,-nbitq), 
to_sfixed(289.0/65536.0,1,-nbitq), 
to_sfixed(-7257.0/65536.0,1,-nbitq), 
to_sfixed(10656.0/65536.0,1,-nbitq), 
to_sfixed(-2312.0/65536.0,1,-nbitq), 
to_sfixed(-1766.0/65536.0,1,-nbitq), 
to_sfixed(-1254.0/65536.0,1,-nbitq), 
to_sfixed(-3145.0/65536.0,1,-nbitq), 
to_sfixed(-1298.0/65536.0,1,-nbitq), 
to_sfixed(-2477.0/65536.0,1,-nbitq), 
to_sfixed(-171.0/65536.0,1,-nbitq), 
to_sfixed(280.0/65536.0,1,-nbitq), 
to_sfixed(1745.0/65536.0,1,-nbitq), 
to_sfixed(7066.0/65536.0,1,-nbitq), 
to_sfixed(6339.0/65536.0,1,-nbitq), 
to_sfixed(1748.0/65536.0,1,-nbitq), 
to_sfixed(-3722.0/65536.0,1,-nbitq), 
to_sfixed(-1050.0/65536.0,1,-nbitq), 
to_sfixed(-1141.0/65536.0,1,-nbitq), 
to_sfixed(2676.0/65536.0,1,-nbitq), 
to_sfixed(426.0/65536.0,1,-nbitq), 
to_sfixed(-109.0/65536.0,1,-nbitq), 
to_sfixed(6459.0/65536.0,1,-nbitq), 
to_sfixed(9773.0/65536.0,1,-nbitq), 
to_sfixed(6782.0/65536.0,1,-nbitq), 
to_sfixed(-1527.0/65536.0,1,-nbitq), 
to_sfixed(471.0/65536.0,1,-nbitq), 
to_sfixed(1999.0/65536.0,1,-nbitq), 
to_sfixed(2585.0/65536.0,1,-nbitq), 
to_sfixed(-473.0/65536.0,1,-nbitq), 
to_sfixed(-3883.0/65536.0,1,-nbitq), 
to_sfixed(-5877.0/65536.0,1,-nbitq), 
to_sfixed(-924.0/65536.0,1,-nbitq), 
to_sfixed(-2758.0/65536.0,1,-nbitq), 
to_sfixed(-433.0/65536.0,1,-nbitq), 
to_sfixed(-4481.0/65536.0,1,-nbitq), 
to_sfixed(7458.0/65536.0,1,-nbitq), 
to_sfixed(7207.0/65536.0,1,-nbitq), 
to_sfixed(3807.0/65536.0,1,-nbitq), 
to_sfixed(-5824.0/65536.0,1,-nbitq), 
to_sfixed(-8857.0/65536.0,1,-nbitq), 
to_sfixed(2775.0/65536.0,1,-nbitq), 
to_sfixed(-4193.0/65536.0,1,-nbitq), 
to_sfixed(6299.0/65536.0,1,-nbitq), 
to_sfixed(-2328.0/65536.0,1,-nbitq), 
to_sfixed(-2750.0/65536.0,1,-nbitq), 
to_sfixed(1338.0/65536.0,1,-nbitq), 
to_sfixed(-4876.0/65536.0,1,-nbitq), 
to_sfixed(261.0/65536.0,1,-nbitq), 
to_sfixed(-1781.0/65536.0,1,-nbitq), 
to_sfixed(-9505.0/65536.0,1,-nbitq)  ), 
( to_sfixed(8064.0/65536.0,1,-nbitq), 
to_sfixed(1076.0/65536.0,1,-nbitq), 
to_sfixed(-2821.0/65536.0,1,-nbitq), 
to_sfixed(1113.0/65536.0,1,-nbitq), 
to_sfixed(2835.0/65536.0,1,-nbitq), 
to_sfixed(1980.0/65536.0,1,-nbitq), 
to_sfixed(1917.0/65536.0,1,-nbitq), 
to_sfixed(5435.0/65536.0,1,-nbitq), 
to_sfixed(-3810.0/65536.0,1,-nbitq), 
to_sfixed(1179.0/65536.0,1,-nbitq), 
to_sfixed(1785.0/65536.0,1,-nbitq), 
to_sfixed(-6653.0/65536.0,1,-nbitq), 
to_sfixed(2084.0/65536.0,1,-nbitq), 
to_sfixed(1658.0/65536.0,1,-nbitq), 
to_sfixed(4.0/65536.0,1,-nbitq), 
to_sfixed(1185.0/65536.0,1,-nbitq), 
to_sfixed(-714.0/65536.0,1,-nbitq), 
to_sfixed(4861.0/65536.0,1,-nbitq), 
to_sfixed(3167.0/65536.0,1,-nbitq), 
to_sfixed(-1715.0/65536.0,1,-nbitq), 
to_sfixed(64.0/65536.0,1,-nbitq), 
to_sfixed(-5136.0/65536.0,1,-nbitq), 
to_sfixed(-1936.0/65536.0,1,-nbitq), 
to_sfixed(1754.0/65536.0,1,-nbitq), 
to_sfixed(-785.0/65536.0,1,-nbitq), 
to_sfixed(3761.0/65536.0,1,-nbitq), 
to_sfixed(839.0/65536.0,1,-nbitq), 
to_sfixed(1426.0/65536.0,1,-nbitq), 
to_sfixed(5335.0/65536.0,1,-nbitq), 
to_sfixed(-1944.0/65536.0,1,-nbitq), 
to_sfixed(3581.0/65536.0,1,-nbitq), 
to_sfixed(-4302.0/65536.0,1,-nbitq), 
to_sfixed(5724.0/65536.0,1,-nbitq), 
to_sfixed(-2962.0/65536.0,1,-nbitq), 
to_sfixed(-3025.0/65536.0,1,-nbitq), 
to_sfixed(2461.0/65536.0,1,-nbitq), 
to_sfixed(792.0/65536.0,1,-nbitq), 
to_sfixed(3596.0/65536.0,1,-nbitq), 
to_sfixed(-2822.0/65536.0,1,-nbitq), 
to_sfixed(3370.0/65536.0,1,-nbitq), 
to_sfixed(2138.0/65536.0,1,-nbitq), 
to_sfixed(-700.0/65536.0,1,-nbitq), 
to_sfixed(3079.0/65536.0,1,-nbitq), 
to_sfixed(6492.0/65536.0,1,-nbitq), 
to_sfixed(2903.0/65536.0,1,-nbitq), 
to_sfixed(-2032.0/65536.0,1,-nbitq), 
to_sfixed(-3108.0/65536.0,1,-nbitq), 
to_sfixed(-4824.0/65536.0,1,-nbitq), 
to_sfixed(2264.0/65536.0,1,-nbitq), 
to_sfixed(2233.0/65536.0,1,-nbitq), 
to_sfixed(596.0/65536.0,1,-nbitq), 
to_sfixed(6832.0/65536.0,1,-nbitq), 
to_sfixed(6561.0/65536.0,1,-nbitq), 
to_sfixed(10656.0/65536.0,1,-nbitq), 
to_sfixed(-2302.0/65536.0,1,-nbitq), 
to_sfixed(1942.0/65536.0,1,-nbitq), 
to_sfixed(-1348.0/65536.0,1,-nbitq), 
to_sfixed(2096.0/65536.0,1,-nbitq), 
to_sfixed(-1579.0/65536.0,1,-nbitq), 
to_sfixed(-6898.0/65536.0,1,-nbitq), 
to_sfixed(-3430.0/65536.0,1,-nbitq), 
to_sfixed(505.0/65536.0,1,-nbitq), 
to_sfixed(-1523.0/65536.0,1,-nbitq), 
to_sfixed(-438.0/65536.0,1,-nbitq), 
to_sfixed(1258.0/65536.0,1,-nbitq), 
to_sfixed(4710.0/65536.0,1,-nbitq), 
to_sfixed(9653.0/65536.0,1,-nbitq), 
to_sfixed(7017.0/65536.0,1,-nbitq), 
to_sfixed(-191.0/65536.0,1,-nbitq), 
to_sfixed(-3311.0/65536.0,1,-nbitq), 
to_sfixed(5130.0/65536.0,1,-nbitq), 
to_sfixed(207.0/65536.0,1,-nbitq), 
to_sfixed(5462.0/65536.0,1,-nbitq), 
to_sfixed(-3242.0/65536.0,1,-nbitq), 
to_sfixed(211.0/65536.0,1,-nbitq), 
to_sfixed(1991.0/65536.0,1,-nbitq), 
to_sfixed(-3741.0/65536.0,1,-nbitq), 
to_sfixed(1214.0/65536.0,1,-nbitq), 
to_sfixed(-2351.0/65536.0,1,-nbitq), 
to_sfixed(-40.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4193.0/65536.0,1,-nbitq), 
to_sfixed(2585.0/65536.0,1,-nbitq), 
to_sfixed(-5269.0/65536.0,1,-nbitq), 
to_sfixed(549.0/65536.0,1,-nbitq), 
to_sfixed(331.0/65536.0,1,-nbitq), 
to_sfixed(-1016.0/65536.0,1,-nbitq), 
to_sfixed(1611.0/65536.0,1,-nbitq), 
to_sfixed(264.0/65536.0,1,-nbitq), 
to_sfixed(-1350.0/65536.0,1,-nbitq), 
to_sfixed(1324.0/65536.0,1,-nbitq), 
to_sfixed(-2666.0/65536.0,1,-nbitq), 
to_sfixed(657.0/65536.0,1,-nbitq), 
to_sfixed(2095.0/65536.0,1,-nbitq), 
to_sfixed(1455.0/65536.0,1,-nbitq), 
to_sfixed(-1361.0/65536.0,1,-nbitq), 
to_sfixed(-2140.0/65536.0,1,-nbitq), 
to_sfixed(2340.0/65536.0,1,-nbitq), 
to_sfixed(2587.0/65536.0,1,-nbitq), 
to_sfixed(-2072.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(3927.0/65536.0,1,-nbitq), 
to_sfixed(-2632.0/65536.0,1,-nbitq), 
to_sfixed(-2654.0/65536.0,1,-nbitq), 
to_sfixed(-997.0/65536.0,1,-nbitq), 
to_sfixed(-788.0/65536.0,1,-nbitq), 
to_sfixed(-376.0/65536.0,1,-nbitq), 
to_sfixed(-1407.0/65536.0,1,-nbitq), 
to_sfixed(-2755.0/65536.0,1,-nbitq), 
to_sfixed(2094.0/65536.0,1,-nbitq), 
to_sfixed(323.0/65536.0,1,-nbitq), 
to_sfixed(646.0/65536.0,1,-nbitq), 
to_sfixed(-1175.0/65536.0,1,-nbitq), 
to_sfixed(4719.0/65536.0,1,-nbitq), 
to_sfixed(-1341.0/65536.0,1,-nbitq), 
to_sfixed(778.0/65536.0,1,-nbitq), 
to_sfixed(-1369.0/65536.0,1,-nbitq), 
to_sfixed(1361.0/65536.0,1,-nbitq), 
to_sfixed(2448.0/65536.0,1,-nbitq), 
to_sfixed(-5049.0/65536.0,1,-nbitq), 
to_sfixed(-1212.0/65536.0,1,-nbitq), 
to_sfixed(175.0/65536.0,1,-nbitq), 
to_sfixed(-208.0/65536.0,1,-nbitq), 
to_sfixed(4242.0/65536.0,1,-nbitq), 
to_sfixed(5295.0/65536.0,1,-nbitq), 
to_sfixed(-1182.0/65536.0,1,-nbitq), 
to_sfixed(-3475.0/65536.0,1,-nbitq), 
to_sfixed(1206.0/65536.0,1,-nbitq), 
to_sfixed(-926.0/65536.0,1,-nbitq), 
to_sfixed(2145.0/65536.0,1,-nbitq), 
to_sfixed(867.0/65536.0,1,-nbitq), 
to_sfixed(-1069.0/65536.0,1,-nbitq), 
to_sfixed(3800.0/65536.0,1,-nbitq), 
to_sfixed(437.0/65536.0,1,-nbitq), 
to_sfixed(6144.0/65536.0,1,-nbitq), 
to_sfixed(-4236.0/65536.0,1,-nbitq), 
to_sfixed(2532.0/65536.0,1,-nbitq), 
to_sfixed(193.0/65536.0,1,-nbitq), 
to_sfixed(-54.0/65536.0,1,-nbitq), 
to_sfixed(31.0/65536.0,1,-nbitq), 
to_sfixed(-3684.0/65536.0,1,-nbitq), 
to_sfixed(-1394.0/65536.0,1,-nbitq), 
to_sfixed(2317.0/65536.0,1,-nbitq), 
to_sfixed(701.0/65536.0,1,-nbitq), 
to_sfixed(-1278.0/65536.0,1,-nbitq), 
to_sfixed(1059.0/65536.0,1,-nbitq), 
to_sfixed(681.0/65536.0,1,-nbitq), 
to_sfixed(2796.0/65536.0,1,-nbitq), 
to_sfixed(109.0/65536.0,1,-nbitq), 
to_sfixed(2401.0/65536.0,1,-nbitq), 
to_sfixed(1281.0/65536.0,1,-nbitq), 
to_sfixed(-1193.0/65536.0,1,-nbitq), 
to_sfixed(-171.0/65536.0,1,-nbitq), 
to_sfixed(6329.0/65536.0,1,-nbitq), 
to_sfixed(925.0/65536.0,1,-nbitq), 
to_sfixed(2612.0/65536.0,1,-nbitq), 
to_sfixed(1647.0/65536.0,1,-nbitq), 
to_sfixed(-2772.0/65536.0,1,-nbitq), 
to_sfixed(3718.0/65536.0,1,-nbitq), 
to_sfixed(2210.0/65536.0,1,-nbitq), 
to_sfixed(462.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1907.0/65536.0,1,-nbitq), 
to_sfixed(-2252.0/65536.0,1,-nbitq), 
to_sfixed(-1782.0/65536.0,1,-nbitq), 
to_sfixed(2772.0/65536.0,1,-nbitq), 
to_sfixed(-4575.0/65536.0,1,-nbitq), 
to_sfixed(-2446.0/65536.0,1,-nbitq), 
to_sfixed(-3183.0/65536.0,1,-nbitq), 
to_sfixed(2776.0/65536.0,1,-nbitq), 
to_sfixed(1226.0/65536.0,1,-nbitq), 
to_sfixed(1715.0/65536.0,1,-nbitq), 
to_sfixed(-460.0/65536.0,1,-nbitq), 
to_sfixed(-2732.0/65536.0,1,-nbitq), 
to_sfixed(2374.0/65536.0,1,-nbitq), 
to_sfixed(1129.0/65536.0,1,-nbitq), 
to_sfixed(3319.0/65536.0,1,-nbitq), 
to_sfixed(2360.0/65536.0,1,-nbitq), 
to_sfixed(1480.0/65536.0,1,-nbitq), 
to_sfixed(3770.0/65536.0,1,-nbitq), 
to_sfixed(2027.0/65536.0,1,-nbitq), 
to_sfixed(-737.0/65536.0,1,-nbitq), 
to_sfixed(737.0/65536.0,1,-nbitq), 
to_sfixed(3186.0/65536.0,1,-nbitq), 
to_sfixed(-3246.0/65536.0,1,-nbitq), 
to_sfixed(71.0/65536.0,1,-nbitq), 
to_sfixed(-993.0/65536.0,1,-nbitq), 
to_sfixed(-815.0/65536.0,1,-nbitq), 
to_sfixed(-1884.0/65536.0,1,-nbitq), 
to_sfixed(-2503.0/65536.0,1,-nbitq), 
to_sfixed(2714.0/65536.0,1,-nbitq), 
to_sfixed(-1304.0/65536.0,1,-nbitq), 
to_sfixed(315.0/65536.0,1,-nbitq), 
to_sfixed(2063.0/65536.0,1,-nbitq), 
to_sfixed(1660.0/65536.0,1,-nbitq), 
to_sfixed(-3947.0/65536.0,1,-nbitq), 
to_sfixed(-1426.0/65536.0,1,-nbitq), 
to_sfixed(1957.0/65536.0,1,-nbitq), 
to_sfixed(-4835.0/65536.0,1,-nbitq), 
to_sfixed(-2425.0/65536.0,1,-nbitq), 
to_sfixed(-3402.0/65536.0,1,-nbitq), 
to_sfixed(1485.0/65536.0,1,-nbitq), 
to_sfixed(-11.0/65536.0,1,-nbitq), 
to_sfixed(467.0/65536.0,1,-nbitq), 
to_sfixed(-2710.0/65536.0,1,-nbitq), 
to_sfixed(-747.0/65536.0,1,-nbitq), 
to_sfixed(-1204.0/65536.0,1,-nbitq), 
to_sfixed(295.0/65536.0,1,-nbitq), 
to_sfixed(1886.0/65536.0,1,-nbitq), 
to_sfixed(1960.0/65536.0,1,-nbitq), 
to_sfixed(1399.0/65536.0,1,-nbitq), 
to_sfixed(94.0/65536.0,1,-nbitq), 
to_sfixed(1072.0/65536.0,1,-nbitq), 
to_sfixed(-28.0/65536.0,1,-nbitq), 
to_sfixed(-256.0/65536.0,1,-nbitq), 
to_sfixed(-468.0/65536.0,1,-nbitq), 
to_sfixed(-1200.0/65536.0,1,-nbitq), 
to_sfixed(-2712.0/65536.0,1,-nbitq), 
to_sfixed(-1214.0/65536.0,1,-nbitq), 
to_sfixed(138.0/65536.0,1,-nbitq), 
to_sfixed(-1125.0/65536.0,1,-nbitq), 
to_sfixed(3032.0/65536.0,1,-nbitq), 
to_sfixed(-4227.0/65536.0,1,-nbitq), 
to_sfixed(-2598.0/65536.0,1,-nbitq), 
to_sfixed(2632.0/65536.0,1,-nbitq), 
to_sfixed(2074.0/65536.0,1,-nbitq), 
to_sfixed(-1491.0/65536.0,1,-nbitq), 
to_sfixed(957.0/65536.0,1,-nbitq), 
to_sfixed(2017.0/65536.0,1,-nbitq), 
to_sfixed(29.0/65536.0,1,-nbitq), 
to_sfixed(1488.0/65536.0,1,-nbitq), 
to_sfixed(1749.0/65536.0,1,-nbitq), 
to_sfixed(2327.0/65536.0,1,-nbitq), 
to_sfixed(-3063.0/65536.0,1,-nbitq), 
to_sfixed(-109.0/65536.0,1,-nbitq), 
to_sfixed(184.0/65536.0,1,-nbitq), 
to_sfixed(1264.0/65536.0,1,-nbitq), 
to_sfixed(-257.0/65536.0,1,-nbitq), 
to_sfixed(750.0/65536.0,1,-nbitq), 
to_sfixed(5231.0/65536.0,1,-nbitq), 
to_sfixed(1709.0/65536.0,1,-nbitq), 
to_sfixed(2411.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2523.0/65536.0,1,-nbitq), 
to_sfixed(1919.0/65536.0,1,-nbitq), 
to_sfixed(-1293.0/65536.0,1,-nbitq), 
to_sfixed(571.0/65536.0,1,-nbitq), 
to_sfixed(-1449.0/65536.0,1,-nbitq), 
to_sfixed(-4400.0/65536.0,1,-nbitq), 
to_sfixed(-2557.0/65536.0,1,-nbitq), 
to_sfixed(1035.0/65536.0,1,-nbitq), 
to_sfixed(2032.0/65536.0,1,-nbitq), 
to_sfixed(925.0/65536.0,1,-nbitq), 
to_sfixed(1497.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(-858.0/65536.0,1,-nbitq), 
to_sfixed(-1661.0/65536.0,1,-nbitq), 
to_sfixed(3294.0/65536.0,1,-nbitq), 
to_sfixed(-383.0/65536.0,1,-nbitq), 
to_sfixed(-3127.0/65536.0,1,-nbitq), 
to_sfixed(-800.0/65536.0,1,-nbitq), 
to_sfixed(2531.0/65536.0,1,-nbitq), 
to_sfixed(2893.0/65536.0,1,-nbitq), 
to_sfixed(735.0/65536.0,1,-nbitq), 
to_sfixed(12.0/65536.0,1,-nbitq), 
to_sfixed(-1481.0/65536.0,1,-nbitq), 
to_sfixed(1399.0/65536.0,1,-nbitq), 
to_sfixed(1269.0/65536.0,1,-nbitq), 
to_sfixed(2884.0/65536.0,1,-nbitq), 
to_sfixed(2345.0/65536.0,1,-nbitq), 
to_sfixed(1510.0/65536.0,1,-nbitq), 
to_sfixed(-697.0/65536.0,1,-nbitq), 
to_sfixed(-724.0/65536.0,1,-nbitq), 
to_sfixed(-1025.0/65536.0,1,-nbitq), 
to_sfixed(-234.0/65536.0,1,-nbitq), 
to_sfixed(-1156.0/65536.0,1,-nbitq), 
to_sfixed(-1068.0/65536.0,1,-nbitq), 
to_sfixed(1342.0/65536.0,1,-nbitq), 
to_sfixed(2339.0/65536.0,1,-nbitq), 
to_sfixed(-1815.0/65536.0,1,-nbitq), 
to_sfixed(-144.0/65536.0,1,-nbitq), 
to_sfixed(773.0/65536.0,1,-nbitq), 
to_sfixed(1284.0/65536.0,1,-nbitq), 
to_sfixed(717.0/65536.0,1,-nbitq), 
to_sfixed(34.0/65536.0,1,-nbitq), 
to_sfixed(-4621.0/65536.0,1,-nbitq), 
to_sfixed(1605.0/65536.0,1,-nbitq), 
to_sfixed(-1446.0/65536.0,1,-nbitq), 
to_sfixed(3277.0/65536.0,1,-nbitq), 
to_sfixed(2811.0/65536.0,1,-nbitq), 
to_sfixed(-1971.0/65536.0,1,-nbitq), 
to_sfixed(3314.0/65536.0,1,-nbitq), 
to_sfixed(3867.0/65536.0,1,-nbitq), 
to_sfixed(-2226.0/65536.0,1,-nbitq), 
to_sfixed(2117.0/65536.0,1,-nbitq), 
to_sfixed(-1174.0/65536.0,1,-nbitq), 
to_sfixed(-3190.0/65536.0,1,-nbitq), 
to_sfixed(207.0/65536.0,1,-nbitq), 
to_sfixed(1094.0/65536.0,1,-nbitq), 
to_sfixed(-749.0/65536.0,1,-nbitq), 
to_sfixed(465.0/65536.0,1,-nbitq), 
to_sfixed(2936.0/65536.0,1,-nbitq), 
to_sfixed(3746.0/65536.0,1,-nbitq), 
to_sfixed(812.0/65536.0,1,-nbitq), 
to_sfixed(-630.0/65536.0,1,-nbitq), 
to_sfixed(-48.0/65536.0,1,-nbitq), 
to_sfixed(-2623.0/65536.0,1,-nbitq), 
to_sfixed(-1880.0/65536.0,1,-nbitq), 
to_sfixed(1036.0/65536.0,1,-nbitq), 
to_sfixed(3080.0/65536.0,1,-nbitq), 
to_sfixed(-1297.0/65536.0,1,-nbitq), 
to_sfixed(-739.0/65536.0,1,-nbitq), 
to_sfixed(-1218.0/65536.0,1,-nbitq), 
to_sfixed(2888.0/65536.0,1,-nbitq), 
to_sfixed(-493.0/65536.0,1,-nbitq), 
to_sfixed(3479.0/65536.0,1,-nbitq), 
to_sfixed(2254.0/65536.0,1,-nbitq), 
to_sfixed(-1151.0/65536.0,1,-nbitq), 
to_sfixed(-316.0/65536.0,1,-nbitq), 
to_sfixed(-496.0/65536.0,1,-nbitq), 
to_sfixed(2988.0/65536.0,1,-nbitq), 
to_sfixed(211.0/65536.0,1,-nbitq), 
to_sfixed(-223.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4.0/65536.0,1,-nbitq), 
to_sfixed(-340.0/65536.0,1,-nbitq), 
to_sfixed(331.0/65536.0,1,-nbitq), 
to_sfixed(2268.0/65536.0,1,-nbitq), 
to_sfixed(-2439.0/65536.0,1,-nbitq), 
to_sfixed(-2937.0/65536.0,1,-nbitq), 
to_sfixed(2616.0/65536.0,1,-nbitq), 
to_sfixed(1672.0/65536.0,1,-nbitq), 
to_sfixed(-1072.0/65536.0,1,-nbitq), 
to_sfixed(-169.0/65536.0,1,-nbitq), 
to_sfixed(-2151.0/65536.0,1,-nbitq), 
to_sfixed(-373.0/65536.0,1,-nbitq), 
to_sfixed(2177.0/65536.0,1,-nbitq), 
to_sfixed(-2642.0/65536.0,1,-nbitq), 
to_sfixed(3452.0/65536.0,1,-nbitq), 
to_sfixed(611.0/65536.0,1,-nbitq), 
to_sfixed(-2582.0/65536.0,1,-nbitq), 
to_sfixed(1019.0/65536.0,1,-nbitq), 
to_sfixed(368.0/65536.0,1,-nbitq), 
to_sfixed(-981.0/65536.0,1,-nbitq), 
to_sfixed(-1067.0/65536.0,1,-nbitq), 
to_sfixed(797.0/65536.0,1,-nbitq), 
to_sfixed(2125.0/65536.0,1,-nbitq), 
to_sfixed(-1052.0/65536.0,1,-nbitq), 
to_sfixed(2174.0/65536.0,1,-nbitq), 
to_sfixed(79.0/65536.0,1,-nbitq), 
to_sfixed(947.0/65536.0,1,-nbitq), 
to_sfixed(1026.0/65536.0,1,-nbitq), 
to_sfixed(-820.0/65536.0,1,-nbitq), 
to_sfixed(-2972.0/65536.0,1,-nbitq), 
to_sfixed(2606.0/65536.0,1,-nbitq), 
to_sfixed(1375.0/65536.0,1,-nbitq), 
to_sfixed(-764.0/65536.0,1,-nbitq), 
to_sfixed(-3550.0/65536.0,1,-nbitq), 
to_sfixed(1003.0/65536.0,1,-nbitq), 
to_sfixed(-694.0/65536.0,1,-nbitq), 
to_sfixed(493.0/65536.0,1,-nbitq), 
to_sfixed(-692.0/65536.0,1,-nbitq), 
to_sfixed(1410.0/65536.0,1,-nbitq), 
to_sfixed(151.0/65536.0,1,-nbitq), 
to_sfixed(-1211.0/65536.0,1,-nbitq), 
to_sfixed(-2738.0/65536.0,1,-nbitq), 
to_sfixed(-2262.0/65536.0,1,-nbitq), 
to_sfixed(1158.0/65536.0,1,-nbitq), 
to_sfixed(-169.0/65536.0,1,-nbitq), 
to_sfixed(4939.0/65536.0,1,-nbitq), 
to_sfixed(-2357.0/65536.0,1,-nbitq), 
to_sfixed(-2023.0/65536.0,1,-nbitq), 
to_sfixed(3485.0/65536.0,1,-nbitq), 
to_sfixed(2618.0/65536.0,1,-nbitq), 
to_sfixed(1209.0/65536.0,1,-nbitq), 
to_sfixed(1760.0/65536.0,1,-nbitq), 
to_sfixed(-1001.0/65536.0,1,-nbitq), 
to_sfixed(582.0/65536.0,1,-nbitq), 
to_sfixed(-1431.0/65536.0,1,-nbitq), 
to_sfixed(-2375.0/65536.0,1,-nbitq), 
to_sfixed(2336.0/65536.0,1,-nbitq), 
to_sfixed(3284.0/65536.0,1,-nbitq), 
to_sfixed(3035.0/65536.0,1,-nbitq), 
to_sfixed(4116.0/65536.0,1,-nbitq), 
to_sfixed(-3339.0/65536.0,1,-nbitq), 
to_sfixed(-2221.0/65536.0,1,-nbitq), 
to_sfixed(2064.0/65536.0,1,-nbitq), 
to_sfixed(-276.0/65536.0,1,-nbitq), 
to_sfixed(2598.0/65536.0,1,-nbitq), 
to_sfixed(2659.0/65536.0,1,-nbitq), 
to_sfixed(2092.0/65536.0,1,-nbitq), 
to_sfixed(900.0/65536.0,1,-nbitq), 
to_sfixed(1205.0/65536.0,1,-nbitq), 
to_sfixed(1452.0/65536.0,1,-nbitq), 
to_sfixed(-1248.0/65536.0,1,-nbitq), 
to_sfixed(-1955.0/65536.0,1,-nbitq), 
to_sfixed(3030.0/65536.0,1,-nbitq), 
to_sfixed(927.0/65536.0,1,-nbitq), 
to_sfixed(1032.0/65536.0,1,-nbitq), 
to_sfixed(-688.0/65536.0,1,-nbitq), 
to_sfixed(2061.0/65536.0,1,-nbitq), 
to_sfixed(2234.0/65536.0,1,-nbitq), 
to_sfixed(207.0/65536.0,1,-nbitq), 
to_sfixed(3107.0/65536.0,1,-nbitq)  ), 
( to_sfixed(788.0/65536.0,1,-nbitq), 
to_sfixed(-2711.0/65536.0,1,-nbitq), 
to_sfixed(4797.0/65536.0,1,-nbitq), 
to_sfixed(-2792.0/65536.0,1,-nbitq), 
to_sfixed(-856.0/65536.0,1,-nbitq), 
to_sfixed(-2277.0/65536.0,1,-nbitq), 
to_sfixed(1402.0/65536.0,1,-nbitq), 
to_sfixed(-1844.0/65536.0,1,-nbitq), 
to_sfixed(-4722.0/65536.0,1,-nbitq), 
to_sfixed(2719.0/65536.0,1,-nbitq), 
to_sfixed(-1144.0/65536.0,1,-nbitq), 
to_sfixed(-2080.0/65536.0,1,-nbitq), 
to_sfixed(1830.0/65536.0,1,-nbitq), 
to_sfixed(1104.0/65536.0,1,-nbitq), 
to_sfixed(2568.0/65536.0,1,-nbitq), 
to_sfixed(2574.0/65536.0,1,-nbitq), 
to_sfixed(1056.0/65536.0,1,-nbitq), 
to_sfixed(1931.0/65536.0,1,-nbitq), 
to_sfixed(1062.0/65536.0,1,-nbitq), 
to_sfixed(388.0/65536.0,1,-nbitq), 
to_sfixed(-1149.0/65536.0,1,-nbitq), 
to_sfixed(181.0/65536.0,1,-nbitq), 
to_sfixed(1352.0/65536.0,1,-nbitq), 
to_sfixed(1763.0/65536.0,1,-nbitq), 
to_sfixed(-667.0/65536.0,1,-nbitq), 
to_sfixed(3078.0/65536.0,1,-nbitq), 
to_sfixed(-1839.0/65536.0,1,-nbitq), 
to_sfixed(-1318.0/65536.0,1,-nbitq), 
to_sfixed(256.0/65536.0,1,-nbitq), 
to_sfixed(-3101.0/65536.0,1,-nbitq), 
to_sfixed(-2416.0/65536.0,1,-nbitq), 
to_sfixed(2144.0/65536.0,1,-nbitq), 
to_sfixed(-1854.0/65536.0,1,-nbitq), 
to_sfixed(-3951.0/65536.0,1,-nbitq), 
to_sfixed(767.0/65536.0,1,-nbitq), 
to_sfixed(-343.0/65536.0,1,-nbitq), 
to_sfixed(1780.0/65536.0,1,-nbitq), 
to_sfixed(24.0/65536.0,1,-nbitq), 
to_sfixed(-1879.0/65536.0,1,-nbitq), 
to_sfixed(2399.0/65536.0,1,-nbitq), 
to_sfixed(750.0/65536.0,1,-nbitq), 
to_sfixed(-2786.0/65536.0,1,-nbitq), 
to_sfixed(-2985.0/65536.0,1,-nbitq), 
to_sfixed(-1874.0/65536.0,1,-nbitq), 
to_sfixed(3263.0/65536.0,1,-nbitq), 
to_sfixed(5595.0/65536.0,1,-nbitq), 
to_sfixed(445.0/65536.0,1,-nbitq), 
to_sfixed(1218.0/65536.0,1,-nbitq), 
to_sfixed(-1786.0/65536.0,1,-nbitq), 
to_sfixed(2687.0/65536.0,1,-nbitq), 
to_sfixed(-2387.0/65536.0,1,-nbitq), 
to_sfixed(157.0/65536.0,1,-nbitq), 
to_sfixed(3426.0/65536.0,1,-nbitq), 
to_sfixed(-1520.0/65536.0,1,-nbitq), 
to_sfixed(-89.0/65536.0,1,-nbitq), 
to_sfixed(3358.0/65536.0,1,-nbitq), 
to_sfixed(1124.0/65536.0,1,-nbitq), 
to_sfixed(-1322.0/65536.0,1,-nbitq), 
to_sfixed(659.0/65536.0,1,-nbitq), 
to_sfixed(2012.0/65536.0,1,-nbitq), 
to_sfixed(-3745.0/65536.0,1,-nbitq), 
to_sfixed(2158.0/65536.0,1,-nbitq), 
to_sfixed(-1354.0/65536.0,1,-nbitq), 
to_sfixed(-3231.0/65536.0,1,-nbitq), 
to_sfixed(-898.0/65536.0,1,-nbitq), 
to_sfixed(456.0/65536.0,1,-nbitq), 
to_sfixed(-1010.0/65536.0,1,-nbitq), 
to_sfixed(-508.0/65536.0,1,-nbitq), 
to_sfixed(-3082.0/65536.0,1,-nbitq), 
to_sfixed(-523.0/65536.0,1,-nbitq), 
to_sfixed(-1688.0/65536.0,1,-nbitq), 
to_sfixed(-2866.0/65536.0,1,-nbitq), 
to_sfixed(3654.0/65536.0,1,-nbitq), 
to_sfixed(2497.0/65536.0,1,-nbitq), 
to_sfixed(312.0/65536.0,1,-nbitq), 
to_sfixed(-715.0/65536.0,1,-nbitq), 
to_sfixed(1785.0/65536.0,1,-nbitq), 
to_sfixed(2065.0/65536.0,1,-nbitq), 
to_sfixed(-366.0/65536.0,1,-nbitq), 
to_sfixed(3880.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2100.0/65536.0,1,-nbitq), 
to_sfixed(1594.0/65536.0,1,-nbitq), 
to_sfixed(4102.0/65536.0,1,-nbitq), 
to_sfixed(3396.0/65536.0,1,-nbitq), 
to_sfixed(2657.0/65536.0,1,-nbitq), 
to_sfixed(224.0/65536.0,1,-nbitq), 
to_sfixed(-14.0/65536.0,1,-nbitq), 
to_sfixed(-2582.0/65536.0,1,-nbitq), 
to_sfixed(-5456.0/65536.0,1,-nbitq), 
to_sfixed(2815.0/65536.0,1,-nbitq), 
to_sfixed(1803.0/65536.0,1,-nbitq), 
to_sfixed(2992.0/65536.0,1,-nbitq), 
to_sfixed(647.0/65536.0,1,-nbitq), 
to_sfixed(1711.0/65536.0,1,-nbitq), 
to_sfixed(2631.0/65536.0,1,-nbitq), 
to_sfixed(-2178.0/65536.0,1,-nbitq), 
to_sfixed(-1829.0/65536.0,1,-nbitq), 
to_sfixed(-4046.0/65536.0,1,-nbitq), 
to_sfixed(4318.0/65536.0,1,-nbitq), 
to_sfixed(286.0/65536.0,1,-nbitq), 
to_sfixed(-522.0/65536.0,1,-nbitq), 
to_sfixed(-2193.0/65536.0,1,-nbitq), 
to_sfixed(-1446.0/65536.0,1,-nbitq), 
to_sfixed(6337.0/65536.0,1,-nbitq), 
to_sfixed(2964.0/65536.0,1,-nbitq), 
to_sfixed(9920.0/65536.0,1,-nbitq), 
to_sfixed(1453.0/65536.0,1,-nbitq), 
to_sfixed(575.0/65536.0,1,-nbitq), 
to_sfixed(-1285.0/65536.0,1,-nbitq), 
to_sfixed(3505.0/65536.0,1,-nbitq), 
to_sfixed(-3751.0/65536.0,1,-nbitq), 
to_sfixed(44.0/65536.0,1,-nbitq), 
to_sfixed(-354.0/65536.0,1,-nbitq), 
to_sfixed(-1593.0/65536.0,1,-nbitq), 
to_sfixed(-2625.0/65536.0,1,-nbitq), 
to_sfixed(-1264.0/65536.0,1,-nbitq), 
to_sfixed(-370.0/65536.0,1,-nbitq), 
to_sfixed(-3674.0/65536.0,1,-nbitq), 
to_sfixed(-429.0/65536.0,1,-nbitq), 
to_sfixed(-4742.0/65536.0,1,-nbitq), 
to_sfixed(-2008.0/65536.0,1,-nbitq), 
to_sfixed(-1416.0/65536.0,1,-nbitq), 
to_sfixed(-3772.0/65536.0,1,-nbitq), 
to_sfixed(-4542.0/65536.0,1,-nbitq), 
to_sfixed(1644.0/65536.0,1,-nbitq), 
to_sfixed(6935.0/65536.0,1,-nbitq), 
to_sfixed(1368.0/65536.0,1,-nbitq), 
to_sfixed(2090.0/65536.0,1,-nbitq), 
to_sfixed(2395.0/65536.0,1,-nbitq), 
to_sfixed(-1162.0/65536.0,1,-nbitq), 
to_sfixed(866.0/65536.0,1,-nbitq), 
to_sfixed(-67.0/65536.0,1,-nbitq), 
to_sfixed(-2030.0/65536.0,1,-nbitq), 
to_sfixed(956.0/65536.0,1,-nbitq), 
to_sfixed(1448.0/65536.0,1,-nbitq), 
to_sfixed(263.0/65536.0,1,-nbitq), 
to_sfixed(-817.0/65536.0,1,-nbitq), 
to_sfixed(-625.0/65536.0,1,-nbitq), 
to_sfixed(2447.0/65536.0,1,-nbitq), 
to_sfixed(7396.0/65536.0,1,-nbitq), 
to_sfixed(-1311.0/65536.0,1,-nbitq), 
to_sfixed(-456.0/65536.0,1,-nbitq), 
to_sfixed(231.0/65536.0,1,-nbitq), 
to_sfixed(2264.0/65536.0,1,-nbitq), 
to_sfixed(-1851.0/65536.0,1,-nbitq), 
to_sfixed(-346.0/65536.0,1,-nbitq), 
to_sfixed(-25.0/65536.0,1,-nbitq), 
to_sfixed(-3909.0/65536.0,1,-nbitq), 
to_sfixed(-1100.0/65536.0,1,-nbitq), 
to_sfixed(-74.0/65536.0,1,-nbitq), 
to_sfixed(-876.0/65536.0,1,-nbitq), 
to_sfixed(-1799.0/65536.0,1,-nbitq), 
to_sfixed(3548.0/65536.0,1,-nbitq), 
to_sfixed(-3266.0/65536.0,1,-nbitq), 
to_sfixed(2371.0/65536.0,1,-nbitq), 
to_sfixed(-1653.0/65536.0,1,-nbitq), 
to_sfixed(-2232.0/65536.0,1,-nbitq), 
to_sfixed(-2283.0/65536.0,1,-nbitq), 
to_sfixed(250.0/65536.0,1,-nbitq), 
to_sfixed(-908.0/65536.0,1,-nbitq)  ), 
( to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(-377.0/65536.0,1,-nbitq), 
to_sfixed(3601.0/65536.0,1,-nbitq), 
to_sfixed(7744.0/65536.0,1,-nbitq), 
to_sfixed(1994.0/65536.0,1,-nbitq), 
to_sfixed(2684.0/65536.0,1,-nbitq), 
to_sfixed(-4102.0/65536.0,1,-nbitq), 
to_sfixed(-671.0/65536.0,1,-nbitq), 
to_sfixed(-3669.0/65536.0,1,-nbitq), 
to_sfixed(1824.0/65536.0,1,-nbitq), 
to_sfixed(2076.0/65536.0,1,-nbitq), 
to_sfixed(8037.0/65536.0,1,-nbitq), 
to_sfixed(-1948.0/65536.0,1,-nbitq), 
to_sfixed(6518.0/65536.0,1,-nbitq), 
to_sfixed(5059.0/65536.0,1,-nbitq), 
to_sfixed(-2641.0/65536.0,1,-nbitq), 
to_sfixed(-2878.0/65536.0,1,-nbitq), 
to_sfixed(-7440.0/65536.0,1,-nbitq), 
to_sfixed(422.0/65536.0,1,-nbitq), 
to_sfixed(-1783.0/65536.0,1,-nbitq), 
to_sfixed(-2134.0/65536.0,1,-nbitq), 
to_sfixed(390.0/65536.0,1,-nbitq), 
to_sfixed(2684.0/65536.0,1,-nbitq), 
to_sfixed(8644.0/65536.0,1,-nbitq), 
to_sfixed(-1363.0/65536.0,1,-nbitq), 
to_sfixed(16748.0/65536.0,1,-nbitq), 
to_sfixed(8889.0/65536.0,1,-nbitq), 
to_sfixed(-1722.0/65536.0,1,-nbitq), 
to_sfixed(-1456.0/65536.0,1,-nbitq), 
to_sfixed(1449.0/65536.0,1,-nbitq), 
to_sfixed(-246.0/65536.0,1,-nbitq), 
to_sfixed(2520.0/65536.0,1,-nbitq), 
to_sfixed(2474.0/65536.0,1,-nbitq), 
to_sfixed(-331.0/65536.0,1,-nbitq), 
to_sfixed(3321.0/65536.0,1,-nbitq), 
to_sfixed(537.0/65536.0,1,-nbitq), 
to_sfixed(-3746.0/65536.0,1,-nbitq), 
to_sfixed(-7714.0/65536.0,1,-nbitq), 
to_sfixed(-556.0/65536.0,1,-nbitq), 
to_sfixed(-5817.0/65536.0,1,-nbitq), 
to_sfixed(554.0/65536.0,1,-nbitq), 
to_sfixed(-2986.0/65536.0,1,-nbitq), 
to_sfixed(-3980.0/65536.0,1,-nbitq), 
to_sfixed(-1079.0/65536.0,1,-nbitq), 
to_sfixed(-2329.0/65536.0,1,-nbitq), 
to_sfixed(3196.0/65536.0,1,-nbitq), 
to_sfixed(16.0/65536.0,1,-nbitq), 
to_sfixed(3454.0/65536.0,1,-nbitq), 
to_sfixed(-972.0/65536.0,1,-nbitq), 
to_sfixed(-856.0/65536.0,1,-nbitq), 
to_sfixed(-1263.0/65536.0,1,-nbitq), 
to_sfixed(-3462.0/65536.0,1,-nbitq), 
to_sfixed(1688.0/65536.0,1,-nbitq), 
to_sfixed(5452.0/65536.0,1,-nbitq), 
to_sfixed(676.0/65536.0,1,-nbitq), 
to_sfixed(5384.0/65536.0,1,-nbitq), 
to_sfixed(-975.0/65536.0,1,-nbitq), 
to_sfixed(-392.0/65536.0,1,-nbitq), 
to_sfixed(-868.0/65536.0,1,-nbitq), 
to_sfixed(3910.0/65536.0,1,-nbitq), 
to_sfixed(-4367.0/65536.0,1,-nbitq), 
to_sfixed(-2465.0/65536.0,1,-nbitq), 
to_sfixed(-1775.0/65536.0,1,-nbitq), 
to_sfixed(-1676.0/65536.0,1,-nbitq), 
to_sfixed(3339.0/65536.0,1,-nbitq), 
to_sfixed(3874.0/65536.0,1,-nbitq), 
to_sfixed(-40.0/65536.0,1,-nbitq), 
to_sfixed(-8135.0/65536.0,1,-nbitq), 
to_sfixed(-7427.0/65536.0,1,-nbitq), 
to_sfixed(1034.0/65536.0,1,-nbitq), 
to_sfixed(3064.0/65536.0,1,-nbitq), 
to_sfixed(-4700.0/65536.0,1,-nbitq), 
to_sfixed(-2347.0/65536.0,1,-nbitq), 
to_sfixed(-1117.0/65536.0,1,-nbitq), 
to_sfixed(-2241.0/65536.0,1,-nbitq), 
to_sfixed(96.0/65536.0,1,-nbitq), 
to_sfixed(309.0/65536.0,1,-nbitq), 
to_sfixed(-2975.0/65536.0,1,-nbitq), 
to_sfixed(-2543.0/65536.0,1,-nbitq), 
to_sfixed(-2619.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1689.0/65536.0,1,-nbitq), 
to_sfixed(1227.0/65536.0,1,-nbitq), 
to_sfixed(4989.0/65536.0,1,-nbitq), 
to_sfixed(8608.0/65536.0,1,-nbitq), 
to_sfixed(1619.0/65536.0,1,-nbitq), 
to_sfixed(3867.0/65536.0,1,-nbitq), 
to_sfixed(-233.0/65536.0,1,-nbitq), 
to_sfixed(-670.0/65536.0,1,-nbitq), 
to_sfixed(-1229.0/65536.0,1,-nbitq), 
to_sfixed(1914.0/65536.0,1,-nbitq), 
to_sfixed(-365.0/65536.0,1,-nbitq), 
to_sfixed(12184.0/65536.0,1,-nbitq), 
to_sfixed(1211.0/65536.0,1,-nbitq), 
to_sfixed(-1931.0/65536.0,1,-nbitq), 
to_sfixed(4443.0/65536.0,1,-nbitq), 
to_sfixed(-2146.0/65536.0,1,-nbitq), 
to_sfixed(955.0/65536.0,1,-nbitq), 
to_sfixed(-2585.0/65536.0,1,-nbitq), 
to_sfixed(1072.0/65536.0,1,-nbitq), 
to_sfixed(706.0/65536.0,1,-nbitq), 
to_sfixed(3343.0/65536.0,1,-nbitq), 
to_sfixed(6592.0/65536.0,1,-nbitq), 
to_sfixed(2973.0/65536.0,1,-nbitq), 
to_sfixed(4085.0/65536.0,1,-nbitq), 
to_sfixed(5483.0/65536.0,1,-nbitq), 
to_sfixed(15816.0/65536.0,1,-nbitq), 
to_sfixed(9545.0/65536.0,1,-nbitq), 
to_sfixed(-1172.0/65536.0,1,-nbitq), 
to_sfixed(-290.0/65536.0,1,-nbitq), 
to_sfixed(3067.0/65536.0,1,-nbitq), 
to_sfixed(-2739.0/65536.0,1,-nbitq), 
to_sfixed(1577.0/65536.0,1,-nbitq), 
to_sfixed(4264.0/65536.0,1,-nbitq), 
to_sfixed(437.0/65536.0,1,-nbitq), 
to_sfixed(1595.0/65536.0,1,-nbitq), 
to_sfixed(-1878.0/65536.0,1,-nbitq), 
to_sfixed(-5386.0/65536.0,1,-nbitq), 
to_sfixed(-2192.0/65536.0,1,-nbitq), 
to_sfixed(-1890.0/65536.0,1,-nbitq), 
to_sfixed(-5028.0/65536.0,1,-nbitq), 
to_sfixed(-2763.0/65536.0,1,-nbitq), 
to_sfixed(1858.0/65536.0,1,-nbitq), 
to_sfixed(-1021.0/65536.0,1,-nbitq), 
to_sfixed(-2382.0/65536.0,1,-nbitq), 
to_sfixed(-570.0/65536.0,1,-nbitq), 
to_sfixed(3104.0/65536.0,1,-nbitq), 
to_sfixed(-1329.0/65536.0,1,-nbitq), 
to_sfixed(-727.0/65536.0,1,-nbitq), 
to_sfixed(1300.0/65536.0,1,-nbitq), 
to_sfixed(1268.0/65536.0,1,-nbitq), 
to_sfixed(1629.0/65536.0,1,-nbitq), 
to_sfixed(345.0/65536.0,1,-nbitq), 
to_sfixed(965.0/65536.0,1,-nbitq), 
to_sfixed(7718.0/65536.0,1,-nbitq), 
to_sfixed(-2181.0/65536.0,1,-nbitq), 
to_sfixed(6043.0/65536.0,1,-nbitq), 
to_sfixed(-1941.0/65536.0,1,-nbitq), 
to_sfixed(-3070.0/65536.0,1,-nbitq), 
to_sfixed(-1721.0/65536.0,1,-nbitq), 
to_sfixed(-2466.0/65536.0,1,-nbitq), 
to_sfixed(-1714.0/65536.0,1,-nbitq), 
to_sfixed(1748.0/65536.0,1,-nbitq), 
to_sfixed(1431.0/65536.0,1,-nbitq), 
to_sfixed(-1394.0/65536.0,1,-nbitq), 
to_sfixed(2139.0/65536.0,1,-nbitq), 
to_sfixed(7704.0/65536.0,1,-nbitq), 
to_sfixed(-86.0/65536.0,1,-nbitq), 
to_sfixed(-13794.0/65536.0,1,-nbitq), 
to_sfixed(-7874.0/65536.0,1,-nbitq), 
to_sfixed(-3219.0/65536.0,1,-nbitq), 
to_sfixed(-517.0/65536.0,1,-nbitq), 
to_sfixed(-1678.0/65536.0,1,-nbitq), 
to_sfixed(-2160.0/65536.0,1,-nbitq), 
to_sfixed(1210.0/65536.0,1,-nbitq), 
to_sfixed(1198.0/65536.0,1,-nbitq), 
to_sfixed(2495.0/65536.0,1,-nbitq), 
to_sfixed(-2210.0/65536.0,1,-nbitq), 
to_sfixed(-5531.0/65536.0,1,-nbitq), 
to_sfixed(-1567.0/65536.0,1,-nbitq), 
to_sfixed(-416.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-451.0/65536.0,1,-nbitq), 
to_sfixed(-3980.0/65536.0,1,-nbitq), 
to_sfixed(5837.0/65536.0,1,-nbitq), 
to_sfixed(5055.0/65536.0,1,-nbitq), 
to_sfixed(2297.0/65536.0,1,-nbitq), 
to_sfixed(7666.0/65536.0,1,-nbitq), 
to_sfixed(-858.0/65536.0,1,-nbitq), 
to_sfixed(1052.0/65536.0,1,-nbitq), 
to_sfixed(-2548.0/65536.0,1,-nbitq), 
to_sfixed(2079.0/65536.0,1,-nbitq), 
to_sfixed(3784.0/65536.0,1,-nbitq), 
to_sfixed(28112.0/65536.0,1,-nbitq), 
to_sfixed(1693.0/65536.0,1,-nbitq), 
to_sfixed(485.0/65536.0,1,-nbitq), 
to_sfixed(793.0/65536.0,1,-nbitq), 
to_sfixed(1042.0/65536.0,1,-nbitq), 
to_sfixed(2586.0/65536.0,1,-nbitq), 
to_sfixed(-3978.0/65536.0,1,-nbitq), 
to_sfixed(-365.0/65536.0,1,-nbitq), 
to_sfixed(-705.0/65536.0,1,-nbitq), 
to_sfixed(1068.0/65536.0,1,-nbitq), 
to_sfixed(1184.0/65536.0,1,-nbitq), 
to_sfixed(-1336.0/65536.0,1,-nbitq), 
to_sfixed(-8121.0/65536.0,1,-nbitq), 
to_sfixed(4592.0/65536.0,1,-nbitq), 
to_sfixed(10868.0/65536.0,1,-nbitq), 
to_sfixed(17300.0/65536.0,1,-nbitq), 
to_sfixed(-2413.0/65536.0,1,-nbitq), 
to_sfixed(915.0/65536.0,1,-nbitq), 
to_sfixed(553.0/65536.0,1,-nbitq), 
to_sfixed(-1177.0/65536.0,1,-nbitq), 
to_sfixed(-1513.0/65536.0,1,-nbitq), 
to_sfixed(1664.0/65536.0,1,-nbitq), 
to_sfixed(-6494.0/65536.0,1,-nbitq), 
to_sfixed(-2326.0/65536.0,1,-nbitq), 
to_sfixed(1936.0/65536.0,1,-nbitq), 
to_sfixed(-7051.0/65536.0,1,-nbitq), 
to_sfixed(1261.0/65536.0,1,-nbitq), 
to_sfixed(-7064.0/65536.0,1,-nbitq), 
to_sfixed(-3547.0/65536.0,1,-nbitq), 
to_sfixed(-10297.0/65536.0,1,-nbitq), 
to_sfixed(-1409.0/65536.0,1,-nbitq), 
to_sfixed(5116.0/65536.0,1,-nbitq), 
to_sfixed(1603.0/65536.0,1,-nbitq), 
to_sfixed(2116.0/65536.0,1,-nbitq), 
to_sfixed(-245.0/65536.0,1,-nbitq), 
to_sfixed(1222.0/65536.0,1,-nbitq), 
to_sfixed(-2727.0/65536.0,1,-nbitq), 
to_sfixed(3601.0/65536.0,1,-nbitq), 
to_sfixed(3316.0/65536.0,1,-nbitq), 
to_sfixed(529.0/65536.0,1,-nbitq), 
to_sfixed(2674.0/65536.0,1,-nbitq), 
to_sfixed(2680.0/65536.0,1,-nbitq), 
to_sfixed(4765.0/65536.0,1,-nbitq), 
to_sfixed(-5341.0/65536.0,1,-nbitq), 
to_sfixed(12725.0/65536.0,1,-nbitq), 
to_sfixed(832.0/65536.0,1,-nbitq), 
to_sfixed(-6421.0/65536.0,1,-nbitq), 
to_sfixed(3730.0/65536.0,1,-nbitq), 
to_sfixed(-5385.0/65536.0,1,-nbitq), 
to_sfixed(-2534.0/65536.0,1,-nbitq), 
to_sfixed(-738.0/65536.0,1,-nbitq), 
to_sfixed(217.0/65536.0,1,-nbitq), 
to_sfixed(-3391.0/65536.0,1,-nbitq), 
to_sfixed(-2513.0/65536.0,1,-nbitq), 
to_sfixed(10205.0/65536.0,1,-nbitq), 
to_sfixed(-4451.0/65536.0,1,-nbitq), 
to_sfixed(-14592.0/65536.0,1,-nbitq), 
to_sfixed(-5449.0/65536.0,1,-nbitq), 
to_sfixed(-1251.0/65536.0,1,-nbitq), 
to_sfixed(-1086.0/65536.0,1,-nbitq), 
to_sfixed(-8408.0/65536.0,1,-nbitq), 
to_sfixed(-41.0/65536.0,1,-nbitq), 
to_sfixed(633.0/65536.0,1,-nbitq), 
to_sfixed(2609.0/65536.0,1,-nbitq), 
to_sfixed(695.0/65536.0,1,-nbitq), 
to_sfixed(-1351.0/65536.0,1,-nbitq), 
to_sfixed(-6324.0/65536.0,1,-nbitq), 
to_sfixed(-948.0/65536.0,1,-nbitq), 
to_sfixed(-3924.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2582.0/65536.0,1,-nbitq), 
to_sfixed(1619.0/65536.0,1,-nbitq), 
to_sfixed(1475.0/65536.0,1,-nbitq), 
to_sfixed(8279.0/65536.0,1,-nbitq), 
to_sfixed(2133.0/65536.0,1,-nbitq), 
to_sfixed(-5183.0/65536.0,1,-nbitq), 
to_sfixed(1112.0/65536.0,1,-nbitq), 
to_sfixed(9586.0/65536.0,1,-nbitq), 
to_sfixed(-381.0/65536.0,1,-nbitq), 
to_sfixed(-1476.0/65536.0,1,-nbitq), 
to_sfixed(2983.0/65536.0,1,-nbitq), 
to_sfixed(21790.0/65536.0,1,-nbitq), 
to_sfixed(-2208.0/65536.0,1,-nbitq), 
to_sfixed(2486.0/65536.0,1,-nbitq), 
to_sfixed(-564.0/65536.0,1,-nbitq), 
to_sfixed(507.0/65536.0,1,-nbitq), 
to_sfixed(-3056.0/65536.0,1,-nbitq), 
to_sfixed(7948.0/65536.0,1,-nbitq), 
to_sfixed(315.0/65536.0,1,-nbitq), 
to_sfixed(-2544.0/65536.0,1,-nbitq), 
to_sfixed(4578.0/65536.0,1,-nbitq), 
to_sfixed(-4366.0/65536.0,1,-nbitq), 
to_sfixed(-9783.0/65536.0,1,-nbitq), 
to_sfixed(-15932.0/65536.0,1,-nbitq), 
to_sfixed(1940.0/65536.0,1,-nbitq), 
to_sfixed(3917.0/65536.0,1,-nbitq), 
to_sfixed(11199.0/65536.0,1,-nbitq), 
to_sfixed(-3403.0/65536.0,1,-nbitq), 
to_sfixed(2227.0/65536.0,1,-nbitq), 
to_sfixed(-1045.0/65536.0,1,-nbitq), 
to_sfixed(1628.0/65536.0,1,-nbitq), 
to_sfixed(934.0/65536.0,1,-nbitq), 
to_sfixed(3061.0/65536.0,1,-nbitq), 
to_sfixed(3685.0/65536.0,1,-nbitq), 
to_sfixed(-3191.0/65536.0,1,-nbitq), 
to_sfixed(2378.0/65536.0,1,-nbitq), 
to_sfixed(-3656.0/65536.0,1,-nbitq), 
to_sfixed(3783.0/65536.0,1,-nbitq), 
to_sfixed(-8621.0/65536.0,1,-nbitq), 
to_sfixed(683.0/65536.0,1,-nbitq), 
to_sfixed(-9480.0/65536.0,1,-nbitq), 
to_sfixed(-579.0/65536.0,1,-nbitq), 
to_sfixed(3941.0/65536.0,1,-nbitq), 
to_sfixed(2677.0/65536.0,1,-nbitq), 
to_sfixed(-1610.0/65536.0,1,-nbitq), 
to_sfixed(-107.0/65536.0,1,-nbitq), 
to_sfixed(-1736.0/65536.0,1,-nbitq), 
to_sfixed(719.0/65536.0,1,-nbitq), 
to_sfixed(234.0/65536.0,1,-nbitq), 
to_sfixed(-89.0/65536.0,1,-nbitq), 
to_sfixed(-2331.0/65536.0,1,-nbitq), 
to_sfixed(10044.0/65536.0,1,-nbitq), 
to_sfixed(1110.0/65536.0,1,-nbitq), 
to_sfixed(5584.0/65536.0,1,-nbitq), 
to_sfixed(-2217.0/65536.0,1,-nbitq), 
to_sfixed(8798.0/65536.0,1,-nbitq), 
to_sfixed(829.0/65536.0,1,-nbitq), 
to_sfixed(-166.0/65536.0,1,-nbitq), 
to_sfixed(-654.0/65536.0,1,-nbitq), 
to_sfixed(-2300.0/65536.0,1,-nbitq), 
to_sfixed(-2730.0/65536.0,1,-nbitq), 
to_sfixed(338.0/65536.0,1,-nbitq), 
to_sfixed(1473.0/65536.0,1,-nbitq), 
to_sfixed(1312.0/65536.0,1,-nbitq), 
to_sfixed(-8393.0/65536.0,1,-nbitq), 
to_sfixed(4676.0/65536.0,1,-nbitq), 
to_sfixed(-1181.0/65536.0,1,-nbitq), 
to_sfixed(-9581.0/65536.0,1,-nbitq), 
to_sfixed(-4623.0/65536.0,1,-nbitq), 
to_sfixed(1662.0/65536.0,1,-nbitq), 
to_sfixed(-478.0/65536.0,1,-nbitq), 
to_sfixed(-1189.0/65536.0,1,-nbitq), 
to_sfixed(198.0/65536.0,1,-nbitq), 
to_sfixed(-2260.0/65536.0,1,-nbitq), 
to_sfixed(2054.0/65536.0,1,-nbitq), 
to_sfixed(-1955.0/65536.0,1,-nbitq), 
to_sfixed(4228.0/65536.0,1,-nbitq), 
to_sfixed(-5802.0/65536.0,1,-nbitq), 
to_sfixed(-1728.0/65536.0,1,-nbitq), 
to_sfixed(-1761.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2980.0/65536.0,1,-nbitq), 
to_sfixed(-2547.0/65536.0,1,-nbitq), 
to_sfixed(4020.0/65536.0,1,-nbitq), 
to_sfixed(7266.0/65536.0,1,-nbitq), 
to_sfixed(7686.0/65536.0,1,-nbitq), 
to_sfixed(-3227.0/65536.0,1,-nbitq), 
to_sfixed(-1594.0/65536.0,1,-nbitq), 
to_sfixed(2476.0/65536.0,1,-nbitq), 
to_sfixed(309.0/65536.0,1,-nbitq), 
to_sfixed(-2043.0/65536.0,1,-nbitq), 
to_sfixed(-1014.0/65536.0,1,-nbitq), 
to_sfixed(6862.0/65536.0,1,-nbitq), 
to_sfixed(-565.0/65536.0,1,-nbitq), 
to_sfixed(15308.0/65536.0,1,-nbitq), 
to_sfixed(4175.0/65536.0,1,-nbitq), 
to_sfixed(-2690.0/65536.0,1,-nbitq), 
to_sfixed(-3020.0/65536.0,1,-nbitq), 
to_sfixed(13426.0/65536.0,1,-nbitq), 
to_sfixed(989.0/65536.0,1,-nbitq), 
to_sfixed(-1602.0/65536.0,1,-nbitq), 
to_sfixed(5021.0/65536.0,1,-nbitq), 
to_sfixed(-7228.0/65536.0,1,-nbitq), 
to_sfixed(-6523.0/65536.0,1,-nbitq), 
to_sfixed(-5946.0/65536.0,1,-nbitq), 
to_sfixed(-1782.0/65536.0,1,-nbitq), 
to_sfixed(11578.0/65536.0,1,-nbitq), 
to_sfixed(19688.0/65536.0,1,-nbitq), 
to_sfixed(1857.0/65536.0,1,-nbitq), 
to_sfixed(-2383.0/65536.0,1,-nbitq), 
to_sfixed(-5737.0/65536.0,1,-nbitq), 
to_sfixed(-2254.0/65536.0,1,-nbitq), 
to_sfixed(3324.0/65536.0,1,-nbitq), 
to_sfixed(1115.0/65536.0,1,-nbitq), 
to_sfixed(-354.0/65536.0,1,-nbitq), 
to_sfixed(33.0/65536.0,1,-nbitq), 
to_sfixed(-630.0/65536.0,1,-nbitq), 
to_sfixed(773.0/65536.0,1,-nbitq), 
to_sfixed(-1549.0/65536.0,1,-nbitq), 
to_sfixed(-8608.0/65536.0,1,-nbitq), 
to_sfixed(73.0/65536.0,1,-nbitq), 
to_sfixed(-7512.0/65536.0,1,-nbitq), 
to_sfixed(-348.0/65536.0,1,-nbitq), 
to_sfixed(1581.0/65536.0,1,-nbitq), 
to_sfixed(5765.0/65536.0,1,-nbitq), 
to_sfixed(2977.0/65536.0,1,-nbitq), 
to_sfixed(-22.0/65536.0,1,-nbitq), 
to_sfixed(2452.0/65536.0,1,-nbitq), 
to_sfixed(6471.0/65536.0,1,-nbitq), 
to_sfixed(-1847.0/65536.0,1,-nbitq), 
to_sfixed(-35.0/65536.0,1,-nbitq), 
to_sfixed(1253.0/65536.0,1,-nbitq), 
to_sfixed(14734.0/65536.0,1,-nbitq), 
to_sfixed(-1547.0/65536.0,1,-nbitq), 
to_sfixed(7483.0/65536.0,1,-nbitq), 
to_sfixed(-2709.0/65536.0,1,-nbitq), 
to_sfixed(10489.0/65536.0,1,-nbitq), 
to_sfixed(1506.0/65536.0,1,-nbitq), 
to_sfixed(1614.0/65536.0,1,-nbitq), 
to_sfixed(-976.0/65536.0,1,-nbitq), 
to_sfixed(4146.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(-1707.0/65536.0,1,-nbitq), 
to_sfixed(-1822.0/65536.0,1,-nbitq), 
to_sfixed(-750.0/65536.0,1,-nbitq), 
to_sfixed(-10142.0/65536.0,1,-nbitq), 
to_sfixed(4361.0/65536.0,1,-nbitq), 
to_sfixed(-359.0/65536.0,1,-nbitq), 
to_sfixed(-6038.0/65536.0,1,-nbitq), 
to_sfixed(-3973.0/65536.0,1,-nbitq), 
to_sfixed(-10949.0/65536.0,1,-nbitq), 
to_sfixed(-1473.0/65536.0,1,-nbitq), 
to_sfixed(-1125.0/65536.0,1,-nbitq), 
to_sfixed(-1990.0/65536.0,1,-nbitq), 
to_sfixed(309.0/65536.0,1,-nbitq), 
to_sfixed(1001.0/65536.0,1,-nbitq), 
to_sfixed(-1440.0/65536.0,1,-nbitq), 
to_sfixed(17155.0/65536.0,1,-nbitq), 
to_sfixed(-3126.0/65536.0,1,-nbitq), 
to_sfixed(1771.0/65536.0,1,-nbitq), 
to_sfixed(-1480.0/65536.0,1,-nbitq)  ), 
( to_sfixed(780.0/65536.0,1,-nbitq), 
to_sfixed(-3514.0/65536.0,1,-nbitq), 
to_sfixed(767.0/65536.0,1,-nbitq), 
to_sfixed(9999.0/65536.0,1,-nbitq), 
to_sfixed(-3538.0/65536.0,1,-nbitq), 
to_sfixed(-3439.0/65536.0,1,-nbitq), 
to_sfixed(-3497.0/65536.0,1,-nbitq), 
to_sfixed(-4674.0/65536.0,1,-nbitq), 
to_sfixed(4395.0/65536.0,1,-nbitq), 
to_sfixed(2080.0/65536.0,1,-nbitq), 
to_sfixed(-499.0/65536.0,1,-nbitq), 
to_sfixed(5649.0/65536.0,1,-nbitq), 
to_sfixed(-1279.0/65536.0,1,-nbitq), 
to_sfixed(17059.0/65536.0,1,-nbitq), 
to_sfixed(4182.0/65536.0,1,-nbitq), 
to_sfixed(1743.0/65536.0,1,-nbitq), 
to_sfixed(2228.0/65536.0,1,-nbitq), 
to_sfixed(9992.0/65536.0,1,-nbitq), 
to_sfixed(8037.0/65536.0,1,-nbitq), 
to_sfixed(1958.0/65536.0,1,-nbitq), 
to_sfixed(4430.0/65536.0,1,-nbitq), 
to_sfixed(2085.0/65536.0,1,-nbitq), 
to_sfixed(1241.0/65536.0,1,-nbitq), 
to_sfixed(1097.0/65536.0,1,-nbitq), 
to_sfixed(-1426.0/65536.0,1,-nbitq), 
to_sfixed(9833.0/65536.0,1,-nbitq), 
to_sfixed(30823.0/65536.0,1,-nbitq), 
to_sfixed(-2679.0/65536.0,1,-nbitq), 
to_sfixed(-3721.0/65536.0,1,-nbitq), 
to_sfixed(-7263.0/65536.0,1,-nbitq), 
to_sfixed(-1834.0/65536.0,1,-nbitq), 
to_sfixed(6309.0/65536.0,1,-nbitq), 
to_sfixed(6404.0/65536.0,1,-nbitq), 
to_sfixed(4613.0/65536.0,1,-nbitq), 
to_sfixed(3504.0/65536.0,1,-nbitq), 
to_sfixed(2566.0/65536.0,1,-nbitq), 
to_sfixed(3971.0/65536.0,1,-nbitq), 
to_sfixed(-1563.0/65536.0,1,-nbitq), 
to_sfixed(-10058.0/65536.0,1,-nbitq), 
to_sfixed(-2554.0/65536.0,1,-nbitq), 
to_sfixed(-1111.0/65536.0,1,-nbitq), 
to_sfixed(-2347.0/65536.0,1,-nbitq), 
to_sfixed(1920.0/65536.0,1,-nbitq), 
to_sfixed(3819.0/65536.0,1,-nbitq), 
to_sfixed(2566.0/65536.0,1,-nbitq), 
to_sfixed(-6249.0/65536.0,1,-nbitq), 
to_sfixed(2643.0/65536.0,1,-nbitq), 
to_sfixed(2892.0/65536.0,1,-nbitq), 
to_sfixed(2455.0/65536.0,1,-nbitq), 
to_sfixed(903.0/65536.0,1,-nbitq), 
to_sfixed(2420.0/65536.0,1,-nbitq), 
to_sfixed(11879.0/65536.0,1,-nbitq), 
to_sfixed(2854.0/65536.0,1,-nbitq), 
to_sfixed(10695.0/65536.0,1,-nbitq), 
to_sfixed(624.0/65536.0,1,-nbitq), 
to_sfixed(9139.0/65536.0,1,-nbitq), 
to_sfixed(1504.0/65536.0,1,-nbitq), 
to_sfixed(-1832.0/65536.0,1,-nbitq), 
to_sfixed(569.0/65536.0,1,-nbitq), 
to_sfixed(2923.0/65536.0,1,-nbitq), 
to_sfixed(3210.0/65536.0,1,-nbitq), 
to_sfixed(-527.0/65536.0,1,-nbitq), 
to_sfixed(-1853.0/65536.0,1,-nbitq), 
to_sfixed(-1349.0/65536.0,1,-nbitq), 
to_sfixed(-7612.0/65536.0,1,-nbitq), 
to_sfixed(6264.0/65536.0,1,-nbitq), 
to_sfixed(-6290.0/65536.0,1,-nbitq), 
to_sfixed(-7358.0/65536.0,1,-nbitq), 
to_sfixed(-5587.0/65536.0,1,-nbitq), 
to_sfixed(-11487.0/65536.0,1,-nbitq), 
to_sfixed(-1312.0/65536.0,1,-nbitq), 
to_sfixed(-6467.0/65536.0,1,-nbitq), 
to_sfixed(-4025.0/65536.0,1,-nbitq), 
to_sfixed(-2538.0/65536.0,1,-nbitq), 
to_sfixed(-2839.0/65536.0,1,-nbitq), 
to_sfixed(3448.0/65536.0,1,-nbitq), 
to_sfixed(9021.0/65536.0,1,-nbitq), 
to_sfixed(-15619.0/65536.0,1,-nbitq), 
to_sfixed(-2017.0/65536.0,1,-nbitq), 
to_sfixed(-2303.0/65536.0,1,-nbitq)  ), 
( to_sfixed(674.0/65536.0,1,-nbitq), 
to_sfixed(-5265.0/65536.0,1,-nbitq), 
to_sfixed(5236.0/65536.0,1,-nbitq), 
to_sfixed(6231.0/65536.0,1,-nbitq), 
to_sfixed(1135.0/65536.0,1,-nbitq), 
to_sfixed(-7926.0/65536.0,1,-nbitq), 
to_sfixed(2058.0/65536.0,1,-nbitq), 
to_sfixed(-11259.0/65536.0,1,-nbitq), 
to_sfixed(5961.0/65536.0,1,-nbitq), 
to_sfixed(-244.0/65536.0,1,-nbitq), 
to_sfixed(839.0/65536.0,1,-nbitq), 
to_sfixed(11218.0/65536.0,1,-nbitq), 
to_sfixed(-2.0/65536.0,1,-nbitq), 
to_sfixed(4362.0/65536.0,1,-nbitq), 
to_sfixed(-4389.0/65536.0,1,-nbitq), 
to_sfixed(-31.0/65536.0,1,-nbitq), 
to_sfixed(-3.0/65536.0,1,-nbitq), 
to_sfixed(11751.0/65536.0,1,-nbitq), 
to_sfixed(-8667.0/65536.0,1,-nbitq), 
to_sfixed(1718.0/65536.0,1,-nbitq), 
to_sfixed(8767.0/65536.0,1,-nbitq), 
to_sfixed(2917.0/65536.0,1,-nbitq), 
to_sfixed(6827.0/65536.0,1,-nbitq), 
to_sfixed(-3115.0/65536.0,1,-nbitq), 
to_sfixed(-2680.0/65536.0,1,-nbitq), 
to_sfixed(-2915.0/65536.0,1,-nbitq), 
to_sfixed(30695.0/65536.0,1,-nbitq), 
to_sfixed(-746.0/65536.0,1,-nbitq), 
to_sfixed(-1661.0/65536.0,1,-nbitq), 
to_sfixed(-5807.0/65536.0,1,-nbitq), 
to_sfixed(-2660.0/65536.0,1,-nbitq), 
to_sfixed(7848.0/65536.0,1,-nbitq), 
to_sfixed(1873.0/65536.0,1,-nbitq), 
to_sfixed(8786.0/65536.0,1,-nbitq), 
to_sfixed(507.0/65536.0,1,-nbitq), 
to_sfixed(-1343.0/65536.0,1,-nbitq), 
to_sfixed(15255.0/65536.0,1,-nbitq), 
to_sfixed(-3787.0/65536.0,1,-nbitq), 
to_sfixed(-5584.0/65536.0,1,-nbitq), 
to_sfixed(-7574.0/65536.0,1,-nbitq), 
to_sfixed(5322.0/65536.0,1,-nbitq), 
to_sfixed(2231.0/65536.0,1,-nbitq), 
to_sfixed(4378.0/65536.0,1,-nbitq), 
to_sfixed(4944.0/65536.0,1,-nbitq), 
to_sfixed(-951.0/65536.0,1,-nbitq), 
to_sfixed(-19034.0/65536.0,1,-nbitq), 
to_sfixed(-291.0/65536.0,1,-nbitq), 
to_sfixed(1118.0/65536.0,1,-nbitq), 
to_sfixed(-1469.0/65536.0,1,-nbitq), 
to_sfixed(3859.0/65536.0,1,-nbitq), 
to_sfixed(1234.0/65536.0,1,-nbitq), 
to_sfixed(8330.0/65536.0,1,-nbitq), 
to_sfixed(3464.0/65536.0,1,-nbitq), 
to_sfixed(4794.0/65536.0,1,-nbitq), 
to_sfixed(-148.0/65536.0,1,-nbitq), 
to_sfixed(12158.0/65536.0,1,-nbitq), 
to_sfixed(508.0/65536.0,1,-nbitq), 
to_sfixed(-4597.0/65536.0,1,-nbitq), 
to_sfixed(274.0/65536.0,1,-nbitq), 
to_sfixed(5466.0/65536.0,1,-nbitq), 
to_sfixed(13017.0/65536.0,1,-nbitq), 
to_sfixed(-667.0/65536.0,1,-nbitq), 
to_sfixed(834.0/65536.0,1,-nbitq), 
to_sfixed(1474.0/65536.0,1,-nbitq), 
to_sfixed(-7000.0/65536.0,1,-nbitq), 
to_sfixed(-1838.0/65536.0,1,-nbitq), 
to_sfixed(-414.0/65536.0,1,-nbitq), 
to_sfixed(-2816.0/65536.0,1,-nbitq), 
to_sfixed(-8264.0/65536.0,1,-nbitq), 
to_sfixed(-4229.0/65536.0,1,-nbitq), 
to_sfixed(-826.0/65536.0,1,-nbitq), 
to_sfixed(-306.0/65536.0,1,-nbitq), 
to_sfixed(-3446.0/65536.0,1,-nbitq), 
to_sfixed(742.0/65536.0,1,-nbitq), 
to_sfixed(-942.0/65536.0,1,-nbitq), 
to_sfixed(9217.0/65536.0,1,-nbitq), 
to_sfixed(-8697.0/65536.0,1,-nbitq), 
to_sfixed(-20234.0/65536.0,1,-nbitq), 
to_sfixed(72.0/65536.0,1,-nbitq), 
to_sfixed(-1221.0/65536.0,1,-nbitq)  ), 
( to_sfixed(862.0/65536.0,1,-nbitq), 
to_sfixed(-4362.0/65536.0,1,-nbitq), 
to_sfixed(8494.0/65536.0,1,-nbitq), 
to_sfixed(11681.0/65536.0,1,-nbitq), 
to_sfixed(4027.0/65536.0,1,-nbitq), 
to_sfixed(-3480.0/65536.0,1,-nbitq), 
to_sfixed(-1092.0/65536.0,1,-nbitq), 
to_sfixed(-16451.0/65536.0,1,-nbitq), 
to_sfixed(688.0/65536.0,1,-nbitq), 
to_sfixed(-1675.0/65536.0,1,-nbitq), 
to_sfixed(2146.0/65536.0,1,-nbitq), 
to_sfixed(11202.0/65536.0,1,-nbitq), 
to_sfixed(-647.0/65536.0,1,-nbitq), 
to_sfixed(-10598.0/65536.0,1,-nbitq), 
to_sfixed(2267.0/65536.0,1,-nbitq), 
to_sfixed(-613.0/65536.0,1,-nbitq), 
to_sfixed(-152.0/65536.0,1,-nbitq), 
to_sfixed(11561.0/65536.0,1,-nbitq), 
to_sfixed(-10173.0/65536.0,1,-nbitq), 
to_sfixed(229.0/65536.0,1,-nbitq), 
to_sfixed(4883.0/65536.0,1,-nbitq), 
to_sfixed(-8162.0/65536.0,1,-nbitq), 
to_sfixed(6370.0/65536.0,1,-nbitq), 
to_sfixed(3001.0/65536.0,1,-nbitq), 
to_sfixed(815.0/65536.0,1,-nbitq), 
to_sfixed(-2131.0/65536.0,1,-nbitq), 
to_sfixed(34279.0/65536.0,1,-nbitq), 
to_sfixed(-1596.0/65536.0,1,-nbitq), 
to_sfixed(1539.0/65536.0,1,-nbitq), 
to_sfixed(-2800.0/65536.0,1,-nbitq), 
to_sfixed(-3447.0/65536.0,1,-nbitq), 
to_sfixed(11046.0/65536.0,1,-nbitq), 
to_sfixed(2518.0/65536.0,1,-nbitq), 
to_sfixed(12660.0/65536.0,1,-nbitq), 
to_sfixed(606.0/65536.0,1,-nbitq), 
to_sfixed(-4795.0/65536.0,1,-nbitq), 
to_sfixed(11172.0/65536.0,1,-nbitq), 
to_sfixed(-4757.0/65536.0,1,-nbitq), 
to_sfixed(-4673.0/65536.0,1,-nbitq), 
to_sfixed(-4550.0/65536.0,1,-nbitq), 
to_sfixed(-1215.0/65536.0,1,-nbitq), 
to_sfixed(-2281.0/65536.0,1,-nbitq), 
to_sfixed(7969.0/65536.0,1,-nbitq), 
to_sfixed(6454.0/65536.0,1,-nbitq), 
to_sfixed(3213.0/65536.0,1,-nbitq), 
to_sfixed(-9506.0/65536.0,1,-nbitq), 
to_sfixed(4154.0/65536.0,1,-nbitq), 
to_sfixed(26.0/65536.0,1,-nbitq), 
to_sfixed(-2615.0/65536.0,1,-nbitq), 
to_sfixed(1634.0/65536.0,1,-nbitq), 
to_sfixed(-895.0/65536.0,1,-nbitq), 
to_sfixed(1992.0/65536.0,1,-nbitq), 
to_sfixed(-8982.0/65536.0,1,-nbitq), 
to_sfixed(417.0/65536.0,1,-nbitq), 
to_sfixed(1896.0/65536.0,1,-nbitq), 
to_sfixed(6936.0/65536.0,1,-nbitq), 
to_sfixed(-851.0/65536.0,1,-nbitq), 
to_sfixed(-2601.0/65536.0,1,-nbitq), 
to_sfixed(790.0/65536.0,1,-nbitq), 
to_sfixed(7803.0/65536.0,1,-nbitq), 
to_sfixed(15648.0/65536.0,1,-nbitq), 
to_sfixed(107.0/65536.0,1,-nbitq), 
to_sfixed(-291.0/65536.0,1,-nbitq), 
to_sfixed(1725.0/65536.0,1,-nbitq), 
to_sfixed(-12368.0/65536.0,1,-nbitq), 
to_sfixed(-5871.0/65536.0,1,-nbitq), 
to_sfixed(623.0/65536.0,1,-nbitq), 
to_sfixed(-4514.0/65536.0,1,-nbitq), 
to_sfixed(-9269.0/65536.0,1,-nbitq), 
to_sfixed(200.0/65536.0,1,-nbitq), 
to_sfixed(2633.0/65536.0,1,-nbitq), 
to_sfixed(10749.0/65536.0,1,-nbitq), 
to_sfixed(-836.0/65536.0,1,-nbitq), 
to_sfixed(-1009.0/65536.0,1,-nbitq), 
to_sfixed(2143.0/65536.0,1,-nbitq), 
to_sfixed(2633.0/65536.0,1,-nbitq), 
to_sfixed(-8580.0/65536.0,1,-nbitq), 
to_sfixed(-11969.0/65536.0,1,-nbitq), 
to_sfixed(2873.0/65536.0,1,-nbitq), 
to_sfixed(-7100.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3191.0/65536.0,1,-nbitq), 
to_sfixed(-4273.0/65536.0,1,-nbitq), 
to_sfixed(-9828.0/65536.0,1,-nbitq), 
to_sfixed(15568.0/65536.0,1,-nbitq), 
to_sfixed(17749.0/65536.0,1,-nbitq), 
to_sfixed(-4289.0/65536.0,1,-nbitq), 
to_sfixed(-448.0/65536.0,1,-nbitq), 
to_sfixed(-3310.0/65536.0,1,-nbitq), 
to_sfixed(-2882.0/65536.0,1,-nbitq), 
to_sfixed(-598.0/65536.0,1,-nbitq), 
to_sfixed(3453.0/65536.0,1,-nbitq), 
to_sfixed(20424.0/65536.0,1,-nbitq), 
to_sfixed(4029.0/65536.0,1,-nbitq), 
to_sfixed(-4898.0/65536.0,1,-nbitq), 
to_sfixed(-2823.0/65536.0,1,-nbitq), 
to_sfixed(2819.0/65536.0,1,-nbitq), 
to_sfixed(-2323.0/65536.0,1,-nbitq), 
to_sfixed(-12605.0/65536.0,1,-nbitq), 
to_sfixed(-9702.0/65536.0,1,-nbitq), 
to_sfixed(105.0/65536.0,1,-nbitq), 
to_sfixed(864.0/65536.0,1,-nbitq), 
to_sfixed(-16309.0/65536.0,1,-nbitq), 
to_sfixed(7358.0/65536.0,1,-nbitq), 
to_sfixed(10628.0/65536.0,1,-nbitq), 
to_sfixed(-1521.0/65536.0,1,-nbitq), 
to_sfixed(-798.0/65536.0,1,-nbitq), 
to_sfixed(29260.0/65536.0,1,-nbitq), 
to_sfixed(1049.0/65536.0,1,-nbitq), 
to_sfixed(4878.0/65536.0,1,-nbitq), 
to_sfixed(-3515.0/65536.0,1,-nbitq), 
to_sfixed(-2543.0/65536.0,1,-nbitq), 
to_sfixed(11807.0/65536.0,1,-nbitq), 
to_sfixed(8892.0/65536.0,1,-nbitq), 
to_sfixed(5923.0/65536.0,1,-nbitq), 
to_sfixed(2070.0/65536.0,1,-nbitq), 
to_sfixed(399.0/65536.0,1,-nbitq), 
to_sfixed(8145.0/65536.0,1,-nbitq), 
to_sfixed(-4919.0/65536.0,1,-nbitq), 
to_sfixed(-18099.0/65536.0,1,-nbitq), 
to_sfixed(-95.0/65536.0,1,-nbitq), 
to_sfixed(-768.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(4744.0/65536.0,1,-nbitq), 
to_sfixed(5307.0/65536.0,1,-nbitq), 
to_sfixed(-37.0/65536.0,1,-nbitq), 
to_sfixed(8610.0/65536.0,1,-nbitq), 
to_sfixed(1143.0/65536.0,1,-nbitq), 
to_sfixed(-10653.0/65536.0,1,-nbitq), 
to_sfixed(-1392.0/65536.0,1,-nbitq), 
to_sfixed(2365.0/65536.0,1,-nbitq), 
to_sfixed(1517.0/65536.0,1,-nbitq), 
to_sfixed(3210.0/65536.0,1,-nbitq), 
to_sfixed(-7183.0/65536.0,1,-nbitq), 
to_sfixed(7245.0/65536.0,1,-nbitq), 
to_sfixed(1624.0/65536.0,1,-nbitq), 
to_sfixed(2841.0/65536.0,1,-nbitq), 
to_sfixed(2772.0/65536.0,1,-nbitq), 
to_sfixed(-5680.0/65536.0,1,-nbitq), 
to_sfixed(2197.0/65536.0,1,-nbitq), 
to_sfixed(-2059.0/65536.0,1,-nbitq), 
to_sfixed(7027.0/65536.0,1,-nbitq), 
to_sfixed(2320.0/65536.0,1,-nbitq), 
to_sfixed(613.0/65536.0,1,-nbitq), 
to_sfixed(47.0/65536.0,1,-nbitq), 
to_sfixed(-13836.0/65536.0,1,-nbitq), 
to_sfixed(-22582.0/65536.0,1,-nbitq), 
to_sfixed(-2089.0/65536.0,1,-nbitq), 
to_sfixed(-8061.0/65536.0,1,-nbitq), 
to_sfixed(-14858.0/65536.0,1,-nbitq), 
to_sfixed(9414.0/65536.0,1,-nbitq), 
to_sfixed(-1111.0/65536.0,1,-nbitq), 
to_sfixed(14849.0/65536.0,1,-nbitq), 
to_sfixed(-5077.0/65536.0,1,-nbitq), 
to_sfixed(1110.0/65536.0,1,-nbitq), 
to_sfixed(-1955.0/65536.0,1,-nbitq), 
to_sfixed(-12210.0/65536.0,1,-nbitq), 
to_sfixed(-8231.0/65536.0,1,-nbitq), 
to_sfixed(7333.0/65536.0,1,-nbitq), 
to_sfixed(2521.0/65536.0,1,-nbitq), 
to_sfixed(-5935.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-5998.0/65536.0,1,-nbitq), 
to_sfixed(-3896.0/65536.0,1,-nbitq), 
to_sfixed(-13678.0/65536.0,1,-nbitq), 
to_sfixed(9226.0/65536.0,1,-nbitq), 
to_sfixed(32955.0/65536.0,1,-nbitq), 
to_sfixed(-10379.0/65536.0,1,-nbitq), 
to_sfixed(2263.0/65536.0,1,-nbitq), 
to_sfixed(3447.0/65536.0,1,-nbitq), 
to_sfixed(4400.0/65536.0,1,-nbitq), 
to_sfixed(2260.0/65536.0,1,-nbitq), 
to_sfixed(2515.0/65536.0,1,-nbitq), 
to_sfixed(20207.0/65536.0,1,-nbitq), 
to_sfixed(3323.0/65536.0,1,-nbitq), 
to_sfixed(-5462.0/65536.0,1,-nbitq), 
to_sfixed(-5305.0/65536.0,1,-nbitq), 
to_sfixed(714.0/65536.0,1,-nbitq), 
to_sfixed(-2480.0/65536.0,1,-nbitq), 
to_sfixed(-7375.0/65536.0,1,-nbitq), 
to_sfixed(-10018.0/65536.0,1,-nbitq), 
to_sfixed(1545.0/65536.0,1,-nbitq), 
to_sfixed(6729.0/65536.0,1,-nbitq), 
to_sfixed(-22686.0/65536.0,1,-nbitq), 
to_sfixed(9096.0/65536.0,1,-nbitq), 
to_sfixed(13872.0/65536.0,1,-nbitq), 
to_sfixed(-1596.0/65536.0,1,-nbitq), 
to_sfixed(-1938.0/65536.0,1,-nbitq), 
to_sfixed(22270.0/65536.0,1,-nbitq), 
to_sfixed(-1561.0/65536.0,1,-nbitq), 
to_sfixed(120.0/65536.0,1,-nbitq), 
to_sfixed(-1084.0/65536.0,1,-nbitq), 
to_sfixed(-705.0/65536.0,1,-nbitq), 
to_sfixed(10114.0/65536.0,1,-nbitq), 
to_sfixed(4138.0/65536.0,1,-nbitq), 
to_sfixed(-6772.0/65536.0,1,-nbitq), 
to_sfixed(2885.0/65536.0,1,-nbitq), 
to_sfixed(2941.0/65536.0,1,-nbitq), 
to_sfixed(243.0/65536.0,1,-nbitq), 
to_sfixed(605.0/65536.0,1,-nbitq), 
to_sfixed(-9116.0/65536.0,1,-nbitq), 
to_sfixed(-3047.0/65536.0,1,-nbitq), 
to_sfixed(2892.0/65536.0,1,-nbitq), 
to_sfixed(1123.0/65536.0,1,-nbitq), 
to_sfixed(5252.0/65536.0,1,-nbitq), 
to_sfixed(6808.0/65536.0,1,-nbitq), 
to_sfixed(-2448.0/65536.0,1,-nbitq), 
to_sfixed(7404.0/65536.0,1,-nbitq), 
to_sfixed(-2276.0/65536.0,1,-nbitq), 
to_sfixed(-8273.0/65536.0,1,-nbitq), 
to_sfixed(137.0/65536.0,1,-nbitq), 
to_sfixed(-1431.0/65536.0,1,-nbitq), 
to_sfixed(1118.0/65536.0,1,-nbitq), 
to_sfixed(4485.0/65536.0,1,-nbitq), 
to_sfixed(-2394.0/65536.0,1,-nbitq), 
to_sfixed(7540.0/65536.0,1,-nbitq), 
to_sfixed(576.0/65536.0,1,-nbitq), 
to_sfixed(8137.0/65536.0,1,-nbitq), 
to_sfixed(2134.0/65536.0,1,-nbitq), 
to_sfixed(67.0/65536.0,1,-nbitq), 
to_sfixed(-1119.0/65536.0,1,-nbitq), 
to_sfixed(955.0/65536.0,1,-nbitq), 
to_sfixed(-2191.0/65536.0,1,-nbitq), 
to_sfixed(978.0/65536.0,1,-nbitq), 
to_sfixed(-129.0/65536.0,1,-nbitq), 
to_sfixed(-1776.0/65536.0,1,-nbitq), 
to_sfixed(-18191.0/65536.0,1,-nbitq), 
to_sfixed(-10941.0/65536.0,1,-nbitq), 
to_sfixed(-12266.0/65536.0,1,-nbitq), 
to_sfixed(-9804.0/65536.0,1,-nbitq), 
to_sfixed(-15318.0/65536.0,1,-nbitq), 
to_sfixed(10184.0/65536.0,1,-nbitq), 
to_sfixed(-1571.0/65536.0,1,-nbitq), 
to_sfixed(7810.0/65536.0,1,-nbitq), 
to_sfixed(-3512.0/65536.0,1,-nbitq), 
to_sfixed(-2960.0/65536.0,1,-nbitq), 
to_sfixed(-1768.0/65536.0,1,-nbitq), 
to_sfixed(-18555.0/65536.0,1,-nbitq), 
to_sfixed(-8353.0/65536.0,1,-nbitq), 
to_sfixed(9937.0/65536.0,1,-nbitq), 
to_sfixed(2471.0/65536.0,1,-nbitq), 
to_sfixed(-5939.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-5955.0/65536.0,1,-nbitq), 
to_sfixed(-30.0/65536.0,1,-nbitq), 
to_sfixed(5947.0/65536.0,1,-nbitq), 
to_sfixed(-297.0/65536.0,1,-nbitq), 
to_sfixed(10024.0/65536.0,1,-nbitq), 
to_sfixed(-14272.0/65536.0,1,-nbitq), 
to_sfixed(-614.0/65536.0,1,-nbitq), 
to_sfixed(9191.0/65536.0,1,-nbitq), 
to_sfixed(2749.0/65536.0,1,-nbitq), 
to_sfixed(2877.0/65536.0,1,-nbitq), 
to_sfixed(4306.0/65536.0,1,-nbitq), 
to_sfixed(14549.0/65536.0,1,-nbitq), 
to_sfixed(-2979.0/65536.0,1,-nbitq), 
to_sfixed(-12277.0/65536.0,1,-nbitq), 
to_sfixed(-3060.0/65536.0,1,-nbitq), 
to_sfixed(-430.0/65536.0,1,-nbitq), 
to_sfixed(-777.0/65536.0,1,-nbitq), 
to_sfixed(2151.0/65536.0,1,-nbitq), 
to_sfixed(-7053.0/65536.0,1,-nbitq), 
to_sfixed(-1795.0/65536.0,1,-nbitq), 
to_sfixed(4139.0/65536.0,1,-nbitq), 
to_sfixed(-17535.0/65536.0,1,-nbitq), 
to_sfixed(-4693.0/65536.0,1,-nbitq), 
to_sfixed(6203.0/65536.0,1,-nbitq), 
to_sfixed(1478.0/65536.0,1,-nbitq), 
to_sfixed(898.0/65536.0,1,-nbitq), 
to_sfixed(17511.0/65536.0,1,-nbitq), 
to_sfixed(1270.0/65536.0,1,-nbitq), 
to_sfixed(-10494.0/65536.0,1,-nbitq), 
to_sfixed(3052.0/65536.0,1,-nbitq), 
to_sfixed(-5993.0/65536.0,1,-nbitq), 
to_sfixed(7196.0/65536.0,1,-nbitq), 
to_sfixed(-1346.0/65536.0,1,-nbitq), 
to_sfixed(-5528.0/65536.0,1,-nbitq), 
to_sfixed(-2314.0/65536.0,1,-nbitq), 
to_sfixed(3166.0/65536.0,1,-nbitq), 
to_sfixed(-1520.0/65536.0,1,-nbitq), 
to_sfixed(-809.0/65536.0,1,-nbitq), 
to_sfixed(9880.0/65536.0,1,-nbitq), 
to_sfixed(2132.0/65536.0,1,-nbitq), 
to_sfixed(2830.0/65536.0,1,-nbitq), 
to_sfixed(-605.0/65536.0,1,-nbitq), 
to_sfixed(6196.0/65536.0,1,-nbitq), 
to_sfixed(731.0/65536.0,1,-nbitq), 
to_sfixed(2155.0/65536.0,1,-nbitq), 
to_sfixed(11682.0/65536.0,1,-nbitq), 
to_sfixed(-123.0/65536.0,1,-nbitq), 
to_sfixed(-4763.0/65536.0,1,-nbitq), 
to_sfixed(1532.0/65536.0,1,-nbitq), 
to_sfixed(2181.0/65536.0,1,-nbitq), 
to_sfixed(-1634.0/65536.0,1,-nbitq), 
to_sfixed(11760.0/65536.0,1,-nbitq), 
to_sfixed(-6419.0/65536.0,1,-nbitq), 
to_sfixed(-3982.0/65536.0,1,-nbitq), 
to_sfixed(-26.0/65536.0,1,-nbitq), 
to_sfixed(6916.0/65536.0,1,-nbitq), 
to_sfixed(1472.0/65536.0,1,-nbitq), 
to_sfixed(-1699.0/65536.0,1,-nbitq), 
to_sfixed(-1990.0/65536.0,1,-nbitq), 
to_sfixed(9050.0/65536.0,1,-nbitq), 
to_sfixed(-1862.0/65536.0,1,-nbitq), 
to_sfixed(-15.0/65536.0,1,-nbitq), 
to_sfixed(111.0/65536.0,1,-nbitq), 
to_sfixed(2270.0/65536.0,1,-nbitq), 
to_sfixed(-14249.0/65536.0,1,-nbitq), 
to_sfixed(4123.0/65536.0,1,-nbitq), 
to_sfixed(-10089.0/65536.0,1,-nbitq), 
to_sfixed(-3880.0/65536.0,1,-nbitq), 
to_sfixed(-4376.0/65536.0,1,-nbitq), 
to_sfixed(5537.0/65536.0,1,-nbitq), 
to_sfixed(453.0/65536.0,1,-nbitq), 
to_sfixed(8072.0/65536.0,1,-nbitq), 
to_sfixed(-9867.0/65536.0,1,-nbitq), 
to_sfixed(1602.0/65536.0,1,-nbitq), 
to_sfixed(-531.0/65536.0,1,-nbitq), 
to_sfixed(-15937.0/65536.0,1,-nbitq), 
to_sfixed(-4746.0/65536.0,1,-nbitq), 
to_sfixed(2966.0/65536.0,1,-nbitq), 
to_sfixed(-1296.0/65536.0,1,-nbitq), 
to_sfixed(1959.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-9343.0/65536.0,1,-nbitq), 
to_sfixed(1146.0/65536.0,1,-nbitq), 
to_sfixed(11762.0/65536.0,1,-nbitq), 
to_sfixed(-5166.0/65536.0,1,-nbitq), 
to_sfixed(-2993.0/65536.0,1,-nbitq), 
to_sfixed(2379.0/65536.0,1,-nbitq), 
to_sfixed(1838.0/65536.0,1,-nbitq), 
to_sfixed(11598.0/65536.0,1,-nbitq), 
to_sfixed(444.0/65536.0,1,-nbitq), 
to_sfixed(-1859.0/65536.0,1,-nbitq), 
to_sfixed(5358.0/65536.0,1,-nbitq), 
to_sfixed(16268.0/65536.0,1,-nbitq), 
to_sfixed(1017.0/65536.0,1,-nbitq), 
to_sfixed(-4994.0/65536.0,1,-nbitq), 
to_sfixed(-1605.0/65536.0,1,-nbitq), 
to_sfixed(3018.0/65536.0,1,-nbitq), 
to_sfixed(1978.0/65536.0,1,-nbitq), 
to_sfixed(522.0/65536.0,1,-nbitq), 
to_sfixed(3818.0/65536.0,1,-nbitq), 
to_sfixed(-2357.0/65536.0,1,-nbitq), 
to_sfixed(-1193.0/65536.0,1,-nbitq), 
to_sfixed(-17483.0/65536.0,1,-nbitq), 
to_sfixed(-13471.0/65536.0,1,-nbitq), 
to_sfixed(-2592.0/65536.0,1,-nbitq), 
to_sfixed(-3329.0/65536.0,1,-nbitq), 
to_sfixed(-2646.0/65536.0,1,-nbitq), 
to_sfixed(17753.0/65536.0,1,-nbitq), 
to_sfixed(-1601.0/65536.0,1,-nbitq), 
to_sfixed(-2631.0/65536.0,1,-nbitq), 
to_sfixed(5409.0/65536.0,1,-nbitq), 
to_sfixed(-4582.0/65536.0,1,-nbitq), 
to_sfixed(-180.0/65536.0,1,-nbitq), 
to_sfixed(-11198.0/65536.0,1,-nbitq), 
to_sfixed(-474.0/65536.0,1,-nbitq), 
to_sfixed(-319.0/65536.0,1,-nbitq), 
to_sfixed(2402.0/65536.0,1,-nbitq), 
to_sfixed(-1086.0/65536.0,1,-nbitq), 
to_sfixed(8656.0/65536.0,1,-nbitq), 
to_sfixed(316.0/65536.0,1,-nbitq), 
to_sfixed(2392.0/65536.0,1,-nbitq), 
to_sfixed(-8326.0/65536.0,1,-nbitq), 
to_sfixed(-3070.0/65536.0,1,-nbitq), 
to_sfixed(-802.0/65536.0,1,-nbitq), 
to_sfixed(-171.0/65536.0,1,-nbitq), 
to_sfixed(-1705.0/65536.0,1,-nbitq), 
to_sfixed(11664.0/65536.0,1,-nbitq), 
to_sfixed(-3639.0/65536.0,1,-nbitq), 
to_sfixed(-1652.0/65536.0,1,-nbitq), 
to_sfixed(2605.0/65536.0,1,-nbitq), 
to_sfixed(275.0/65536.0,1,-nbitq), 
to_sfixed(-1310.0/65536.0,1,-nbitq), 
to_sfixed(7312.0/65536.0,1,-nbitq), 
to_sfixed(-1399.0/65536.0,1,-nbitq), 
to_sfixed(3024.0/65536.0,1,-nbitq), 
to_sfixed(3095.0/65536.0,1,-nbitq), 
to_sfixed(-21146.0/65536.0,1,-nbitq), 
to_sfixed(3864.0/65536.0,1,-nbitq), 
to_sfixed(1677.0/65536.0,1,-nbitq), 
to_sfixed(830.0/65536.0,1,-nbitq), 
to_sfixed(5500.0/65536.0,1,-nbitq), 
to_sfixed(3507.0/65536.0,1,-nbitq), 
to_sfixed(276.0/65536.0,1,-nbitq), 
to_sfixed(-830.0/65536.0,1,-nbitq), 
to_sfixed(496.0/65536.0,1,-nbitq), 
to_sfixed(-14316.0/65536.0,1,-nbitq), 
to_sfixed(4710.0/65536.0,1,-nbitq), 
to_sfixed(-1339.0/65536.0,1,-nbitq), 
to_sfixed(-4058.0/65536.0,1,-nbitq), 
to_sfixed(-1843.0/65536.0,1,-nbitq), 
to_sfixed(8877.0/65536.0,1,-nbitq), 
to_sfixed(1758.0/65536.0,1,-nbitq), 
to_sfixed(6781.0/65536.0,1,-nbitq), 
to_sfixed(-9728.0/65536.0,1,-nbitq), 
to_sfixed(596.0/65536.0,1,-nbitq), 
to_sfixed(-2736.0/65536.0,1,-nbitq), 
to_sfixed(-9142.0/65536.0,1,-nbitq), 
to_sfixed(-927.0/65536.0,1,-nbitq), 
to_sfixed(5203.0/65536.0,1,-nbitq), 
to_sfixed(734.0/65536.0,1,-nbitq), 
to_sfixed(10699.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-8860.0/65536.0,1,-nbitq), 
to_sfixed(779.0/65536.0,1,-nbitq), 
to_sfixed(8092.0/65536.0,1,-nbitq), 
to_sfixed(-2563.0/65536.0,1,-nbitq), 
to_sfixed(-5777.0/65536.0,1,-nbitq), 
to_sfixed(16904.0/65536.0,1,-nbitq), 
to_sfixed(2099.0/65536.0,1,-nbitq), 
to_sfixed(9102.0/65536.0,1,-nbitq), 
to_sfixed(5539.0/65536.0,1,-nbitq), 
to_sfixed(318.0/65536.0,1,-nbitq), 
to_sfixed(3392.0/65536.0,1,-nbitq), 
to_sfixed(5286.0/65536.0,1,-nbitq), 
to_sfixed(629.0/65536.0,1,-nbitq), 
to_sfixed(233.0/65536.0,1,-nbitq), 
to_sfixed(2216.0/65536.0,1,-nbitq), 
to_sfixed(1087.0/65536.0,1,-nbitq), 
to_sfixed(2879.0/65536.0,1,-nbitq), 
to_sfixed(-6734.0/65536.0,1,-nbitq), 
to_sfixed(4553.0/65536.0,1,-nbitq), 
to_sfixed(1490.0/65536.0,1,-nbitq), 
to_sfixed(-3685.0/65536.0,1,-nbitq), 
to_sfixed(-11951.0/65536.0,1,-nbitq), 
to_sfixed(-15710.0/65536.0,1,-nbitq), 
to_sfixed(589.0/65536.0,1,-nbitq), 
to_sfixed(-3199.0/65536.0,1,-nbitq), 
to_sfixed(2284.0/65536.0,1,-nbitq), 
to_sfixed(15421.0/65536.0,1,-nbitq), 
to_sfixed(1314.0/65536.0,1,-nbitq), 
to_sfixed(5508.0/65536.0,1,-nbitq), 
to_sfixed(7752.0/65536.0,1,-nbitq), 
to_sfixed(-4369.0/65536.0,1,-nbitq), 
to_sfixed(-1351.0/65536.0,1,-nbitq), 
to_sfixed(-14877.0/65536.0,1,-nbitq), 
to_sfixed(-3450.0/65536.0,1,-nbitq), 
to_sfixed(734.0/65536.0,1,-nbitq), 
to_sfixed(738.0/65536.0,1,-nbitq), 
to_sfixed(11026.0/65536.0,1,-nbitq), 
to_sfixed(9063.0/65536.0,1,-nbitq), 
to_sfixed(1536.0/65536.0,1,-nbitq), 
to_sfixed(1474.0/65536.0,1,-nbitq), 
to_sfixed(3860.0/65536.0,1,-nbitq), 
to_sfixed(1331.0/65536.0,1,-nbitq), 
to_sfixed(-1227.0/65536.0,1,-nbitq), 
to_sfixed(134.0/65536.0,1,-nbitq), 
to_sfixed(779.0/65536.0,1,-nbitq), 
to_sfixed(-3452.0/65536.0,1,-nbitq), 
to_sfixed(-1660.0/65536.0,1,-nbitq), 
to_sfixed(4112.0/65536.0,1,-nbitq), 
to_sfixed(-1697.0/65536.0,1,-nbitq), 
to_sfixed(-770.0/65536.0,1,-nbitq), 
to_sfixed(1815.0/65536.0,1,-nbitq), 
to_sfixed(1978.0/65536.0,1,-nbitq), 
to_sfixed(-9089.0/65536.0,1,-nbitq), 
to_sfixed(-5756.0/65536.0,1,-nbitq), 
to_sfixed(8276.0/65536.0,1,-nbitq), 
to_sfixed(-17632.0/65536.0,1,-nbitq), 
to_sfixed(-1294.0/65536.0,1,-nbitq), 
to_sfixed(540.0/65536.0,1,-nbitq), 
to_sfixed(-2031.0/65536.0,1,-nbitq), 
to_sfixed(-163.0/65536.0,1,-nbitq), 
to_sfixed(-177.0/65536.0,1,-nbitq), 
to_sfixed(-2465.0/65536.0,1,-nbitq), 
to_sfixed(-2288.0/65536.0,1,-nbitq), 
to_sfixed(-2342.0/65536.0,1,-nbitq), 
to_sfixed(-7986.0/65536.0,1,-nbitq), 
to_sfixed(5301.0/65536.0,1,-nbitq), 
to_sfixed(4843.0/65536.0,1,-nbitq), 
to_sfixed(-6079.0/65536.0,1,-nbitq), 
to_sfixed(910.0/65536.0,1,-nbitq), 
to_sfixed(7242.0/65536.0,1,-nbitq), 
to_sfixed(-321.0/65536.0,1,-nbitq), 
to_sfixed(2481.0/65536.0,1,-nbitq), 
to_sfixed(11149.0/65536.0,1,-nbitq), 
to_sfixed(-2934.0/65536.0,1,-nbitq), 
to_sfixed(-1597.0/65536.0,1,-nbitq), 
to_sfixed(-4495.0/65536.0,1,-nbitq), 
to_sfixed(-5462.0/65536.0,1,-nbitq), 
to_sfixed(13657.0/65536.0,1,-nbitq), 
to_sfixed(-1999.0/65536.0,1,-nbitq), 
to_sfixed(9037.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-5473.0/65536.0,1,-nbitq), 
to_sfixed(3491.0/65536.0,1,-nbitq), 
to_sfixed(2117.0/65536.0,1,-nbitq), 
to_sfixed(-2198.0/65536.0,1,-nbitq), 
to_sfixed(357.0/65536.0,1,-nbitq), 
to_sfixed(20393.0/65536.0,1,-nbitq), 
to_sfixed(2378.0/65536.0,1,-nbitq), 
to_sfixed(9167.0/65536.0,1,-nbitq), 
to_sfixed(8779.0/65536.0,1,-nbitq), 
to_sfixed(96.0/65536.0,1,-nbitq), 
to_sfixed(5917.0/65536.0,1,-nbitq), 
to_sfixed(-5325.0/65536.0,1,-nbitq), 
to_sfixed(-1941.0/65536.0,1,-nbitq), 
to_sfixed(4488.0/65536.0,1,-nbitq), 
to_sfixed(2748.0/65536.0,1,-nbitq), 
to_sfixed(911.0/65536.0,1,-nbitq), 
to_sfixed(-598.0/65536.0,1,-nbitq), 
to_sfixed(1507.0/65536.0,1,-nbitq), 
to_sfixed(3419.0/65536.0,1,-nbitq), 
to_sfixed(1682.0/65536.0,1,-nbitq), 
to_sfixed(2392.0/65536.0,1,-nbitq), 
to_sfixed(-14636.0/65536.0,1,-nbitq), 
to_sfixed(-13896.0/65536.0,1,-nbitq), 
to_sfixed(-39.0/65536.0,1,-nbitq), 
to_sfixed(246.0/65536.0,1,-nbitq), 
to_sfixed(15481.0/65536.0,1,-nbitq), 
to_sfixed(4177.0/65536.0,1,-nbitq), 
to_sfixed(2194.0/65536.0,1,-nbitq), 
to_sfixed(9239.0/65536.0,1,-nbitq), 
to_sfixed(2556.0/65536.0,1,-nbitq), 
to_sfixed(-6367.0/65536.0,1,-nbitq), 
to_sfixed(-3084.0/65536.0,1,-nbitq), 
to_sfixed(-16003.0/65536.0,1,-nbitq), 
to_sfixed(236.0/65536.0,1,-nbitq), 
to_sfixed(752.0/65536.0,1,-nbitq), 
to_sfixed(808.0/65536.0,1,-nbitq), 
to_sfixed(8857.0/65536.0,1,-nbitq), 
to_sfixed(-3194.0/65536.0,1,-nbitq), 
to_sfixed(1494.0/65536.0,1,-nbitq), 
to_sfixed(237.0/65536.0,1,-nbitq), 
to_sfixed(10134.0/65536.0,1,-nbitq), 
to_sfixed(1297.0/65536.0,1,-nbitq), 
to_sfixed(8978.0/65536.0,1,-nbitq), 
to_sfixed(-784.0/65536.0,1,-nbitq), 
to_sfixed(2888.0/65536.0,1,-nbitq), 
to_sfixed(-15236.0/65536.0,1,-nbitq), 
to_sfixed(391.0/65536.0,1,-nbitq), 
to_sfixed(6823.0/65536.0,1,-nbitq), 
to_sfixed(-1609.0/65536.0,1,-nbitq), 
to_sfixed(1258.0/65536.0,1,-nbitq), 
to_sfixed(-2537.0/65536.0,1,-nbitq), 
to_sfixed(-3404.0/65536.0,1,-nbitq), 
to_sfixed(-4315.0/65536.0,1,-nbitq), 
to_sfixed(-469.0/65536.0,1,-nbitq), 
to_sfixed(12878.0/65536.0,1,-nbitq), 
to_sfixed(-3152.0/65536.0,1,-nbitq), 
to_sfixed(2071.0/65536.0,1,-nbitq), 
to_sfixed(-4090.0/65536.0,1,-nbitq), 
to_sfixed(1489.0/65536.0,1,-nbitq), 
to_sfixed(4605.0/65536.0,1,-nbitq), 
to_sfixed(-3811.0/65536.0,1,-nbitq), 
to_sfixed(-1757.0/65536.0,1,-nbitq), 
to_sfixed(2075.0/65536.0,1,-nbitq), 
to_sfixed(1972.0/65536.0,1,-nbitq), 
to_sfixed(-3600.0/65536.0,1,-nbitq), 
to_sfixed(15564.0/65536.0,1,-nbitq), 
to_sfixed(-2795.0/65536.0,1,-nbitq), 
to_sfixed(-439.0/65536.0,1,-nbitq), 
to_sfixed(-10185.0/65536.0,1,-nbitq), 
to_sfixed(668.0/65536.0,1,-nbitq), 
to_sfixed(1626.0/65536.0,1,-nbitq), 
to_sfixed(-732.0/65536.0,1,-nbitq), 
to_sfixed(24141.0/65536.0,1,-nbitq), 
to_sfixed(2386.0/65536.0,1,-nbitq), 
to_sfixed(256.0/65536.0,1,-nbitq), 
to_sfixed(394.0/65536.0,1,-nbitq), 
to_sfixed(-11755.0/65536.0,1,-nbitq), 
to_sfixed(-4255.0/65536.0,1,-nbitq), 
to_sfixed(-3529.0/65536.0,1,-nbitq), 
to_sfixed(8864.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3010.0/65536.0,1,-nbitq), 
to_sfixed(4965.0/65536.0,1,-nbitq), 
to_sfixed(4418.0/65536.0,1,-nbitq), 
to_sfixed(7207.0/65536.0,1,-nbitq), 
to_sfixed(-4592.0/65536.0,1,-nbitq), 
to_sfixed(14658.0/65536.0,1,-nbitq), 
to_sfixed(-76.0/65536.0,1,-nbitq), 
to_sfixed(6264.0/65536.0,1,-nbitq), 
to_sfixed(5661.0/65536.0,1,-nbitq), 
to_sfixed(2631.0/65536.0,1,-nbitq), 
to_sfixed(663.0/65536.0,1,-nbitq), 
to_sfixed(3208.0/65536.0,1,-nbitq), 
to_sfixed(-315.0/65536.0,1,-nbitq), 
to_sfixed(9316.0/65536.0,1,-nbitq), 
to_sfixed(413.0/65536.0,1,-nbitq), 
to_sfixed(2671.0/65536.0,1,-nbitq), 
to_sfixed(1977.0/65536.0,1,-nbitq), 
to_sfixed(2350.0/65536.0,1,-nbitq), 
to_sfixed(-38.0/65536.0,1,-nbitq), 
to_sfixed(2479.0/65536.0,1,-nbitq), 
to_sfixed(1647.0/65536.0,1,-nbitq), 
to_sfixed(-5918.0/65536.0,1,-nbitq), 
to_sfixed(-10719.0/65536.0,1,-nbitq), 
to_sfixed(117.0/65536.0,1,-nbitq), 
to_sfixed(-4474.0/65536.0,1,-nbitq), 
to_sfixed(16348.0/65536.0,1,-nbitq), 
to_sfixed(-648.0/65536.0,1,-nbitq), 
to_sfixed(-1343.0/65536.0,1,-nbitq), 
to_sfixed(9513.0/65536.0,1,-nbitq), 
to_sfixed(-1338.0/65536.0,1,-nbitq), 
to_sfixed(-2285.0/65536.0,1,-nbitq), 
to_sfixed(-7717.0/65536.0,1,-nbitq), 
to_sfixed(-14862.0/65536.0,1,-nbitq), 
to_sfixed(5094.0/65536.0,1,-nbitq), 
to_sfixed(-2702.0/65536.0,1,-nbitq), 
to_sfixed(2593.0/65536.0,1,-nbitq), 
to_sfixed(4816.0/65536.0,1,-nbitq), 
to_sfixed(-3696.0/65536.0,1,-nbitq), 
to_sfixed(2843.0/65536.0,1,-nbitq), 
to_sfixed(-2116.0/65536.0,1,-nbitq), 
to_sfixed(7694.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(7746.0/65536.0,1,-nbitq), 
to_sfixed(-5201.0/65536.0,1,-nbitq), 
to_sfixed(-2903.0/65536.0,1,-nbitq), 
to_sfixed(-21270.0/65536.0,1,-nbitq), 
to_sfixed(1865.0/65536.0,1,-nbitq), 
to_sfixed(3388.0/65536.0,1,-nbitq), 
to_sfixed(2021.0/65536.0,1,-nbitq), 
to_sfixed(-1101.0/65536.0,1,-nbitq), 
to_sfixed(2141.0/65536.0,1,-nbitq), 
to_sfixed(81.0/65536.0,1,-nbitq), 
to_sfixed(1623.0/65536.0,1,-nbitq), 
to_sfixed(-1602.0/65536.0,1,-nbitq), 
to_sfixed(13479.0/65536.0,1,-nbitq), 
to_sfixed(-2790.0/65536.0,1,-nbitq), 
to_sfixed(-2747.0/65536.0,1,-nbitq), 
to_sfixed(-4228.0/65536.0,1,-nbitq), 
to_sfixed(-2610.0/65536.0,1,-nbitq), 
to_sfixed(1740.0/65536.0,1,-nbitq), 
to_sfixed(-7900.0/65536.0,1,-nbitq), 
to_sfixed(2537.0/65536.0,1,-nbitq), 
to_sfixed(2828.0/65536.0,1,-nbitq), 
to_sfixed(-1061.0/65536.0,1,-nbitq), 
to_sfixed(298.0/65536.0,1,-nbitq), 
to_sfixed(7565.0/65536.0,1,-nbitq), 
to_sfixed(-1375.0/65536.0,1,-nbitq), 
to_sfixed(3149.0/65536.0,1,-nbitq), 
to_sfixed(-4666.0/65536.0,1,-nbitq), 
to_sfixed(-1332.0/65536.0,1,-nbitq), 
to_sfixed(4926.0/65536.0,1,-nbitq), 
to_sfixed(-3758.0/65536.0,1,-nbitq), 
to_sfixed(11897.0/65536.0,1,-nbitq), 
to_sfixed(2339.0/65536.0,1,-nbitq), 
to_sfixed(-1961.0/65536.0,1,-nbitq), 
to_sfixed(2189.0/65536.0,1,-nbitq), 
to_sfixed(-5202.0/65536.0,1,-nbitq), 
to_sfixed(-15089.0/65536.0,1,-nbitq), 
to_sfixed(1582.0/65536.0,1,-nbitq), 
to_sfixed(-591.0/65536.0,1,-nbitq)  ), 
( to_sfixed(184.0/65536.0,1,-nbitq), 
to_sfixed(-815.0/65536.0,1,-nbitq), 
to_sfixed(5477.0/65536.0,1,-nbitq), 
to_sfixed(8833.0/65536.0,1,-nbitq), 
to_sfixed(3853.0/65536.0,1,-nbitq), 
to_sfixed(13383.0/65536.0,1,-nbitq), 
to_sfixed(3096.0/65536.0,1,-nbitq), 
to_sfixed(4692.0/65536.0,1,-nbitq), 
to_sfixed(6975.0/65536.0,1,-nbitq), 
to_sfixed(1074.0/65536.0,1,-nbitq), 
to_sfixed(3058.0/65536.0,1,-nbitq), 
to_sfixed(5052.0/65536.0,1,-nbitq), 
to_sfixed(-891.0/65536.0,1,-nbitq), 
to_sfixed(9230.0/65536.0,1,-nbitq), 
to_sfixed(462.0/65536.0,1,-nbitq), 
to_sfixed(-2293.0/65536.0,1,-nbitq), 
to_sfixed(1657.0/65536.0,1,-nbitq), 
to_sfixed(-67.0/65536.0,1,-nbitq), 
to_sfixed(-57.0/65536.0,1,-nbitq), 
to_sfixed(-182.0/65536.0,1,-nbitq), 
to_sfixed(6276.0/65536.0,1,-nbitq), 
to_sfixed(-6014.0/65536.0,1,-nbitq), 
to_sfixed(-7327.0/65536.0,1,-nbitq), 
to_sfixed(1218.0/65536.0,1,-nbitq), 
to_sfixed(-1821.0/65536.0,1,-nbitq), 
to_sfixed(16508.0/65536.0,1,-nbitq), 
to_sfixed(3870.0/65536.0,1,-nbitq), 
to_sfixed(993.0/65536.0,1,-nbitq), 
to_sfixed(7717.0/65536.0,1,-nbitq), 
to_sfixed(-2590.0/65536.0,1,-nbitq), 
to_sfixed(3705.0/65536.0,1,-nbitq), 
to_sfixed(-12222.0/65536.0,1,-nbitq), 
to_sfixed(-7541.0/65536.0,1,-nbitq), 
to_sfixed(6596.0/65536.0,1,-nbitq), 
to_sfixed(-406.0/65536.0,1,-nbitq), 
to_sfixed(-664.0/65536.0,1,-nbitq), 
to_sfixed(81.0/65536.0,1,-nbitq), 
to_sfixed(-3408.0/65536.0,1,-nbitq), 
to_sfixed(-1646.0/65536.0,1,-nbitq), 
to_sfixed(-1917.0/65536.0,1,-nbitq), 
to_sfixed(6364.0/65536.0,1,-nbitq), 
to_sfixed(-2039.0/65536.0,1,-nbitq), 
to_sfixed(4655.0/65536.0,1,-nbitq), 
to_sfixed(-6699.0/65536.0,1,-nbitq), 
to_sfixed(-928.0/65536.0,1,-nbitq), 
to_sfixed(-5041.0/65536.0,1,-nbitq), 
to_sfixed(1397.0/65536.0,1,-nbitq), 
to_sfixed(1400.0/65536.0,1,-nbitq), 
to_sfixed(122.0/65536.0,1,-nbitq), 
to_sfixed(98.0/65536.0,1,-nbitq), 
to_sfixed(377.0/65536.0,1,-nbitq), 
to_sfixed(428.0/65536.0,1,-nbitq), 
to_sfixed(-2709.0/65536.0,1,-nbitq), 
to_sfixed(-1158.0/65536.0,1,-nbitq), 
to_sfixed(6030.0/65536.0,1,-nbitq), 
to_sfixed(364.0/65536.0,1,-nbitq), 
to_sfixed(-1707.0/65536.0,1,-nbitq), 
to_sfixed(1835.0/65536.0,1,-nbitq), 
to_sfixed(-1990.0/65536.0,1,-nbitq), 
to_sfixed(4066.0/65536.0,1,-nbitq), 
to_sfixed(-3564.0/65536.0,1,-nbitq), 
to_sfixed(-2430.0/65536.0,1,-nbitq), 
to_sfixed(-1741.0/65536.0,1,-nbitq), 
to_sfixed(1071.0/65536.0,1,-nbitq), 
to_sfixed(268.0/65536.0,1,-nbitq), 
to_sfixed(5198.0/65536.0,1,-nbitq), 
to_sfixed(-1614.0/65536.0,1,-nbitq), 
to_sfixed(8123.0/65536.0,1,-nbitq), 
to_sfixed(-3434.0/65536.0,1,-nbitq), 
to_sfixed(-13837.0/65536.0,1,-nbitq), 
to_sfixed(5521.0/65536.0,1,-nbitq), 
to_sfixed(-632.0/65536.0,1,-nbitq), 
to_sfixed(15287.0/65536.0,1,-nbitq), 
to_sfixed(-300.0/65536.0,1,-nbitq), 
to_sfixed(-378.0/65536.0,1,-nbitq), 
to_sfixed(-1844.0/65536.0,1,-nbitq), 
to_sfixed(-8360.0/65536.0,1,-nbitq), 
to_sfixed(-15880.0/65536.0,1,-nbitq), 
to_sfixed(-2929.0/65536.0,1,-nbitq), 
to_sfixed(-6422.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5063.0/65536.0,1,-nbitq), 
to_sfixed(3208.0/65536.0,1,-nbitq), 
to_sfixed(-3660.0/65536.0,1,-nbitq), 
to_sfixed(-388.0/65536.0,1,-nbitq), 
to_sfixed(4651.0/65536.0,1,-nbitq), 
to_sfixed(9452.0/65536.0,1,-nbitq), 
to_sfixed(104.0/65536.0,1,-nbitq), 
to_sfixed(887.0/65536.0,1,-nbitq), 
to_sfixed(-582.0/65536.0,1,-nbitq), 
to_sfixed(-2080.0/65536.0,1,-nbitq), 
to_sfixed(5034.0/65536.0,1,-nbitq), 
to_sfixed(-3158.0/65536.0,1,-nbitq), 
to_sfixed(-1084.0/65536.0,1,-nbitq), 
to_sfixed(534.0/65536.0,1,-nbitq), 
to_sfixed(-3911.0/65536.0,1,-nbitq), 
to_sfixed(-2478.0/65536.0,1,-nbitq), 
to_sfixed(2464.0/65536.0,1,-nbitq), 
to_sfixed(936.0/65536.0,1,-nbitq), 
to_sfixed(3325.0/65536.0,1,-nbitq), 
to_sfixed(1410.0/65536.0,1,-nbitq), 
to_sfixed(6587.0/65536.0,1,-nbitq), 
to_sfixed(-9926.0/65536.0,1,-nbitq), 
to_sfixed(-7188.0/65536.0,1,-nbitq), 
to_sfixed(2479.0/65536.0,1,-nbitq), 
to_sfixed(2392.0/65536.0,1,-nbitq), 
to_sfixed(8212.0/65536.0,1,-nbitq), 
to_sfixed(2974.0/65536.0,1,-nbitq), 
to_sfixed(1798.0/65536.0,1,-nbitq), 
to_sfixed(7958.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(3549.0/65536.0,1,-nbitq), 
to_sfixed(-8506.0/65536.0,1,-nbitq), 
to_sfixed(-551.0/65536.0,1,-nbitq), 
to_sfixed(17760.0/65536.0,1,-nbitq), 
to_sfixed(1227.0/65536.0,1,-nbitq), 
to_sfixed(76.0/65536.0,1,-nbitq), 
to_sfixed(460.0/65536.0,1,-nbitq), 
to_sfixed(-5859.0/65536.0,1,-nbitq), 
to_sfixed(165.0/65536.0,1,-nbitq), 
to_sfixed(3408.0/65536.0,1,-nbitq), 
to_sfixed(5345.0/65536.0,1,-nbitq), 
to_sfixed(-2247.0/65536.0,1,-nbitq), 
to_sfixed(9156.0/65536.0,1,-nbitq), 
to_sfixed(-2202.0/65536.0,1,-nbitq), 
to_sfixed(-1065.0/65536.0,1,-nbitq), 
to_sfixed(115.0/65536.0,1,-nbitq), 
to_sfixed(2600.0/65536.0,1,-nbitq), 
to_sfixed(-1228.0/65536.0,1,-nbitq), 
to_sfixed(1690.0/65536.0,1,-nbitq), 
to_sfixed(-2281.0/65536.0,1,-nbitq), 
to_sfixed(-644.0/65536.0,1,-nbitq), 
to_sfixed(5622.0/65536.0,1,-nbitq), 
to_sfixed(1696.0/65536.0,1,-nbitq), 
to_sfixed(-1545.0/65536.0,1,-nbitq), 
to_sfixed(5417.0/65536.0,1,-nbitq), 
to_sfixed(-1164.0/65536.0,1,-nbitq), 
to_sfixed(-2595.0/65536.0,1,-nbitq), 
to_sfixed(-1791.0/65536.0,1,-nbitq), 
to_sfixed(1597.0/65536.0,1,-nbitq), 
to_sfixed(2103.0/65536.0,1,-nbitq), 
to_sfixed(1856.0/65536.0,1,-nbitq), 
to_sfixed(1153.0/65536.0,1,-nbitq), 
to_sfixed(-2619.0/65536.0,1,-nbitq), 
to_sfixed(2589.0/65536.0,1,-nbitq), 
to_sfixed(2057.0/65536.0,1,-nbitq), 
to_sfixed(-2782.0/65536.0,1,-nbitq), 
to_sfixed(4284.0/65536.0,1,-nbitq), 
to_sfixed(3523.0/65536.0,1,-nbitq), 
to_sfixed(-1732.0/65536.0,1,-nbitq), 
to_sfixed(-14673.0/65536.0,1,-nbitq), 
to_sfixed(7621.0/65536.0,1,-nbitq), 
to_sfixed(-3064.0/65536.0,1,-nbitq), 
to_sfixed(8136.0/65536.0,1,-nbitq), 
to_sfixed(-1369.0/65536.0,1,-nbitq), 
to_sfixed(1052.0/65536.0,1,-nbitq), 
to_sfixed(1285.0/65536.0,1,-nbitq), 
to_sfixed(-5132.0/65536.0,1,-nbitq), 
to_sfixed(-10040.0/65536.0,1,-nbitq), 
to_sfixed(-1817.0/65536.0,1,-nbitq), 
to_sfixed(-11085.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2423.0/65536.0,1,-nbitq), 
to_sfixed(6362.0/65536.0,1,-nbitq), 
to_sfixed(-2814.0/65536.0,1,-nbitq), 
to_sfixed(2318.0/65536.0,1,-nbitq), 
to_sfixed(-4908.0/65536.0,1,-nbitq), 
to_sfixed(9393.0/65536.0,1,-nbitq), 
to_sfixed(-4303.0/65536.0,1,-nbitq), 
to_sfixed(8134.0/65536.0,1,-nbitq), 
to_sfixed(1234.0/65536.0,1,-nbitq), 
to_sfixed(-137.0/65536.0,1,-nbitq), 
to_sfixed(7817.0/65536.0,1,-nbitq), 
to_sfixed(-3083.0/65536.0,1,-nbitq), 
to_sfixed(691.0/65536.0,1,-nbitq), 
to_sfixed(7916.0/65536.0,1,-nbitq), 
to_sfixed(-4688.0/65536.0,1,-nbitq), 
to_sfixed(-1968.0/65536.0,1,-nbitq), 
to_sfixed(546.0/65536.0,1,-nbitq), 
to_sfixed(7547.0/65536.0,1,-nbitq), 
to_sfixed(1854.0/65536.0,1,-nbitq), 
to_sfixed(384.0/65536.0,1,-nbitq), 
to_sfixed(6926.0/65536.0,1,-nbitq), 
to_sfixed(-17350.0/65536.0,1,-nbitq), 
to_sfixed(-3591.0/65536.0,1,-nbitq), 
to_sfixed(3274.0/65536.0,1,-nbitq), 
to_sfixed(-435.0/65536.0,1,-nbitq), 
to_sfixed(7541.0/65536.0,1,-nbitq), 
to_sfixed(948.0/65536.0,1,-nbitq), 
to_sfixed(2600.0/65536.0,1,-nbitq), 
to_sfixed(5142.0/65536.0,1,-nbitq), 
to_sfixed(-4947.0/65536.0,1,-nbitq), 
to_sfixed(476.0/65536.0,1,-nbitq), 
to_sfixed(-9219.0/65536.0,1,-nbitq), 
to_sfixed(9365.0/65536.0,1,-nbitq), 
to_sfixed(11026.0/65536.0,1,-nbitq), 
to_sfixed(1298.0/65536.0,1,-nbitq), 
to_sfixed(1778.0/65536.0,1,-nbitq), 
to_sfixed(-2798.0/65536.0,1,-nbitq), 
to_sfixed(-2.0/65536.0,1,-nbitq), 
to_sfixed(3594.0/65536.0,1,-nbitq), 
to_sfixed(-2335.0/65536.0,1,-nbitq), 
to_sfixed(6389.0/65536.0,1,-nbitq), 
to_sfixed(-1177.0/65536.0,1,-nbitq), 
to_sfixed(11518.0/65536.0,1,-nbitq), 
to_sfixed(1521.0/65536.0,1,-nbitq), 
to_sfixed(-1653.0/65536.0,1,-nbitq), 
to_sfixed(828.0/65536.0,1,-nbitq), 
to_sfixed(-3041.0/65536.0,1,-nbitq), 
to_sfixed(-3009.0/65536.0,1,-nbitq), 
to_sfixed(1096.0/65536.0,1,-nbitq), 
to_sfixed(-27.0/65536.0,1,-nbitq), 
to_sfixed(3035.0/65536.0,1,-nbitq), 
to_sfixed(5423.0/65536.0,1,-nbitq), 
to_sfixed(8023.0/65536.0,1,-nbitq), 
to_sfixed(4264.0/65536.0,1,-nbitq), 
to_sfixed(-1323.0/65536.0,1,-nbitq), 
to_sfixed(-898.0/65536.0,1,-nbitq), 
to_sfixed(-2061.0/65536.0,1,-nbitq), 
to_sfixed(3034.0/65536.0,1,-nbitq), 
to_sfixed(908.0/65536.0,1,-nbitq), 
to_sfixed(-2027.0/65536.0,1,-nbitq), 
to_sfixed(2364.0/65536.0,1,-nbitq), 
to_sfixed(-137.0/65536.0,1,-nbitq), 
to_sfixed(-589.0/65536.0,1,-nbitq), 
to_sfixed(-543.0/65536.0,1,-nbitq), 
to_sfixed(-2256.0/65536.0,1,-nbitq), 
to_sfixed(-3071.0/65536.0,1,-nbitq), 
to_sfixed(5212.0/65536.0,1,-nbitq), 
to_sfixed(5214.0/65536.0,1,-nbitq), 
to_sfixed(-2615.0/65536.0,1,-nbitq), 
to_sfixed(-4675.0/65536.0,1,-nbitq), 
to_sfixed(1851.0/65536.0,1,-nbitq), 
to_sfixed(-1575.0/65536.0,1,-nbitq), 
to_sfixed(2716.0/65536.0,1,-nbitq), 
to_sfixed(-350.0/65536.0,1,-nbitq), 
to_sfixed(-2040.0/65536.0,1,-nbitq), 
to_sfixed(3448.0/65536.0,1,-nbitq), 
to_sfixed(-5176.0/65536.0,1,-nbitq), 
to_sfixed(-3980.0/65536.0,1,-nbitq), 
to_sfixed(2228.0/65536.0,1,-nbitq), 
to_sfixed(-13010.0/65536.0,1,-nbitq)  ), 
( to_sfixed(8531.0/65536.0,1,-nbitq), 
to_sfixed(4772.0/65536.0,1,-nbitq), 
to_sfixed(-1507.0/65536.0,1,-nbitq), 
to_sfixed(-3242.0/65536.0,1,-nbitq), 
to_sfixed(-2599.0/65536.0,1,-nbitq), 
to_sfixed(5334.0/65536.0,1,-nbitq), 
to_sfixed(-3239.0/65536.0,1,-nbitq), 
to_sfixed(12013.0/65536.0,1,-nbitq), 
to_sfixed(-4942.0/65536.0,1,-nbitq), 
to_sfixed(-2237.0/65536.0,1,-nbitq), 
to_sfixed(5272.0/65536.0,1,-nbitq), 
to_sfixed(-12817.0/65536.0,1,-nbitq), 
to_sfixed(2732.0/65536.0,1,-nbitq), 
to_sfixed(9850.0/65536.0,1,-nbitq), 
to_sfixed(-1645.0/65536.0,1,-nbitq), 
to_sfixed(912.0/65536.0,1,-nbitq), 
to_sfixed(-1337.0/65536.0,1,-nbitq), 
to_sfixed(8191.0/65536.0,1,-nbitq), 
to_sfixed(4120.0/65536.0,1,-nbitq), 
to_sfixed(-2301.0/65536.0,1,-nbitq), 
to_sfixed(5396.0/65536.0,1,-nbitq), 
to_sfixed(-9996.0/65536.0,1,-nbitq), 
to_sfixed(-7952.0/65536.0,1,-nbitq), 
to_sfixed(1614.0/65536.0,1,-nbitq), 
to_sfixed(3174.0/65536.0,1,-nbitq), 
to_sfixed(5081.0/65536.0,1,-nbitq), 
to_sfixed(689.0/65536.0,1,-nbitq), 
to_sfixed(678.0/65536.0,1,-nbitq), 
to_sfixed(1017.0/65536.0,1,-nbitq), 
to_sfixed(-322.0/65536.0,1,-nbitq), 
to_sfixed(1937.0/65536.0,1,-nbitq), 
to_sfixed(-10657.0/65536.0,1,-nbitq), 
to_sfixed(5746.0/65536.0,1,-nbitq), 
to_sfixed(83.0/65536.0,1,-nbitq), 
to_sfixed(2242.0/65536.0,1,-nbitq), 
to_sfixed(494.0/65536.0,1,-nbitq), 
to_sfixed(-939.0/65536.0,1,-nbitq), 
to_sfixed(5370.0/65536.0,1,-nbitq), 
to_sfixed(-625.0/65536.0,1,-nbitq), 
to_sfixed(2889.0/65536.0,1,-nbitq), 
to_sfixed(1548.0/65536.0,1,-nbitq), 
to_sfixed(-665.0/65536.0,1,-nbitq), 
to_sfixed(14229.0/65536.0,1,-nbitq), 
to_sfixed(5342.0/65536.0,1,-nbitq), 
to_sfixed(-94.0/65536.0,1,-nbitq), 
to_sfixed(-5889.0/65536.0,1,-nbitq), 
to_sfixed(305.0/65536.0,1,-nbitq), 
to_sfixed(-5711.0/65536.0,1,-nbitq), 
to_sfixed(-2555.0/65536.0,1,-nbitq), 
to_sfixed(4048.0/65536.0,1,-nbitq), 
to_sfixed(-1453.0/65536.0,1,-nbitq), 
to_sfixed(6913.0/65536.0,1,-nbitq), 
to_sfixed(7298.0/65536.0,1,-nbitq), 
to_sfixed(1548.0/65536.0,1,-nbitq), 
to_sfixed(-3496.0/65536.0,1,-nbitq), 
to_sfixed(376.0/65536.0,1,-nbitq), 
to_sfixed(-686.0/65536.0,1,-nbitq), 
to_sfixed(-941.0/65536.0,1,-nbitq), 
to_sfixed(-311.0/65536.0,1,-nbitq), 
to_sfixed(660.0/65536.0,1,-nbitq), 
to_sfixed(-2892.0/65536.0,1,-nbitq), 
to_sfixed(2432.0/65536.0,1,-nbitq), 
to_sfixed(-1382.0/65536.0,1,-nbitq), 
to_sfixed(2795.0/65536.0,1,-nbitq), 
to_sfixed(-6943.0/65536.0,1,-nbitq), 
to_sfixed(5134.0/65536.0,1,-nbitq), 
to_sfixed(4548.0/65536.0,1,-nbitq), 
to_sfixed(2702.0/65536.0,1,-nbitq), 
to_sfixed(-5481.0/65536.0,1,-nbitq), 
to_sfixed(-2447.0/65536.0,1,-nbitq), 
to_sfixed(1887.0/65536.0,1,-nbitq), 
to_sfixed(-140.0/65536.0,1,-nbitq), 
to_sfixed(5766.0/65536.0,1,-nbitq), 
to_sfixed(345.0/65536.0,1,-nbitq), 
to_sfixed(688.0/65536.0,1,-nbitq), 
to_sfixed(4627.0/65536.0,1,-nbitq), 
to_sfixed(871.0/65536.0,1,-nbitq), 
to_sfixed(1699.0/65536.0,1,-nbitq), 
to_sfixed(-998.0/65536.0,1,-nbitq), 
to_sfixed(-9849.0/65536.0,1,-nbitq)  ), 
( to_sfixed(6430.0/65536.0,1,-nbitq), 
to_sfixed(-2888.0/65536.0,1,-nbitq), 
to_sfixed(-2164.0/65536.0,1,-nbitq), 
to_sfixed(403.0/65536.0,1,-nbitq), 
to_sfixed(-312.0/65536.0,1,-nbitq), 
to_sfixed(8687.0/65536.0,1,-nbitq), 
to_sfixed(981.0/65536.0,1,-nbitq), 
to_sfixed(8396.0/65536.0,1,-nbitq), 
to_sfixed(-4252.0/65536.0,1,-nbitq), 
to_sfixed(-672.0/65536.0,1,-nbitq), 
to_sfixed(2812.0/65536.0,1,-nbitq), 
to_sfixed(-5324.0/65536.0,1,-nbitq), 
to_sfixed(438.0/65536.0,1,-nbitq), 
to_sfixed(3151.0/65536.0,1,-nbitq), 
to_sfixed(2822.0/65536.0,1,-nbitq), 
to_sfixed(-1979.0/65536.0,1,-nbitq), 
to_sfixed(-2107.0/65536.0,1,-nbitq), 
to_sfixed(8946.0/65536.0,1,-nbitq), 
to_sfixed(1031.0/65536.0,1,-nbitq), 
to_sfixed(3014.0/65536.0,1,-nbitq), 
to_sfixed(4803.0/65536.0,1,-nbitq), 
to_sfixed(-3420.0/65536.0,1,-nbitq), 
to_sfixed(-6634.0/65536.0,1,-nbitq), 
to_sfixed(1139.0/65536.0,1,-nbitq), 
to_sfixed(2977.0/65536.0,1,-nbitq), 
to_sfixed(6439.0/65536.0,1,-nbitq), 
to_sfixed(-2561.0/65536.0,1,-nbitq), 
to_sfixed(1497.0/65536.0,1,-nbitq), 
to_sfixed(4769.0/65536.0,1,-nbitq), 
to_sfixed(-610.0/65536.0,1,-nbitq), 
to_sfixed(889.0/65536.0,1,-nbitq), 
to_sfixed(-7198.0/65536.0,1,-nbitq), 
to_sfixed(6399.0/65536.0,1,-nbitq), 
to_sfixed(-216.0/65536.0,1,-nbitq), 
to_sfixed(-1457.0/65536.0,1,-nbitq), 
to_sfixed(2367.0/65536.0,1,-nbitq), 
to_sfixed(-223.0/65536.0,1,-nbitq), 
to_sfixed(636.0/65536.0,1,-nbitq), 
to_sfixed(-1685.0/65536.0,1,-nbitq), 
to_sfixed(-435.0/65536.0,1,-nbitq), 
to_sfixed(6249.0/65536.0,1,-nbitq), 
to_sfixed(-2107.0/65536.0,1,-nbitq), 
to_sfixed(8809.0/65536.0,1,-nbitq), 
to_sfixed(4266.0/65536.0,1,-nbitq), 
to_sfixed(2994.0/65536.0,1,-nbitq), 
to_sfixed(-4256.0/65536.0,1,-nbitq), 
to_sfixed(976.0/65536.0,1,-nbitq), 
to_sfixed(-2297.0/65536.0,1,-nbitq), 
to_sfixed(-2813.0/65536.0,1,-nbitq), 
to_sfixed(4293.0/65536.0,1,-nbitq), 
to_sfixed(-1799.0/65536.0,1,-nbitq), 
to_sfixed(5522.0/65536.0,1,-nbitq), 
to_sfixed(9762.0/65536.0,1,-nbitq), 
to_sfixed(4654.0/65536.0,1,-nbitq), 
to_sfixed(-2191.0/65536.0,1,-nbitq), 
to_sfixed(2450.0/65536.0,1,-nbitq), 
to_sfixed(-2267.0/65536.0,1,-nbitq), 
to_sfixed(2418.0/65536.0,1,-nbitq), 
to_sfixed(706.0/65536.0,1,-nbitq), 
to_sfixed(1706.0/65536.0,1,-nbitq), 
to_sfixed(171.0/65536.0,1,-nbitq), 
to_sfixed(-2353.0/65536.0,1,-nbitq), 
to_sfixed(-2367.0/65536.0,1,-nbitq), 
to_sfixed(-23.0/65536.0,1,-nbitq), 
to_sfixed(1499.0/65536.0,1,-nbitq), 
to_sfixed(2336.0/65536.0,1,-nbitq), 
to_sfixed(5984.0/65536.0,1,-nbitq), 
to_sfixed(3579.0/65536.0,1,-nbitq), 
to_sfixed(-6827.0/65536.0,1,-nbitq), 
to_sfixed(-8073.0/65536.0,1,-nbitq), 
to_sfixed(5821.0/65536.0,1,-nbitq), 
to_sfixed(-3014.0/65536.0,1,-nbitq), 
to_sfixed(4878.0/65536.0,1,-nbitq), 
to_sfixed(1498.0/65536.0,1,-nbitq), 
to_sfixed(-1061.0/65536.0,1,-nbitq), 
to_sfixed(4659.0/65536.0,1,-nbitq), 
to_sfixed(1062.0/65536.0,1,-nbitq), 
to_sfixed(1118.0/65536.0,1,-nbitq), 
to_sfixed(-735.0/65536.0,1,-nbitq), 
to_sfixed(-10094.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3983.0/65536.0,1,-nbitq), 
to_sfixed(-4086.0/65536.0,1,-nbitq), 
to_sfixed(-1683.0/65536.0,1,-nbitq), 
to_sfixed(-407.0/65536.0,1,-nbitq), 
to_sfixed(380.0/65536.0,1,-nbitq), 
to_sfixed(6510.0/65536.0,1,-nbitq), 
to_sfixed(-1084.0/65536.0,1,-nbitq), 
to_sfixed(3665.0/65536.0,1,-nbitq), 
to_sfixed(1335.0/65536.0,1,-nbitq), 
to_sfixed(-2529.0/65536.0,1,-nbitq), 
to_sfixed(618.0/65536.0,1,-nbitq), 
to_sfixed(-4966.0/65536.0,1,-nbitq), 
to_sfixed(2084.0/65536.0,1,-nbitq), 
to_sfixed(-1333.0/65536.0,1,-nbitq), 
to_sfixed(814.0/65536.0,1,-nbitq), 
to_sfixed(1406.0/65536.0,1,-nbitq), 
to_sfixed(1401.0/65536.0,1,-nbitq), 
to_sfixed(3584.0/65536.0,1,-nbitq), 
to_sfixed(-1973.0/65536.0,1,-nbitq), 
to_sfixed(450.0/65536.0,1,-nbitq), 
to_sfixed(109.0/65536.0,1,-nbitq), 
to_sfixed(-3577.0/65536.0,1,-nbitq), 
to_sfixed(-4848.0/65536.0,1,-nbitq), 
to_sfixed(-2926.0/65536.0,1,-nbitq), 
to_sfixed(2179.0/65536.0,1,-nbitq), 
to_sfixed(7316.0/65536.0,1,-nbitq), 
to_sfixed(-3328.0/65536.0,1,-nbitq), 
to_sfixed(-3064.0/65536.0,1,-nbitq), 
to_sfixed(2505.0/65536.0,1,-nbitq), 
to_sfixed(-2617.0/65536.0,1,-nbitq), 
to_sfixed(-956.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(7736.0/65536.0,1,-nbitq), 
to_sfixed(3.0/65536.0,1,-nbitq), 
to_sfixed(-897.0/65536.0,1,-nbitq), 
to_sfixed(-331.0/65536.0,1,-nbitq), 
to_sfixed(-3212.0/65536.0,1,-nbitq), 
to_sfixed(238.0/65536.0,1,-nbitq), 
to_sfixed(-3341.0/65536.0,1,-nbitq), 
to_sfixed(-270.0/65536.0,1,-nbitq), 
to_sfixed(2533.0/65536.0,1,-nbitq), 
to_sfixed(-1239.0/65536.0,1,-nbitq), 
to_sfixed(4081.0/65536.0,1,-nbitq), 
to_sfixed(1436.0/65536.0,1,-nbitq), 
to_sfixed(-1869.0/65536.0,1,-nbitq), 
to_sfixed(-5322.0/65536.0,1,-nbitq), 
to_sfixed(-2865.0/65536.0,1,-nbitq), 
to_sfixed(-3191.0/65536.0,1,-nbitq), 
to_sfixed(2076.0/65536.0,1,-nbitq), 
to_sfixed(3523.0/65536.0,1,-nbitq), 
to_sfixed(3232.0/65536.0,1,-nbitq), 
to_sfixed(8208.0/65536.0,1,-nbitq), 
to_sfixed(3354.0/65536.0,1,-nbitq), 
to_sfixed(4493.0/65536.0,1,-nbitq), 
to_sfixed(-1073.0/65536.0,1,-nbitq), 
to_sfixed(-823.0/65536.0,1,-nbitq), 
to_sfixed(1578.0/65536.0,1,-nbitq), 
to_sfixed(3313.0/65536.0,1,-nbitq), 
to_sfixed(-1073.0/65536.0,1,-nbitq), 
to_sfixed(-3281.0/65536.0,1,-nbitq), 
to_sfixed(-6117.0/65536.0,1,-nbitq), 
to_sfixed(1830.0/65536.0,1,-nbitq), 
to_sfixed(-1033.0/65536.0,1,-nbitq), 
to_sfixed(2130.0/65536.0,1,-nbitq), 
to_sfixed(-1985.0/65536.0,1,-nbitq), 
to_sfixed(3042.0/65536.0,1,-nbitq), 
to_sfixed(7441.0/65536.0,1,-nbitq), 
to_sfixed(5762.0/65536.0,1,-nbitq), 
to_sfixed(-3041.0/65536.0,1,-nbitq), 
to_sfixed(-4555.0/65536.0,1,-nbitq), 
to_sfixed(2017.0/65536.0,1,-nbitq), 
to_sfixed(429.0/65536.0,1,-nbitq), 
to_sfixed(7505.0/65536.0,1,-nbitq), 
to_sfixed(1175.0/65536.0,1,-nbitq), 
to_sfixed(2419.0/65536.0,1,-nbitq), 
to_sfixed(2462.0/65536.0,1,-nbitq), 
to_sfixed(-2450.0/65536.0,1,-nbitq), 
to_sfixed(4074.0/65536.0,1,-nbitq), 
to_sfixed(1661.0/65536.0,1,-nbitq), 
to_sfixed(-6472.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5035.0/65536.0,1,-nbitq), 
to_sfixed(3073.0/65536.0,1,-nbitq), 
to_sfixed(-4861.0/65536.0,1,-nbitq), 
to_sfixed(2626.0/65536.0,1,-nbitq), 
to_sfixed(914.0/65536.0,1,-nbitq), 
to_sfixed(1799.0/65536.0,1,-nbitq), 
to_sfixed(839.0/65536.0,1,-nbitq), 
to_sfixed(4268.0/65536.0,1,-nbitq), 
to_sfixed(-328.0/65536.0,1,-nbitq), 
to_sfixed(1582.0/65536.0,1,-nbitq), 
to_sfixed(-2100.0/65536.0,1,-nbitq), 
to_sfixed(2561.0/65536.0,1,-nbitq), 
to_sfixed(-3072.0/65536.0,1,-nbitq), 
to_sfixed(-880.0/65536.0,1,-nbitq), 
to_sfixed(2212.0/65536.0,1,-nbitq), 
to_sfixed(1842.0/65536.0,1,-nbitq), 
to_sfixed(-136.0/65536.0,1,-nbitq), 
to_sfixed(5493.0/65536.0,1,-nbitq), 
to_sfixed(779.0/65536.0,1,-nbitq), 
to_sfixed(-1964.0/65536.0,1,-nbitq), 
to_sfixed(1971.0/65536.0,1,-nbitq), 
to_sfixed(985.0/65536.0,1,-nbitq), 
to_sfixed(-3941.0/65536.0,1,-nbitq), 
to_sfixed(-3065.0/65536.0,1,-nbitq), 
to_sfixed(3727.0/65536.0,1,-nbitq), 
to_sfixed(-942.0/65536.0,1,-nbitq), 
to_sfixed(-4890.0/65536.0,1,-nbitq), 
to_sfixed(-439.0/65536.0,1,-nbitq), 
to_sfixed(1622.0/65536.0,1,-nbitq), 
to_sfixed(-323.0/65536.0,1,-nbitq), 
to_sfixed(2775.0/65536.0,1,-nbitq), 
to_sfixed(-3654.0/65536.0,1,-nbitq), 
to_sfixed(511.0/65536.0,1,-nbitq), 
to_sfixed(-921.0/65536.0,1,-nbitq), 
to_sfixed(558.0/65536.0,1,-nbitq), 
to_sfixed(-822.0/65536.0,1,-nbitq), 
to_sfixed(-2144.0/65536.0,1,-nbitq), 
to_sfixed(1431.0/65536.0,1,-nbitq), 
to_sfixed(-2938.0/65536.0,1,-nbitq), 
to_sfixed(1562.0/65536.0,1,-nbitq), 
to_sfixed(1232.0/65536.0,1,-nbitq), 
to_sfixed(2464.0/65536.0,1,-nbitq), 
to_sfixed(2474.0/65536.0,1,-nbitq), 
to_sfixed(1685.0/65536.0,1,-nbitq), 
to_sfixed(-58.0/65536.0,1,-nbitq), 
to_sfixed(-2708.0/65536.0,1,-nbitq), 
to_sfixed(819.0/65536.0,1,-nbitq), 
to_sfixed(-4086.0/65536.0,1,-nbitq), 
to_sfixed(-2403.0/65536.0,1,-nbitq), 
to_sfixed(-64.0/65536.0,1,-nbitq), 
to_sfixed(-1321.0/65536.0,1,-nbitq), 
to_sfixed(850.0/65536.0,1,-nbitq), 
to_sfixed(146.0/65536.0,1,-nbitq), 
to_sfixed(5582.0/65536.0,1,-nbitq), 
to_sfixed(54.0/65536.0,1,-nbitq), 
to_sfixed(3097.0/65536.0,1,-nbitq), 
to_sfixed(29.0/65536.0,1,-nbitq), 
to_sfixed(-388.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(1553.0/65536.0,1,-nbitq), 
to_sfixed(-1571.0/65536.0,1,-nbitq), 
to_sfixed(-683.0/65536.0,1,-nbitq), 
to_sfixed(-1472.0/65536.0,1,-nbitq), 
to_sfixed(-996.0/65536.0,1,-nbitq), 
to_sfixed(-2529.0/65536.0,1,-nbitq), 
to_sfixed(-1950.0/65536.0,1,-nbitq), 
to_sfixed(5679.0/65536.0,1,-nbitq), 
to_sfixed(-466.0/65536.0,1,-nbitq), 
to_sfixed(1325.0/65536.0,1,-nbitq), 
to_sfixed(1532.0/65536.0,1,-nbitq), 
to_sfixed(-205.0/65536.0,1,-nbitq), 
to_sfixed(-2119.0/65536.0,1,-nbitq), 
to_sfixed(2442.0/65536.0,1,-nbitq), 
to_sfixed(2002.0/65536.0,1,-nbitq), 
to_sfixed(294.0/65536.0,1,-nbitq), 
to_sfixed(2222.0/65536.0,1,-nbitq), 
to_sfixed(-1555.0/65536.0,1,-nbitq), 
to_sfixed(1530.0/65536.0,1,-nbitq), 
to_sfixed(2115.0/65536.0,1,-nbitq), 
to_sfixed(-2063.0/65536.0,1,-nbitq)  ), 
( to_sfixed(372.0/65536.0,1,-nbitq), 
to_sfixed(-1859.0/65536.0,1,-nbitq), 
to_sfixed(-3812.0/65536.0,1,-nbitq), 
to_sfixed(-1826.0/65536.0,1,-nbitq), 
to_sfixed(-1369.0/65536.0,1,-nbitq), 
to_sfixed(-72.0/65536.0,1,-nbitq), 
to_sfixed(-958.0/65536.0,1,-nbitq), 
to_sfixed(2316.0/65536.0,1,-nbitq), 
to_sfixed(-2452.0/65536.0,1,-nbitq), 
to_sfixed(-2382.0/65536.0,1,-nbitq), 
to_sfixed(-2485.0/65536.0,1,-nbitq), 
to_sfixed(-2439.0/65536.0,1,-nbitq), 
to_sfixed(1588.0/65536.0,1,-nbitq), 
to_sfixed(1904.0/65536.0,1,-nbitq), 
to_sfixed(-50.0/65536.0,1,-nbitq), 
to_sfixed(-3041.0/65536.0,1,-nbitq), 
to_sfixed(648.0/65536.0,1,-nbitq), 
to_sfixed(417.0/65536.0,1,-nbitq), 
to_sfixed(553.0/65536.0,1,-nbitq), 
to_sfixed(664.0/65536.0,1,-nbitq), 
to_sfixed(-1780.0/65536.0,1,-nbitq), 
to_sfixed(2114.0/65536.0,1,-nbitq), 
to_sfixed(-1369.0/65536.0,1,-nbitq), 
to_sfixed(1819.0/65536.0,1,-nbitq), 
to_sfixed(851.0/65536.0,1,-nbitq), 
to_sfixed(-1430.0/65536.0,1,-nbitq), 
to_sfixed(-2832.0/65536.0,1,-nbitq), 
to_sfixed(1608.0/65536.0,1,-nbitq), 
to_sfixed(-483.0/65536.0,1,-nbitq), 
to_sfixed(-2491.0/65536.0,1,-nbitq), 
to_sfixed(-2667.0/65536.0,1,-nbitq), 
to_sfixed(-686.0/65536.0,1,-nbitq), 
to_sfixed(-355.0/65536.0,1,-nbitq), 
to_sfixed(-1011.0/65536.0,1,-nbitq), 
to_sfixed(-2842.0/65536.0,1,-nbitq), 
to_sfixed(-2407.0/65536.0,1,-nbitq), 
to_sfixed(390.0/65536.0,1,-nbitq), 
to_sfixed(1041.0/65536.0,1,-nbitq), 
to_sfixed(-2656.0/65536.0,1,-nbitq), 
to_sfixed(3032.0/65536.0,1,-nbitq), 
to_sfixed(32.0/65536.0,1,-nbitq), 
to_sfixed(-1130.0/65536.0,1,-nbitq), 
to_sfixed(477.0/65536.0,1,-nbitq), 
to_sfixed(2771.0/65536.0,1,-nbitq), 
to_sfixed(474.0/65536.0,1,-nbitq), 
to_sfixed(238.0/65536.0,1,-nbitq), 
to_sfixed(-2742.0/65536.0,1,-nbitq), 
to_sfixed(-2440.0/65536.0,1,-nbitq), 
to_sfixed(1559.0/65536.0,1,-nbitq), 
to_sfixed(2779.0/65536.0,1,-nbitq), 
to_sfixed(2439.0/65536.0,1,-nbitq), 
to_sfixed(1021.0/65536.0,1,-nbitq), 
to_sfixed(2737.0/65536.0,1,-nbitq), 
to_sfixed(1911.0/65536.0,1,-nbitq), 
to_sfixed(-1231.0/65536.0,1,-nbitq), 
to_sfixed(-949.0/65536.0,1,-nbitq), 
to_sfixed(-1117.0/65536.0,1,-nbitq), 
to_sfixed(-1120.0/65536.0,1,-nbitq), 
to_sfixed(2397.0/65536.0,1,-nbitq), 
to_sfixed(-1113.0/65536.0,1,-nbitq), 
to_sfixed(-888.0/65536.0,1,-nbitq), 
to_sfixed(-180.0/65536.0,1,-nbitq), 
to_sfixed(266.0/65536.0,1,-nbitq), 
to_sfixed(-692.0/65536.0,1,-nbitq), 
to_sfixed(1878.0/65536.0,1,-nbitq), 
to_sfixed(967.0/65536.0,1,-nbitq), 
to_sfixed(2607.0/65536.0,1,-nbitq), 
to_sfixed(-814.0/65536.0,1,-nbitq), 
to_sfixed(-2475.0/65536.0,1,-nbitq), 
to_sfixed(490.0/65536.0,1,-nbitq), 
to_sfixed(311.0/65536.0,1,-nbitq), 
to_sfixed(635.0/65536.0,1,-nbitq), 
to_sfixed(-1404.0/65536.0,1,-nbitq), 
to_sfixed(-1925.0/65536.0,1,-nbitq), 
to_sfixed(1794.0/65536.0,1,-nbitq), 
to_sfixed(-282.0/65536.0,1,-nbitq), 
to_sfixed(-2386.0/65536.0,1,-nbitq), 
to_sfixed(1839.0/65536.0,1,-nbitq), 
to_sfixed(350.0/65536.0,1,-nbitq), 
to_sfixed(664.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2570.0/65536.0,1,-nbitq), 
to_sfixed(1880.0/65536.0,1,-nbitq), 
to_sfixed(1180.0/65536.0,1,-nbitq), 
to_sfixed(-397.0/65536.0,1,-nbitq), 
to_sfixed(-3538.0/65536.0,1,-nbitq), 
to_sfixed(-2050.0/65536.0,1,-nbitq), 
to_sfixed(-2985.0/65536.0,1,-nbitq), 
to_sfixed(-1464.0/65536.0,1,-nbitq), 
to_sfixed(2133.0/65536.0,1,-nbitq), 
to_sfixed(1930.0/65536.0,1,-nbitq), 
to_sfixed(-3105.0/65536.0,1,-nbitq), 
to_sfixed(2942.0/65536.0,1,-nbitq), 
to_sfixed(1120.0/65536.0,1,-nbitq), 
to_sfixed(-170.0/65536.0,1,-nbitq), 
to_sfixed(-938.0/65536.0,1,-nbitq), 
to_sfixed(2614.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(-1272.0/65536.0,1,-nbitq), 
to_sfixed(3193.0/65536.0,1,-nbitq), 
to_sfixed(2777.0/65536.0,1,-nbitq), 
to_sfixed(-308.0/65536.0,1,-nbitq), 
to_sfixed(-1978.0/65536.0,1,-nbitq), 
to_sfixed(720.0/65536.0,1,-nbitq), 
to_sfixed(-1017.0/65536.0,1,-nbitq), 
to_sfixed(-650.0/65536.0,1,-nbitq), 
to_sfixed(2011.0/65536.0,1,-nbitq), 
to_sfixed(-3180.0/65536.0,1,-nbitq), 
to_sfixed(-1406.0/65536.0,1,-nbitq), 
to_sfixed(888.0/65536.0,1,-nbitq), 
to_sfixed(-732.0/65536.0,1,-nbitq), 
to_sfixed(-2000.0/65536.0,1,-nbitq), 
to_sfixed(2628.0/65536.0,1,-nbitq), 
to_sfixed(-2555.0/65536.0,1,-nbitq), 
to_sfixed(-3207.0/65536.0,1,-nbitq), 
to_sfixed(-2277.0/65536.0,1,-nbitq), 
to_sfixed(-923.0/65536.0,1,-nbitq), 
to_sfixed(528.0/65536.0,1,-nbitq), 
to_sfixed(-3897.0/65536.0,1,-nbitq), 
to_sfixed(-1205.0/65536.0,1,-nbitq), 
to_sfixed(-1727.0/65536.0,1,-nbitq), 
to_sfixed(1605.0/65536.0,1,-nbitq), 
to_sfixed(-178.0/65536.0,1,-nbitq), 
to_sfixed(-3808.0/65536.0,1,-nbitq), 
to_sfixed(2768.0/65536.0,1,-nbitq), 
to_sfixed(1867.0/65536.0,1,-nbitq), 
to_sfixed(2180.0/65536.0,1,-nbitq), 
to_sfixed(387.0/65536.0,1,-nbitq), 
to_sfixed(1089.0/65536.0,1,-nbitq), 
to_sfixed(1227.0/65536.0,1,-nbitq), 
to_sfixed(2296.0/65536.0,1,-nbitq), 
to_sfixed(-2404.0/65536.0,1,-nbitq), 
to_sfixed(-1031.0/65536.0,1,-nbitq), 
to_sfixed(2891.0/65536.0,1,-nbitq), 
to_sfixed(508.0/65536.0,1,-nbitq), 
to_sfixed(3700.0/65536.0,1,-nbitq), 
to_sfixed(2536.0/65536.0,1,-nbitq), 
to_sfixed(1336.0/65536.0,1,-nbitq), 
to_sfixed(-315.0/65536.0,1,-nbitq), 
to_sfixed(1804.0/65536.0,1,-nbitq), 
to_sfixed(5038.0/65536.0,1,-nbitq), 
to_sfixed(-3232.0/65536.0,1,-nbitq), 
to_sfixed(-1060.0/65536.0,1,-nbitq), 
to_sfixed(568.0/65536.0,1,-nbitq), 
to_sfixed(-2319.0/65536.0,1,-nbitq), 
to_sfixed(-63.0/65536.0,1,-nbitq), 
to_sfixed(-806.0/65536.0,1,-nbitq), 
to_sfixed(736.0/65536.0,1,-nbitq), 
to_sfixed(909.0/65536.0,1,-nbitq), 
to_sfixed(890.0/65536.0,1,-nbitq), 
to_sfixed(-1801.0/65536.0,1,-nbitq), 
to_sfixed(1325.0/65536.0,1,-nbitq), 
to_sfixed(273.0/65536.0,1,-nbitq), 
to_sfixed(-1587.0/65536.0,1,-nbitq), 
to_sfixed(1262.0/65536.0,1,-nbitq), 
to_sfixed(-2963.0/65536.0,1,-nbitq), 
to_sfixed(3720.0/65536.0,1,-nbitq), 
to_sfixed(523.0/65536.0,1,-nbitq), 
to_sfixed(-172.0/65536.0,1,-nbitq), 
to_sfixed(-1118.0/65536.0,1,-nbitq), 
to_sfixed(-460.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2003.0/65536.0,1,-nbitq), 
to_sfixed(3141.0/65536.0,1,-nbitq), 
to_sfixed(4353.0/65536.0,1,-nbitq), 
to_sfixed(770.0/65536.0,1,-nbitq), 
to_sfixed(1643.0/65536.0,1,-nbitq), 
to_sfixed(-496.0/65536.0,1,-nbitq), 
to_sfixed(1031.0/65536.0,1,-nbitq), 
to_sfixed(213.0/65536.0,1,-nbitq), 
to_sfixed(2059.0/65536.0,1,-nbitq), 
to_sfixed(1419.0/65536.0,1,-nbitq), 
to_sfixed(-1725.0/65536.0,1,-nbitq), 
to_sfixed(-1429.0/65536.0,1,-nbitq), 
to_sfixed(1150.0/65536.0,1,-nbitq), 
to_sfixed(-2068.0/65536.0,1,-nbitq), 
to_sfixed(308.0/65536.0,1,-nbitq), 
to_sfixed(2109.0/65536.0,1,-nbitq), 
to_sfixed(1923.0/65536.0,1,-nbitq), 
to_sfixed(3645.0/65536.0,1,-nbitq), 
to_sfixed(1432.0/65536.0,1,-nbitq), 
to_sfixed(-1458.0/65536.0,1,-nbitq), 
to_sfixed(-2858.0/65536.0,1,-nbitq), 
to_sfixed(804.0/65536.0,1,-nbitq), 
to_sfixed(4016.0/65536.0,1,-nbitq), 
to_sfixed(2735.0/65536.0,1,-nbitq), 
to_sfixed(1015.0/65536.0,1,-nbitq), 
to_sfixed(-590.0/65536.0,1,-nbitq), 
to_sfixed(-4709.0/65536.0,1,-nbitq), 
to_sfixed(1529.0/65536.0,1,-nbitq), 
to_sfixed(-1264.0/65536.0,1,-nbitq), 
to_sfixed(-1603.0/65536.0,1,-nbitq), 
to_sfixed(-1151.0/65536.0,1,-nbitq), 
to_sfixed(-1944.0/65536.0,1,-nbitq), 
to_sfixed(-1008.0/65536.0,1,-nbitq), 
to_sfixed(-5002.0/65536.0,1,-nbitq), 
to_sfixed(-1664.0/65536.0,1,-nbitq), 
to_sfixed(2135.0/65536.0,1,-nbitq), 
to_sfixed(2839.0/65536.0,1,-nbitq), 
to_sfixed(441.0/65536.0,1,-nbitq), 
to_sfixed(-1558.0/65536.0,1,-nbitq), 
to_sfixed(-1042.0/65536.0,1,-nbitq), 
to_sfixed(316.0/65536.0,1,-nbitq), 
to_sfixed(334.0/65536.0,1,-nbitq), 
to_sfixed(-1584.0/65536.0,1,-nbitq), 
to_sfixed(1783.0/65536.0,1,-nbitq), 
to_sfixed(380.0/65536.0,1,-nbitq), 
to_sfixed(5408.0/65536.0,1,-nbitq), 
to_sfixed(1951.0/65536.0,1,-nbitq), 
to_sfixed(787.0/65536.0,1,-nbitq), 
to_sfixed(1175.0/65536.0,1,-nbitq), 
to_sfixed(477.0/65536.0,1,-nbitq), 
to_sfixed(3157.0/65536.0,1,-nbitq), 
to_sfixed(2169.0/65536.0,1,-nbitq), 
to_sfixed(1253.0/65536.0,1,-nbitq), 
to_sfixed(-1903.0/65536.0,1,-nbitq), 
to_sfixed(-802.0/65536.0,1,-nbitq), 
to_sfixed(-853.0/65536.0,1,-nbitq), 
to_sfixed(954.0/65536.0,1,-nbitq), 
to_sfixed(-422.0/65536.0,1,-nbitq), 
to_sfixed(-957.0/65536.0,1,-nbitq), 
to_sfixed(4029.0/65536.0,1,-nbitq), 
to_sfixed(1796.0/65536.0,1,-nbitq), 
to_sfixed(1860.0/65536.0,1,-nbitq), 
to_sfixed(144.0/65536.0,1,-nbitq), 
to_sfixed(1884.0/65536.0,1,-nbitq), 
to_sfixed(2678.0/65536.0,1,-nbitq), 
to_sfixed(4134.0/65536.0,1,-nbitq), 
to_sfixed(-900.0/65536.0,1,-nbitq), 
to_sfixed(-1507.0/65536.0,1,-nbitq), 
to_sfixed(1831.0/65536.0,1,-nbitq), 
to_sfixed(1472.0/65536.0,1,-nbitq), 
to_sfixed(-1454.0/65536.0,1,-nbitq), 
to_sfixed(1689.0/65536.0,1,-nbitq), 
to_sfixed(897.0/65536.0,1,-nbitq), 
to_sfixed(-960.0/65536.0,1,-nbitq), 
to_sfixed(-316.0/65536.0,1,-nbitq), 
to_sfixed(-2007.0/65536.0,1,-nbitq), 
to_sfixed(191.0/65536.0,1,-nbitq), 
to_sfixed(4963.0/65536.0,1,-nbitq), 
to_sfixed(2110.0/65536.0,1,-nbitq), 
to_sfixed(5143.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-271.0/65536.0,1,-nbitq), 
to_sfixed(500.0/65536.0,1,-nbitq), 
to_sfixed(1738.0/65536.0,1,-nbitq), 
to_sfixed(1791.0/65536.0,1,-nbitq), 
to_sfixed(1953.0/65536.0,1,-nbitq), 
to_sfixed(-4042.0/65536.0,1,-nbitq), 
to_sfixed(-1249.0/65536.0,1,-nbitq), 
to_sfixed(-880.0/65536.0,1,-nbitq), 
to_sfixed(-218.0/65536.0,1,-nbitq), 
to_sfixed(1266.0/65536.0,1,-nbitq), 
to_sfixed(-1471.0/65536.0,1,-nbitq), 
to_sfixed(1682.0/65536.0,1,-nbitq), 
to_sfixed(-1147.0/65536.0,1,-nbitq), 
to_sfixed(-1373.0/65536.0,1,-nbitq), 
to_sfixed(2472.0/65536.0,1,-nbitq), 
to_sfixed(2955.0/65536.0,1,-nbitq), 
to_sfixed(245.0/65536.0,1,-nbitq), 
to_sfixed(3024.0/65536.0,1,-nbitq), 
to_sfixed(3089.0/65536.0,1,-nbitq), 
to_sfixed(-953.0/65536.0,1,-nbitq), 
to_sfixed(-1732.0/65536.0,1,-nbitq), 
to_sfixed(-2416.0/65536.0,1,-nbitq), 
to_sfixed(3521.0/65536.0,1,-nbitq), 
to_sfixed(-169.0/65536.0,1,-nbitq), 
to_sfixed(2718.0/65536.0,1,-nbitq), 
to_sfixed(5174.0/65536.0,1,-nbitq), 
to_sfixed(-611.0/65536.0,1,-nbitq), 
to_sfixed(-901.0/65536.0,1,-nbitq), 
to_sfixed(-2136.0/65536.0,1,-nbitq), 
to_sfixed(828.0/65536.0,1,-nbitq), 
to_sfixed(226.0/65536.0,1,-nbitq), 
to_sfixed(-472.0/65536.0,1,-nbitq), 
to_sfixed(-889.0/65536.0,1,-nbitq), 
to_sfixed(-732.0/65536.0,1,-nbitq), 
to_sfixed(1435.0/65536.0,1,-nbitq), 
to_sfixed(1102.0/65536.0,1,-nbitq), 
to_sfixed(-702.0/65536.0,1,-nbitq), 
to_sfixed(-3747.0/65536.0,1,-nbitq), 
to_sfixed(-1316.0/65536.0,1,-nbitq), 
to_sfixed(2599.0/65536.0,1,-nbitq), 
to_sfixed(-1641.0/65536.0,1,-nbitq), 
to_sfixed(1282.0/65536.0,1,-nbitq), 
to_sfixed(-2695.0/65536.0,1,-nbitq), 
to_sfixed(-49.0/65536.0,1,-nbitq), 
to_sfixed(1354.0/65536.0,1,-nbitq), 
to_sfixed(6214.0/65536.0,1,-nbitq), 
to_sfixed(1537.0/65536.0,1,-nbitq), 
to_sfixed(-1050.0/65536.0,1,-nbitq), 
to_sfixed(2973.0/65536.0,1,-nbitq), 
to_sfixed(437.0/65536.0,1,-nbitq), 
to_sfixed(2874.0/65536.0,1,-nbitq), 
to_sfixed(2539.0/65536.0,1,-nbitq), 
to_sfixed(214.0/65536.0,1,-nbitq), 
to_sfixed(2242.0/65536.0,1,-nbitq), 
to_sfixed(-37.0/65536.0,1,-nbitq), 
to_sfixed(-2115.0/65536.0,1,-nbitq), 
to_sfixed(3115.0/65536.0,1,-nbitq), 
to_sfixed(-677.0/65536.0,1,-nbitq), 
to_sfixed(1001.0/65536.0,1,-nbitq), 
to_sfixed(4728.0/65536.0,1,-nbitq), 
to_sfixed(-2289.0/65536.0,1,-nbitq), 
to_sfixed(-1074.0/65536.0,1,-nbitq), 
to_sfixed(1793.0/65536.0,1,-nbitq), 
to_sfixed(-272.0/65536.0,1,-nbitq), 
to_sfixed(142.0/65536.0,1,-nbitq), 
to_sfixed(544.0/65536.0,1,-nbitq), 
to_sfixed(1249.0/65536.0,1,-nbitq), 
to_sfixed(-6771.0/65536.0,1,-nbitq), 
to_sfixed(-2538.0/65536.0,1,-nbitq), 
to_sfixed(3762.0/65536.0,1,-nbitq), 
to_sfixed(2700.0/65536.0,1,-nbitq), 
to_sfixed(-1756.0/65536.0,1,-nbitq), 
to_sfixed(-1155.0/65536.0,1,-nbitq), 
to_sfixed(-1095.0/65536.0,1,-nbitq), 
to_sfixed(964.0/65536.0,1,-nbitq), 
to_sfixed(2027.0/65536.0,1,-nbitq), 
to_sfixed(-463.0/65536.0,1,-nbitq), 
to_sfixed(1744.0/65536.0,1,-nbitq), 
to_sfixed(-1086.0/65536.0,1,-nbitq), 
to_sfixed(77.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3281.0/65536.0,1,-nbitq), 
to_sfixed(-269.0/65536.0,1,-nbitq), 
to_sfixed(4387.0/65536.0,1,-nbitq), 
to_sfixed(1038.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(-1951.0/65536.0,1,-nbitq), 
to_sfixed(-893.0/65536.0,1,-nbitq), 
to_sfixed(531.0/65536.0,1,-nbitq), 
to_sfixed(1025.0/65536.0,1,-nbitq), 
to_sfixed(-1427.0/65536.0,1,-nbitq), 
to_sfixed(2960.0/65536.0,1,-nbitq), 
to_sfixed(2838.0/65536.0,1,-nbitq), 
to_sfixed(1500.0/65536.0,1,-nbitq), 
to_sfixed(712.0/65536.0,1,-nbitq), 
to_sfixed(4844.0/65536.0,1,-nbitq), 
to_sfixed(-131.0/65536.0,1,-nbitq), 
to_sfixed(2235.0/65536.0,1,-nbitq), 
to_sfixed(-2203.0/65536.0,1,-nbitq), 
to_sfixed(2562.0/65536.0,1,-nbitq), 
to_sfixed(865.0/65536.0,1,-nbitq), 
to_sfixed(1465.0/65536.0,1,-nbitq), 
to_sfixed(-3819.0/65536.0,1,-nbitq), 
to_sfixed(-1726.0/65536.0,1,-nbitq), 
to_sfixed(3705.0/65536.0,1,-nbitq), 
to_sfixed(274.0/65536.0,1,-nbitq), 
to_sfixed(11920.0/65536.0,1,-nbitq), 
to_sfixed(1115.0/65536.0,1,-nbitq), 
to_sfixed(19.0/65536.0,1,-nbitq), 
to_sfixed(-416.0/65536.0,1,-nbitq), 
to_sfixed(413.0/65536.0,1,-nbitq), 
to_sfixed(1174.0/65536.0,1,-nbitq), 
to_sfixed(1931.0/65536.0,1,-nbitq), 
to_sfixed(-85.0/65536.0,1,-nbitq), 
to_sfixed(2071.0/65536.0,1,-nbitq), 
to_sfixed(1101.0/65536.0,1,-nbitq), 
to_sfixed(2489.0/65536.0,1,-nbitq), 
to_sfixed(-1282.0/65536.0,1,-nbitq), 
to_sfixed(-3721.0/65536.0,1,-nbitq), 
to_sfixed(435.0/65536.0,1,-nbitq), 
to_sfixed(-944.0/65536.0,1,-nbitq), 
to_sfixed(-140.0/65536.0,1,-nbitq), 
to_sfixed(2254.0/65536.0,1,-nbitq), 
to_sfixed(-1836.0/65536.0,1,-nbitq), 
to_sfixed(-3325.0/65536.0,1,-nbitq), 
to_sfixed(3029.0/65536.0,1,-nbitq), 
to_sfixed(7287.0/65536.0,1,-nbitq), 
to_sfixed(510.0/65536.0,1,-nbitq), 
to_sfixed(-1241.0/65536.0,1,-nbitq), 
to_sfixed(2490.0/65536.0,1,-nbitq), 
to_sfixed(2251.0/65536.0,1,-nbitq), 
to_sfixed(1896.0/65536.0,1,-nbitq), 
to_sfixed(-3370.0/65536.0,1,-nbitq), 
to_sfixed(111.0/65536.0,1,-nbitq), 
to_sfixed(3485.0/65536.0,1,-nbitq), 
to_sfixed(1850.0/65536.0,1,-nbitq), 
to_sfixed(5260.0/65536.0,1,-nbitq), 
to_sfixed(-1095.0/65536.0,1,-nbitq), 
to_sfixed(-2952.0/65536.0,1,-nbitq), 
to_sfixed(323.0/65536.0,1,-nbitq), 
to_sfixed(2414.0/65536.0,1,-nbitq), 
to_sfixed(1385.0/65536.0,1,-nbitq), 
to_sfixed(-2598.0/65536.0,1,-nbitq), 
to_sfixed(1008.0/65536.0,1,-nbitq), 
to_sfixed(-1414.0/65536.0,1,-nbitq), 
to_sfixed(-1700.0/65536.0,1,-nbitq), 
to_sfixed(3589.0/65536.0,1,-nbitq), 
to_sfixed(-1288.0/65536.0,1,-nbitq), 
to_sfixed(-5333.0/65536.0,1,-nbitq), 
to_sfixed(-306.0/65536.0,1,-nbitq), 
to_sfixed(-1833.0/65536.0,1,-nbitq), 
to_sfixed(-2435.0/65536.0,1,-nbitq), 
to_sfixed(-1322.0/65536.0,1,-nbitq), 
to_sfixed(1271.0/65536.0,1,-nbitq), 
to_sfixed(-2372.0/65536.0,1,-nbitq), 
to_sfixed(-2381.0/65536.0,1,-nbitq), 
to_sfixed(2367.0/65536.0,1,-nbitq), 
to_sfixed(-2112.0/65536.0,1,-nbitq), 
to_sfixed(-2259.0/65536.0,1,-nbitq), 
to_sfixed(-1565.0/65536.0,1,-nbitq), 
to_sfixed(860.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3154.0/65536.0,1,-nbitq), 
to_sfixed(-3044.0/65536.0,1,-nbitq), 
to_sfixed(-390.0/65536.0,1,-nbitq), 
to_sfixed(3629.0/65536.0,1,-nbitq), 
to_sfixed(4073.0/65536.0,1,-nbitq), 
to_sfixed(-1379.0/65536.0,1,-nbitq), 
to_sfixed(520.0/65536.0,1,-nbitq), 
to_sfixed(-1782.0/65536.0,1,-nbitq), 
to_sfixed(1815.0/65536.0,1,-nbitq), 
to_sfixed(-1425.0/65536.0,1,-nbitq), 
to_sfixed(-785.0/65536.0,1,-nbitq), 
to_sfixed(6744.0/65536.0,1,-nbitq), 
to_sfixed(-2940.0/65536.0,1,-nbitq), 
to_sfixed(209.0/65536.0,1,-nbitq), 
to_sfixed(5326.0/65536.0,1,-nbitq), 
to_sfixed(-2441.0/65536.0,1,-nbitq), 
to_sfixed(347.0/65536.0,1,-nbitq), 
to_sfixed(-4162.0/65536.0,1,-nbitq), 
to_sfixed(4345.0/65536.0,1,-nbitq), 
to_sfixed(1295.0/65536.0,1,-nbitq), 
to_sfixed(-761.0/65536.0,1,-nbitq), 
to_sfixed(-2410.0/65536.0,1,-nbitq), 
to_sfixed(-154.0/65536.0,1,-nbitq), 
to_sfixed(6832.0/65536.0,1,-nbitq), 
to_sfixed(-3002.0/65536.0,1,-nbitq), 
to_sfixed(15481.0/65536.0,1,-nbitq), 
to_sfixed(4605.0/65536.0,1,-nbitq), 
to_sfixed(869.0/65536.0,1,-nbitq), 
to_sfixed(1107.0/65536.0,1,-nbitq), 
to_sfixed(732.0/65536.0,1,-nbitq), 
to_sfixed(-2351.0/65536.0,1,-nbitq), 
to_sfixed(-48.0/65536.0,1,-nbitq), 
to_sfixed(77.0/65536.0,1,-nbitq), 
to_sfixed(4606.0/65536.0,1,-nbitq), 
to_sfixed(1695.0/65536.0,1,-nbitq), 
to_sfixed(-3506.0/65536.0,1,-nbitq), 
to_sfixed(-5131.0/65536.0,1,-nbitq), 
to_sfixed(-4532.0/65536.0,1,-nbitq), 
to_sfixed(-4284.0/65536.0,1,-nbitq), 
to_sfixed(-6090.0/65536.0,1,-nbitq), 
to_sfixed(-5122.0/65536.0,1,-nbitq), 
to_sfixed(-2065.0/65536.0,1,-nbitq), 
to_sfixed(-2510.0/65536.0,1,-nbitq), 
to_sfixed(-61.0/65536.0,1,-nbitq), 
to_sfixed(1974.0/65536.0,1,-nbitq), 
to_sfixed(2735.0/65536.0,1,-nbitq), 
to_sfixed(-3113.0/65536.0,1,-nbitq), 
to_sfixed(-893.0/65536.0,1,-nbitq), 
to_sfixed(148.0/65536.0,1,-nbitq), 
to_sfixed(2110.0/65536.0,1,-nbitq), 
to_sfixed(-795.0/65536.0,1,-nbitq), 
to_sfixed(-1191.0/65536.0,1,-nbitq), 
to_sfixed(219.0/65536.0,1,-nbitq), 
to_sfixed(5950.0/65536.0,1,-nbitq), 
to_sfixed(-3818.0/65536.0,1,-nbitq), 
to_sfixed(3470.0/65536.0,1,-nbitq), 
to_sfixed(1272.0/65536.0,1,-nbitq), 
to_sfixed(1540.0/65536.0,1,-nbitq), 
to_sfixed(994.0/65536.0,1,-nbitq), 
to_sfixed(1365.0/65536.0,1,-nbitq), 
to_sfixed(-3276.0/65536.0,1,-nbitq), 
to_sfixed(137.0/65536.0,1,-nbitq), 
to_sfixed(-2207.0/65536.0,1,-nbitq), 
to_sfixed(1517.0/65536.0,1,-nbitq), 
to_sfixed(-330.0/65536.0,1,-nbitq), 
to_sfixed(3465.0/65536.0,1,-nbitq), 
to_sfixed(-728.0/65536.0,1,-nbitq), 
to_sfixed(-6546.0/65536.0,1,-nbitq), 
to_sfixed(-3954.0/65536.0,1,-nbitq), 
to_sfixed(2240.0/65536.0,1,-nbitq), 
to_sfixed(-652.0/65536.0,1,-nbitq), 
to_sfixed(642.0/65536.0,1,-nbitq), 
to_sfixed(-2342.0/65536.0,1,-nbitq), 
to_sfixed(2371.0/65536.0,1,-nbitq), 
to_sfixed(-2156.0/65536.0,1,-nbitq), 
to_sfixed(-1040.0/65536.0,1,-nbitq), 
to_sfixed(-2722.0/65536.0,1,-nbitq), 
to_sfixed(-3663.0/65536.0,1,-nbitq), 
to_sfixed(-1072.0/65536.0,1,-nbitq), 
to_sfixed(-191.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-664.0/65536.0,1,-nbitq), 
to_sfixed(797.0/65536.0,1,-nbitq), 
to_sfixed(5358.0/65536.0,1,-nbitq), 
to_sfixed(7486.0/65536.0,1,-nbitq), 
to_sfixed(3463.0/65536.0,1,-nbitq), 
to_sfixed(902.0/65536.0,1,-nbitq), 
to_sfixed(-3383.0/65536.0,1,-nbitq), 
to_sfixed(-222.0/65536.0,1,-nbitq), 
to_sfixed(-281.0/65536.0,1,-nbitq), 
to_sfixed(1485.0/65536.0,1,-nbitq), 
to_sfixed(2893.0/65536.0,1,-nbitq), 
to_sfixed(12146.0/65536.0,1,-nbitq), 
to_sfixed(-2073.0/65536.0,1,-nbitq), 
to_sfixed(2488.0/65536.0,1,-nbitq), 
to_sfixed(1616.0/65536.0,1,-nbitq), 
to_sfixed(-674.0/65536.0,1,-nbitq), 
to_sfixed(2563.0/65536.0,1,-nbitq), 
to_sfixed(-5657.0/65536.0,1,-nbitq), 
to_sfixed(2159.0/65536.0,1,-nbitq), 
to_sfixed(1912.0/65536.0,1,-nbitq), 
to_sfixed(1281.0/65536.0,1,-nbitq), 
to_sfixed(-1268.0/65536.0,1,-nbitq), 
to_sfixed(6175.0/65536.0,1,-nbitq), 
to_sfixed(6338.0/65536.0,1,-nbitq), 
to_sfixed(-176.0/65536.0,1,-nbitq), 
to_sfixed(15304.0/65536.0,1,-nbitq), 
to_sfixed(3836.0/65536.0,1,-nbitq), 
to_sfixed(-2657.0/65536.0,1,-nbitq), 
to_sfixed(233.0/65536.0,1,-nbitq), 
to_sfixed(2913.0/65536.0,1,-nbitq), 
to_sfixed(-3110.0/65536.0,1,-nbitq), 
to_sfixed(-1167.0/65536.0,1,-nbitq), 
to_sfixed(6233.0/65536.0,1,-nbitq), 
to_sfixed(2489.0/65536.0,1,-nbitq), 
to_sfixed(-2456.0/65536.0,1,-nbitq), 
to_sfixed(-452.0/65536.0,1,-nbitq), 
to_sfixed(-1288.0/65536.0,1,-nbitq), 
to_sfixed(-744.0/65536.0,1,-nbitq), 
to_sfixed(-5699.0/65536.0,1,-nbitq), 
to_sfixed(-5565.0/65536.0,1,-nbitq), 
to_sfixed(-8309.0/65536.0,1,-nbitq), 
to_sfixed(-1016.0/65536.0,1,-nbitq), 
to_sfixed(3439.0/65536.0,1,-nbitq), 
to_sfixed(457.0/65536.0,1,-nbitq), 
to_sfixed(-1342.0/65536.0,1,-nbitq), 
to_sfixed(-2130.0/65536.0,1,-nbitq), 
to_sfixed(-1578.0/65536.0,1,-nbitq), 
to_sfixed(-2945.0/65536.0,1,-nbitq), 
to_sfixed(901.0/65536.0,1,-nbitq), 
to_sfixed(3876.0/65536.0,1,-nbitq), 
to_sfixed(-210.0/65536.0,1,-nbitq), 
to_sfixed(-3298.0/65536.0,1,-nbitq), 
to_sfixed(939.0/65536.0,1,-nbitq), 
to_sfixed(7514.0/65536.0,1,-nbitq), 
to_sfixed(-6600.0/65536.0,1,-nbitq), 
to_sfixed(6422.0/65536.0,1,-nbitq), 
to_sfixed(1630.0/65536.0,1,-nbitq), 
to_sfixed(-5633.0/65536.0,1,-nbitq), 
to_sfixed(1977.0/65536.0,1,-nbitq), 
to_sfixed(-500.0/65536.0,1,-nbitq), 
to_sfixed(-3884.0/65536.0,1,-nbitq), 
to_sfixed(-1222.0/65536.0,1,-nbitq), 
to_sfixed(910.0/65536.0,1,-nbitq), 
to_sfixed(-2702.0/65536.0,1,-nbitq), 
to_sfixed(-3687.0/65536.0,1,-nbitq), 
to_sfixed(3668.0/65536.0,1,-nbitq), 
to_sfixed(-5337.0/65536.0,1,-nbitq), 
to_sfixed(-11739.0/65536.0,1,-nbitq), 
to_sfixed(-2782.0/65536.0,1,-nbitq), 
to_sfixed(-4361.0/65536.0,1,-nbitq), 
to_sfixed(2304.0/65536.0,1,-nbitq), 
to_sfixed(-6864.0/65536.0,1,-nbitq), 
to_sfixed(-2635.0/65536.0,1,-nbitq), 
to_sfixed(-1943.0/65536.0,1,-nbitq), 
to_sfixed(-2929.0/65536.0,1,-nbitq), 
to_sfixed(-764.0/65536.0,1,-nbitq), 
to_sfixed(-163.0/65536.0,1,-nbitq), 
to_sfixed(-3042.0/65536.0,1,-nbitq), 
to_sfixed(2350.0/65536.0,1,-nbitq), 
to_sfixed(-1694.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-628.0/65536.0,1,-nbitq), 
to_sfixed(-2798.0/65536.0,1,-nbitq), 
to_sfixed(7949.0/65536.0,1,-nbitq), 
to_sfixed(11072.0/65536.0,1,-nbitq), 
to_sfixed(2639.0/65536.0,1,-nbitq), 
to_sfixed(8297.0/65536.0,1,-nbitq), 
to_sfixed(-186.0/65536.0,1,-nbitq), 
to_sfixed(4094.0/65536.0,1,-nbitq), 
to_sfixed(732.0/65536.0,1,-nbitq), 
to_sfixed(2898.0/65536.0,1,-nbitq), 
to_sfixed(120.0/65536.0,1,-nbitq), 
to_sfixed(17893.0/65536.0,1,-nbitq), 
to_sfixed(-2070.0/65536.0,1,-nbitq), 
to_sfixed(6035.0/65536.0,1,-nbitq), 
to_sfixed(-1594.0/65536.0,1,-nbitq), 
to_sfixed(646.0/65536.0,1,-nbitq), 
to_sfixed(-3115.0/65536.0,1,-nbitq), 
to_sfixed(2415.0/65536.0,1,-nbitq), 
to_sfixed(2154.0/65536.0,1,-nbitq), 
to_sfixed(-2510.0/65536.0,1,-nbitq), 
to_sfixed(3767.0/65536.0,1,-nbitq), 
to_sfixed(2658.0/65536.0,1,-nbitq), 
to_sfixed(656.0/65536.0,1,-nbitq), 
to_sfixed(-6480.0/65536.0,1,-nbitq), 
to_sfixed(3652.0/65536.0,1,-nbitq), 
to_sfixed(13796.0/65536.0,1,-nbitq), 
to_sfixed(6628.0/65536.0,1,-nbitq), 
to_sfixed(-3952.0/65536.0,1,-nbitq), 
to_sfixed(3953.0/65536.0,1,-nbitq), 
to_sfixed(4153.0/65536.0,1,-nbitq), 
to_sfixed(-2086.0/65536.0,1,-nbitq), 
to_sfixed(-2826.0/65536.0,1,-nbitq), 
to_sfixed(3473.0/65536.0,1,-nbitq), 
to_sfixed(-2863.0/65536.0,1,-nbitq), 
to_sfixed(-3867.0/65536.0,1,-nbitq), 
to_sfixed(-1434.0/65536.0,1,-nbitq), 
to_sfixed(-4579.0/65536.0,1,-nbitq), 
to_sfixed(2030.0/65536.0,1,-nbitq), 
to_sfixed(-3521.0/65536.0,1,-nbitq), 
to_sfixed(-6865.0/65536.0,1,-nbitq), 
to_sfixed(-9838.0/65536.0,1,-nbitq), 
to_sfixed(2481.0/65536.0,1,-nbitq), 
to_sfixed(231.0/65536.0,1,-nbitq), 
to_sfixed(-2560.0/65536.0,1,-nbitq), 
to_sfixed(1711.0/65536.0,1,-nbitq), 
to_sfixed(-899.0/65536.0,1,-nbitq), 
to_sfixed(-1698.0/65536.0,1,-nbitq), 
to_sfixed(-1931.0/65536.0,1,-nbitq), 
to_sfixed(-26.0/65536.0,1,-nbitq), 
to_sfixed(2478.0/65536.0,1,-nbitq), 
to_sfixed(157.0/65536.0,1,-nbitq), 
to_sfixed(728.0/65536.0,1,-nbitq), 
to_sfixed(-1653.0/65536.0,1,-nbitq), 
to_sfixed(9060.0/65536.0,1,-nbitq), 
to_sfixed(-3073.0/65536.0,1,-nbitq), 
to_sfixed(8534.0/65536.0,1,-nbitq), 
to_sfixed(1743.0/65536.0,1,-nbitq), 
to_sfixed(-3994.0/65536.0,1,-nbitq), 
to_sfixed(-1737.0/65536.0,1,-nbitq), 
to_sfixed(853.0/65536.0,1,-nbitq), 
to_sfixed(-3217.0/65536.0,1,-nbitq), 
to_sfixed(2560.0/65536.0,1,-nbitq), 
to_sfixed(2005.0/65536.0,1,-nbitq), 
to_sfixed(2020.0/65536.0,1,-nbitq), 
to_sfixed(-1858.0/65536.0,1,-nbitq), 
to_sfixed(9269.0/65536.0,1,-nbitq), 
to_sfixed(-2012.0/65536.0,1,-nbitq), 
to_sfixed(-6007.0/65536.0,1,-nbitq), 
to_sfixed(-7333.0/65536.0,1,-nbitq), 
to_sfixed(-10463.0/65536.0,1,-nbitq), 
to_sfixed(-2203.0/65536.0,1,-nbitq), 
to_sfixed(-4121.0/65536.0,1,-nbitq), 
to_sfixed(-2970.0/65536.0,1,-nbitq), 
to_sfixed(-2853.0/65536.0,1,-nbitq), 
to_sfixed(832.0/65536.0,1,-nbitq), 
to_sfixed(-2033.0/65536.0,1,-nbitq), 
to_sfixed(-2803.0/65536.0,1,-nbitq), 
to_sfixed(-2689.0/65536.0,1,-nbitq), 
to_sfixed(-2149.0/65536.0,1,-nbitq), 
to_sfixed(-4693.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5853.0/65536.0,1,-nbitq), 
to_sfixed(-552.0/65536.0,1,-nbitq), 
to_sfixed(7543.0/65536.0,1,-nbitq), 
to_sfixed(4713.0/65536.0,1,-nbitq), 
to_sfixed(454.0/65536.0,1,-nbitq), 
to_sfixed(3498.0/65536.0,1,-nbitq), 
to_sfixed(1486.0/65536.0,1,-nbitq), 
to_sfixed(2171.0/65536.0,1,-nbitq), 
to_sfixed(1060.0/65536.0,1,-nbitq), 
to_sfixed(-2540.0/65536.0,1,-nbitq), 
to_sfixed(-1282.0/65536.0,1,-nbitq), 
to_sfixed(21836.0/65536.0,1,-nbitq), 
to_sfixed(3006.0/65536.0,1,-nbitq), 
to_sfixed(8472.0/65536.0,1,-nbitq), 
to_sfixed(-8451.0/65536.0,1,-nbitq), 
to_sfixed(2119.0/65536.0,1,-nbitq), 
to_sfixed(-3220.0/65536.0,1,-nbitq), 
to_sfixed(6652.0/65536.0,1,-nbitq), 
to_sfixed(195.0/65536.0,1,-nbitq), 
to_sfixed(2609.0/65536.0,1,-nbitq), 
to_sfixed(4762.0/65536.0,1,-nbitq), 
to_sfixed(-793.0/65536.0,1,-nbitq), 
to_sfixed(504.0/65536.0,1,-nbitq), 
to_sfixed(-13713.0/65536.0,1,-nbitq), 
to_sfixed(1882.0/65536.0,1,-nbitq), 
to_sfixed(6356.0/65536.0,1,-nbitq), 
to_sfixed(5473.0/65536.0,1,-nbitq), 
to_sfixed(-3393.0/65536.0,1,-nbitq), 
to_sfixed(-3771.0/65536.0,1,-nbitq), 
to_sfixed(6701.0/65536.0,1,-nbitq), 
to_sfixed(441.0/65536.0,1,-nbitq), 
to_sfixed(1475.0/65536.0,1,-nbitq), 
to_sfixed(4154.0/65536.0,1,-nbitq), 
to_sfixed(-97.0/65536.0,1,-nbitq), 
to_sfixed(-607.0/65536.0,1,-nbitq), 
to_sfixed(2301.0/65536.0,1,-nbitq), 
to_sfixed(-1632.0/65536.0,1,-nbitq), 
to_sfixed(186.0/65536.0,1,-nbitq), 
to_sfixed(-9528.0/65536.0,1,-nbitq), 
to_sfixed(2300.0/65536.0,1,-nbitq), 
to_sfixed(-13570.0/65536.0,1,-nbitq), 
to_sfixed(-708.0/65536.0,1,-nbitq), 
to_sfixed(4565.0/65536.0,1,-nbitq), 
to_sfixed(2250.0/65536.0,1,-nbitq), 
to_sfixed(1913.0/65536.0,1,-nbitq), 
to_sfixed(-2735.0/65536.0,1,-nbitq), 
to_sfixed(-1271.0/65536.0,1,-nbitq), 
to_sfixed(5636.0/65536.0,1,-nbitq), 
to_sfixed(3189.0/65536.0,1,-nbitq), 
to_sfixed(-1647.0/65536.0,1,-nbitq), 
to_sfixed(898.0/65536.0,1,-nbitq), 
to_sfixed(8150.0/65536.0,1,-nbitq), 
to_sfixed(-1736.0/65536.0,1,-nbitq), 
to_sfixed(6785.0/65536.0,1,-nbitq), 
to_sfixed(-1566.0/65536.0,1,-nbitq), 
to_sfixed(7269.0/65536.0,1,-nbitq), 
to_sfixed(-257.0/65536.0,1,-nbitq), 
to_sfixed(711.0/65536.0,1,-nbitq), 
to_sfixed(1796.0/65536.0,1,-nbitq), 
to_sfixed(-1181.0/65536.0,1,-nbitq), 
to_sfixed(-3825.0/65536.0,1,-nbitq), 
to_sfixed(925.0/65536.0,1,-nbitq), 
to_sfixed(1372.0/65536.0,1,-nbitq), 
to_sfixed(-1112.0/65536.0,1,-nbitq), 
to_sfixed(-1786.0/65536.0,1,-nbitq), 
to_sfixed(5307.0/65536.0,1,-nbitq), 
to_sfixed(-2326.0/65536.0,1,-nbitq), 
to_sfixed(-6164.0/65536.0,1,-nbitq), 
to_sfixed(-2561.0/65536.0,1,-nbitq), 
to_sfixed(-5307.0/65536.0,1,-nbitq), 
to_sfixed(1981.0/65536.0,1,-nbitq), 
to_sfixed(-3986.0/65536.0,1,-nbitq), 
to_sfixed(1031.0/65536.0,1,-nbitq), 
to_sfixed(330.0/65536.0,1,-nbitq), 
to_sfixed(2822.0/65536.0,1,-nbitq), 
to_sfixed(-5069.0/65536.0,1,-nbitq), 
to_sfixed(1744.0/65536.0,1,-nbitq), 
to_sfixed(-6295.0/65536.0,1,-nbitq), 
to_sfixed(-2486.0/65536.0,1,-nbitq), 
to_sfixed(-4609.0/65536.0,1,-nbitq)  ), 
( to_sfixed(6782.0/65536.0,1,-nbitq), 
to_sfixed(-3221.0/65536.0,1,-nbitq), 
to_sfixed(7072.0/65536.0,1,-nbitq), 
to_sfixed(7355.0/65536.0,1,-nbitq), 
to_sfixed(-2920.0/65536.0,1,-nbitq), 
to_sfixed(-3471.0/65536.0,1,-nbitq), 
to_sfixed(3472.0/65536.0,1,-nbitq), 
to_sfixed(9805.0/65536.0,1,-nbitq), 
to_sfixed(-3343.0/65536.0,1,-nbitq), 
to_sfixed(-2076.0/65536.0,1,-nbitq), 
to_sfixed(-20.0/65536.0,1,-nbitq), 
to_sfixed(9042.0/65536.0,1,-nbitq), 
to_sfixed(2101.0/65536.0,1,-nbitq), 
to_sfixed(13726.0/65536.0,1,-nbitq), 
to_sfixed(-1997.0/65536.0,1,-nbitq), 
to_sfixed(-588.0/65536.0,1,-nbitq), 
to_sfixed(1451.0/65536.0,1,-nbitq), 
to_sfixed(4431.0/65536.0,1,-nbitq), 
to_sfixed(3320.0/65536.0,1,-nbitq), 
to_sfixed(2337.0/65536.0,1,-nbitq), 
to_sfixed(6344.0/65536.0,1,-nbitq), 
to_sfixed(-5702.0/65536.0,1,-nbitq), 
to_sfixed(-2251.0/65536.0,1,-nbitq), 
to_sfixed(-11637.0/65536.0,1,-nbitq), 
to_sfixed(585.0/65536.0,1,-nbitq), 
to_sfixed(4093.0/65536.0,1,-nbitq), 
to_sfixed(10290.0/65536.0,1,-nbitq), 
to_sfixed(-2656.0/65536.0,1,-nbitq), 
to_sfixed(-5612.0/65536.0,1,-nbitq), 
to_sfixed(3608.0/65536.0,1,-nbitq), 
to_sfixed(1914.0/65536.0,1,-nbitq), 
to_sfixed(4905.0/65536.0,1,-nbitq), 
to_sfixed(3553.0/65536.0,1,-nbitq), 
to_sfixed(5401.0/65536.0,1,-nbitq), 
to_sfixed(-1861.0/65536.0,1,-nbitq), 
to_sfixed(2757.0/65536.0,1,-nbitq), 
to_sfixed(5802.0/65536.0,1,-nbitq), 
to_sfixed(-5439.0/65536.0,1,-nbitq), 
to_sfixed(-5328.0/65536.0,1,-nbitq), 
to_sfixed(7470.0/65536.0,1,-nbitq), 
to_sfixed(-11701.0/65536.0,1,-nbitq), 
to_sfixed(293.0/65536.0,1,-nbitq), 
to_sfixed(6967.0/65536.0,1,-nbitq), 
to_sfixed(718.0/65536.0,1,-nbitq), 
to_sfixed(-160.0/65536.0,1,-nbitq), 
to_sfixed(-2513.0/65536.0,1,-nbitq), 
to_sfixed(-1651.0/65536.0,1,-nbitq), 
to_sfixed(5772.0/65536.0,1,-nbitq), 
to_sfixed(-509.0/65536.0,1,-nbitq), 
to_sfixed(-1882.0/65536.0,1,-nbitq), 
to_sfixed(-1668.0/65536.0,1,-nbitq), 
to_sfixed(11139.0/65536.0,1,-nbitq), 
to_sfixed(4775.0/65536.0,1,-nbitq), 
to_sfixed(11720.0/65536.0,1,-nbitq), 
to_sfixed(3439.0/65536.0,1,-nbitq), 
to_sfixed(8808.0/65536.0,1,-nbitq), 
to_sfixed(2212.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(2386.0/65536.0,1,-nbitq), 
to_sfixed(-2282.0/65536.0,1,-nbitq), 
to_sfixed(-1753.0/65536.0,1,-nbitq), 
to_sfixed(2870.0/65536.0,1,-nbitq), 
to_sfixed(-780.0/65536.0,1,-nbitq), 
to_sfixed(1636.0/65536.0,1,-nbitq), 
to_sfixed(-3204.0/65536.0,1,-nbitq), 
to_sfixed(3049.0/65536.0,1,-nbitq), 
to_sfixed(-2158.0/65536.0,1,-nbitq), 
to_sfixed(-9432.0/65536.0,1,-nbitq), 
to_sfixed(-7784.0/65536.0,1,-nbitq), 
to_sfixed(-7081.0/65536.0,1,-nbitq), 
to_sfixed(-1192.0/65536.0,1,-nbitq), 
to_sfixed(1897.0/65536.0,1,-nbitq), 
to_sfixed(-1246.0/65536.0,1,-nbitq), 
to_sfixed(-1855.0/65536.0,1,-nbitq), 
to_sfixed(813.0/65536.0,1,-nbitq), 
to_sfixed(-3948.0/65536.0,1,-nbitq), 
to_sfixed(6227.0/65536.0,1,-nbitq), 
to_sfixed(1269.0/65536.0,1,-nbitq), 
to_sfixed(2550.0/65536.0,1,-nbitq), 
to_sfixed(-761.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3627.0/65536.0,1,-nbitq), 
to_sfixed(-1611.0/65536.0,1,-nbitq), 
to_sfixed(2529.0/65536.0,1,-nbitq), 
to_sfixed(5181.0/65536.0,1,-nbitq), 
to_sfixed(-7509.0/65536.0,1,-nbitq), 
to_sfixed(-4461.0/65536.0,1,-nbitq), 
to_sfixed(1140.0/65536.0,1,-nbitq), 
to_sfixed(5335.0/65536.0,1,-nbitq), 
to_sfixed(1232.0/65536.0,1,-nbitq), 
to_sfixed(1704.0/65536.0,1,-nbitq), 
to_sfixed(2995.0/65536.0,1,-nbitq), 
to_sfixed(11497.0/65536.0,1,-nbitq), 
to_sfixed(1926.0/65536.0,1,-nbitq), 
to_sfixed(15822.0/65536.0,1,-nbitq), 
to_sfixed(5784.0/65536.0,1,-nbitq), 
to_sfixed(-664.0/65536.0,1,-nbitq), 
to_sfixed(-2234.0/65536.0,1,-nbitq), 
to_sfixed(5564.0/65536.0,1,-nbitq), 
to_sfixed(3733.0/65536.0,1,-nbitq), 
to_sfixed(-2665.0/65536.0,1,-nbitq), 
to_sfixed(8353.0/65536.0,1,-nbitq), 
to_sfixed(5911.0/65536.0,1,-nbitq), 
to_sfixed(-3277.0/65536.0,1,-nbitq), 
to_sfixed(-4993.0/65536.0,1,-nbitq), 
to_sfixed(-827.0/65536.0,1,-nbitq), 
to_sfixed(-4266.0/65536.0,1,-nbitq), 
to_sfixed(18043.0/65536.0,1,-nbitq), 
to_sfixed(-4148.0/65536.0,1,-nbitq), 
to_sfixed(-2885.0/65536.0,1,-nbitq), 
to_sfixed(-1955.0/65536.0,1,-nbitq), 
to_sfixed(-1560.0/65536.0,1,-nbitq), 
to_sfixed(4205.0/65536.0,1,-nbitq), 
to_sfixed(7471.0/65536.0,1,-nbitq), 
to_sfixed(6106.0/65536.0,1,-nbitq), 
to_sfixed(-1901.0/65536.0,1,-nbitq), 
to_sfixed(2026.0/65536.0,1,-nbitq), 
to_sfixed(7645.0/65536.0,1,-nbitq), 
to_sfixed(2282.0/65536.0,1,-nbitq), 
to_sfixed(-216.0/65536.0,1,-nbitq), 
to_sfixed(5068.0/65536.0,1,-nbitq), 
to_sfixed(-10678.0/65536.0,1,-nbitq), 
to_sfixed(1988.0/65536.0,1,-nbitq), 
to_sfixed(14367.0/65536.0,1,-nbitq), 
to_sfixed(4098.0/65536.0,1,-nbitq), 
to_sfixed(-2434.0/65536.0,1,-nbitq), 
to_sfixed(-12624.0/65536.0,1,-nbitq), 
to_sfixed(40.0/65536.0,1,-nbitq), 
to_sfixed(3636.0/65536.0,1,-nbitq), 
to_sfixed(1549.0/65536.0,1,-nbitq), 
to_sfixed(5018.0/65536.0,1,-nbitq), 
to_sfixed(-1233.0/65536.0,1,-nbitq), 
to_sfixed(6278.0/65536.0,1,-nbitq), 
to_sfixed(4554.0/65536.0,1,-nbitq), 
to_sfixed(15485.0/65536.0,1,-nbitq), 
to_sfixed(3162.0/65536.0,1,-nbitq), 
to_sfixed(4114.0/65536.0,1,-nbitq), 
to_sfixed(-72.0/65536.0,1,-nbitq), 
to_sfixed(-3921.0/65536.0,1,-nbitq), 
to_sfixed(-1983.0/65536.0,1,-nbitq), 
to_sfixed(-1374.0/65536.0,1,-nbitq), 
to_sfixed(5509.0/65536.0,1,-nbitq), 
to_sfixed(1612.0/65536.0,1,-nbitq), 
to_sfixed(-1907.0/65536.0,1,-nbitq), 
to_sfixed(1790.0/65536.0,1,-nbitq), 
to_sfixed(-4708.0/65536.0,1,-nbitq), 
to_sfixed(1835.0/65536.0,1,-nbitq), 
to_sfixed(-9701.0/65536.0,1,-nbitq), 
to_sfixed(929.0/65536.0,1,-nbitq), 
to_sfixed(-6376.0/65536.0,1,-nbitq), 
to_sfixed(-5058.0/65536.0,1,-nbitq), 
to_sfixed(-1433.0/65536.0,1,-nbitq), 
to_sfixed(5389.0/65536.0,1,-nbitq), 
to_sfixed(-2746.0/65536.0,1,-nbitq), 
to_sfixed(1638.0/65536.0,1,-nbitq), 
to_sfixed(-2649.0/65536.0,1,-nbitq), 
to_sfixed(6322.0/65536.0,1,-nbitq), 
to_sfixed(3445.0/65536.0,1,-nbitq), 
to_sfixed(-6023.0/65536.0,1,-nbitq), 
to_sfixed(77.0/65536.0,1,-nbitq), 
to_sfixed(-1191.0/65536.0,1,-nbitq)  ), 
( to_sfixed(6630.0/65536.0,1,-nbitq), 
to_sfixed(-1601.0/65536.0,1,-nbitq), 
to_sfixed(2989.0/65536.0,1,-nbitq), 
to_sfixed(2944.0/65536.0,1,-nbitq), 
to_sfixed(-1587.0/65536.0,1,-nbitq), 
to_sfixed(-8901.0/65536.0,1,-nbitq), 
to_sfixed(3081.0/65536.0,1,-nbitq), 
to_sfixed(151.0/65536.0,1,-nbitq), 
to_sfixed(820.0/65536.0,1,-nbitq), 
to_sfixed(-2422.0/65536.0,1,-nbitq), 
to_sfixed(2907.0/65536.0,1,-nbitq), 
to_sfixed(3160.0/65536.0,1,-nbitq), 
to_sfixed(5131.0/65536.0,1,-nbitq), 
to_sfixed(1228.0/65536.0,1,-nbitq), 
to_sfixed(-1666.0/65536.0,1,-nbitq), 
to_sfixed(-3200.0/65536.0,1,-nbitq), 
to_sfixed(-1931.0/65536.0,1,-nbitq), 
to_sfixed(7660.0/65536.0,1,-nbitq), 
to_sfixed(-1118.0/65536.0,1,-nbitq), 
to_sfixed(865.0/65536.0,1,-nbitq), 
to_sfixed(10685.0/65536.0,1,-nbitq), 
to_sfixed(1016.0/65536.0,1,-nbitq), 
to_sfixed(2783.0/65536.0,1,-nbitq), 
to_sfixed(1308.0/65536.0,1,-nbitq), 
to_sfixed(3993.0/65536.0,1,-nbitq), 
to_sfixed(-280.0/65536.0,1,-nbitq), 
to_sfixed(20250.0/65536.0,1,-nbitq), 
to_sfixed(87.0/65536.0,1,-nbitq), 
to_sfixed(-8565.0/65536.0,1,-nbitq), 
to_sfixed(-5541.0/65536.0,1,-nbitq), 
to_sfixed(-3795.0/65536.0,1,-nbitq), 
to_sfixed(3537.0/65536.0,1,-nbitq), 
to_sfixed(3582.0/65536.0,1,-nbitq), 
to_sfixed(1511.0/65536.0,1,-nbitq), 
to_sfixed(1978.0/65536.0,1,-nbitq), 
to_sfixed(586.0/65536.0,1,-nbitq), 
to_sfixed(19566.0/65536.0,1,-nbitq), 
to_sfixed(-5864.0/65536.0,1,-nbitq), 
to_sfixed(-969.0/65536.0,1,-nbitq), 
to_sfixed(-1565.0/65536.0,1,-nbitq), 
to_sfixed(-5410.0/65536.0,1,-nbitq), 
to_sfixed(581.0/65536.0,1,-nbitq), 
to_sfixed(6843.0/65536.0,1,-nbitq), 
to_sfixed(-43.0/65536.0,1,-nbitq), 
to_sfixed(-786.0/65536.0,1,-nbitq), 
to_sfixed(-13463.0/65536.0,1,-nbitq), 
to_sfixed(-3167.0/65536.0,1,-nbitq), 
to_sfixed(5567.0/65536.0,1,-nbitq), 
to_sfixed(-158.0/65536.0,1,-nbitq), 
to_sfixed(1473.0/65536.0,1,-nbitq), 
to_sfixed(207.0/65536.0,1,-nbitq), 
to_sfixed(6063.0/65536.0,1,-nbitq), 
to_sfixed(997.0/65536.0,1,-nbitq), 
to_sfixed(8896.0/65536.0,1,-nbitq), 
to_sfixed(1415.0/65536.0,1,-nbitq), 
to_sfixed(9974.0/65536.0,1,-nbitq), 
to_sfixed(1601.0/65536.0,1,-nbitq), 
to_sfixed(-2389.0/65536.0,1,-nbitq), 
to_sfixed(-2953.0/65536.0,1,-nbitq), 
to_sfixed(3780.0/65536.0,1,-nbitq), 
to_sfixed(11698.0/65536.0,1,-nbitq), 
to_sfixed(2322.0/65536.0,1,-nbitq), 
to_sfixed(-2269.0/65536.0,1,-nbitq), 
to_sfixed(-1859.0/65536.0,1,-nbitq), 
to_sfixed(-6397.0/65536.0,1,-nbitq), 
to_sfixed(-5307.0/65536.0,1,-nbitq), 
to_sfixed(-4858.0/65536.0,1,-nbitq), 
to_sfixed(-4153.0/65536.0,1,-nbitq), 
to_sfixed(-6840.0/65536.0,1,-nbitq), 
to_sfixed(-2604.0/65536.0,1,-nbitq), 
to_sfixed(-778.0/65536.0,1,-nbitq), 
to_sfixed(9983.0/65536.0,1,-nbitq), 
to_sfixed(-7601.0/65536.0,1,-nbitq), 
to_sfixed(112.0/65536.0,1,-nbitq), 
to_sfixed(-2745.0/65536.0,1,-nbitq), 
to_sfixed(4007.0/65536.0,1,-nbitq), 
to_sfixed(148.0/65536.0,1,-nbitq), 
to_sfixed(-19411.0/65536.0,1,-nbitq), 
to_sfixed(2629.0/65536.0,1,-nbitq), 
to_sfixed(-3111.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3822.0/65536.0,1,-nbitq), 
to_sfixed(-8434.0/65536.0,1,-nbitq), 
to_sfixed(-7425.0/65536.0,1,-nbitq), 
to_sfixed(5437.0/65536.0,1,-nbitq), 
to_sfixed(10471.0/65536.0,1,-nbitq), 
to_sfixed(-11932.0/65536.0,1,-nbitq), 
to_sfixed(3288.0/65536.0,1,-nbitq), 
to_sfixed(-9450.0/65536.0,1,-nbitq), 
to_sfixed(-1460.0/65536.0,1,-nbitq), 
to_sfixed(553.0/65536.0,1,-nbitq), 
to_sfixed(1142.0/65536.0,1,-nbitq), 
to_sfixed(8523.0/65536.0,1,-nbitq), 
to_sfixed(1898.0/65536.0,1,-nbitq), 
to_sfixed(-10462.0/65536.0,1,-nbitq), 
to_sfixed(-3343.0/65536.0,1,-nbitq), 
to_sfixed(1393.0/65536.0,1,-nbitq), 
to_sfixed(2373.0/65536.0,1,-nbitq), 
to_sfixed(6479.0/65536.0,1,-nbitq), 
to_sfixed(-13231.0/65536.0,1,-nbitq), 
to_sfixed(1743.0/65536.0,1,-nbitq), 
to_sfixed(498.0/65536.0,1,-nbitq), 
to_sfixed(-3254.0/65536.0,1,-nbitq), 
to_sfixed(3241.0/65536.0,1,-nbitq), 
to_sfixed(5702.0/65536.0,1,-nbitq), 
to_sfixed(2425.0/65536.0,1,-nbitq), 
to_sfixed(-4946.0/65536.0,1,-nbitq), 
to_sfixed(24100.0/65536.0,1,-nbitq), 
to_sfixed(1413.0/65536.0,1,-nbitq), 
to_sfixed(-6644.0/65536.0,1,-nbitq), 
to_sfixed(-2897.0/65536.0,1,-nbitq), 
to_sfixed(-2873.0/65536.0,1,-nbitq), 
to_sfixed(10942.0/65536.0,1,-nbitq), 
to_sfixed(3094.0/65536.0,1,-nbitq), 
to_sfixed(7340.0/65536.0,1,-nbitq), 
to_sfixed(-1411.0/65536.0,1,-nbitq), 
to_sfixed(-4415.0/65536.0,1,-nbitq), 
to_sfixed(14748.0/65536.0,1,-nbitq), 
to_sfixed(-4878.0/65536.0,1,-nbitq), 
to_sfixed(-4961.0/65536.0,1,-nbitq), 
to_sfixed(-299.0/65536.0,1,-nbitq), 
to_sfixed(-5906.0/65536.0,1,-nbitq), 
to_sfixed(613.0/65536.0,1,-nbitq), 
to_sfixed(-2326.0/65536.0,1,-nbitq), 
to_sfixed(2547.0/65536.0,1,-nbitq), 
to_sfixed(1988.0/65536.0,1,-nbitq), 
to_sfixed(-9797.0/65536.0,1,-nbitq), 
to_sfixed(1903.0/65536.0,1,-nbitq), 
to_sfixed(2728.0/65536.0,1,-nbitq), 
to_sfixed(-741.0/65536.0,1,-nbitq), 
to_sfixed(-464.0/65536.0,1,-nbitq), 
to_sfixed(-1478.0/65536.0,1,-nbitq), 
to_sfixed(5177.0/65536.0,1,-nbitq), 
to_sfixed(-3634.0/65536.0,1,-nbitq), 
to_sfixed(4651.0/65536.0,1,-nbitq), 
to_sfixed(-6224.0/65536.0,1,-nbitq), 
to_sfixed(9769.0/65536.0,1,-nbitq), 
to_sfixed(-1051.0/65536.0,1,-nbitq), 
to_sfixed(426.0/65536.0,1,-nbitq), 
to_sfixed(-1795.0/65536.0,1,-nbitq), 
to_sfixed(4238.0/65536.0,1,-nbitq), 
to_sfixed(12404.0/65536.0,1,-nbitq), 
to_sfixed(-1501.0/65536.0,1,-nbitq), 
to_sfixed(1310.0/65536.0,1,-nbitq), 
to_sfixed(-3094.0/65536.0,1,-nbitq), 
to_sfixed(-8967.0/65536.0,1,-nbitq), 
to_sfixed(-5721.0/65536.0,1,-nbitq), 
to_sfixed(-2076.0/65536.0,1,-nbitq), 
to_sfixed(-3239.0/65536.0,1,-nbitq), 
to_sfixed(-9136.0/65536.0,1,-nbitq), 
to_sfixed(2732.0/65536.0,1,-nbitq), 
to_sfixed(371.0/65536.0,1,-nbitq), 
to_sfixed(11121.0/65536.0,1,-nbitq), 
to_sfixed(-4697.0/65536.0,1,-nbitq), 
to_sfixed(-2595.0/65536.0,1,-nbitq), 
to_sfixed(-38.0/65536.0,1,-nbitq), 
to_sfixed(-4604.0/65536.0,1,-nbitq), 
to_sfixed(-1657.0/65536.0,1,-nbitq), 
to_sfixed(-10770.0/65536.0,1,-nbitq), 
to_sfixed(-680.0/65536.0,1,-nbitq), 
to_sfixed(-6254.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3911.0/65536.0,1,-nbitq), 
to_sfixed(-10705.0/65536.0,1,-nbitq), 
to_sfixed(-16988.0/65536.0,1,-nbitq), 
to_sfixed(9870.0/65536.0,1,-nbitq), 
to_sfixed(14006.0/65536.0,1,-nbitq), 
to_sfixed(-16340.0/65536.0,1,-nbitq), 
to_sfixed(1947.0/65536.0,1,-nbitq), 
to_sfixed(-15893.0/65536.0,1,-nbitq), 
to_sfixed(-4723.0/65536.0,1,-nbitq), 
to_sfixed(2875.0/65536.0,1,-nbitq), 
to_sfixed(1360.0/65536.0,1,-nbitq), 
to_sfixed(11729.0/65536.0,1,-nbitq), 
to_sfixed(1585.0/65536.0,1,-nbitq), 
to_sfixed(-1584.0/65536.0,1,-nbitq), 
to_sfixed(-6131.0/65536.0,1,-nbitq), 
to_sfixed(159.0/65536.0,1,-nbitq), 
to_sfixed(1814.0/65536.0,1,-nbitq), 
to_sfixed(-16595.0/65536.0,1,-nbitq), 
to_sfixed(-11617.0/65536.0,1,-nbitq), 
to_sfixed(-496.0/65536.0,1,-nbitq), 
to_sfixed(3190.0/65536.0,1,-nbitq), 
to_sfixed(-12661.0/65536.0,1,-nbitq), 
to_sfixed(15266.0/65536.0,1,-nbitq), 
to_sfixed(6693.0/65536.0,1,-nbitq), 
to_sfixed(510.0/65536.0,1,-nbitq), 
to_sfixed(-4417.0/65536.0,1,-nbitq), 
to_sfixed(18397.0/65536.0,1,-nbitq), 
to_sfixed(-669.0/65536.0,1,-nbitq), 
to_sfixed(-5092.0/65536.0,1,-nbitq), 
to_sfixed(-3079.0/65536.0,1,-nbitq), 
to_sfixed(-3247.0/65536.0,1,-nbitq), 
to_sfixed(5511.0/65536.0,1,-nbitq), 
to_sfixed(2350.0/65536.0,1,-nbitq), 
to_sfixed(-5267.0/65536.0,1,-nbitq), 
to_sfixed(-217.0/65536.0,1,-nbitq), 
to_sfixed(1865.0/65536.0,1,-nbitq), 
to_sfixed(9011.0/65536.0,1,-nbitq), 
to_sfixed(-9864.0/65536.0,1,-nbitq), 
to_sfixed(-14731.0/65536.0,1,-nbitq), 
to_sfixed(-3584.0/65536.0,1,-nbitq), 
to_sfixed(-8723.0/65536.0,1,-nbitq), 
to_sfixed(1915.0/65536.0,1,-nbitq), 
to_sfixed(-6343.0/65536.0,1,-nbitq), 
to_sfixed(4213.0/65536.0,1,-nbitq), 
to_sfixed(1243.0/65536.0,1,-nbitq), 
to_sfixed(10640.0/65536.0,1,-nbitq), 
to_sfixed(1392.0/65536.0,1,-nbitq), 
to_sfixed(-8932.0/65536.0,1,-nbitq), 
to_sfixed(2360.0/65536.0,1,-nbitq), 
to_sfixed(-164.0/65536.0,1,-nbitq), 
to_sfixed(2293.0/65536.0,1,-nbitq), 
to_sfixed(7392.0/65536.0,1,-nbitq), 
to_sfixed(-743.0/65536.0,1,-nbitq), 
to_sfixed(-959.0/65536.0,1,-nbitq), 
to_sfixed(-4229.0/65536.0,1,-nbitq), 
to_sfixed(7241.0/65536.0,1,-nbitq), 
to_sfixed(-2020.0/65536.0,1,-nbitq), 
to_sfixed(-488.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(-1125.0/65536.0,1,-nbitq), 
to_sfixed(10967.0/65536.0,1,-nbitq), 
to_sfixed(-1336.0/65536.0,1,-nbitq), 
to_sfixed(232.0/65536.0,1,-nbitq), 
to_sfixed(1590.0/65536.0,1,-nbitq), 
to_sfixed(-8324.0/65536.0,1,-nbitq), 
to_sfixed(-16011.0/65536.0,1,-nbitq), 
to_sfixed(-10658.0/65536.0,1,-nbitq), 
to_sfixed(-13336.0/65536.0,1,-nbitq), 
to_sfixed(-16594.0/65536.0,1,-nbitq), 
to_sfixed(6500.0/65536.0,1,-nbitq), 
to_sfixed(2006.0/65536.0,1,-nbitq), 
to_sfixed(15762.0/65536.0,1,-nbitq), 
to_sfixed(-3984.0/65536.0,1,-nbitq), 
to_sfixed(-19.0/65536.0,1,-nbitq), 
to_sfixed(-107.0/65536.0,1,-nbitq), 
to_sfixed(-12941.0/65536.0,1,-nbitq), 
to_sfixed(-5013.0/65536.0,1,-nbitq), 
to_sfixed(4327.0/65536.0,1,-nbitq), 
to_sfixed(-2729.0/65536.0,1,-nbitq), 
to_sfixed(-9460.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1905.0/65536.0,1,-nbitq), 
to_sfixed(-6316.0/65536.0,1,-nbitq), 
to_sfixed(-15734.0/65536.0,1,-nbitq), 
to_sfixed(8159.0/65536.0,1,-nbitq), 
to_sfixed(17929.0/65536.0,1,-nbitq), 
to_sfixed(-15193.0/65536.0,1,-nbitq), 
to_sfixed(-1283.0/65536.0,1,-nbitq), 
to_sfixed(-8543.0/65536.0,1,-nbitq), 
to_sfixed(425.0/65536.0,1,-nbitq), 
to_sfixed(-1108.0/65536.0,1,-nbitq), 
to_sfixed(8801.0/65536.0,1,-nbitq), 
to_sfixed(12173.0/65536.0,1,-nbitq), 
to_sfixed(-336.0/65536.0,1,-nbitq), 
to_sfixed(-13757.0/65536.0,1,-nbitq), 
to_sfixed(-7362.0/65536.0,1,-nbitq), 
to_sfixed(3214.0/65536.0,1,-nbitq), 
to_sfixed(-1860.0/65536.0,1,-nbitq), 
to_sfixed(-7548.0/65536.0,1,-nbitq), 
to_sfixed(-9078.0/65536.0,1,-nbitq), 
to_sfixed(-1947.0/65536.0,1,-nbitq), 
to_sfixed(13425.0/65536.0,1,-nbitq), 
to_sfixed(-12656.0/65536.0,1,-nbitq), 
to_sfixed(11678.0/65536.0,1,-nbitq), 
to_sfixed(8245.0/65536.0,1,-nbitq), 
to_sfixed(-399.0/65536.0,1,-nbitq), 
to_sfixed(-7170.0/65536.0,1,-nbitq), 
to_sfixed(15606.0/65536.0,1,-nbitq), 
to_sfixed(-20.0/65536.0,1,-nbitq), 
to_sfixed(-5439.0/65536.0,1,-nbitq), 
to_sfixed(-4845.0/65536.0,1,-nbitq), 
to_sfixed(-833.0/65536.0,1,-nbitq), 
to_sfixed(4066.0/65536.0,1,-nbitq), 
to_sfixed(11329.0/65536.0,1,-nbitq), 
to_sfixed(-11264.0/65536.0,1,-nbitq), 
to_sfixed(1987.0/65536.0,1,-nbitq), 
to_sfixed(2746.0/65536.0,1,-nbitq), 
to_sfixed(-2081.0/65536.0,1,-nbitq), 
to_sfixed(2222.0/65536.0,1,-nbitq), 
to_sfixed(-8584.0/65536.0,1,-nbitq), 
to_sfixed(-8125.0/65536.0,1,-nbitq), 
to_sfixed(-4216.0/65536.0,1,-nbitq), 
to_sfixed(-1987.0/65536.0,1,-nbitq), 
to_sfixed(2480.0/65536.0,1,-nbitq), 
to_sfixed(8562.0/65536.0,1,-nbitq), 
to_sfixed(-1520.0/65536.0,1,-nbitq), 
to_sfixed(7441.0/65536.0,1,-nbitq), 
to_sfixed(768.0/65536.0,1,-nbitq), 
to_sfixed(-4506.0/65536.0,1,-nbitq), 
to_sfixed(3770.0/65536.0,1,-nbitq), 
to_sfixed(500.0/65536.0,1,-nbitq), 
to_sfixed(-379.0/65536.0,1,-nbitq), 
to_sfixed(10318.0/65536.0,1,-nbitq), 
to_sfixed(-7514.0/65536.0,1,-nbitq), 
to_sfixed(1321.0/65536.0,1,-nbitq), 
to_sfixed(-3915.0/65536.0,1,-nbitq), 
to_sfixed(9969.0/65536.0,1,-nbitq), 
to_sfixed(-149.0/65536.0,1,-nbitq), 
to_sfixed(4063.0/65536.0,1,-nbitq), 
to_sfixed(1648.0/65536.0,1,-nbitq), 
to_sfixed(-534.0/65536.0,1,-nbitq), 
to_sfixed(-847.0/65536.0,1,-nbitq), 
to_sfixed(2008.0/65536.0,1,-nbitq), 
to_sfixed(914.0/65536.0,1,-nbitq), 
to_sfixed(2594.0/65536.0,1,-nbitq), 
to_sfixed(-16934.0/65536.0,1,-nbitq), 
to_sfixed(-9138.0/65536.0,1,-nbitq), 
to_sfixed(-13739.0/65536.0,1,-nbitq), 
to_sfixed(-4239.0/65536.0,1,-nbitq), 
to_sfixed(-15485.0/65536.0,1,-nbitq), 
to_sfixed(9867.0/65536.0,1,-nbitq), 
to_sfixed(-3553.0/65536.0,1,-nbitq), 
to_sfixed(9447.0/65536.0,1,-nbitq), 
to_sfixed(-9236.0/65536.0,1,-nbitq), 
to_sfixed(-1034.0/65536.0,1,-nbitq), 
to_sfixed(-2671.0/65536.0,1,-nbitq), 
to_sfixed(-15673.0/65536.0,1,-nbitq), 
to_sfixed(-14341.0/65536.0,1,-nbitq), 
to_sfixed(10943.0/65536.0,1,-nbitq), 
to_sfixed(1604.0/65536.0,1,-nbitq), 
to_sfixed(-4875.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1256.0/65536.0,1,-nbitq), 
to_sfixed(-5194.0/65536.0,1,-nbitq), 
to_sfixed(11946.0/65536.0,1,-nbitq), 
to_sfixed(-1164.0/65536.0,1,-nbitq), 
to_sfixed(98.0/65536.0,1,-nbitq), 
to_sfixed(-10663.0/65536.0,1,-nbitq), 
to_sfixed(-1034.0/65536.0,1,-nbitq), 
to_sfixed(3236.0/65536.0,1,-nbitq), 
to_sfixed(-3217.0/65536.0,1,-nbitq), 
to_sfixed(137.0/65536.0,1,-nbitq), 
to_sfixed(6842.0/65536.0,1,-nbitq), 
to_sfixed(15329.0/65536.0,1,-nbitq), 
to_sfixed(-1492.0/65536.0,1,-nbitq), 
to_sfixed(-9473.0/65536.0,1,-nbitq), 
to_sfixed(-5687.0/65536.0,1,-nbitq), 
to_sfixed(-1807.0/65536.0,1,-nbitq), 
to_sfixed(1867.0/65536.0,1,-nbitq), 
to_sfixed(1918.0/65536.0,1,-nbitq), 
to_sfixed(735.0/65536.0,1,-nbitq), 
to_sfixed(-176.0/65536.0,1,-nbitq), 
to_sfixed(5394.0/65536.0,1,-nbitq), 
to_sfixed(-10308.0/65536.0,1,-nbitq), 
to_sfixed(-3019.0/65536.0,1,-nbitq), 
to_sfixed(7749.0/65536.0,1,-nbitq), 
to_sfixed(1603.0/65536.0,1,-nbitq), 
to_sfixed(1579.0/65536.0,1,-nbitq), 
to_sfixed(11483.0/65536.0,1,-nbitq), 
to_sfixed(-1473.0/65536.0,1,-nbitq), 
to_sfixed(-7009.0/65536.0,1,-nbitq), 
to_sfixed(4739.0/65536.0,1,-nbitq), 
to_sfixed(4400.0/65536.0,1,-nbitq), 
to_sfixed(8106.0/65536.0,1,-nbitq), 
to_sfixed(976.0/65536.0,1,-nbitq), 
to_sfixed(-1161.0/65536.0,1,-nbitq), 
to_sfixed(-27.0/65536.0,1,-nbitq), 
to_sfixed(576.0/65536.0,1,-nbitq), 
to_sfixed(756.0/65536.0,1,-nbitq), 
to_sfixed(3692.0/65536.0,1,-nbitq), 
to_sfixed(12058.0/65536.0,1,-nbitq), 
to_sfixed(-3688.0/65536.0,1,-nbitq), 
to_sfixed(-8723.0/65536.0,1,-nbitq), 
to_sfixed(-1066.0/65536.0,1,-nbitq), 
to_sfixed(-3627.0/65536.0,1,-nbitq), 
to_sfixed(7120.0/65536.0,1,-nbitq), 
to_sfixed(2168.0/65536.0,1,-nbitq), 
to_sfixed(8327.0/65536.0,1,-nbitq), 
to_sfixed(2474.0/65536.0,1,-nbitq), 
to_sfixed(-4930.0/65536.0,1,-nbitq), 
to_sfixed(655.0/65536.0,1,-nbitq), 
to_sfixed(-3193.0/65536.0,1,-nbitq), 
to_sfixed(-2568.0/65536.0,1,-nbitq), 
to_sfixed(14399.0/65536.0,1,-nbitq), 
to_sfixed(-3989.0/65536.0,1,-nbitq), 
to_sfixed(3276.0/65536.0,1,-nbitq), 
to_sfixed(-7506.0/65536.0,1,-nbitq), 
to_sfixed(4134.0/65536.0,1,-nbitq), 
to_sfixed(1902.0/65536.0,1,-nbitq), 
to_sfixed(-68.0/65536.0,1,-nbitq), 
to_sfixed(2314.0/65536.0,1,-nbitq), 
to_sfixed(-413.0/65536.0,1,-nbitq), 
to_sfixed(-3793.0/65536.0,1,-nbitq), 
to_sfixed(54.0/65536.0,1,-nbitq), 
to_sfixed(-88.0/65536.0,1,-nbitq), 
to_sfixed(317.0/65536.0,1,-nbitq), 
to_sfixed(-6716.0/65536.0,1,-nbitq), 
to_sfixed(-2337.0/65536.0,1,-nbitq), 
to_sfixed(-12485.0/65536.0,1,-nbitq), 
to_sfixed(-4396.0/65536.0,1,-nbitq), 
to_sfixed(-702.0/65536.0,1,-nbitq), 
to_sfixed(-1976.0/65536.0,1,-nbitq), 
to_sfixed(-2627.0/65536.0,1,-nbitq), 
to_sfixed(75.0/65536.0,1,-nbitq), 
to_sfixed(-22778.0/65536.0,1,-nbitq), 
to_sfixed(537.0/65536.0,1,-nbitq), 
to_sfixed(-2165.0/65536.0,1,-nbitq), 
to_sfixed(-11630.0/65536.0,1,-nbitq), 
to_sfixed(-12123.0/65536.0,1,-nbitq), 
to_sfixed(5112.0/65536.0,1,-nbitq), 
to_sfixed(-1772.0/65536.0,1,-nbitq), 
to_sfixed(10183.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2789.0/65536.0,1,-nbitq), 
to_sfixed(-1171.0/65536.0,1,-nbitq), 
to_sfixed(12136.0/65536.0,1,-nbitq), 
to_sfixed(-11161.0/65536.0,1,-nbitq), 
to_sfixed(-1607.0/65536.0,1,-nbitq), 
to_sfixed(16184.0/65536.0,1,-nbitq), 
to_sfixed(-3057.0/65536.0,1,-nbitq), 
to_sfixed(9699.0/65536.0,1,-nbitq), 
to_sfixed(4012.0/65536.0,1,-nbitq), 
to_sfixed(1330.0/65536.0,1,-nbitq), 
to_sfixed(10192.0/65536.0,1,-nbitq), 
to_sfixed(6680.0/65536.0,1,-nbitq), 
to_sfixed(-2189.0/65536.0,1,-nbitq), 
to_sfixed(-6455.0/65536.0,1,-nbitq), 
to_sfixed(1037.0/65536.0,1,-nbitq), 
to_sfixed(604.0/65536.0,1,-nbitq), 
to_sfixed(-2718.0/65536.0,1,-nbitq), 
to_sfixed(1977.0/65536.0,1,-nbitq), 
to_sfixed(3310.0/65536.0,1,-nbitq), 
to_sfixed(-571.0/65536.0,1,-nbitq), 
to_sfixed(4582.0/65536.0,1,-nbitq), 
to_sfixed(-13354.0/65536.0,1,-nbitq), 
to_sfixed(-14576.0/65536.0,1,-nbitq), 
to_sfixed(12143.0/65536.0,1,-nbitq), 
to_sfixed(-1829.0/65536.0,1,-nbitq), 
to_sfixed(7638.0/65536.0,1,-nbitq), 
to_sfixed(12114.0/65536.0,1,-nbitq), 
to_sfixed(3761.0/65536.0,1,-nbitq), 
to_sfixed(-806.0/65536.0,1,-nbitq), 
to_sfixed(6681.0/65536.0,1,-nbitq), 
to_sfixed(3601.0/65536.0,1,-nbitq), 
to_sfixed(5582.0/65536.0,1,-nbitq), 
to_sfixed(-10649.0/65536.0,1,-nbitq), 
to_sfixed(1024.0/65536.0,1,-nbitq), 
to_sfixed(-2094.0/65536.0,1,-nbitq), 
to_sfixed(-80.0/65536.0,1,-nbitq), 
to_sfixed(10359.0/65536.0,1,-nbitq), 
to_sfixed(9847.0/65536.0,1,-nbitq), 
to_sfixed(963.0/65536.0,1,-nbitq), 
to_sfixed(953.0/65536.0,1,-nbitq), 
to_sfixed(-9842.0/65536.0,1,-nbitq), 
to_sfixed(-1082.0/65536.0,1,-nbitq), 
to_sfixed(-3597.0/65536.0,1,-nbitq), 
to_sfixed(1733.0/65536.0,1,-nbitq), 
to_sfixed(-681.0/65536.0,1,-nbitq), 
to_sfixed(6396.0/65536.0,1,-nbitq), 
to_sfixed(-46.0/65536.0,1,-nbitq), 
to_sfixed(-111.0/65536.0,1,-nbitq), 
to_sfixed(-2486.0/65536.0,1,-nbitq), 
to_sfixed(1579.0/65536.0,1,-nbitq), 
to_sfixed(246.0/65536.0,1,-nbitq), 
to_sfixed(11977.0/65536.0,1,-nbitq), 
to_sfixed(-4907.0/65536.0,1,-nbitq), 
to_sfixed(10261.0/65536.0,1,-nbitq), 
to_sfixed(-480.0/65536.0,1,-nbitq), 
to_sfixed(-19777.0/65536.0,1,-nbitq), 
to_sfixed(2663.0/65536.0,1,-nbitq), 
to_sfixed(123.0/65536.0,1,-nbitq), 
to_sfixed(794.0/65536.0,1,-nbitq), 
to_sfixed(-7825.0/65536.0,1,-nbitq), 
to_sfixed(1027.0/65536.0,1,-nbitq), 
to_sfixed(-385.0/65536.0,1,-nbitq), 
to_sfixed(-1533.0/65536.0,1,-nbitq), 
to_sfixed(-705.0/65536.0,1,-nbitq), 
to_sfixed(-6796.0/65536.0,1,-nbitq), 
to_sfixed(-4027.0/65536.0,1,-nbitq), 
to_sfixed(-3549.0/65536.0,1,-nbitq), 
to_sfixed(2028.0/65536.0,1,-nbitq), 
to_sfixed(1450.0/65536.0,1,-nbitq), 
to_sfixed(-8860.0/65536.0,1,-nbitq), 
to_sfixed(-2707.0/65536.0,1,-nbitq), 
to_sfixed(-6753.0/65536.0,1,-nbitq), 
to_sfixed(-12220.0/65536.0,1,-nbitq), 
to_sfixed(1531.0/65536.0,1,-nbitq), 
to_sfixed(974.0/65536.0,1,-nbitq), 
to_sfixed(-8233.0/65536.0,1,-nbitq), 
to_sfixed(-6789.0/65536.0,1,-nbitq), 
to_sfixed(9456.0/65536.0,1,-nbitq), 
to_sfixed(-2776.0/65536.0,1,-nbitq), 
to_sfixed(11568.0/65536.0,1,-nbitq)  ), 
( to_sfixed(58.0/65536.0,1,-nbitq), 
to_sfixed(5330.0/65536.0,1,-nbitq), 
to_sfixed(5968.0/65536.0,1,-nbitq), 
to_sfixed(-5122.0/65536.0,1,-nbitq), 
to_sfixed(3477.0/65536.0,1,-nbitq), 
to_sfixed(13390.0/65536.0,1,-nbitq), 
to_sfixed(-1858.0/65536.0,1,-nbitq), 
to_sfixed(4971.0/65536.0,1,-nbitq), 
to_sfixed(11762.0/65536.0,1,-nbitq), 
to_sfixed(3186.0/65536.0,1,-nbitq), 
to_sfixed(14029.0/65536.0,1,-nbitq), 
to_sfixed(-1018.0/65536.0,1,-nbitq), 
to_sfixed(-227.0/65536.0,1,-nbitq), 
to_sfixed(-1000.0/65536.0,1,-nbitq), 
to_sfixed(-1112.0/65536.0,1,-nbitq), 
to_sfixed(-1562.0/65536.0,1,-nbitq), 
to_sfixed(-370.0/65536.0,1,-nbitq), 
to_sfixed(-2857.0/65536.0,1,-nbitq), 
to_sfixed(1392.0/65536.0,1,-nbitq), 
to_sfixed(-2563.0/65536.0,1,-nbitq), 
to_sfixed(-225.0/65536.0,1,-nbitq), 
to_sfixed(-18237.0/65536.0,1,-nbitq), 
to_sfixed(-3828.0/65536.0,1,-nbitq), 
to_sfixed(13463.0/65536.0,1,-nbitq), 
to_sfixed(-3826.0/65536.0,1,-nbitq), 
to_sfixed(6765.0/65536.0,1,-nbitq), 
to_sfixed(10414.0/65536.0,1,-nbitq), 
to_sfixed(-337.0/65536.0,1,-nbitq), 
to_sfixed(-550.0/65536.0,1,-nbitq), 
to_sfixed(5125.0/65536.0,1,-nbitq), 
to_sfixed(-1083.0/65536.0,1,-nbitq), 
to_sfixed(-4663.0/65536.0,1,-nbitq), 
to_sfixed(-19813.0/65536.0,1,-nbitq), 
to_sfixed(-1590.0/65536.0,1,-nbitq), 
to_sfixed(14.0/65536.0,1,-nbitq), 
to_sfixed(33.0/65536.0,1,-nbitq), 
to_sfixed(13580.0/65536.0,1,-nbitq), 
to_sfixed(8000.0/65536.0,1,-nbitq), 
to_sfixed(3430.0/65536.0,1,-nbitq), 
to_sfixed(-1063.0/65536.0,1,-nbitq), 
to_sfixed(-9392.0/65536.0,1,-nbitq), 
to_sfixed(-2985.0/65536.0,1,-nbitq), 
to_sfixed(2045.0/65536.0,1,-nbitq), 
to_sfixed(-5362.0/65536.0,1,-nbitq), 
to_sfixed(-1099.0/65536.0,1,-nbitq), 
to_sfixed(-3910.0/65536.0,1,-nbitq), 
to_sfixed(-2203.0/65536.0,1,-nbitq), 
to_sfixed(10166.0/65536.0,1,-nbitq), 
to_sfixed(-844.0/65536.0,1,-nbitq), 
to_sfixed(2800.0/65536.0,1,-nbitq), 
to_sfixed(947.0/65536.0,1,-nbitq), 
to_sfixed(247.0/65536.0,1,-nbitq), 
to_sfixed(-10048.0/65536.0,1,-nbitq), 
to_sfixed(8299.0/65536.0,1,-nbitq), 
to_sfixed(6722.0/65536.0,1,-nbitq), 
to_sfixed(-14845.0/65536.0,1,-nbitq), 
to_sfixed(-1421.0/65536.0,1,-nbitq), 
to_sfixed(-2291.0/65536.0,1,-nbitq), 
to_sfixed(-1580.0/65536.0,1,-nbitq), 
to_sfixed(-7893.0/65536.0,1,-nbitq), 
to_sfixed(1036.0/65536.0,1,-nbitq), 
to_sfixed(-2764.0/65536.0,1,-nbitq), 
to_sfixed(-1578.0/65536.0,1,-nbitq), 
to_sfixed(2762.0/65536.0,1,-nbitq), 
to_sfixed(1377.0/65536.0,1,-nbitq), 
to_sfixed(6153.0/65536.0,1,-nbitq), 
to_sfixed(-4020.0/65536.0,1,-nbitq), 
to_sfixed(-977.0/65536.0,1,-nbitq), 
to_sfixed(822.0/65536.0,1,-nbitq), 
to_sfixed(-7556.0/65536.0,1,-nbitq), 
to_sfixed(508.0/65536.0,1,-nbitq), 
to_sfixed(-2853.0/65536.0,1,-nbitq), 
to_sfixed(15232.0/65536.0,1,-nbitq), 
to_sfixed(714.0/65536.0,1,-nbitq), 
to_sfixed(2419.0/65536.0,1,-nbitq), 
to_sfixed(-3732.0/65536.0,1,-nbitq), 
to_sfixed(-4798.0/65536.0,1,-nbitq), 
to_sfixed(17994.0/65536.0,1,-nbitq), 
to_sfixed(-1138.0/65536.0,1,-nbitq), 
to_sfixed(9865.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5485.0/65536.0,1,-nbitq), 
to_sfixed(7591.0/65536.0,1,-nbitq), 
to_sfixed(-8489.0/65536.0,1,-nbitq), 
to_sfixed(-3528.0/65536.0,1,-nbitq), 
to_sfixed(-881.0/65536.0,1,-nbitq), 
to_sfixed(11845.0/65536.0,1,-nbitq), 
to_sfixed(1685.0/65536.0,1,-nbitq), 
to_sfixed(1954.0/65536.0,1,-nbitq), 
to_sfixed(16036.0/65536.0,1,-nbitq), 
to_sfixed(1466.0/65536.0,1,-nbitq), 
to_sfixed(9720.0/65536.0,1,-nbitq), 
to_sfixed(-924.0/65536.0,1,-nbitq), 
to_sfixed(-177.0/65536.0,1,-nbitq), 
to_sfixed(773.0/65536.0,1,-nbitq), 
to_sfixed(2402.0/65536.0,1,-nbitq), 
to_sfixed(3627.0/65536.0,1,-nbitq), 
to_sfixed(2614.0/65536.0,1,-nbitq), 
to_sfixed(5870.0/65536.0,1,-nbitq), 
to_sfixed(-4604.0/65536.0,1,-nbitq), 
to_sfixed(-2961.0/65536.0,1,-nbitq), 
to_sfixed(4509.0/65536.0,1,-nbitq), 
to_sfixed(-14605.0/65536.0,1,-nbitq), 
to_sfixed(-5619.0/65536.0,1,-nbitq), 
to_sfixed(6440.0/65536.0,1,-nbitq), 
to_sfixed(-1494.0/65536.0,1,-nbitq), 
to_sfixed(4825.0/65536.0,1,-nbitq), 
to_sfixed(7494.0/65536.0,1,-nbitq), 
to_sfixed(801.0/65536.0,1,-nbitq), 
to_sfixed(98.0/65536.0,1,-nbitq), 
to_sfixed(1358.0/65536.0,1,-nbitq), 
to_sfixed(-4826.0/65536.0,1,-nbitq), 
to_sfixed(-12101.0/65536.0,1,-nbitq), 
to_sfixed(-11310.0/65536.0,1,-nbitq), 
to_sfixed(4786.0/65536.0,1,-nbitq), 
to_sfixed(38.0/65536.0,1,-nbitq), 
to_sfixed(30.0/65536.0,1,-nbitq), 
to_sfixed(10796.0/65536.0,1,-nbitq), 
to_sfixed(35.0/65536.0,1,-nbitq), 
to_sfixed(6259.0/65536.0,1,-nbitq), 
to_sfixed(-577.0/65536.0,1,-nbitq), 
to_sfixed(4516.0/65536.0,1,-nbitq), 
to_sfixed(-2138.0/65536.0,1,-nbitq), 
to_sfixed(1793.0/65536.0,1,-nbitq), 
to_sfixed(-2493.0/65536.0,1,-nbitq), 
to_sfixed(-1113.0/65536.0,1,-nbitq), 
to_sfixed(-9346.0/65536.0,1,-nbitq), 
to_sfixed(-889.0/65536.0,1,-nbitq), 
to_sfixed(4910.0/65536.0,1,-nbitq), 
to_sfixed(-1765.0/65536.0,1,-nbitq), 
to_sfixed(-1979.0/65536.0,1,-nbitq), 
to_sfixed(2309.0/65536.0,1,-nbitq), 
to_sfixed(-3476.0/65536.0,1,-nbitq), 
to_sfixed(-6832.0/65536.0,1,-nbitq), 
to_sfixed(-5262.0/65536.0,1,-nbitq), 
to_sfixed(10675.0/65536.0,1,-nbitq), 
to_sfixed(-5254.0/65536.0,1,-nbitq), 
to_sfixed(2650.0/65536.0,1,-nbitq), 
to_sfixed(-2461.0/65536.0,1,-nbitq), 
to_sfixed(-1170.0/65536.0,1,-nbitq), 
to_sfixed(-867.0/65536.0,1,-nbitq), 
to_sfixed(-4117.0/65536.0,1,-nbitq), 
to_sfixed(-2200.0/65536.0,1,-nbitq), 
to_sfixed(1641.0/65536.0,1,-nbitq), 
to_sfixed(-953.0/65536.0,1,-nbitq), 
to_sfixed(-2477.0/65536.0,1,-nbitq), 
to_sfixed(4714.0/65536.0,1,-nbitq), 
to_sfixed(-2066.0/65536.0,1,-nbitq), 
to_sfixed(7995.0/65536.0,1,-nbitq), 
to_sfixed(-4412.0/65536.0,1,-nbitq), 
to_sfixed(-6965.0/65536.0,1,-nbitq), 
to_sfixed(2162.0/65536.0,1,-nbitq), 
to_sfixed(-2073.0/65536.0,1,-nbitq), 
to_sfixed(20459.0/65536.0,1,-nbitq), 
to_sfixed(2018.0/65536.0,1,-nbitq), 
to_sfixed(1292.0/65536.0,1,-nbitq), 
to_sfixed(4641.0/65536.0,1,-nbitq), 
to_sfixed(-8111.0/65536.0,1,-nbitq), 
to_sfixed(2394.0/65536.0,1,-nbitq), 
to_sfixed(50.0/65536.0,1,-nbitq), 
to_sfixed(8458.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5926.0/65536.0,1,-nbitq), 
to_sfixed(3587.0/65536.0,1,-nbitq), 
to_sfixed(-746.0/65536.0,1,-nbitq), 
to_sfixed(-2753.0/65536.0,1,-nbitq), 
to_sfixed(-1244.0/65536.0,1,-nbitq), 
to_sfixed(10472.0/65536.0,1,-nbitq), 
to_sfixed(1462.0/65536.0,1,-nbitq), 
to_sfixed(4613.0/65536.0,1,-nbitq), 
to_sfixed(9994.0/65536.0,1,-nbitq), 
to_sfixed(-1135.0/65536.0,1,-nbitq), 
to_sfixed(8086.0/65536.0,1,-nbitq), 
to_sfixed(-4243.0/65536.0,1,-nbitq), 
to_sfixed(-3739.0/65536.0,1,-nbitq), 
to_sfixed(8684.0/65536.0,1,-nbitq), 
to_sfixed(4239.0/65536.0,1,-nbitq), 
to_sfixed(2841.0/65536.0,1,-nbitq), 
to_sfixed(2779.0/65536.0,1,-nbitq), 
to_sfixed(7912.0/65536.0,1,-nbitq), 
to_sfixed(-1247.0/65536.0,1,-nbitq), 
to_sfixed(2372.0/65536.0,1,-nbitq), 
to_sfixed(4921.0/65536.0,1,-nbitq), 
to_sfixed(-6057.0/65536.0,1,-nbitq), 
to_sfixed(-3756.0/65536.0,1,-nbitq), 
to_sfixed(6101.0/65536.0,1,-nbitq), 
to_sfixed(-4057.0/65536.0,1,-nbitq), 
to_sfixed(6547.0/65536.0,1,-nbitq), 
to_sfixed(5471.0/65536.0,1,-nbitq), 
to_sfixed(633.0/65536.0,1,-nbitq), 
to_sfixed(117.0/65536.0,1,-nbitq), 
to_sfixed(-2775.0/65536.0,1,-nbitq), 
to_sfixed(-3469.0/65536.0,1,-nbitq), 
to_sfixed(-8225.0/65536.0,1,-nbitq), 
to_sfixed(-8017.0/65536.0,1,-nbitq), 
to_sfixed(11138.0/65536.0,1,-nbitq), 
to_sfixed(-370.0/65536.0,1,-nbitq), 
to_sfixed(-4141.0/65536.0,1,-nbitq), 
to_sfixed(6705.0/65536.0,1,-nbitq), 
to_sfixed(-5708.0/65536.0,1,-nbitq), 
to_sfixed(7138.0/65536.0,1,-nbitq), 
to_sfixed(-384.0/65536.0,1,-nbitq), 
to_sfixed(8096.0/65536.0,1,-nbitq), 
to_sfixed(1583.0/65536.0,1,-nbitq), 
to_sfixed(6962.0/65536.0,1,-nbitq), 
to_sfixed(-2618.0/65536.0,1,-nbitq), 
to_sfixed(-744.0/65536.0,1,-nbitq), 
to_sfixed(-20619.0/65536.0,1,-nbitq), 
to_sfixed(-919.0/65536.0,1,-nbitq), 
to_sfixed(3482.0/65536.0,1,-nbitq), 
to_sfixed(-3979.0/65536.0,1,-nbitq), 
to_sfixed(1320.0/65536.0,1,-nbitq), 
to_sfixed(-2714.0/65536.0,1,-nbitq), 
to_sfixed(-923.0/65536.0,1,-nbitq), 
to_sfixed(-5907.0/65536.0,1,-nbitq), 
to_sfixed(-1192.0/65536.0,1,-nbitq), 
to_sfixed(9434.0/65536.0,1,-nbitq), 
to_sfixed(2276.0/65536.0,1,-nbitq), 
to_sfixed(873.0/65536.0,1,-nbitq), 
to_sfixed(-63.0/65536.0,1,-nbitq), 
to_sfixed(-182.0/65536.0,1,-nbitq), 
to_sfixed(-5557.0/65536.0,1,-nbitq), 
to_sfixed(-9310.0/65536.0,1,-nbitq), 
to_sfixed(90.0/65536.0,1,-nbitq), 
to_sfixed(-2339.0/65536.0,1,-nbitq), 
to_sfixed(2802.0/65536.0,1,-nbitq), 
to_sfixed(-1432.0/65536.0,1,-nbitq), 
to_sfixed(3031.0/65536.0,1,-nbitq), 
to_sfixed(1662.0/65536.0,1,-nbitq), 
to_sfixed(7301.0/65536.0,1,-nbitq), 
to_sfixed(-173.0/65536.0,1,-nbitq), 
to_sfixed(-13601.0/65536.0,1,-nbitq), 
to_sfixed(1246.0/65536.0,1,-nbitq), 
to_sfixed(2183.0/65536.0,1,-nbitq), 
to_sfixed(6695.0/65536.0,1,-nbitq), 
to_sfixed(1912.0/65536.0,1,-nbitq), 
to_sfixed(143.0/65536.0,1,-nbitq), 
to_sfixed(2081.0/65536.0,1,-nbitq), 
to_sfixed(-6469.0/65536.0,1,-nbitq), 
to_sfixed(-10761.0/65536.0,1,-nbitq), 
to_sfixed(-2744.0/65536.0,1,-nbitq), 
to_sfixed(5513.0/65536.0,1,-nbitq)  ), 
( to_sfixed(659.0/65536.0,1,-nbitq), 
to_sfixed(480.0/65536.0,1,-nbitq), 
to_sfixed(-4798.0/65536.0,1,-nbitq), 
to_sfixed(123.0/65536.0,1,-nbitq), 
to_sfixed(12718.0/65536.0,1,-nbitq), 
to_sfixed(13350.0/65536.0,1,-nbitq), 
to_sfixed(-2024.0/65536.0,1,-nbitq), 
to_sfixed(4360.0/65536.0,1,-nbitq), 
to_sfixed(6187.0/65536.0,1,-nbitq), 
to_sfixed(-681.0/65536.0,1,-nbitq), 
to_sfixed(8157.0/65536.0,1,-nbitq), 
to_sfixed(-2617.0/65536.0,1,-nbitq), 
to_sfixed(-322.0/65536.0,1,-nbitq), 
to_sfixed(13261.0/65536.0,1,-nbitq), 
to_sfixed(-362.0/65536.0,1,-nbitq), 
to_sfixed(2671.0/65536.0,1,-nbitq), 
to_sfixed(-1.0/65536.0,1,-nbitq), 
to_sfixed(7066.0/65536.0,1,-nbitq), 
to_sfixed(3240.0/65536.0,1,-nbitq), 
to_sfixed(1577.0/65536.0,1,-nbitq), 
to_sfixed(9983.0/65536.0,1,-nbitq), 
to_sfixed(-10986.0/65536.0,1,-nbitq), 
to_sfixed(-10650.0/65536.0,1,-nbitq), 
to_sfixed(8058.0/65536.0,1,-nbitq), 
to_sfixed(1361.0/65536.0,1,-nbitq), 
to_sfixed(7339.0/65536.0,1,-nbitq), 
to_sfixed(2622.0/65536.0,1,-nbitq), 
to_sfixed(3342.0/65536.0,1,-nbitq), 
to_sfixed(-265.0/65536.0,1,-nbitq), 
to_sfixed(-2020.0/65536.0,1,-nbitq), 
to_sfixed(1798.0/65536.0,1,-nbitq), 
to_sfixed(-8793.0/65536.0,1,-nbitq), 
to_sfixed(-3299.0/65536.0,1,-nbitq), 
to_sfixed(10638.0/65536.0,1,-nbitq), 
to_sfixed(136.0/65536.0,1,-nbitq), 
to_sfixed(-3253.0/65536.0,1,-nbitq), 
to_sfixed(2081.0/65536.0,1,-nbitq), 
to_sfixed(-2671.0/65536.0,1,-nbitq), 
to_sfixed(-820.0/65536.0,1,-nbitq), 
to_sfixed(-3608.0/65536.0,1,-nbitq), 
to_sfixed(2330.0/65536.0,1,-nbitq), 
to_sfixed(-3032.0/65536.0,1,-nbitq), 
to_sfixed(12365.0/65536.0,1,-nbitq), 
to_sfixed(58.0/65536.0,1,-nbitq), 
to_sfixed(-1250.0/65536.0,1,-nbitq), 
to_sfixed(-10715.0/65536.0,1,-nbitq), 
to_sfixed(-2442.0/65536.0,1,-nbitq), 
to_sfixed(-683.0/65536.0,1,-nbitq), 
to_sfixed(-3218.0/65536.0,1,-nbitq), 
to_sfixed(588.0/65536.0,1,-nbitq), 
to_sfixed(-2514.0/65536.0,1,-nbitq), 
to_sfixed(2323.0/65536.0,1,-nbitq), 
to_sfixed(-4724.0/65536.0,1,-nbitq), 
to_sfixed(-4405.0/65536.0,1,-nbitq), 
to_sfixed(1199.0/65536.0,1,-nbitq), 
to_sfixed(751.0/65536.0,1,-nbitq), 
to_sfixed(-1773.0/65536.0,1,-nbitq), 
to_sfixed(2967.0/65536.0,1,-nbitq), 
to_sfixed(1887.0/65536.0,1,-nbitq), 
to_sfixed(-7217.0/65536.0,1,-nbitq), 
to_sfixed(711.0/65536.0,1,-nbitq), 
to_sfixed(1481.0/65536.0,1,-nbitq), 
to_sfixed(1919.0/65536.0,1,-nbitq), 
to_sfixed(2135.0/65536.0,1,-nbitq), 
to_sfixed(-4144.0/65536.0,1,-nbitq), 
to_sfixed(-307.0/65536.0,1,-nbitq), 
to_sfixed(816.0/65536.0,1,-nbitq), 
to_sfixed(7208.0/65536.0,1,-nbitq), 
to_sfixed(-1141.0/65536.0,1,-nbitq), 
to_sfixed(-9861.0/65536.0,1,-nbitq), 
to_sfixed(1426.0/65536.0,1,-nbitq), 
to_sfixed(4226.0/65536.0,1,-nbitq), 
to_sfixed(7604.0/65536.0,1,-nbitq), 
to_sfixed(1660.0/65536.0,1,-nbitq), 
to_sfixed(1361.0/65536.0,1,-nbitq), 
to_sfixed(-3341.0/65536.0,1,-nbitq), 
to_sfixed(-6554.0/65536.0,1,-nbitq), 
to_sfixed(-15366.0/65536.0,1,-nbitq), 
to_sfixed(907.0/65536.0,1,-nbitq), 
to_sfixed(-5315.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1324.0/65536.0,1,-nbitq), 
to_sfixed(2437.0/65536.0,1,-nbitq), 
to_sfixed(-4414.0/65536.0,1,-nbitq), 
to_sfixed(-1492.0/65536.0,1,-nbitq), 
to_sfixed(5727.0/65536.0,1,-nbitq), 
to_sfixed(5072.0/65536.0,1,-nbitq), 
to_sfixed(-720.0/65536.0,1,-nbitq), 
to_sfixed(3403.0/65536.0,1,-nbitq), 
to_sfixed(1263.0/65536.0,1,-nbitq), 
to_sfixed(2749.0/65536.0,1,-nbitq), 
to_sfixed(3675.0/65536.0,1,-nbitq), 
to_sfixed(-6077.0/65536.0,1,-nbitq), 
to_sfixed(-3068.0/65536.0,1,-nbitq), 
to_sfixed(842.0/65536.0,1,-nbitq), 
to_sfixed(-496.0/65536.0,1,-nbitq), 
to_sfixed(2286.0/65536.0,1,-nbitq), 
to_sfixed(-1615.0/65536.0,1,-nbitq), 
to_sfixed(3775.0/65536.0,1,-nbitq), 
to_sfixed(1447.0/65536.0,1,-nbitq), 
to_sfixed(-1380.0/65536.0,1,-nbitq), 
to_sfixed(10258.0/65536.0,1,-nbitq), 
to_sfixed(-12139.0/65536.0,1,-nbitq), 
to_sfixed(-4926.0/65536.0,1,-nbitq), 
to_sfixed(7810.0/65536.0,1,-nbitq), 
to_sfixed(2486.0/65536.0,1,-nbitq), 
to_sfixed(4442.0/65536.0,1,-nbitq), 
to_sfixed(1256.0/65536.0,1,-nbitq), 
to_sfixed(3751.0/65536.0,1,-nbitq), 
to_sfixed(4841.0/65536.0,1,-nbitq), 
to_sfixed(-6412.0/65536.0,1,-nbitq), 
to_sfixed(-2859.0/65536.0,1,-nbitq), 
to_sfixed(-7673.0/65536.0,1,-nbitq), 
to_sfixed(2277.0/65536.0,1,-nbitq), 
to_sfixed(11022.0/65536.0,1,-nbitq), 
to_sfixed(-4110.0/65536.0,1,-nbitq), 
to_sfixed(1861.0/65536.0,1,-nbitq), 
to_sfixed(389.0/65536.0,1,-nbitq), 
to_sfixed(-3341.0/65536.0,1,-nbitq), 
to_sfixed(5635.0/65536.0,1,-nbitq), 
to_sfixed(373.0/65536.0,1,-nbitq), 
to_sfixed(3140.0/65536.0,1,-nbitq), 
to_sfixed(2183.0/65536.0,1,-nbitq), 
to_sfixed(7926.0/65536.0,1,-nbitq), 
to_sfixed(-1287.0/65536.0,1,-nbitq), 
to_sfixed(-69.0/65536.0,1,-nbitq), 
to_sfixed(-2129.0/65536.0,1,-nbitq), 
to_sfixed(-3772.0/65536.0,1,-nbitq), 
to_sfixed(-2419.0/65536.0,1,-nbitq), 
to_sfixed(-2814.0/65536.0,1,-nbitq), 
to_sfixed(128.0/65536.0,1,-nbitq), 
to_sfixed(2148.0/65536.0,1,-nbitq), 
to_sfixed(6545.0/65536.0,1,-nbitq), 
to_sfixed(-2804.0/65536.0,1,-nbitq), 
to_sfixed(-3490.0/65536.0,1,-nbitq), 
to_sfixed(3809.0/65536.0,1,-nbitq), 
to_sfixed(-2050.0/65536.0,1,-nbitq), 
to_sfixed(-3046.0/65536.0,1,-nbitq), 
to_sfixed(-809.0/65536.0,1,-nbitq), 
to_sfixed(2204.0/65536.0,1,-nbitq), 
to_sfixed(-3197.0/65536.0,1,-nbitq), 
to_sfixed(795.0/65536.0,1,-nbitq), 
to_sfixed(-2451.0/65536.0,1,-nbitq), 
to_sfixed(-1746.0/65536.0,1,-nbitq), 
to_sfixed(2744.0/65536.0,1,-nbitq), 
to_sfixed(-2426.0/65536.0,1,-nbitq), 
to_sfixed(-3692.0/65536.0,1,-nbitq), 
to_sfixed(-2251.0/65536.0,1,-nbitq), 
to_sfixed(1428.0/65536.0,1,-nbitq), 
to_sfixed(-2232.0/65536.0,1,-nbitq), 
to_sfixed(-5930.0/65536.0,1,-nbitq), 
to_sfixed(693.0/65536.0,1,-nbitq), 
to_sfixed(1697.0/65536.0,1,-nbitq), 
to_sfixed(4850.0/65536.0,1,-nbitq), 
to_sfixed(-1187.0/65536.0,1,-nbitq), 
to_sfixed(-2281.0/65536.0,1,-nbitq), 
to_sfixed(247.0/65536.0,1,-nbitq), 
to_sfixed(-3412.0/65536.0,1,-nbitq), 
to_sfixed(-7428.0/65536.0,1,-nbitq), 
to_sfixed(-846.0/65536.0,1,-nbitq), 
to_sfixed(-7648.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3666.0/65536.0,1,-nbitq), 
to_sfixed(7068.0/65536.0,1,-nbitq), 
to_sfixed(-4216.0/65536.0,1,-nbitq), 
to_sfixed(-5893.0/65536.0,1,-nbitq), 
to_sfixed(-6489.0/65536.0,1,-nbitq), 
to_sfixed(7127.0/65536.0,1,-nbitq), 
to_sfixed(-4448.0/65536.0,1,-nbitq), 
to_sfixed(6323.0/65536.0,1,-nbitq), 
to_sfixed(-2093.0/65536.0,1,-nbitq), 
to_sfixed(206.0/65536.0,1,-nbitq), 
to_sfixed(6596.0/65536.0,1,-nbitq), 
to_sfixed(-6004.0/65536.0,1,-nbitq), 
to_sfixed(1575.0/65536.0,1,-nbitq), 
to_sfixed(960.0/65536.0,1,-nbitq), 
to_sfixed(711.0/65536.0,1,-nbitq), 
to_sfixed(2642.0/65536.0,1,-nbitq), 
to_sfixed(1823.0/65536.0,1,-nbitq), 
to_sfixed(7572.0/65536.0,1,-nbitq), 
to_sfixed(1588.0/65536.0,1,-nbitq), 
to_sfixed(1856.0/65536.0,1,-nbitq), 
to_sfixed(8116.0/65536.0,1,-nbitq), 
to_sfixed(-11052.0/65536.0,1,-nbitq), 
to_sfixed(-6573.0/65536.0,1,-nbitq), 
to_sfixed(3895.0/65536.0,1,-nbitq), 
to_sfixed(-291.0/65536.0,1,-nbitq), 
to_sfixed(2425.0/65536.0,1,-nbitq), 
to_sfixed(4021.0/65536.0,1,-nbitq), 
to_sfixed(1904.0/65536.0,1,-nbitq), 
to_sfixed(3221.0/65536.0,1,-nbitq), 
to_sfixed(-570.0/65536.0,1,-nbitq), 
to_sfixed(1020.0/65536.0,1,-nbitq), 
to_sfixed(-3548.0/65536.0,1,-nbitq), 
to_sfixed(6924.0/65536.0,1,-nbitq), 
to_sfixed(6185.0/65536.0,1,-nbitq), 
to_sfixed(39.0/65536.0,1,-nbitq), 
to_sfixed(-2958.0/65536.0,1,-nbitq), 
to_sfixed(542.0/65536.0,1,-nbitq), 
to_sfixed(-1751.0/65536.0,1,-nbitq), 
to_sfixed(2917.0/65536.0,1,-nbitq), 
to_sfixed(-1787.0/65536.0,1,-nbitq), 
to_sfixed(2497.0/65536.0,1,-nbitq), 
to_sfixed(-821.0/65536.0,1,-nbitq), 
to_sfixed(12409.0/65536.0,1,-nbitq), 
to_sfixed(-819.0/65536.0,1,-nbitq), 
to_sfixed(461.0/65536.0,1,-nbitq), 
to_sfixed(-86.0/65536.0,1,-nbitq), 
to_sfixed(-623.0/65536.0,1,-nbitq), 
to_sfixed(-7455.0/65536.0,1,-nbitq), 
to_sfixed(-298.0/65536.0,1,-nbitq), 
to_sfixed(1371.0/65536.0,1,-nbitq), 
to_sfixed(2787.0/65536.0,1,-nbitq), 
to_sfixed(7017.0/65536.0,1,-nbitq), 
to_sfixed(5161.0/65536.0,1,-nbitq), 
to_sfixed(-1043.0/65536.0,1,-nbitq), 
to_sfixed(-4252.0/65536.0,1,-nbitq), 
to_sfixed(-657.0/65536.0,1,-nbitq), 
to_sfixed(394.0/65536.0,1,-nbitq), 
to_sfixed(648.0/65536.0,1,-nbitq), 
to_sfixed(1397.0/65536.0,1,-nbitq), 
to_sfixed(1175.0/65536.0,1,-nbitq), 
to_sfixed(-4763.0/65536.0,1,-nbitq), 
to_sfixed(-1448.0/65536.0,1,-nbitq), 
to_sfixed(552.0/65536.0,1,-nbitq), 
to_sfixed(1503.0/65536.0,1,-nbitq), 
to_sfixed(-3918.0/65536.0,1,-nbitq), 
to_sfixed(-869.0/65536.0,1,-nbitq), 
to_sfixed(2552.0/65536.0,1,-nbitq), 
to_sfixed(2083.0/65536.0,1,-nbitq), 
to_sfixed(-6921.0/65536.0,1,-nbitq), 
to_sfixed(-2482.0/65536.0,1,-nbitq), 
to_sfixed(3276.0/65536.0,1,-nbitq), 
to_sfixed(132.0/65536.0,1,-nbitq), 
to_sfixed(571.0/65536.0,1,-nbitq), 
to_sfixed(210.0/65536.0,1,-nbitq), 
to_sfixed(-1107.0/65536.0,1,-nbitq), 
to_sfixed(3444.0/65536.0,1,-nbitq), 
to_sfixed(1702.0/65536.0,1,-nbitq), 
to_sfixed(-4464.0/65536.0,1,-nbitq), 
to_sfixed(1532.0/65536.0,1,-nbitq), 
to_sfixed(-8558.0/65536.0,1,-nbitq)  ), 
( to_sfixed(9583.0/65536.0,1,-nbitq), 
to_sfixed(5297.0/65536.0,1,-nbitq), 
to_sfixed(-571.0/65536.0,1,-nbitq), 
to_sfixed(-5412.0/65536.0,1,-nbitq), 
to_sfixed(174.0/65536.0,1,-nbitq), 
to_sfixed(8394.0/65536.0,1,-nbitq), 
to_sfixed(-479.0/65536.0,1,-nbitq), 
to_sfixed(5305.0/65536.0,1,-nbitq), 
to_sfixed(-6021.0/65536.0,1,-nbitq), 
to_sfixed(-986.0/65536.0,1,-nbitq), 
to_sfixed(1275.0/65536.0,1,-nbitq), 
to_sfixed(-4649.0/65536.0,1,-nbitq), 
to_sfixed(-2003.0/65536.0,1,-nbitq), 
to_sfixed(2619.0/65536.0,1,-nbitq), 
to_sfixed(-18.0/65536.0,1,-nbitq), 
to_sfixed(-1196.0/65536.0,1,-nbitq), 
to_sfixed(-1890.0/65536.0,1,-nbitq), 
to_sfixed(6656.0/65536.0,1,-nbitq), 
to_sfixed(1381.0/65536.0,1,-nbitq), 
to_sfixed(2836.0/65536.0,1,-nbitq), 
to_sfixed(5461.0/65536.0,1,-nbitq), 
to_sfixed(-5859.0/65536.0,1,-nbitq), 
to_sfixed(-5967.0/65536.0,1,-nbitq), 
to_sfixed(1249.0/65536.0,1,-nbitq), 
to_sfixed(-2867.0/65536.0,1,-nbitq), 
to_sfixed(2539.0/65536.0,1,-nbitq), 
to_sfixed(3982.0/65536.0,1,-nbitq), 
to_sfixed(-1166.0/65536.0,1,-nbitq), 
to_sfixed(3150.0/65536.0,1,-nbitq), 
to_sfixed(863.0/65536.0,1,-nbitq), 
to_sfixed(-3558.0/65536.0,1,-nbitq), 
to_sfixed(-4902.0/65536.0,1,-nbitq), 
to_sfixed(10677.0/65536.0,1,-nbitq), 
to_sfixed(-128.0/65536.0,1,-nbitq), 
to_sfixed(-372.0/65536.0,1,-nbitq), 
to_sfixed(-2290.0/65536.0,1,-nbitq), 
to_sfixed(2651.0/65536.0,1,-nbitq), 
to_sfixed(1836.0/65536.0,1,-nbitq), 
to_sfixed(2960.0/65536.0,1,-nbitq), 
to_sfixed(-1652.0/65536.0,1,-nbitq), 
to_sfixed(5112.0/65536.0,1,-nbitq), 
to_sfixed(-1591.0/65536.0,1,-nbitq), 
to_sfixed(9380.0/65536.0,1,-nbitq), 
to_sfixed(3024.0/65536.0,1,-nbitq), 
to_sfixed(1758.0/65536.0,1,-nbitq), 
to_sfixed(-5929.0/65536.0,1,-nbitq), 
to_sfixed(-2826.0/65536.0,1,-nbitq), 
to_sfixed(-3656.0/65536.0,1,-nbitq), 
to_sfixed(-158.0/65536.0,1,-nbitq), 
to_sfixed(-1246.0/65536.0,1,-nbitq), 
to_sfixed(691.0/65536.0,1,-nbitq), 
to_sfixed(5981.0/65536.0,1,-nbitq), 
to_sfixed(5606.0/65536.0,1,-nbitq), 
to_sfixed(-664.0/65536.0,1,-nbitq), 
to_sfixed(-489.0/65536.0,1,-nbitq), 
to_sfixed(-542.0/65536.0,1,-nbitq), 
to_sfixed(-805.0/65536.0,1,-nbitq), 
to_sfixed(3467.0/65536.0,1,-nbitq), 
to_sfixed(-1146.0/65536.0,1,-nbitq), 
to_sfixed(3751.0/65536.0,1,-nbitq), 
to_sfixed(-4710.0/65536.0,1,-nbitq), 
to_sfixed(2449.0/65536.0,1,-nbitq), 
to_sfixed(459.0/65536.0,1,-nbitq), 
to_sfixed(1828.0/65536.0,1,-nbitq), 
to_sfixed(-2416.0/65536.0,1,-nbitq), 
to_sfixed(1850.0/65536.0,1,-nbitq), 
to_sfixed(3280.0/65536.0,1,-nbitq), 
to_sfixed(1506.0/65536.0,1,-nbitq), 
to_sfixed(-4670.0/65536.0,1,-nbitq), 
to_sfixed(-3138.0/65536.0,1,-nbitq), 
to_sfixed(5723.0/65536.0,1,-nbitq), 
to_sfixed(182.0/65536.0,1,-nbitq), 
to_sfixed(651.0/65536.0,1,-nbitq), 
to_sfixed(689.0/65536.0,1,-nbitq), 
to_sfixed(-388.0/65536.0,1,-nbitq), 
to_sfixed(6776.0/65536.0,1,-nbitq), 
to_sfixed(-1619.0/65536.0,1,-nbitq), 
to_sfixed(-2155.0/65536.0,1,-nbitq), 
to_sfixed(-406.0/65536.0,1,-nbitq), 
to_sfixed(-8851.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3937.0/65536.0,1,-nbitq), 
to_sfixed(-2475.0/65536.0,1,-nbitq), 
to_sfixed(1333.0/65536.0,1,-nbitq), 
to_sfixed(583.0/65536.0,1,-nbitq), 
to_sfixed(1598.0/65536.0,1,-nbitq), 
to_sfixed(4691.0/65536.0,1,-nbitq), 
to_sfixed(1265.0/65536.0,1,-nbitq), 
to_sfixed(2444.0/65536.0,1,-nbitq), 
to_sfixed(-2061.0/65536.0,1,-nbitq), 
to_sfixed(-1734.0/65536.0,1,-nbitq), 
to_sfixed(3243.0/65536.0,1,-nbitq), 
to_sfixed(-5112.0/65536.0,1,-nbitq), 
to_sfixed(2758.0/65536.0,1,-nbitq), 
to_sfixed(4559.0/65536.0,1,-nbitq), 
to_sfixed(2360.0/65536.0,1,-nbitq), 
to_sfixed(2103.0/65536.0,1,-nbitq), 
to_sfixed(-3304.0/65536.0,1,-nbitq), 
to_sfixed(1462.0/65536.0,1,-nbitq), 
to_sfixed(-2046.0/65536.0,1,-nbitq), 
to_sfixed(-1951.0/65536.0,1,-nbitq), 
to_sfixed(5790.0/65536.0,1,-nbitq), 
to_sfixed(-152.0/65536.0,1,-nbitq), 
to_sfixed(-6308.0/65536.0,1,-nbitq), 
to_sfixed(1606.0/65536.0,1,-nbitq), 
to_sfixed(782.0/65536.0,1,-nbitq), 
to_sfixed(4937.0/65536.0,1,-nbitq), 
to_sfixed(2388.0/65536.0,1,-nbitq), 
to_sfixed(-2171.0/65536.0,1,-nbitq), 
to_sfixed(3117.0/65536.0,1,-nbitq), 
to_sfixed(-1846.0/65536.0,1,-nbitq), 
to_sfixed(857.0/65536.0,1,-nbitq), 
to_sfixed(-2398.0/65536.0,1,-nbitq), 
to_sfixed(9201.0/65536.0,1,-nbitq), 
to_sfixed(-2046.0/65536.0,1,-nbitq), 
to_sfixed(-1978.0/65536.0,1,-nbitq), 
to_sfixed(1950.0/65536.0,1,-nbitq), 
to_sfixed(3512.0/65536.0,1,-nbitq), 
to_sfixed(2148.0/65536.0,1,-nbitq), 
to_sfixed(-2231.0/65536.0,1,-nbitq), 
to_sfixed(1127.0/65536.0,1,-nbitq), 
to_sfixed(1316.0/65536.0,1,-nbitq), 
to_sfixed(74.0/65536.0,1,-nbitq), 
to_sfixed(9838.0/65536.0,1,-nbitq), 
to_sfixed(1627.0/65536.0,1,-nbitq), 
to_sfixed(700.0/65536.0,1,-nbitq), 
to_sfixed(-6100.0/65536.0,1,-nbitq), 
to_sfixed(1924.0/65536.0,1,-nbitq), 
to_sfixed(-1901.0/65536.0,1,-nbitq), 
to_sfixed(-2302.0/65536.0,1,-nbitq), 
to_sfixed(2354.0/65536.0,1,-nbitq), 
to_sfixed(-1596.0/65536.0,1,-nbitq), 
to_sfixed(4286.0/65536.0,1,-nbitq), 
to_sfixed(9339.0/65536.0,1,-nbitq), 
to_sfixed(-1575.0/65536.0,1,-nbitq), 
to_sfixed(-717.0/65536.0,1,-nbitq), 
to_sfixed(6430.0/65536.0,1,-nbitq), 
to_sfixed(1286.0/65536.0,1,-nbitq), 
to_sfixed(540.0/65536.0,1,-nbitq), 
to_sfixed(751.0/65536.0,1,-nbitq), 
to_sfixed(2020.0/65536.0,1,-nbitq), 
to_sfixed(1868.0/65536.0,1,-nbitq), 
to_sfixed(2577.0/65536.0,1,-nbitq), 
to_sfixed(666.0/65536.0,1,-nbitq), 
to_sfixed(-1261.0/65536.0,1,-nbitq), 
to_sfixed(920.0/65536.0,1,-nbitq), 
to_sfixed(6775.0/65536.0,1,-nbitq), 
to_sfixed(6002.0/65536.0,1,-nbitq), 
to_sfixed(6252.0/65536.0,1,-nbitq), 
to_sfixed(-8233.0/65536.0,1,-nbitq), 
to_sfixed(-8443.0/65536.0,1,-nbitq), 
to_sfixed(2653.0/65536.0,1,-nbitq), 
to_sfixed(-651.0/65536.0,1,-nbitq), 
to_sfixed(2273.0/65536.0,1,-nbitq), 
to_sfixed(-567.0/65536.0,1,-nbitq), 
to_sfixed(1318.0/65536.0,1,-nbitq), 
to_sfixed(2249.0/65536.0,1,-nbitq), 
to_sfixed(-1207.0/65536.0,1,-nbitq), 
to_sfixed(1832.0/65536.0,1,-nbitq), 
to_sfixed(1554.0/65536.0,1,-nbitq), 
to_sfixed(-7009.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2216.0/65536.0,1,-nbitq), 
to_sfixed(-2313.0/65536.0,1,-nbitq), 
to_sfixed(-3117.0/65536.0,1,-nbitq), 
to_sfixed(428.0/65536.0,1,-nbitq), 
to_sfixed(1184.0/65536.0,1,-nbitq), 
to_sfixed(2440.0/65536.0,1,-nbitq), 
to_sfixed(100.0/65536.0,1,-nbitq), 
to_sfixed(6203.0/65536.0,1,-nbitq), 
to_sfixed(-3697.0/65536.0,1,-nbitq), 
to_sfixed(1241.0/65536.0,1,-nbitq), 
to_sfixed(3820.0/65536.0,1,-nbitq), 
to_sfixed(1498.0/65536.0,1,-nbitq), 
to_sfixed(2815.0/65536.0,1,-nbitq), 
to_sfixed(3390.0/65536.0,1,-nbitq), 
to_sfixed(1304.0/65536.0,1,-nbitq), 
to_sfixed(-2044.0/65536.0,1,-nbitq), 
to_sfixed(-1275.0/65536.0,1,-nbitq), 
to_sfixed(4415.0/65536.0,1,-nbitq), 
to_sfixed(-3256.0/65536.0,1,-nbitq), 
to_sfixed(-2330.0/65536.0,1,-nbitq), 
to_sfixed(5637.0/65536.0,1,-nbitq), 
to_sfixed(-2334.0/65536.0,1,-nbitq), 
to_sfixed(-3532.0/65536.0,1,-nbitq), 
to_sfixed(817.0/65536.0,1,-nbitq), 
to_sfixed(-203.0/65536.0,1,-nbitq), 
to_sfixed(2257.0/65536.0,1,-nbitq), 
to_sfixed(2738.0/65536.0,1,-nbitq), 
to_sfixed(1440.0/65536.0,1,-nbitq), 
to_sfixed(79.0/65536.0,1,-nbitq), 
to_sfixed(-2523.0/65536.0,1,-nbitq), 
to_sfixed(1994.0/65536.0,1,-nbitq), 
to_sfixed(-246.0/65536.0,1,-nbitq), 
to_sfixed(6540.0/65536.0,1,-nbitq), 
to_sfixed(-1729.0/65536.0,1,-nbitq), 
to_sfixed(1490.0/65536.0,1,-nbitq), 
to_sfixed(-2812.0/65536.0,1,-nbitq), 
to_sfixed(-224.0/65536.0,1,-nbitq), 
to_sfixed(5812.0/65536.0,1,-nbitq), 
to_sfixed(731.0/65536.0,1,-nbitq), 
to_sfixed(-1102.0/65536.0,1,-nbitq), 
to_sfixed(1565.0/65536.0,1,-nbitq), 
to_sfixed(172.0/65536.0,1,-nbitq), 
to_sfixed(8398.0/65536.0,1,-nbitq), 
to_sfixed(5304.0/65536.0,1,-nbitq), 
to_sfixed(-1702.0/65536.0,1,-nbitq), 
to_sfixed(-4820.0/65536.0,1,-nbitq), 
to_sfixed(-3149.0/65536.0,1,-nbitq), 
to_sfixed(-1396.0/65536.0,1,-nbitq), 
to_sfixed(1944.0/65536.0,1,-nbitq), 
to_sfixed(1573.0/65536.0,1,-nbitq), 
to_sfixed(-1014.0/65536.0,1,-nbitq), 
to_sfixed(761.0/65536.0,1,-nbitq), 
to_sfixed(7265.0/65536.0,1,-nbitq), 
to_sfixed(4569.0/65536.0,1,-nbitq), 
to_sfixed(-1869.0/65536.0,1,-nbitq), 
to_sfixed(3136.0/65536.0,1,-nbitq), 
to_sfixed(44.0/65536.0,1,-nbitq), 
to_sfixed(3871.0/65536.0,1,-nbitq), 
to_sfixed(2761.0/65536.0,1,-nbitq), 
to_sfixed(2045.0/65536.0,1,-nbitq), 
to_sfixed(-2494.0/65536.0,1,-nbitq), 
to_sfixed(-13.0/65536.0,1,-nbitq), 
to_sfixed(1140.0/65536.0,1,-nbitq), 
to_sfixed(-2415.0/65536.0,1,-nbitq), 
to_sfixed(-4019.0/65536.0,1,-nbitq), 
to_sfixed(-182.0/65536.0,1,-nbitq), 
to_sfixed(1055.0/65536.0,1,-nbitq), 
to_sfixed(4923.0/65536.0,1,-nbitq), 
to_sfixed(-7341.0/65536.0,1,-nbitq), 
to_sfixed(-5203.0/65536.0,1,-nbitq), 
to_sfixed(5713.0/65536.0,1,-nbitq), 
to_sfixed(-631.0/65536.0,1,-nbitq), 
to_sfixed(4480.0/65536.0,1,-nbitq), 
to_sfixed(-2381.0/65536.0,1,-nbitq), 
to_sfixed(805.0/65536.0,1,-nbitq), 
to_sfixed(2091.0/65536.0,1,-nbitq), 
to_sfixed(-1439.0/65536.0,1,-nbitq), 
to_sfixed(1131.0/65536.0,1,-nbitq), 
to_sfixed(-2908.0/65536.0,1,-nbitq), 
to_sfixed(-4463.0/65536.0,1,-nbitq)  ), 
( to_sfixed(719.0/65536.0,1,-nbitq), 
to_sfixed(-2326.0/65536.0,1,-nbitq), 
to_sfixed(-2956.0/65536.0,1,-nbitq), 
to_sfixed(-2012.0/65536.0,1,-nbitq), 
to_sfixed(-2326.0/65536.0,1,-nbitq), 
to_sfixed(-279.0/65536.0,1,-nbitq), 
to_sfixed(449.0/65536.0,1,-nbitq), 
to_sfixed(2125.0/65536.0,1,-nbitq), 
to_sfixed(851.0/65536.0,1,-nbitq), 
to_sfixed(2402.0/65536.0,1,-nbitq), 
to_sfixed(577.0/65536.0,1,-nbitq), 
to_sfixed(1608.0/65536.0,1,-nbitq), 
to_sfixed(785.0/65536.0,1,-nbitq), 
to_sfixed(469.0/65536.0,1,-nbitq), 
to_sfixed(-1249.0/65536.0,1,-nbitq), 
to_sfixed(-2312.0/65536.0,1,-nbitq), 
to_sfixed(-1845.0/65536.0,1,-nbitq), 
to_sfixed(-932.0/65536.0,1,-nbitq), 
to_sfixed(-2452.0/65536.0,1,-nbitq), 
to_sfixed(-2162.0/65536.0,1,-nbitq), 
to_sfixed(2787.0/65536.0,1,-nbitq), 
to_sfixed(4227.0/65536.0,1,-nbitq), 
to_sfixed(-3708.0/65536.0,1,-nbitq), 
to_sfixed(455.0/65536.0,1,-nbitq), 
to_sfixed(1076.0/65536.0,1,-nbitq), 
to_sfixed(1953.0/65536.0,1,-nbitq), 
to_sfixed(-1380.0/65536.0,1,-nbitq), 
to_sfixed(-1369.0/65536.0,1,-nbitq), 
to_sfixed(-1257.0/65536.0,1,-nbitq), 
to_sfixed(1630.0/65536.0,1,-nbitq), 
to_sfixed(-1119.0/65536.0,1,-nbitq), 
to_sfixed(887.0/65536.0,1,-nbitq), 
to_sfixed(1945.0/65536.0,1,-nbitq), 
to_sfixed(3117.0/65536.0,1,-nbitq), 
to_sfixed(1841.0/65536.0,1,-nbitq), 
to_sfixed(-321.0/65536.0,1,-nbitq), 
to_sfixed(-407.0/65536.0,1,-nbitq), 
to_sfixed(1211.0/65536.0,1,-nbitq), 
to_sfixed(-3807.0/65536.0,1,-nbitq), 
to_sfixed(2589.0/65536.0,1,-nbitq), 
to_sfixed(-2584.0/65536.0,1,-nbitq), 
to_sfixed(1114.0/65536.0,1,-nbitq), 
to_sfixed(1035.0/65536.0,1,-nbitq), 
to_sfixed(4010.0/65536.0,1,-nbitq), 
to_sfixed(1994.0/65536.0,1,-nbitq), 
to_sfixed(1009.0/65536.0,1,-nbitq), 
to_sfixed(-1906.0/65536.0,1,-nbitq), 
to_sfixed(-1937.0/65536.0,1,-nbitq), 
to_sfixed(-2989.0/65536.0,1,-nbitq), 
to_sfixed(1555.0/65536.0,1,-nbitq), 
to_sfixed(1167.0/65536.0,1,-nbitq), 
to_sfixed(-232.0/65536.0,1,-nbitq), 
to_sfixed(3431.0/65536.0,1,-nbitq), 
to_sfixed(2301.0/65536.0,1,-nbitq), 
to_sfixed(2408.0/65536.0,1,-nbitq), 
to_sfixed(1581.0/65536.0,1,-nbitq), 
to_sfixed(1400.0/65536.0,1,-nbitq), 
to_sfixed(-1229.0/65536.0,1,-nbitq), 
to_sfixed(974.0/65536.0,1,-nbitq), 
to_sfixed(1997.0/65536.0,1,-nbitq), 
to_sfixed(-3358.0/65536.0,1,-nbitq), 
to_sfixed(1377.0/65536.0,1,-nbitq), 
to_sfixed(69.0/65536.0,1,-nbitq), 
to_sfixed(-2380.0/65536.0,1,-nbitq), 
to_sfixed(-415.0/65536.0,1,-nbitq), 
to_sfixed(3312.0/65536.0,1,-nbitq), 
to_sfixed(-69.0/65536.0,1,-nbitq), 
to_sfixed(-989.0/65536.0,1,-nbitq), 
to_sfixed(-5580.0/65536.0,1,-nbitq), 
to_sfixed(289.0/65536.0,1,-nbitq), 
to_sfixed(1112.0/65536.0,1,-nbitq), 
to_sfixed(252.0/65536.0,1,-nbitq), 
to_sfixed(-310.0/65536.0,1,-nbitq), 
to_sfixed(-272.0/65536.0,1,-nbitq), 
to_sfixed(2486.0/65536.0,1,-nbitq), 
to_sfixed(1845.0/65536.0,1,-nbitq), 
to_sfixed(-968.0/65536.0,1,-nbitq), 
to_sfixed(2042.0/65536.0,1,-nbitq), 
to_sfixed(-924.0/65536.0,1,-nbitq), 
to_sfixed(-6233.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1199.0/65536.0,1,-nbitq), 
to_sfixed(-873.0/65536.0,1,-nbitq), 
to_sfixed(1849.0/65536.0,1,-nbitq), 
to_sfixed(-486.0/65536.0,1,-nbitq), 
to_sfixed(-2400.0/65536.0,1,-nbitq), 
to_sfixed(-1657.0/65536.0,1,-nbitq), 
to_sfixed(-2441.0/65536.0,1,-nbitq), 
to_sfixed(227.0/65536.0,1,-nbitq), 
to_sfixed(-652.0/65536.0,1,-nbitq), 
to_sfixed(-1190.0/65536.0,1,-nbitq), 
to_sfixed(-3.0/65536.0,1,-nbitq), 
to_sfixed(947.0/65536.0,1,-nbitq), 
to_sfixed(1653.0/65536.0,1,-nbitq), 
to_sfixed(-2200.0/65536.0,1,-nbitq), 
to_sfixed(-143.0/65536.0,1,-nbitq), 
to_sfixed(-1230.0/65536.0,1,-nbitq), 
to_sfixed(761.0/65536.0,1,-nbitq), 
to_sfixed(4532.0/65536.0,1,-nbitq), 
to_sfixed(1604.0/65536.0,1,-nbitq), 
to_sfixed(-165.0/65536.0,1,-nbitq), 
to_sfixed(-1546.0/65536.0,1,-nbitq), 
to_sfixed(859.0/65536.0,1,-nbitq), 
to_sfixed(984.0/65536.0,1,-nbitq), 
to_sfixed(3121.0/65536.0,1,-nbitq), 
to_sfixed(774.0/65536.0,1,-nbitq), 
to_sfixed(1931.0/65536.0,1,-nbitq), 
to_sfixed(-2712.0/65536.0,1,-nbitq), 
to_sfixed(-1450.0/65536.0,1,-nbitq), 
to_sfixed(-3105.0/65536.0,1,-nbitq), 
to_sfixed(-3498.0/65536.0,1,-nbitq), 
to_sfixed(-1914.0/65536.0,1,-nbitq), 
to_sfixed(1681.0/65536.0,1,-nbitq), 
to_sfixed(282.0/65536.0,1,-nbitq), 
to_sfixed(-2294.0/65536.0,1,-nbitq), 
to_sfixed(-1351.0/65536.0,1,-nbitq), 
to_sfixed(-2239.0/65536.0,1,-nbitq), 
to_sfixed(1295.0/65536.0,1,-nbitq), 
to_sfixed(410.0/65536.0,1,-nbitq), 
to_sfixed(-4256.0/65536.0,1,-nbitq), 
to_sfixed(2778.0/65536.0,1,-nbitq), 
to_sfixed(1987.0/65536.0,1,-nbitq), 
to_sfixed(-1658.0/65536.0,1,-nbitq), 
to_sfixed(949.0/65536.0,1,-nbitq), 
to_sfixed(3741.0/65536.0,1,-nbitq), 
to_sfixed(1119.0/65536.0,1,-nbitq), 
to_sfixed(2315.0/65536.0,1,-nbitq), 
to_sfixed(751.0/65536.0,1,-nbitq), 
to_sfixed(-1879.0/65536.0,1,-nbitq), 
to_sfixed(490.0/65536.0,1,-nbitq), 
to_sfixed(722.0/65536.0,1,-nbitq), 
to_sfixed(709.0/65536.0,1,-nbitq), 
to_sfixed(849.0/65536.0,1,-nbitq), 
to_sfixed(-16.0/65536.0,1,-nbitq), 
to_sfixed(-1712.0/65536.0,1,-nbitq), 
to_sfixed(2529.0/65536.0,1,-nbitq), 
to_sfixed(-88.0/65536.0,1,-nbitq), 
to_sfixed(141.0/65536.0,1,-nbitq), 
to_sfixed(1002.0/65536.0,1,-nbitq), 
to_sfixed(938.0/65536.0,1,-nbitq), 
to_sfixed(4366.0/65536.0,1,-nbitq), 
to_sfixed(-4276.0/65536.0,1,-nbitq), 
to_sfixed(-132.0/65536.0,1,-nbitq), 
to_sfixed(762.0/65536.0,1,-nbitq), 
to_sfixed(1053.0/65536.0,1,-nbitq), 
to_sfixed(-2338.0/65536.0,1,-nbitq), 
to_sfixed(680.0/65536.0,1,-nbitq), 
to_sfixed(1505.0/65536.0,1,-nbitq), 
to_sfixed(-2947.0/65536.0,1,-nbitq), 
to_sfixed(491.0/65536.0,1,-nbitq), 
to_sfixed(-105.0/65536.0,1,-nbitq), 
to_sfixed(3076.0/65536.0,1,-nbitq), 
to_sfixed(-143.0/65536.0,1,-nbitq), 
to_sfixed(409.0/65536.0,1,-nbitq), 
to_sfixed(-1121.0/65536.0,1,-nbitq), 
to_sfixed(-2947.0/65536.0,1,-nbitq), 
to_sfixed(-1689.0/65536.0,1,-nbitq), 
to_sfixed(-1207.0/65536.0,1,-nbitq), 
to_sfixed(700.0/65536.0,1,-nbitq), 
to_sfixed(-2221.0/65536.0,1,-nbitq), 
to_sfixed(462.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2158.0/65536.0,1,-nbitq), 
to_sfixed(80.0/65536.0,1,-nbitq), 
to_sfixed(558.0/65536.0,1,-nbitq), 
to_sfixed(-761.0/65536.0,1,-nbitq), 
to_sfixed(-539.0/65536.0,1,-nbitq), 
to_sfixed(-2391.0/65536.0,1,-nbitq), 
to_sfixed(-3185.0/65536.0,1,-nbitq), 
to_sfixed(107.0/65536.0,1,-nbitq), 
to_sfixed(692.0/65536.0,1,-nbitq), 
to_sfixed(1342.0/65536.0,1,-nbitq), 
to_sfixed(-319.0/65536.0,1,-nbitq), 
to_sfixed(-172.0/65536.0,1,-nbitq), 
to_sfixed(-1897.0/65536.0,1,-nbitq), 
to_sfixed(-884.0/65536.0,1,-nbitq), 
to_sfixed(-828.0/65536.0,1,-nbitq), 
to_sfixed(-1293.0/65536.0,1,-nbitq), 
to_sfixed(-46.0/65536.0,1,-nbitq), 
to_sfixed(497.0/65536.0,1,-nbitq), 
to_sfixed(1720.0/65536.0,1,-nbitq), 
to_sfixed(2090.0/65536.0,1,-nbitq), 
to_sfixed(-2627.0/65536.0,1,-nbitq), 
to_sfixed(-314.0/65536.0,1,-nbitq), 
to_sfixed(-1511.0/65536.0,1,-nbitq), 
to_sfixed(1448.0/65536.0,1,-nbitq), 
to_sfixed(420.0/65536.0,1,-nbitq), 
to_sfixed(3604.0/65536.0,1,-nbitq), 
to_sfixed(1261.0/65536.0,1,-nbitq), 
to_sfixed(1528.0/65536.0,1,-nbitq), 
to_sfixed(-763.0/65536.0,1,-nbitq), 
to_sfixed(-2116.0/65536.0,1,-nbitq), 
to_sfixed(2266.0/65536.0,1,-nbitq), 
to_sfixed(1171.0/65536.0,1,-nbitq), 
to_sfixed(798.0/65536.0,1,-nbitq), 
to_sfixed(-3691.0/65536.0,1,-nbitq), 
to_sfixed(1748.0/65536.0,1,-nbitq), 
to_sfixed(961.0/65536.0,1,-nbitq), 
to_sfixed(626.0/65536.0,1,-nbitq), 
to_sfixed(417.0/65536.0,1,-nbitq), 
to_sfixed(-1315.0/65536.0,1,-nbitq), 
to_sfixed(-2857.0/65536.0,1,-nbitq), 
to_sfixed(-1188.0/65536.0,1,-nbitq), 
to_sfixed(880.0/65536.0,1,-nbitq), 
to_sfixed(128.0/65536.0,1,-nbitq), 
to_sfixed(408.0/65536.0,1,-nbitq), 
to_sfixed(-2144.0/65536.0,1,-nbitq), 
to_sfixed(3998.0/65536.0,1,-nbitq), 
to_sfixed(1425.0/65536.0,1,-nbitq), 
to_sfixed(3125.0/65536.0,1,-nbitq), 
to_sfixed(-1683.0/65536.0,1,-nbitq), 
to_sfixed(4292.0/65536.0,1,-nbitq), 
to_sfixed(1739.0/65536.0,1,-nbitq), 
to_sfixed(-1707.0/65536.0,1,-nbitq), 
to_sfixed(570.0/65536.0,1,-nbitq), 
to_sfixed(441.0/65536.0,1,-nbitq), 
to_sfixed(432.0/65536.0,1,-nbitq), 
to_sfixed(1679.0/65536.0,1,-nbitq), 
to_sfixed(2785.0/65536.0,1,-nbitq), 
to_sfixed(2240.0/65536.0,1,-nbitq), 
to_sfixed(2883.0/65536.0,1,-nbitq), 
to_sfixed(1657.0/65536.0,1,-nbitq), 
to_sfixed(-3307.0/65536.0,1,-nbitq), 
to_sfixed(-858.0/65536.0,1,-nbitq), 
to_sfixed(-2397.0/65536.0,1,-nbitq), 
to_sfixed(-327.0/65536.0,1,-nbitq), 
to_sfixed(-2549.0/65536.0,1,-nbitq), 
to_sfixed(3561.0/65536.0,1,-nbitq), 
to_sfixed(1.0/65536.0,1,-nbitq), 
to_sfixed(-2906.0/65536.0,1,-nbitq), 
to_sfixed(325.0/65536.0,1,-nbitq), 
to_sfixed(-1439.0/65536.0,1,-nbitq), 
to_sfixed(1965.0/65536.0,1,-nbitq), 
to_sfixed(-2239.0/65536.0,1,-nbitq), 
to_sfixed(-92.0/65536.0,1,-nbitq), 
to_sfixed(-1030.0/65536.0,1,-nbitq), 
to_sfixed(-1027.0/65536.0,1,-nbitq), 
to_sfixed(2307.0/65536.0,1,-nbitq), 
to_sfixed(-1164.0/65536.0,1,-nbitq), 
to_sfixed(2322.0/65536.0,1,-nbitq), 
to_sfixed(2480.0/65536.0,1,-nbitq), 
to_sfixed(1282.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1338.0/65536.0,1,-nbitq), 
to_sfixed(-210.0/65536.0,1,-nbitq), 
to_sfixed(2765.0/65536.0,1,-nbitq), 
to_sfixed(2906.0/65536.0,1,-nbitq), 
to_sfixed(-1146.0/65536.0,1,-nbitq), 
to_sfixed(-399.0/65536.0,1,-nbitq), 
to_sfixed(1121.0/65536.0,1,-nbitq), 
to_sfixed(-738.0/65536.0,1,-nbitq), 
to_sfixed(280.0/65536.0,1,-nbitq), 
to_sfixed(-1838.0/65536.0,1,-nbitq), 
to_sfixed(-2177.0/65536.0,1,-nbitq), 
to_sfixed(-1134.0/65536.0,1,-nbitq), 
to_sfixed(289.0/65536.0,1,-nbitq), 
to_sfixed(-2679.0/65536.0,1,-nbitq), 
to_sfixed(153.0/65536.0,1,-nbitq), 
to_sfixed(1394.0/65536.0,1,-nbitq), 
to_sfixed(-1814.0/65536.0,1,-nbitq), 
to_sfixed(-1250.0/65536.0,1,-nbitq), 
to_sfixed(-2691.0/65536.0,1,-nbitq), 
to_sfixed(-1092.0/65536.0,1,-nbitq), 
to_sfixed(679.0/65536.0,1,-nbitq), 
to_sfixed(3008.0/65536.0,1,-nbitq), 
to_sfixed(-1067.0/65536.0,1,-nbitq), 
to_sfixed(1037.0/65536.0,1,-nbitq), 
to_sfixed(606.0/65536.0,1,-nbitq), 
to_sfixed(3229.0/65536.0,1,-nbitq), 
to_sfixed(371.0/65536.0,1,-nbitq), 
to_sfixed(736.0/65536.0,1,-nbitq), 
to_sfixed(1428.0/65536.0,1,-nbitq), 
to_sfixed(-1078.0/65536.0,1,-nbitq), 
to_sfixed(-2806.0/65536.0,1,-nbitq), 
to_sfixed(727.0/65536.0,1,-nbitq), 
to_sfixed(-569.0/65536.0,1,-nbitq), 
to_sfixed(679.0/65536.0,1,-nbitq), 
to_sfixed(-3181.0/65536.0,1,-nbitq), 
to_sfixed(2578.0/65536.0,1,-nbitq), 
to_sfixed(1328.0/65536.0,1,-nbitq), 
to_sfixed(471.0/65536.0,1,-nbitq), 
to_sfixed(63.0/65536.0,1,-nbitq), 
to_sfixed(-1992.0/65536.0,1,-nbitq), 
to_sfixed(-2140.0/65536.0,1,-nbitq), 
to_sfixed(2368.0/65536.0,1,-nbitq), 
to_sfixed(-3057.0/65536.0,1,-nbitq), 
to_sfixed(2798.0/65536.0,1,-nbitq), 
to_sfixed(305.0/65536.0,1,-nbitq), 
to_sfixed(594.0/65536.0,1,-nbitq), 
to_sfixed(143.0/65536.0,1,-nbitq), 
to_sfixed(1730.0/65536.0,1,-nbitq), 
to_sfixed(1124.0/65536.0,1,-nbitq), 
to_sfixed(2692.0/65536.0,1,-nbitq), 
to_sfixed(2543.0/65536.0,1,-nbitq), 
to_sfixed(-474.0/65536.0,1,-nbitq), 
to_sfixed(-872.0/65536.0,1,-nbitq), 
to_sfixed(2202.0/65536.0,1,-nbitq), 
to_sfixed(1139.0/65536.0,1,-nbitq), 
to_sfixed(2171.0/65536.0,1,-nbitq), 
to_sfixed(1598.0/65536.0,1,-nbitq), 
to_sfixed(-58.0/65536.0,1,-nbitq), 
to_sfixed(2688.0/65536.0,1,-nbitq), 
to_sfixed(687.0/65536.0,1,-nbitq), 
to_sfixed(-3451.0/65536.0,1,-nbitq), 
to_sfixed(1220.0/65536.0,1,-nbitq), 
to_sfixed(-2298.0/65536.0,1,-nbitq), 
to_sfixed(398.0/65536.0,1,-nbitq), 
to_sfixed(-120.0/65536.0,1,-nbitq), 
to_sfixed(911.0/65536.0,1,-nbitq), 
to_sfixed(-499.0/65536.0,1,-nbitq), 
to_sfixed(-374.0/65536.0,1,-nbitq), 
to_sfixed(1517.0/65536.0,1,-nbitq), 
to_sfixed(-1391.0/65536.0,1,-nbitq), 
to_sfixed(64.0/65536.0,1,-nbitq), 
to_sfixed(-3521.0/65536.0,1,-nbitq), 
to_sfixed(-996.0/65536.0,1,-nbitq), 
to_sfixed(-1266.0/65536.0,1,-nbitq), 
to_sfixed(-2627.0/65536.0,1,-nbitq), 
to_sfixed(3914.0/65536.0,1,-nbitq), 
to_sfixed(542.0/65536.0,1,-nbitq), 
to_sfixed(2835.0/65536.0,1,-nbitq), 
to_sfixed(-2176.0/65536.0,1,-nbitq), 
to_sfixed(2319.0/65536.0,1,-nbitq)  ), 
( to_sfixed(379.0/65536.0,1,-nbitq), 
to_sfixed(-870.0/65536.0,1,-nbitq), 
to_sfixed(-501.0/65536.0,1,-nbitq), 
to_sfixed(-603.0/65536.0,1,-nbitq), 
to_sfixed(-2116.0/65536.0,1,-nbitq), 
to_sfixed(-4485.0/65536.0,1,-nbitq), 
to_sfixed(-2757.0/65536.0,1,-nbitq), 
to_sfixed(-2497.0/65536.0,1,-nbitq), 
to_sfixed(-777.0/65536.0,1,-nbitq), 
to_sfixed(322.0/65536.0,1,-nbitq), 
to_sfixed(1141.0/65536.0,1,-nbitq), 
to_sfixed(-1823.0/65536.0,1,-nbitq), 
to_sfixed(-3090.0/65536.0,1,-nbitq), 
to_sfixed(-1041.0/65536.0,1,-nbitq), 
to_sfixed(1207.0/65536.0,1,-nbitq), 
to_sfixed(-587.0/65536.0,1,-nbitq), 
to_sfixed(-342.0/65536.0,1,-nbitq), 
to_sfixed(2941.0/65536.0,1,-nbitq), 
to_sfixed(-1158.0/65536.0,1,-nbitq), 
to_sfixed(-2141.0/65536.0,1,-nbitq), 
to_sfixed(651.0/65536.0,1,-nbitq), 
to_sfixed(-1463.0/65536.0,1,-nbitq), 
to_sfixed(-910.0/65536.0,1,-nbitq), 
to_sfixed(343.0/65536.0,1,-nbitq), 
to_sfixed(-2777.0/65536.0,1,-nbitq), 
to_sfixed(308.0/65536.0,1,-nbitq), 
to_sfixed(428.0/65536.0,1,-nbitq), 
to_sfixed(1618.0/65536.0,1,-nbitq), 
to_sfixed(-1442.0/65536.0,1,-nbitq), 
to_sfixed(902.0/65536.0,1,-nbitq), 
to_sfixed(-492.0/65536.0,1,-nbitq), 
to_sfixed(-1914.0/65536.0,1,-nbitq), 
to_sfixed(-1215.0/65536.0,1,-nbitq), 
to_sfixed(-2981.0/65536.0,1,-nbitq), 
to_sfixed(-2737.0/65536.0,1,-nbitq), 
to_sfixed(-1090.0/65536.0,1,-nbitq), 
to_sfixed(-318.0/65536.0,1,-nbitq), 
to_sfixed(-1134.0/65536.0,1,-nbitq), 
to_sfixed(-2181.0/65536.0,1,-nbitq), 
to_sfixed(260.0/65536.0,1,-nbitq), 
to_sfixed(-1624.0/65536.0,1,-nbitq), 
to_sfixed(2495.0/65536.0,1,-nbitq), 
to_sfixed(-1435.0/65536.0,1,-nbitq), 
to_sfixed(590.0/65536.0,1,-nbitq), 
to_sfixed(-1300.0/65536.0,1,-nbitq), 
to_sfixed(3706.0/65536.0,1,-nbitq), 
to_sfixed(-827.0/65536.0,1,-nbitq), 
to_sfixed(1302.0/65536.0,1,-nbitq), 
to_sfixed(2936.0/65536.0,1,-nbitq), 
to_sfixed(618.0/65536.0,1,-nbitq), 
to_sfixed(-777.0/65536.0,1,-nbitq), 
to_sfixed(-2520.0/65536.0,1,-nbitq), 
to_sfixed(-1812.0/65536.0,1,-nbitq), 
to_sfixed(2656.0/65536.0,1,-nbitq), 
to_sfixed(2025.0/65536.0,1,-nbitq), 
to_sfixed(-347.0/65536.0,1,-nbitq), 
to_sfixed(-1472.0/65536.0,1,-nbitq), 
to_sfixed(1464.0/65536.0,1,-nbitq), 
to_sfixed(2140.0/65536.0,1,-nbitq), 
to_sfixed(3867.0/65536.0,1,-nbitq), 
to_sfixed(-515.0/65536.0,1,-nbitq), 
to_sfixed(755.0/65536.0,1,-nbitq), 
to_sfixed(-165.0/65536.0,1,-nbitq), 
to_sfixed(-2553.0/65536.0,1,-nbitq), 
to_sfixed(1164.0/65536.0,1,-nbitq), 
to_sfixed(4126.0/65536.0,1,-nbitq), 
to_sfixed(-381.0/65536.0,1,-nbitq), 
to_sfixed(-1488.0/65536.0,1,-nbitq), 
to_sfixed(-322.0/65536.0,1,-nbitq), 
to_sfixed(-2301.0/65536.0,1,-nbitq), 
to_sfixed(-134.0/65536.0,1,-nbitq), 
to_sfixed(-1456.0/65536.0,1,-nbitq), 
to_sfixed(2321.0/65536.0,1,-nbitq), 
to_sfixed(-912.0/65536.0,1,-nbitq), 
to_sfixed(2293.0/65536.0,1,-nbitq), 
to_sfixed(67.0/65536.0,1,-nbitq), 
to_sfixed(-630.0/65536.0,1,-nbitq), 
to_sfixed(325.0/65536.0,1,-nbitq), 
to_sfixed(-188.0/65536.0,1,-nbitq), 
to_sfixed(1602.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1611.0/65536.0,1,-nbitq), 
to_sfixed(2309.0/65536.0,1,-nbitq), 
to_sfixed(-1372.0/65536.0,1,-nbitq), 
to_sfixed(197.0/65536.0,1,-nbitq), 
to_sfixed(1324.0/65536.0,1,-nbitq), 
to_sfixed(-2231.0/65536.0,1,-nbitq), 
to_sfixed(-270.0/65536.0,1,-nbitq), 
to_sfixed(2919.0/65536.0,1,-nbitq), 
to_sfixed(-2037.0/65536.0,1,-nbitq), 
to_sfixed(-1347.0/65536.0,1,-nbitq), 
to_sfixed(2140.0/65536.0,1,-nbitq), 
to_sfixed(2095.0/65536.0,1,-nbitq), 
to_sfixed(-752.0/65536.0,1,-nbitq), 
to_sfixed(-2193.0/65536.0,1,-nbitq), 
to_sfixed(1272.0/65536.0,1,-nbitq), 
to_sfixed(-845.0/65536.0,1,-nbitq), 
to_sfixed(2698.0/65536.0,1,-nbitq), 
to_sfixed(2969.0/65536.0,1,-nbitq), 
to_sfixed(551.0/65536.0,1,-nbitq), 
to_sfixed(-1919.0/65536.0,1,-nbitq), 
to_sfixed(-33.0/65536.0,1,-nbitq), 
to_sfixed(-1005.0/65536.0,1,-nbitq), 
to_sfixed(897.0/65536.0,1,-nbitq), 
to_sfixed(-1940.0/65536.0,1,-nbitq), 
to_sfixed(1798.0/65536.0,1,-nbitq), 
to_sfixed(3873.0/65536.0,1,-nbitq), 
to_sfixed(976.0/65536.0,1,-nbitq), 
to_sfixed(2299.0/65536.0,1,-nbitq), 
to_sfixed(1754.0/65536.0,1,-nbitq), 
to_sfixed(1220.0/65536.0,1,-nbitq), 
to_sfixed(1713.0/65536.0,1,-nbitq), 
to_sfixed(799.0/65536.0,1,-nbitq), 
to_sfixed(-2075.0/65536.0,1,-nbitq), 
to_sfixed(-2015.0/65536.0,1,-nbitq), 
to_sfixed(-2772.0/65536.0,1,-nbitq), 
to_sfixed(-2498.0/65536.0,1,-nbitq), 
to_sfixed(-163.0/65536.0,1,-nbitq), 
to_sfixed(1210.0/65536.0,1,-nbitq), 
to_sfixed(-1779.0/65536.0,1,-nbitq), 
to_sfixed(2878.0/65536.0,1,-nbitq), 
to_sfixed(-2249.0/65536.0,1,-nbitq), 
to_sfixed(-590.0/65536.0,1,-nbitq), 
to_sfixed(997.0/65536.0,1,-nbitq), 
to_sfixed(173.0/65536.0,1,-nbitq), 
to_sfixed(2484.0/65536.0,1,-nbitq), 
to_sfixed(2625.0/65536.0,1,-nbitq), 
to_sfixed(375.0/65536.0,1,-nbitq), 
to_sfixed(1000.0/65536.0,1,-nbitq), 
to_sfixed(2475.0/65536.0,1,-nbitq), 
to_sfixed(1320.0/65536.0,1,-nbitq), 
to_sfixed(-2291.0/65536.0,1,-nbitq), 
to_sfixed(1175.0/65536.0,1,-nbitq), 
to_sfixed(1901.0/65536.0,1,-nbitq), 
to_sfixed(988.0/65536.0,1,-nbitq), 
to_sfixed(3700.0/65536.0,1,-nbitq), 
to_sfixed(-353.0/65536.0,1,-nbitq), 
to_sfixed(-2075.0/65536.0,1,-nbitq), 
to_sfixed(1988.0/65536.0,1,-nbitq), 
to_sfixed(2500.0/65536.0,1,-nbitq), 
to_sfixed(-1176.0/65536.0,1,-nbitq), 
to_sfixed(-707.0/65536.0,1,-nbitq), 
to_sfixed(-407.0/65536.0,1,-nbitq), 
to_sfixed(-1182.0/65536.0,1,-nbitq), 
to_sfixed(1451.0/65536.0,1,-nbitq), 
to_sfixed(-776.0/65536.0,1,-nbitq), 
to_sfixed(-1132.0/65536.0,1,-nbitq), 
to_sfixed(-2308.0/65536.0,1,-nbitq), 
to_sfixed(-2092.0/65536.0,1,-nbitq), 
to_sfixed(-1000.0/65536.0,1,-nbitq), 
to_sfixed(1190.0/65536.0,1,-nbitq), 
to_sfixed(2013.0/65536.0,1,-nbitq), 
to_sfixed(914.0/65536.0,1,-nbitq), 
to_sfixed(1798.0/65536.0,1,-nbitq), 
to_sfixed(1366.0/65536.0,1,-nbitq), 
to_sfixed(-1042.0/65536.0,1,-nbitq), 
to_sfixed(-2006.0/65536.0,1,-nbitq), 
to_sfixed(1090.0/65536.0,1,-nbitq), 
to_sfixed(750.0/65536.0,1,-nbitq), 
to_sfixed(-809.0/65536.0,1,-nbitq), 
to_sfixed(2640.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2289.0/65536.0,1,-nbitq), 
to_sfixed(-1177.0/65536.0,1,-nbitq), 
to_sfixed(1595.0/65536.0,1,-nbitq), 
to_sfixed(-17.0/65536.0,1,-nbitq), 
to_sfixed(-1454.0/65536.0,1,-nbitq), 
to_sfixed(4171.0/65536.0,1,-nbitq), 
to_sfixed(-115.0/65536.0,1,-nbitq), 
to_sfixed(-2212.0/65536.0,1,-nbitq), 
to_sfixed(-879.0/65536.0,1,-nbitq), 
to_sfixed(1546.0/65536.0,1,-nbitq), 
to_sfixed(3576.0/65536.0,1,-nbitq), 
to_sfixed(3037.0/65536.0,1,-nbitq), 
to_sfixed(-591.0/65536.0,1,-nbitq), 
to_sfixed(3329.0/65536.0,1,-nbitq), 
to_sfixed(98.0/65536.0,1,-nbitq), 
to_sfixed(-226.0/65536.0,1,-nbitq), 
to_sfixed(469.0/65536.0,1,-nbitq), 
to_sfixed(2043.0/65536.0,1,-nbitq), 
to_sfixed(637.0/65536.0,1,-nbitq), 
to_sfixed(1854.0/65536.0,1,-nbitq), 
to_sfixed(675.0/65536.0,1,-nbitq), 
to_sfixed(-314.0/65536.0,1,-nbitq), 
to_sfixed(-479.0/65536.0,1,-nbitq), 
to_sfixed(1330.0/65536.0,1,-nbitq), 
to_sfixed(-2413.0/65536.0,1,-nbitq), 
to_sfixed(8101.0/65536.0,1,-nbitq), 
to_sfixed(-142.0/65536.0,1,-nbitq), 
to_sfixed(-1562.0/65536.0,1,-nbitq), 
to_sfixed(1596.0/65536.0,1,-nbitq), 
to_sfixed(1691.0/65536.0,1,-nbitq), 
to_sfixed(-2112.0/65536.0,1,-nbitq), 
to_sfixed(2876.0/65536.0,1,-nbitq), 
to_sfixed(2659.0/65536.0,1,-nbitq), 
to_sfixed(-340.0/65536.0,1,-nbitq), 
to_sfixed(-1354.0/65536.0,1,-nbitq), 
to_sfixed(1229.0/65536.0,1,-nbitq), 
to_sfixed(-2963.0/65536.0,1,-nbitq), 
to_sfixed(-1842.0/65536.0,1,-nbitq), 
to_sfixed(-3523.0/65536.0,1,-nbitq), 
to_sfixed(-2369.0/65536.0,1,-nbitq), 
to_sfixed(-1101.0/65536.0,1,-nbitq), 
to_sfixed(-2542.0/65536.0,1,-nbitq), 
to_sfixed(-2150.0/65536.0,1,-nbitq), 
to_sfixed(-2065.0/65536.0,1,-nbitq), 
to_sfixed(-1047.0/65536.0,1,-nbitq), 
to_sfixed(2197.0/65536.0,1,-nbitq), 
to_sfixed(-2346.0/65536.0,1,-nbitq), 
to_sfixed(1127.0/65536.0,1,-nbitq), 
to_sfixed(2053.0/65536.0,1,-nbitq), 
to_sfixed(4682.0/65536.0,1,-nbitq), 
to_sfixed(2547.0/65536.0,1,-nbitq), 
to_sfixed(-3053.0/65536.0,1,-nbitq), 
to_sfixed(2039.0/65536.0,1,-nbitq), 
to_sfixed(-2368.0/65536.0,1,-nbitq), 
to_sfixed(1781.0/65536.0,1,-nbitq), 
to_sfixed(-163.0/65536.0,1,-nbitq), 
to_sfixed(793.0/65536.0,1,-nbitq), 
to_sfixed(1154.0/65536.0,1,-nbitq), 
to_sfixed(1372.0/65536.0,1,-nbitq), 
to_sfixed(2200.0/65536.0,1,-nbitq), 
to_sfixed(-2344.0/65536.0,1,-nbitq), 
to_sfixed(1433.0/65536.0,1,-nbitq), 
to_sfixed(2053.0/65536.0,1,-nbitq), 
to_sfixed(384.0/65536.0,1,-nbitq), 
to_sfixed(-2556.0/65536.0,1,-nbitq), 
to_sfixed(1631.0/65536.0,1,-nbitq), 
to_sfixed(-3840.0/65536.0,1,-nbitq), 
to_sfixed(-4422.0/65536.0,1,-nbitq), 
to_sfixed(293.0/65536.0,1,-nbitq), 
to_sfixed(3752.0/65536.0,1,-nbitq), 
to_sfixed(-2569.0/65536.0,1,-nbitq), 
to_sfixed(-618.0/65536.0,1,-nbitq), 
to_sfixed(2454.0/65536.0,1,-nbitq), 
to_sfixed(-2621.0/65536.0,1,-nbitq), 
to_sfixed(2397.0/65536.0,1,-nbitq), 
to_sfixed(-607.0/65536.0,1,-nbitq), 
to_sfixed(-5368.0/65536.0,1,-nbitq), 
to_sfixed(762.0/65536.0,1,-nbitq), 
to_sfixed(-2598.0/65536.0,1,-nbitq), 
to_sfixed(-3782.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3466.0/65536.0,1,-nbitq), 
to_sfixed(2165.0/65536.0,1,-nbitq), 
to_sfixed(2710.0/65536.0,1,-nbitq), 
to_sfixed(1544.0/65536.0,1,-nbitq), 
to_sfixed(-3565.0/65536.0,1,-nbitq), 
to_sfixed(4082.0/65536.0,1,-nbitq), 
to_sfixed(-3110.0/65536.0,1,-nbitq), 
to_sfixed(-1889.0/65536.0,1,-nbitq), 
to_sfixed(-86.0/65536.0,1,-nbitq), 
to_sfixed(2649.0/65536.0,1,-nbitq), 
to_sfixed(-782.0/65536.0,1,-nbitq), 
to_sfixed(9626.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(3653.0/65536.0,1,-nbitq), 
to_sfixed(7882.0/65536.0,1,-nbitq), 
to_sfixed(-1813.0/65536.0,1,-nbitq), 
to_sfixed(-1988.0/65536.0,1,-nbitq), 
to_sfixed(-1253.0/65536.0,1,-nbitq), 
to_sfixed(2651.0/65536.0,1,-nbitq), 
to_sfixed(-755.0/65536.0,1,-nbitq), 
to_sfixed(1063.0/65536.0,1,-nbitq), 
to_sfixed(1065.0/65536.0,1,-nbitq), 
to_sfixed(2300.0/65536.0,1,-nbitq), 
to_sfixed(-2948.0/65536.0,1,-nbitq), 
to_sfixed(-2445.0/65536.0,1,-nbitq), 
to_sfixed(6812.0/65536.0,1,-nbitq), 
to_sfixed(1000.0/65536.0,1,-nbitq), 
to_sfixed(-1660.0/65536.0,1,-nbitq), 
to_sfixed(5424.0/65536.0,1,-nbitq), 
to_sfixed(1930.0/65536.0,1,-nbitq), 
to_sfixed(-815.0/65536.0,1,-nbitq), 
to_sfixed(1949.0/65536.0,1,-nbitq), 
to_sfixed(516.0/65536.0,1,-nbitq), 
to_sfixed(528.0/65536.0,1,-nbitq), 
to_sfixed(-1711.0/65536.0,1,-nbitq), 
to_sfixed(-1273.0/65536.0,1,-nbitq), 
to_sfixed(-3293.0/65536.0,1,-nbitq), 
to_sfixed(-2198.0/65536.0,1,-nbitq), 
to_sfixed(-1526.0/65536.0,1,-nbitq), 
to_sfixed(1074.0/65536.0,1,-nbitq), 
to_sfixed(-7495.0/65536.0,1,-nbitq), 
to_sfixed(-2040.0/65536.0,1,-nbitq), 
to_sfixed(2214.0/65536.0,1,-nbitq), 
to_sfixed(-3208.0/65536.0,1,-nbitq), 
to_sfixed(2285.0/65536.0,1,-nbitq), 
to_sfixed(7199.0/65536.0,1,-nbitq), 
to_sfixed(-46.0/65536.0,1,-nbitq), 
to_sfixed(412.0/65536.0,1,-nbitq), 
to_sfixed(107.0/65536.0,1,-nbitq), 
to_sfixed(684.0/65536.0,1,-nbitq), 
to_sfixed(-1248.0/65536.0,1,-nbitq), 
to_sfixed(-1210.0/65536.0,1,-nbitq), 
to_sfixed(2628.0/65536.0,1,-nbitq), 
to_sfixed(1866.0/65536.0,1,-nbitq), 
to_sfixed(-4219.0/65536.0,1,-nbitq), 
to_sfixed(3264.0/65536.0,1,-nbitq), 
to_sfixed(274.0/65536.0,1,-nbitq), 
to_sfixed(-2386.0/65536.0,1,-nbitq), 
to_sfixed(-2464.0/65536.0,1,-nbitq), 
to_sfixed(-1273.0/65536.0,1,-nbitq), 
to_sfixed(-3000.0/65536.0,1,-nbitq), 
to_sfixed(-521.0/65536.0,1,-nbitq), 
to_sfixed(-2251.0/65536.0,1,-nbitq), 
to_sfixed(799.0/65536.0,1,-nbitq), 
to_sfixed(-3798.0/65536.0,1,-nbitq), 
to_sfixed(3681.0/65536.0,1,-nbitq), 
to_sfixed(-1691.0/65536.0,1,-nbitq), 
to_sfixed(-4958.0/65536.0,1,-nbitq), 
to_sfixed(-4164.0/65536.0,1,-nbitq), 
to_sfixed(-2449.0/65536.0,1,-nbitq), 
to_sfixed(-2007.0/65536.0,1,-nbitq), 
to_sfixed(607.0/65536.0,1,-nbitq), 
to_sfixed(-1780.0/65536.0,1,-nbitq), 
to_sfixed(-2676.0/65536.0,1,-nbitq), 
to_sfixed(942.0/65536.0,1,-nbitq), 
to_sfixed(100.0/65536.0,1,-nbitq), 
to_sfixed(-4730.0/65536.0,1,-nbitq), 
to_sfixed(559.0/65536.0,1,-nbitq), 
to_sfixed(-2538.0/65536.0,1,-nbitq), 
to_sfixed(-573.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-502.0/65536.0,1,-nbitq), 
to_sfixed(346.0/65536.0,1,-nbitq), 
to_sfixed(1306.0/65536.0,1,-nbitq), 
to_sfixed(5538.0/65536.0,1,-nbitq), 
to_sfixed(1491.0/65536.0,1,-nbitq), 
to_sfixed(2392.0/65536.0,1,-nbitq), 
to_sfixed(-4822.0/65536.0,1,-nbitq), 
to_sfixed(-1249.0/65536.0,1,-nbitq), 
to_sfixed(3409.0/65536.0,1,-nbitq), 
to_sfixed(93.0/65536.0,1,-nbitq), 
to_sfixed(204.0/65536.0,1,-nbitq), 
to_sfixed(13830.0/65536.0,1,-nbitq), 
to_sfixed(2225.0/65536.0,1,-nbitq), 
to_sfixed(1823.0/65536.0,1,-nbitq), 
to_sfixed(6097.0/65536.0,1,-nbitq), 
to_sfixed(-2844.0/65536.0,1,-nbitq), 
to_sfixed(-1830.0/65536.0,1,-nbitq), 
to_sfixed(-3967.0/65536.0,1,-nbitq), 
to_sfixed(3645.0/65536.0,1,-nbitq), 
to_sfixed(-198.0/65536.0,1,-nbitq), 
to_sfixed(5796.0/65536.0,1,-nbitq), 
to_sfixed(142.0/65536.0,1,-nbitq), 
to_sfixed(779.0/65536.0,1,-nbitq), 
to_sfixed(-978.0/65536.0,1,-nbitq), 
to_sfixed(2590.0/65536.0,1,-nbitq), 
to_sfixed(6469.0/65536.0,1,-nbitq), 
to_sfixed(842.0/65536.0,1,-nbitq), 
to_sfixed(401.0/65536.0,1,-nbitq), 
to_sfixed(2907.0/65536.0,1,-nbitq), 
to_sfixed(2067.0/65536.0,1,-nbitq), 
to_sfixed(-2140.0/65536.0,1,-nbitq), 
to_sfixed(1237.0/65536.0,1,-nbitq), 
to_sfixed(2219.0/65536.0,1,-nbitq), 
to_sfixed(79.0/65536.0,1,-nbitq), 
to_sfixed(-2404.0/65536.0,1,-nbitq), 
to_sfixed(1287.0/65536.0,1,-nbitq), 
to_sfixed(-5278.0/65536.0,1,-nbitq), 
to_sfixed(2767.0/65536.0,1,-nbitq), 
to_sfixed(-2554.0/65536.0,1,-nbitq), 
to_sfixed(-6062.0/65536.0,1,-nbitq), 
to_sfixed(-11698.0/65536.0,1,-nbitq), 
to_sfixed(-376.0/65536.0,1,-nbitq), 
to_sfixed(3983.0/65536.0,1,-nbitq), 
to_sfixed(-278.0/65536.0,1,-nbitq), 
to_sfixed(-1473.0/65536.0,1,-nbitq), 
to_sfixed(-571.0/65536.0,1,-nbitq), 
to_sfixed(-909.0/65536.0,1,-nbitq), 
to_sfixed(-2202.0/65536.0,1,-nbitq), 
to_sfixed(2644.0/65536.0,1,-nbitq), 
to_sfixed(3375.0/65536.0,1,-nbitq), 
to_sfixed(-232.0/65536.0,1,-nbitq), 
to_sfixed(-441.0/65536.0,1,-nbitq), 
to_sfixed(2162.0/65536.0,1,-nbitq), 
to_sfixed(4653.0/65536.0,1,-nbitq), 
to_sfixed(-1879.0/65536.0,1,-nbitq), 
to_sfixed(7067.0/65536.0,1,-nbitq), 
to_sfixed(1922.0/65536.0,1,-nbitq), 
to_sfixed(-2294.0/65536.0,1,-nbitq), 
to_sfixed(-101.0/65536.0,1,-nbitq), 
to_sfixed(-2359.0/65536.0,1,-nbitq), 
to_sfixed(-125.0/65536.0,1,-nbitq), 
to_sfixed(-633.0/65536.0,1,-nbitq), 
to_sfixed(-1148.0/65536.0,1,-nbitq), 
to_sfixed(-2059.0/65536.0,1,-nbitq), 
to_sfixed(-1356.0/65536.0,1,-nbitq), 
to_sfixed(3293.0/65536.0,1,-nbitq), 
to_sfixed(-3116.0/65536.0,1,-nbitq), 
to_sfixed(-5265.0/65536.0,1,-nbitq), 
to_sfixed(-2165.0/65536.0,1,-nbitq), 
to_sfixed(-3881.0/65536.0,1,-nbitq), 
to_sfixed(-906.0/65536.0,1,-nbitq), 
to_sfixed(-4540.0/65536.0,1,-nbitq), 
to_sfixed(-1839.0/65536.0,1,-nbitq), 
to_sfixed(-2187.0/65536.0,1,-nbitq), 
to_sfixed(-246.0/65536.0,1,-nbitq), 
to_sfixed(4808.0/65536.0,1,-nbitq), 
to_sfixed(-410.0/65536.0,1,-nbitq), 
to_sfixed(1029.0/65536.0,1,-nbitq), 
to_sfixed(2435.0/65536.0,1,-nbitq), 
to_sfixed(-1166.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-892.0/65536.0,1,-nbitq), 
to_sfixed(351.0/65536.0,1,-nbitq), 
to_sfixed(8225.0/65536.0,1,-nbitq), 
to_sfixed(7262.0/65536.0,1,-nbitq), 
to_sfixed(-2451.0/65536.0,1,-nbitq), 
to_sfixed(3926.0/65536.0,1,-nbitq), 
to_sfixed(-929.0/65536.0,1,-nbitq), 
to_sfixed(1337.0/65536.0,1,-nbitq), 
to_sfixed(2237.0/65536.0,1,-nbitq), 
to_sfixed(84.0/65536.0,1,-nbitq), 
to_sfixed(2603.0/65536.0,1,-nbitq), 
to_sfixed(16157.0/65536.0,1,-nbitq), 
to_sfixed(-565.0/65536.0,1,-nbitq), 
to_sfixed(-738.0/65536.0,1,-nbitq), 
to_sfixed(-303.0/65536.0,1,-nbitq), 
to_sfixed(-2979.0/65536.0,1,-nbitq), 
to_sfixed(-2031.0/65536.0,1,-nbitq), 
to_sfixed(-5392.0/65536.0,1,-nbitq), 
to_sfixed(4306.0/65536.0,1,-nbitq), 
to_sfixed(2169.0/65536.0,1,-nbitq), 
to_sfixed(3515.0/65536.0,1,-nbitq), 
to_sfixed(1389.0/65536.0,1,-nbitq), 
to_sfixed(3138.0/65536.0,1,-nbitq), 
to_sfixed(-5702.0/65536.0,1,-nbitq), 
to_sfixed(5470.0/65536.0,1,-nbitq), 
to_sfixed(5124.0/65536.0,1,-nbitq), 
to_sfixed(-2354.0/65536.0,1,-nbitq), 
to_sfixed(857.0/65536.0,1,-nbitq), 
to_sfixed(-2962.0/65536.0,1,-nbitq), 
to_sfixed(5747.0/65536.0,1,-nbitq), 
to_sfixed(1337.0/65536.0,1,-nbitq), 
to_sfixed(-2135.0/65536.0,1,-nbitq), 
to_sfixed(6962.0/65536.0,1,-nbitq), 
to_sfixed(1051.0/65536.0,1,-nbitq), 
to_sfixed(-4177.0/65536.0,1,-nbitq), 
to_sfixed(-572.0/65536.0,1,-nbitq), 
to_sfixed(-5581.0/65536.0,1,-nbitq), 
to_sfixed(1604.0/65536.0,1,-nbitq), 
to_sfixed(2332.0/65536.0,1,-nbitq), 
to_sfixed(-6875.0/65536.0,1,-nbitq), 
to_sfixed(-12058.0/65536.0,1,-nbitq), 
to_sfixed(1219.0/65536.0,1,-nbitq), 
to_sfixed(469.0/65536.0,1,-nbitq), 
to_sfixed(-1736.0/65536.0,1,-nbitq), 
to_sfixed(2385.0/65536.0,1,-nbitq), 
to_sfixed(-7457.0/65536.0,1,-nbitq), 
to_sfixed(-1022.0/65536.0,1,-nbitq), 
to_sfixed(-4040.0/65536.0,1,-nbitq), 
to_sfixed(1964.0/65536.0,1,-nbitq), 
to_sfixed(2331.0/65536.0,1,-nbitq), 
to_sfixed(-331.0/65536.0,1,-nbitq), 
to_sfixed(350.0/65536.0,1,-nbitq), 
to_sfixed(1666.0/65536.0,1,-nbitq), 
to_sfixed(3813.0/65536.0,1,-nbitq), 
to_sfixed(-7009.0/65536.0,1,-nbitq), 
to_sfixed(10095.0/65536.0,1,-nbitq), 
to_sfixed(663.0/65536.0,1,-nbitq), 
to_sfixed(-1586.0/65536.0,1,-nbitq), 
to_sfixed(1524.0/65536.0,1,-nbitq), 
to_sfixed(-1712.0/65536.0,1,-nbitq), 
to_sfixed(-2736.0/65536.0,1,-nbitq), 
to_sfixed(-2602.0/65536.0,1,-nbitq), 
to_sfixed(2509.0/65536.0,1,-nbitq), 
to_sfixed(-3274.0/65536.0,1,-nbitq), 
to_sfixed(754.0/65536.0,1,-nbitq), 
to_sfixed(6775.0/65536.0,1,-nbitq), 
to_sfixed(-1909.0/65536.0,1,-nbitq), 
to_sfixed(-9819.0/65536.0,1,-nbitq), 
to_sfixed(-3497.0/65536.0,1,-nbitq), 
to_sfixed(-7934.0/65536.0,1,-nbitq), 
to_sfixed(-2350.0/65536.0,1,-nbitq), 
to_sfixed(-7434.0/65536.0,1,-nbitq), 
to_sfixed(-384.0/65536.0,1,-nbitq), 
to_sfixed(-2515.0/65536.0,1,-nbitq), 
to_sfixed(1672.0/65536.0,1,-nbitq), 
to_sfixed(-3834.0/65536.0,1,-nbitq), 
to_sfixed(-444.0/65536.0,1,-nbitq), 
to_sfixed(-280.0/65536.0,1,-nbitq), 
to_sfixed(1676.0/65536.0,1,-nbitq), 
to_sfixed(779.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1598.0/65536.0,1,-nbitq), 
to_sfixed(748.0/65536.0,1,-nbitq), 
to_sfixed(1591.0/65536.0,1,-nbitq), 
to_sfixed(9011.0/65536.0,1,-nbitq), 
to_sfixed(-3844.0/65536.0,1,-nbitq), 
to_sfixed(4531.0/65536.0,1,-nbitq), 
to_sfixed(2630.0/65536.0,1,-nbitq), 
to_sfixed(2532.0/65536.0,1,-nbitq), 
to_sfixed(-628.0/65536.0,1,-nbitq), 
to_sfixed(-2312.0/65536.0,1,-nbitq), 
to_sfixed(3859.0/65536.0,1,-nbitq), 
to_sfixed(14671.0/65536.0,1,-nbitq), 
to_sfixed(-160.0/65536.0,1,-nbitq), 
to_sfixed(3307.0/65536.0,1,-nbitq), 
to_sfixed(-6250.0/65536.0,1,-nbitq), 
to_sfixed(306.0/65536.0,1,-nbitq), 
to_sfixed(1905.0/65536.0,1,-nbitq), 
to_sfixed(-2052.0/65536.0,1,-nbitq), 
to_sfixed(-1767.0/65536.0,1,-nbitq), 
to_sfixed(1353.0/65536.0,1,-nbitq), 
to_sfixed(6312.0/65536.0,1,-nbitq), 
to_sfixed(-4631.0/65536.0,1,-nbitq), 
to_sfixed(-1229.0/65536.0,1,-nbitq), 
to_sfixed(-3853.0/65536.0,1,-nbitq), 
to_sfixed(5174.0/65536.0,1,-nbitq), 
to_sfixed(7063.0/65536.0,1,-nbitq), 
to_sfixed(-5064.0/65536.0,1,-nbitq), 
to_sfixed(-462.0/65536.0,1,-nbitq), 
to_sfixed(618.0/65536.0,1,-nbitq), 
to_sfixed(4641.0/65536.0,1,-nbitq), 
to_sfixed(-630.0/65536.0,1,-nbitq), 
to_sfixed(1515.0/65536.0,1,-nbitq), 
to_sfixed(11651.0/65536.0,1,-nbitq), 
to_sfixed(-1681.0/65536.0,1,-nbitq), 
to_sfixed(-3415.0/65536.0,1,-nbitq), 
to_sfixed(2541.0/65536.0,1,-nbitq), 
to_sfixed(-5775.0/65536.0,1,-nbitq), 
to_sfixed(-3628.0/65536.0,1,-nbitq), 
to_sfixed(-4801.0/65536.0,1,-nbitq), 
to_sfixed(607.0/65536.0,1,-nbitq), 
to_sfixed(-10128.0/65536.0,1,-nbitq), 
to_sfixed(307.0/65536.0,1,-nbitq), 
to_sfixed(5499.0/65536.0,1,-nbitq), 
to_sfixed(-378.0/65536.0,1,-nbitq), 
to_sfixed(1641.0/65536.0,1,-nbitq), 
to_sfixed(-5561.0/65536.0,1,-nbitq), 
to_sfixed(-1315.0/65536.0,1,-nbitq), 
to_sfixed(-255.0/65536.0,1,-nbitq), 
to_sfixed(2786.0/65536.0,1,-nbitq), 
to_sfixed(-2607.0/65536.0,1,-nbitq), 
to_sfixed(1781.0/65536.0,1,-nbitq), 
to_sfixed(6050.0/65536.0,1,-nbitq), 
to_sfixed(-1962.0/65536.0,1,-nbitq), 
to_sfixed(-337.0/65536.0,1,-nbitq), 
to_sfixed(-422.0/65536.0,1,-nbitq), 
to_sfixed(9231.0/65536.0,1,-nbitq), 
to_sfixed(-3005.0/65536.0,1,-nbitq), 
to_sfixed(-1964.0/65536.0,1,-nbitq), 
to_sfixed(-2925.0/65536.0,1,-nbitq), 
to_sfixed(2784.0/65536.0,1,-nbitq), 
to_sfixed(130.0/65536.0,1,-nbitq), 
to_sfixed(504.0/65536.0,1,-nbitq), 
to_sfixed(-1816.0/65536.0,1,-nbitq), 
to_sfixed(1785.0/65536.0,1,-nbitq), 
to_sfixed(-2771.0/65536.0,1,-nbitq), 
to_sfixed(7590.0/65536.0,1,-nbitq), 
to_sfixed(-3467.0/65536.0,1,-nbitq), 
to_sfixed(-7997.0/65536.0,1,-nbitq), 
to_sfixed(-695.0/65536.0,1,-nbitq), 
to_sfixed(-4665.0/65536.0,1,-nbitq), 
to_sfixed(-2871.0/65536.0,1,-nbitq), 
to_sfixed(-3816.0/65536.0,1,-nbitq), 
to_sfixed(-4455.0/65536.0,1,-nbitq), 
to_sfixed(1474.0/65536.0,1,-nbitq), 
to_sfixed(473.0/65536.0,1,-nbitq), 
to_sfixed(192.0/65536.0,1,-nbitq), 
to_sfixed(-427.0/65536.0,1,-nbitq), 
to_sfixed(822.0/65536.0,1,-nbitq), 
to_sfixed(-1154.0/65536.0,1,-nbitq), 
to_sfixed(-3351.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-334.0/65536.0,1,-nbitq), 
to_sfixed(971.0/65536.0,1,-nbitq), 
to_sfixed(2305.0/65536.0,1,-nbitq), 
to_sfixed(4925.0/65536.0,1,-nbitq), 
to_sfixed(-10245.0/65536.0,1,-nbitq), 
to_sfixed(-1092.0/65536.0,1,-nbitq), 
to_sfixed(-126.0/65536.0,1,-nbitq), 
to_sfixed(3214.0/65536.0,1,-nbitq), 
to_sfixed(5209.0/65536.0,1,-nbitq), 
to_sfixed(-2422.0/65536.0,1,-nbitq), 
to_sfixed(5274.0/65536.0,1,-nbitq), 
to_sfixed(10513.0/65536.0,1,-nbitq), 
to_sfixed(-761.0/65536.0,1,-nbitq), 
to_sfixed(6955.0/65536.0,1,-nbitq), 
to_sfixed(-249.0/65536.0,1,-nbitq), 
to_sfixed(-1139.0/65536.0,1,-nbitq), 
to_sfixed(-268.0/65536.0,1,-nbitq), 
to_sfixed(3304.0/65536.0,1,-nbitq), 
to_sfixed(2622.0/65536.0,1,-nbitq), 
to_sfixed(2001.0/65536.0,1,-nbitq), 
to_sfixed(8349.0/65536.0,1,-nbitq), 
to_sfixed(4509.0/65536.0,1,-nbitq), 
to_sfixed(4390.0/65536.0,1,-nbitq), 
to_sfixed(-9195.0/65536.0,1,-nbitq), 
to_sfixed(4267.0/65536.0,1,-nbitq), 
to_sfixed(-1832.0/65536.0,1,-nbitq), 
to_sfixed(742.0/65536.0,1,-nbitq), 
to_sfixed(-1595.0/65536.0,1,-nbitq), 
to_sfixed(-3607.0/65536.0,1,-nbitq), 
to_sfixed(4119.0/65536.0,1,-nbitq), 
to_sfixed(-2766.0/65536.0,1,-nbitq), 
to_sfixed(3996.0/65536.0,1,-nbitq), 
to_sfixed(6404.0/65536.0,1,-nbitq), 
to_sfixed(4186.0/65536.0,1,-nbitq), 
to_sfixed(-4520.0/65536.0,1,-nbitq), 
to_sfixed(2011.0/65536.0,1,-nbitq), 
to_sfixed(2729.0/65536.0,1,-nbitq), 
to_sfixed(-1323.0/65536.0,1,-nbitq), 
to_sfixed(-3726.0/65536.0,1,-nbitq), 
to_sfixed(6127.0/65536.0,1,-nbitq), 
to_sfixed(-11495.0/65536.0,1,-nbitq), 
to_sfixed(1644.0/65536.0,1,-nbitq), 
to_sfixed(13732.0/65536.0,1,-nbitq), 
to_sfixed(-2861.0/65536.0,1,-nbitq), 
to_sfixed(2183.0/65536.0,1,-nbitq), 
to_sfixed(-9657.0/65536.0,1,-nbitq), 
to_sfixed(-1935.0/65536.0,1,-nbitq), 
to_sfixed(4106.0/65536.0,1,-nbitq), 
to_sfixed(-361.0/65536.0,1,-nbitq), 
to_sfixed(-18.0/65536.0,1,-nbitq), 
to_sfixed(-237.0/65536.0,1,-nbitq), 
to_sfixed(6555.0/65536.0,1,-nbitq), 
to_sfixed(2987.0/65536.0,1,-nbitq), 
to_sfixed(10107.0/65536.0,1,-nbitq), 
to_sfixed(-1702.0/65536.0,1,-nbitq), 
to_sfixed(6355.0/65536.0,1,-nbitq), 
to_sfixed(1885.0/65536.0,1,-nbitq), 
to_sfixed(2463.0/65536.0,1,-nbitq), 
to_sfixed(-1706.0/65536.0,1,-nbitq), 
to_sfixed(2089.0/65536.0,1,-nbitq), 
to_sfixed(-2053.0/65536.0,1,-nbitq), 
to_sfixed(-2063.0/65536.0,1,-nbitq), 
to_sfixed(2366.0/65536.0,1,-nbitq), 
to_sfixed(-1656.0/65536.0,1,-nbitq), 
to_sfixed(-5060.0/65536.0,1,-nbitq), 
to_sfixed(9521.0/65536.0,1,-nbitq), 
to_sfixed(-4698.0/65536.0,1,-nbitq), 
to_sfixed(-1736.0/65536.0,1,-nbitq), 
to_sfixed(1259.0/65536.0,1,-nbitq), 
to_sfixed(-4177.0/65536.0,1,-nbitq), 
to_sfixed(-1088.0/65536.0,1,-nbitq), 
to_sfixed(3875.0/65536.0,1,-nbitq), 
to_sfixed(-4907.0/65536.0,1,-nbitq), 
to_sfixed(367.0/65536.0,1,-nbitq), 
to_sfixed(626.0/65536.0,1,-nbitq), 
to_sfixed(1987.0/65536.0,1,-nbitq), 
to_sfixed(-648.0/65536.0,1,-nbitq), 
to_sfixed(1534.0/65536.0,1,-nbitq), 
to_sfixed(971.0/65536.0,1,-nbitq), 
to_sfixed(-4916.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5359.0/65536.0,1,-nbitq), 
to_sfixed(273.0/65536.0,1,-nbitq), 
to_sfixed(10372.0/65536.0,1,-nbitq), 
to_sfixed(3793.0/65536.0,1,-nbitq), 
to_sfixed(-6952.0/65536.0,1,-nbitq), 
to_sfixed(-1406.0/65536.0,1,-nbitq), 
to_sfixed(-1836.0/65536.0,1,-nbitq), 
to_sfixed(6009.0/65536.0,1,-nbitq), 
to_sfixed(1471.0/65536.0,1,-nbitq), 
to_sfixed(293.0/65536.0,1,-nbitq), 
to_sfixed(3708.0/65536.0,1,-nbitq), 
to_sfixed(9648.0/65536.0,1,-nbitq), 
to_sfixed(71.0/65536.0,1,-nbitq), 
to_sfixed(12606.0/65536.0,1,-nbitq), 
to_sfixed(4538.0/65536.0,1,-nbitq), 
to_sfixed(-502.0/65536.0,1,-nbitq), 
to_sfixed(1103.0/65536.0,1,-nbitq), 
to_sfixed(1201.0/65536.0,1,-nbitq), 
to_sfixed(5361.0/65536.0,1,-nbitq), 
to_sfixed(-1919.0/65536.0,1,-nbitq), 
to_sfixed(6400.0/65536.0,1,-nbitq), 
to_sfixed(-3114.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(-7570.0/65536.0,1,-nbitq), 
to_sfixed(-1466.0/65536.0,1,-nbitq), 
to_sfixed(-6902.0/65536.0,1,-nbitq), 
to_sfixed(1939.0/65536.0,1,-nbitq), 
to_sfixed(-2323.0/65536.0,1,-nbitq), 
to_sfixed(-5669.0/65536.0,1,-nbitq), 
to_sfixed(11027.0/65536.0,1,-nbitq), 
to_sfixed(-843.0/65536.0,1,-nbitq), 
to_sfixed(7530.0/65536.0,1,-nbitq), 
to_sfixed(2146.0/65536.0,1,-nbitq), 
to_sfixed(8056.0/65536.0,1,-nbitq), 
to_sfixed(-2017.0/65536.0,1,-nbitq), 
to_sfixed(-704.0/65536.0,1,-nbitq), 
to_sfixed(11437.0/65536.0,1,-nbitq), 
to_sfixed(-7140.0/65536.0,1,-nbitq), 
to_sfixed(-6150.0/65536.0,1,-nbitq), 
to_sfixed(7997.0/65536.0,1,-nbitq), 
to_sfixed(-8716.0/65536.0,1,-nbitq), 
to_sfixed(1500.0/65536.0,1,-nbitq), 
to_sfixed(10369.0/65536.0,1,-nbitq), 
to_sfixed(-2043.0/65536.0,1,-nbitq), 
to_sfixed(2466.0/65536.0,1,-nbitq), 
to_sfixed(-13410.0/65536.0,1,-nbitq), 
to_sfixed(-4542.0/65536.0,1,-nbitq), 
to_sfixed(2880.0/65536.0,1,-nbitq), 
to_sfixed(-561.0/65536.0,1,-nbitq), 
to_sfixed(2017.0/65536.0,1,-nbitq), 
to_sfixed(1887.0/65536.0,1,-nbitq), 
to_sfixed(3886.0/65536.0,1,-nbitq), 
to_sfixed(4838.0/65536.0,1,-nbitq), 
to_sfixed(17571.0/65536.0,1,-nbitq), 
to_sfixed(1979.0/65536.0,1,-nbitq), 
to_sfixed(5084.0/65536.0,1,-nbitq), 
to_sfixed(1593.0/65536.0,1,-nbitq), 
to_sfixed(1458.0/65536.0,1,-nbitq), 
to_sfixed(-2372.0/65536.0,1,-nbitq), 
to_sfixed(1213.0/65536.0,1,-nbitq), 
to_sfixed(3655.0/65536.0,1,-nbitq), 
to_sfixed(814.0/65536.0,1,-nbitq), 
to_sfixed(-2101.0/65536.0,1,-nbitq), 
to_sfixed(1648.0/65536.0,1,-nbitq), 
to_sfixed(170.0/65536.0,1,-nbitq), 
to_sfixed(1333.0/65536.0,1,-nbitq), 
to_sfixed(-5162.0/65536.0,1,-nbitq), 
to_sfixed(-2067.0/65536.0,1,-nbitq), 
to_sfixed(-2070.0/65536.0,1,-nbitq), 
to_sfixed(-133.0/65536.0,1,-nbitq), 
to_sfixed(633.0/65536.0,1,-nbitq), 
to_sfixed(10855.0/65536.0,1,-nbitq), 
to_sfixed(-3218.0/65536.0,1,-nbitq), 
to_sfixed(-2532.0/65536.0,1,-nbitq), 
to_sfixed(-1761.0/65536.0,1,-nbitq), 
to_sfixed(7495.0/65536.0,1,-nbitq), 
to_sfixed(-226.0/65536.0,1,-nbitq), 
to_sfixed(-3405.0/65536.0,1,-nbitq), 
to_sfixed(-2575.0/65536.0,1,-nbitq), 
to_sfixed(-2941.0/65536.0,1,-nbitq)  ), 
( to_sfixed(7952.0/65536.0,1,-nbitq), 
to_sfixed(-342.0/65536.0,1,-nbitq), 
to_sfixed(-6182.0/65536.0,1,-nbitq), 
to_sfixed(3369.0/65536.0,1,-nbitq), 
to_sfixed(5486.0/65536.0,1,-nbitq), 
to_sfixed(-7392.0/65536.0,1,-nbitq), 
to_sfixed(4048.0/65536.0,1,-nbitq), 
to_sfixed(4531.0/65536.0,1,-nbitq), 
to_sfixed(-5271.0/65536.0,1,-nbitq), 
to_sfixed(948.0/65536.0,1,-nbitq), 
to_sfixed(9178.0/65536.0,1,-nbitq), 
to_sfixed(2830.0/65536.0,1,-nbitq), 
to_sfixed(10.0/65536.0,1,-nbitq), 
to_sfixed(-933.0/65536.0,1,-nbitq), 
to_sfixed(2502.0/65536.0,1,-nbitq), 
to_sfixed(1375.0/65536.0,1,-nbitq), 
to_sfixed(-2912.0/65536.0,1,-nbitq), 
to_sfixed(4726.0/65536.0,1,-nbitq), 
to_sfixed(2236.0/65536.0,1,-nbitq), 
to_sfixed(1844.0/65536.0,1,-nbitq), 
to_sfixed(5999.0/65536.0,1,-nbitq), 
to_sfixed(-7952.0/65536.0,1,-nbitq), 
to_sfixed(6092.0/65536.0,1,-nbitq), 
to_sfixed(-3669.0/65536.0,1,-nbitq), 
to_sfixed(3512.0/65536.0,1,-nbitq), 
to_sfixed(-8777.0/65536.0,1,-nbitq), 
to_sfixed(-274.0/65536.0,1,-nbitq), 
to_sfixed(-2577.0/65536.0,1,-nbitq), 
to_sfixed(-6400.0/65536.0,1,-nbitq), 
to_sfixed(7728.0/65536.0,1,-nbitq), 
to_sfixed(1078.0/65536.0,1,-nbitq), 
to_sfixed(5707.0/65536.0,1,-nbitq), 
to_sfixed(4717.0/65536.0,1,-nbitq), 
to_sfixed(3298.0/65536.0,1,-nbitq), 
to_sfixed(-3277.0/65536.0,1,-nbitq), 
to_sfixed(3379.0/65536.0,1,-nbitq), 
to_sfixed(14362.0/65536.0,1,-nbitq), 
to_sfixed(-11602.0/65536.0,1,-nbitq), 
to_sfixed(-15389.0/65536.0,1,-nbitq), 
to_sfixed(6594.0/65536.0,1,-nbitq), 
to_sfixed(21.0/65536.0,1,-nbitq), 
to_sfixed(886.0/65536.0,1,-nbitq), 
to_sfixed(3376.0/65536.0,1,-nbitq), 
to_sfixed(-2739.0/65536.0,1,-nbitq), 
to_sfixed(2610.0/65536.0,1,-nbitq), 
to_sfixed(-18449.0/65536.0,1,-nbitq), 
to_sfixed(-3111.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(1095.0/65536.0,1,-nbitq), 
to_sfixed(1638.0/65536.0,1,-nbitq), 
to_sfixed(-692.0/65536.0,1,-nbitq), 
to_sfixed(3545.0/65536.0,1,-nbitq), 
to_sfixed(1381.0/65536.0,1,-nbitq), 
to_sfixed(10055.0/65536.0,1,-nbitq), 
to_sfixed(-1566.0/65536.0,1,-nbitq), 
to_sfixed(5783.0/65536.0,1,-nbitq), 
to_sfixed(-1990.0/65536.0,1,-nbitq), 
to_sfixed(-2535.0/65536.0,1,-nbitq), 
to_sfixed(-1387.0/65536.0,1,-nbitq), 
to_sfixed(1673.0/65536.0,1,-nbitq), 
to_sfixed(4855.0/65536.0,1,-nbitq), 
to_sfixed(80.0/65536.0,1,-nbitq), 
to_sfixed(-516.0/65536.0,1,-nbitq), 
to_sfixed(2216.0/65536.0,1,-nbitq), 
to_sfixed(-2241.0/65536.0,1,-nbitq), 
to_sfixed(6488.0/65536.0,1,-nbitq), 
to_sfixed(-5257.0/65536.0,1,-nbitq), 
to_sfixed(-8594.0/65536.0,1,-nbitq), 
to_sfixed(-51.0/65536.0,1,-nbitq), 
to_sfixed(4057.0/65536.0,1,-nbitq), 
to_sfixed(-1184.0/65536.0,1,-nbitq), 
to_sfixed(11005.0/65536.0,1,-nbitq), 
to_sfixed(-5337.0/65536.0,1,-nbitq), 
to_sfixed(2290.0/65536.0,1,-nbitq), 
to_sfixed(1192.0/65536.0,1,-nbitq), 
to_sfixed(1370.0/65536.0,1,-nbitq), 
to_sfixed(-33.0/65536.0,1,-nbitq), 
to_sfixed(-15939.0/65536.0,1,-nbitq), 
to_sfixed(-2538.0/65536.0,1,-nbitq), 
to_sfixed(-9713.0/65536.0,1,-nbitq)  ), 
( to_sfixed(7595.0/65536.0,1,-nbitq), 
to_sfixed(-1918.0/65536.0,1,-nbitq), 
to_sfixed(-6346.0/65536.0,1,-nbitq), 
to_sfixed(7015.0/65536.0,1,-nbitq), 
to_sfixed(13108.0/65536.0,1,-nbitq), 
to_sfixed(-7676.0/65536.0,1,-nbitq), 
to_sfixed(6223.0/65536.0,1,-nbitq), 
to_sfixed(3495.0/65536.0,1,-nbitq), 
to_sfixed(2513.0/65536.0,1,-nbitq), 
to_sfixed(2317.0/65536.0,1,-nbitq), 
to_sfixed(5293.0/65536.0,1,-nbitq), 
to_sfixed(4894.0/65536.0,1,-nbitq), 
to_sfixed(40.0/65536.0,1,-nbitq), 
to_sfixed(-5268.0/65536.0,1,-nbitq), 
to_sfixed(2696.0/65536.0,1,-nbitq), 
to_sfixed(-794.0/65536.0,1,-nbitq), 
to_sfixed(1251.0/65536.0,1,-nbitq), 
to_sfixed(6077.0/65536.0,1,-nbitq), 
to_sfixed(-6081.0/65536.0,1,-nbitq), 
to_sfixed(-562.0/65536.0,1,-nbitq), 
to_sfixed(3322.0/65536.0,1,-nbitq), 
to_sfixed(2590.0/65536.0,1,-nbitq), 
to_sfixed(11800.0/65536.0,1,-nbitq), 
to_sfixed(2982.0/65536.0,1,-nbitq), 
to_sfixed(6737.0/65536.0,1,-nbitq), 
to_sfixed(-1390.0/65536.0,1,-nbitq), 
to_sfixed(780.0/65536.0,1,-nbitq), 
to_sfixed(-3069.0/65536.0,1,-nbitq), 
to_sfixed(-4491.0/65536.0,1,-nbitq), 
to_sfixed(1754.0/65536.0,1,-nbitq), 
to_sfixed(-3581.0/65536.0,1,-nbitq), 
to_sfixed(7299.0/65536.0,1,-nbitq), 
to_sfixed(4412.0/65536.0,1,-nbitq), 
to_sfixed(2418.0/65536.0,1,-nbitq), 
to_sfixed(2911.0/65536.0,1,-nbitq), 
to_sfixed(-3459.0/65536.0,1,-nbitq), 
to_sfixed(20826.0/65536.0,1,-nbitq), 
to_sfixed(-7714.0/65536.0,1,-nbitq), 
to_sfixed(-17357.0/65536.0,1,-nbitq), 
to_sfixed(-1306.0/65536.0,1,-nbitq), 
to_sfixed(-4984.0/65536.0,1,-nbitq), 
to_sfixed(-1105.0/65536.0,1,-nbitq), 
to_sfixed(-1586.0/65536.0,1,-nbitq), 
to_sfixed(-4773.0/65536.0,1,-nbitq), 
to_sfixed(-1833.0/65536.0,1,-nbitq), 
to_sfixed(-7987.0/65536.0,1,-nbitq), 
to_sfixed(225.0/65536.0,1,-nbitq), 
to_sfixed(330.0/65536.0,1,-nbitq), 
to_sfixed(336.0/65536.0,1,-nbitq), 
to_sfixed(-3269.0/65536.0,1,-nbitq), 
to_sfixed(2716.0/65536.0,1,-nbitq), 
to_sfixed(293.0/65536.0,1,-nbitq), 
to_sfixed(4557.0/65536.0,1,-nbitq), 
to_sfixed(7268.0/65536.0,1,-nbitq), 
to_sfixed(-5309.0/65536.0,1,-nbitq), 
to_sfixed(8686.0/65536.0,1,-nbitq), 
to_sfixed(-2170.0/65536.0,1,-nbitq), 
to_sfixed(-3786.0/65536.0,1,-nbitq), 
to_sfixed(-3219.0/65536.0,1,-nbitq), 
to_sfixed(-2199.0/65536.0,1,-nbitq), 
to_sfixed(9057.0/65536.0,1,-nbitq), 
to_sfixed(-2101.0/65536.0,1,-nbitq), 
to_sfixed(1562.0/65536.0,1,-nbitq), 
to_sfixed(-2118.0/65536.0,1,-nbitq), 
to_sfixed(-16459.0/65536.0,1,-nbitq), 
to_sfixed(2178.0/65536.0,1,-nbitq), 
to_sfixed(-7089.0/65536.0,1,-nbitq), 
to_sfixed(-9297.0/65536.0,1,-nbitq), 
to_sfixed(-2616.0/65536.0,1,-nbitq), 
to_sfixed(1372.0/65536.0,1,-nbitq), 
to_sfixed(-455.0/65536.0,1,-nbitq), 
to_sfixed(12464.0/65536.0,1,-nbitq), 
to_sfixed(-4602.0/65536.0,1,-nbitq), 
to_sfixed(784.0/65536.0,1,-nbitq), 
to_sfixed(-1835.0/65536.0,1,-nbitq), 
to_sfixed(-5109.0/65536.0,1,-nbitq), 
to_sfixed(2495.0/65536.0,1,-nbitq), 
to_sfixed(-9976.0/65536.0,1,-nbitq), 
to_sfixed(-79.0/65536.0,1,-nbitq), 
to_sfixed(-9868.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4262.0/65536.0,1,-nbitq), 
to_sfixed(-6605.0/65536.0,1,-nbitq), 
to_sfixed(-15973.0/65536.0,1,-nbitq), 
to_sfixed(6054.0/65536.0,1,-nbitq), 
to_sfixed(17023.0/65536.0,1,-nbitq), 
to_sfixed(-7563.0/65536.0,1,-nbitq), 
to_sfixed(2544.0/65536.0,1,-nbitq), 
to_sfixed(717.0/65536.0,1,-nbitq), 
to_sfixed(-3206.0/65536.0,1,-nbitq), 
to_sfixed(1804.0/65536.0,1,-nbitq), 
to_sfixed(7438.0/65536.0,1,-nbitq), 
to_sfixed(8323.0/65536.0,1,-nbitq), 
to_sfixed(3799.0/65536.0,1,-nbitq), 
to_sfixed(-3450.0/65536.0,1,-nbitq), 
to_sfixed(-4794.0/65536.0,1,-nbitq), 
to_sfixed(1819.0/65536.0,1,-nbitq), 
to_sfixed(132.0/65536.0,1,-nbitq), 
to_sfixed(-3303.0/65536.0,1,-nbitq), 
to_sfixed(-10552.0/65536.0,1,-nbitq), 
to_sfixed(-1381.0/65536.0,1,-nbitq), 
to_sfixed(5003.0/65536.0,1,-nbitq), 
to_sfixed(3033.0/65536.0,1,-nbitq), 
to_sfixed(17591.0/65536.0,1,-nbitq), 
to_sfixed(1309.0/65536.0,1,-nbitq), 
to_sfixed(4329.0/65536.0,1,-nbitq), 
to_sfixed(-5778.0/65536.0,1,-nbitq), 
to_sfixed(-4901.0/65536.0,1,-nbitq), 
to_sfixed(1847.0/65536.0,1,-nbitq), 
to_sfixed(1969.0/65536.0,1,-nbitq), 
to_sfixed(-2199.0/65536.0,1,-nbitq), 
to_sfixed(1520.0/65536.0,1,-nbitq), 
to_sfixed(2342.0/65536.0,1,-nbitq), 
to_sfixed(7018.0/65536.0,1,-nbitq), 
to_sfixed(4601.0/65536.0,1,-nbitq), 
to_sfixed(1726.0/65536.0,1,-nbitq), 
to_sfixed(-2197.0/65536.0,1,-nbitq), 
to_sfixed(8170.0/65536.0,1,-nbitq), 
to_sfixed(-6418.0/65536.0,1,-nbitq), 
to_sfixed(-19983.0/65536.0,1,-nbitq), 
to_sfixed(-5874.0/65536.0,1,-nbitq), 
to_sfixed(-5094.0/65536.0,1,-nbitq), 
to_sfixed(-2671.0/65536.0,1,-nbitq), 
to_sfixed(-8317.0/65536.0,1,-nbitq), 
to_sfixed(-4333.0/65536.0,1,-nbitq), 
to_sfixed(-1194.0/65536.0,1,-nbitq), 
to_sfixed(11285.0/65536.0,1,-nbitq), 
to_sfixed(-3465.0/65536.0,1,-nbitq), 
to_sfixed(-1927.0/65536.0,1,-nbitq), 
to_sfixed(1381.0/65536.0,1,-nbitq), 
to_sfixed(-3334.0/65536.0,1,-nbitq), 
to_sfixed(1708.0/65536.0,1,-nbitq), 
to_sfixed(-1761.0/65536.0,1,-nbitq), 
to_sfixed(1653.0/65536.0,1,-nbitq), 
to_sfixed(-1888.0/65536.0,1,-nbitq), 
to_sfixed(-1317.0/65536.0,1,-nbitq), 
to_sfixed(1952.0/65536.0,1,-nbitq), 
to_sfixed(2209.0/65536.0,1,-nbitq), 
to_sfixed(-3428.0/65536.0,1,-nbitq), 
to_sfixed(-350.0/65536.0,1,-nbitq), 
to_sfixed(-5003.0/65536.0,1,-nbitq), 
to_sfixed(3961.0/65536.0,1,-nbitq), 
to_sfixed(-2375.0/65536.0,1,-nbitq), 
to_sfixed(1096.0/65536.0,1,-nbitq), 
to_sfixed(1425.0/65536.0,1,-nbitq), 
to_sfixed(-16107.0/65536.0,1,-nbitq), 
to_sfixed(-8383.0/65536.0,1,-nbitq), 
to_sfixed(-5431.0/65536.0,1,-nbitq), 
to_sfixed(-5982.0/65536.0,1,-nbitq), 
to_sfixed(-12027.0/65536.0,1,-nbitq), 
to_sfixed(1794.0/65536.0,1,-nbitq), 
to_sfixed(97.0/65536.0,1,-nbitq), 
to_sfixed(5136.0/65536.0,1,-nbitq), 
to_sfixed(-5835.0/65536.0,1,-nbitq), 
to_sfixed(254.0/65536.0,1,-nbitq), 
to_sfixed(1453.0/65536.0,1,-nbitq), 
to_sfixed(-7894.0/65536.0,1,-nbitq), 
to_sfixed(1343.0/65536.0,1,-nbitq), 
to_sfixed(8936.0/65536.0,1,-nbitq), 
to_sfixed(-2082.0/65536.0,1,-nbitq), 
to_sfixed(-10057.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5159.0/65536.0,1,-nbitq), 
to_sfixed(-2936.0/65536.0,1,-nbitq), 
to_sfixed(-12868.0/65536.0,1,-nbitq), 
to_sfixed(8264.0/65536.0,1,-nbitq), 
to_sfixed(-933.0/65536.0,1,-nbitq), 
to_sfixed(-10536.0/65536.0,1,-nbitq), 
to_sfixed(2138.0/65536.0,1,-nbitq), 
to_sfixed(-5507.0/65536.0,1,-nbitq), 
to_sfixed(-4006.0/65536.0,1,-nbitq), 
to_sfixed(263.0/65536.0,1,-nbitq), 
to_sfixed(9700.0/65536.0,1,-nbitq), 
to_sfixed(10780.0/65536.0,1,-nbitq), 
to_sfixed(1061.0/65536.0,1,-nbitq), 
to_sfixed(-8576.0/65536.0,1,-nbitq), 
to_sfixed(-8058.0/65536.0,1,-nbitq), 
to_sfixed(-1882.0/65536.0,1,-nbitq), 
to_sfixed(9.0/65536.0,1,-nbitq), 
to_sfixed(-2012.0/65536.0,1,-nbitq), 
to_sfixed(1642.0/65536.0,1,-nbitq), 
to_sfixed(-1870.0/65536.0,1,-nbitq), 
to_sfixed(5655.0/65536.0,1,-nbitq), 
to_sfixed(5077.0/65536.0,1,-nbitq), 
to_sfixed(10727.0/65536.0,1,-nbitq), 
to_sfixed(666.0/65536.0,1,-nbitq), 
to_sfixed(2550.0/65536.0,1,-nbitq), 
to_sfixed(-8097.0/65536.0,1,-nbitq), 
to_sfixed(-7987.0/65536.0,1,-nbitq), 
to_sfixed(-1066.0/65536.0,1,-nbitq), 
to_sfixed(293.0/65536.0,1,-nbitq), 
to_sfixed(399.0/65536.0,1,-nbitq), 
to_sfixed(251.0/65536.0,1,-nbitq), 
to_sfixed(-393.0/65536.0,1,-nbitq), 
to_sfixed(10868.0/65536.0,1,-nbitq), 
to_sfixed(6089.0/65536.0,1,-nbitq), 
to_sfixed(-2319.0/65536.0,1,-nbitq), 
to_sfixed(2760.0/65536.0,1,-nbitq), 
to_sfixed(-480.0/65536.0,1,-nbitq), 
to_sfixed(600.0/65536.0,1,-nbitq), 
to_sfixed(-12009.0/65536.0,1,-nbitq), 
to_sfixed(-6133.0/65536.0,1,-nbitq), 
to_sfixed(-6310.0/65536.0,1,-nbitq), 
to_sfixed(1484.0/65536.0,1,-nbitq), 
to_sfixed(-8715.0/65536.0,1,-nbitq), 
to_sfixed(1059.0/65536.0,1,-nbitq), 
to_sfixed(-1368.0/65536.0,1,-nbitq), 
to_sfixed(8220.0/65536.0,1,-nbitq), 
to_sfixed(953.0/65536.0,1,-nbitq), 
to_sfixed(2613.0/65536.0,1,-nbitq), 
to_sfixed(931.0/65536.0,1,-nbitq), 
to_sfixed(2695.0/65536.0,1,-nbitq), 
to_sfixed(-2356.0/65536.0,1,-nbitq), 
to_sfixed(10488.0/65536.0,1,-nbitq), 
to_sfixed(621.0/65536.0,1,-nbitq), 
to_sfixed(9602.0/65536.0,1,-nbitq), 
to_sfixed(-1482.0/65536.0,1,-nbitq), 
to_sfixed(-277.0/65536.0,1,-nbitq), 
to_sfixed(405.0/65536.0,1,-nbitq), 
to_sfixed(-5109.0/65536.0,1,-nbitq), 
to_sfixed(167.0/65536.0,1,-nbitq), 
to_sfixed(-952.0/65536.0,1,-nbitq), 
to_sfixed(-2158.0/65536.0,1,-nbitq), 
to_sfixed(80.0/65536.0,1,-nbitq), 
to_sfixed(-1879.0/65536.0,1,-nbitq), 
to_sfixed(1736.0/65536.0,1,-nbitq), 
to_sfixed(-12732.0/65536.0,1,-nbitq), 
to_sfixed(-5994.0/65536.0,1,-nbitq), 
to_sfixed(-10799.0/65536.0,1,-nbitq), 
to_sfixed(-3142.0/65536.0,1,-nbitq), 
to_sfixed(-11030.0/65536.0,1,-nbitq), 
to_sfixed(6377.0/65536.0,1,-nbitq), 
to_sfixed(-1107.0/65536.0,1,-nbitq), 
to_sfixed(-1175.0/65536.0,1,-nbitq), 
to_sfixed(-10605.0/65536.0,1,-nbitq), 
to_sfixed(2204.0/65536.0,1,-nbitq), 
to_sfixed(2426.0/65536.0,1,-nbitq), 
to_sfixed(-9239.0/65536.0,1,-nbitq), 
to_sfixed(-8013.0/65536.0,1,-nbitq), 
to_sfixed(5561.0/65536.0,1,-nbitq), 
to_sfixed(-1416.0/65536.0,1,-nbitq), 
to_sfixed(-910.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4868.0/65536.0,1,-nbitq), 
to_sfixed(-3407.0/65536.0,1,-nbitq), 
to_sfixed(2522.0/65536.0,1,-nbitq), 
to_sfixed(-5878.0/65536.0,1,-nbitq), 
to_sfixed(-8137.0/65536.0,1,-nbitq), 
to_sfixed(-4167.0/65536.0,1,-nbitq), 
to_sfixed(1089.0/65536.0,1,-nbitq), 
to_sfixed(-10612.0/65536.0,1,-nbitq), 
to_sfixed(-3756.0/65536.0,1,-nbitq), 
to_sfixed(-1767.0/65536.0,1,-nbitq), 
to_sfixed(5789.0/65536.0,1,-nbitq), 
to_sfixed(7525.0/65536.0,1,-nbitq), 
to_sfixed(-1584.0/65536.0,1,-nbitq), 
to_sfixed(-14616.0/65536.0,1,-nbitq), 
to_sfixed(-986.0/65536.0,1,-nbitq), 
to_sfixed(23.0/65536.0,1,-nbitq), 
to_sfixed(2654.0/65536.0,1,-nbitq), 
to_sfixed(-3645.0/65536.0,1,-nbitq), 
to_sfixed(5587.0/65536.0,1,-nbitq), 
to_sfixed(1624.0/65536.0,1,-nbitq), 
to_sfixed(11497.0/65536.0,1,-nbitq), 
to_sfixed(-8734.0/65536.0,1,-nbitq), 
to_sfixed(-9013.0/65536.0,1,-nbitq), 
to_sfixed(-1416.0/65536.0,1,-nbitq), 
to_sfixed(-460.0/65536.0,1,-nbitq), 
to_sfixed(1940.0/65536.0,1,-nbitq), 
to_sfixed(-1385.0/65536.0,1,-nbitq), 
to_sfixed(2436.0/65536.0,1,-nbitq), 
to_sfixed(6378.0/65536.0,1,-nbitq), 
to_sfixed(-2197.0/65536.0,1,-nbitq), 
to_sfixed(-1985.0/65536.0,1,-nbitq), 
to_sfixed(6692.0/65536.0,1,-nbitq), 
to_sfixed(-2271.0/65536.0,1,-nbitq), 
to_sfixed(2656.0/65536.0,1,-nbitq), 
to_sfixed(959.0/65536.0,1,-nbitq), 
to_sfixed(-1059.0/65536.0,1,-nbitq), 
to_sfixed(1611.0/65536.0,1,-nbitq), 
to_sfixed(3521.0/65536.0,1,-nbitq), 
to_sfixed(13253.0/65536.0,1,-nbitq), 
to_sfixed(-1438.0/65536.0,1,-nbitq), 
to_sfixed(-3583.0/65536.0,1,-nbitq), 
to_sfixed(1918.0/65536.0,1,-nbitq), 
to_sfixed(-9331.0/65536.0,1,-nbitq), 
to_sfixed(1694.0/65536.0,1,-nbitq), 
to_sfixed(396.0/65536.0,1,-nbitq), 
to_sfixed(1276.0/65536.0,1,-nbitq), 
to_sfixed(-1880.0/65536.0,1,-nbitq), 
to_sfixed(1012.0/65536.0,1,-nbitq), 
to_sfixed(-1846.0/65536.0,1,-nbitq), 
to_sfixed(-1096.0/65536.0,1,-nbitq), 
to_sfixed(292.0/65536.0,1,-nbitq), 
to_sfixed(23096.0/65536.0,1,-nbitq), 
to_sfixed(-4979.0/65536.0,1,-nbitq), 
to_sfixed(1422.0/65536.0,1,-nbitq), 
to_sfixed(-6135.0/65536.0,1,-nbitq), 
to_sfixed(2576.0/65536.0,1,-nbitq), 
to_sfixed(363.0/65536.0,1,-nbitq), 
to_sfixed(-64.0/65536.0,1,-nbitq), 
to_sfixed(-2600.0/65536.0,1,-nbitq), 
to_sfixed(130.0/65536.0,1,-nbitq), 
to_sfixed(-5674.0/65536.0,1,-nbitq), 
to_sfixed(1293.0/65536.0,1,-nbitq), 
to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(-787.0/65536.0,1,-nbitq), 
to_sfixed(-9304.0/65536.0,1,-nbitq), 
to_sfixed(-5113.0/65536.0,1,-nbitq), 
to_sfixed(-8643.0/65536.0,1,-nbitq), 
to_sfixed(-2401.0/65536.0,1,-nbitq), 
to_sfixed(-9456.0/65536.0,1,-nbitq), 
to_sfixed(-2189.0/65536.0,1,-nbitq), 
to_sfixed(-1759.0/65536.0,1,-nbitq), 
to_sfixed(-4438.0/65536.0,1,-nbitq), 
to_sfixed(-13564.0/65536.0,1,-nbitq), 
to_sfixed(-3047.0/65536.0,1,-nbitq), 
to_sfixed(-364.0/65536.0,1,-nbitq), 
to_sfixed(-7016.0/65536.0,1,-nbitq), 
to_sfixed(-5574.0/65536.0,1,-nbitq), 
to_sfixed(1967.0/65536.0,1,-nbitq), 
to_sfixed(2633.0/65536.0,1,-nbitq), 
to_sfixed(12704.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2064.0/65536.0,1,-nbitq), 
to_sfixed(-2401.0/65536.0,1,-nbitq), 
to_sfixed(14599.0/65536.0,1,-nbitq), 
to_sfixed(-9372.0/65536.0,1,-nbitq), 
to_sfixed(-2936.0/65536.0,1,-nbitq), 
to_sfixed(13771.0/65536.0,1,-nbitq), 
to_sfixed(-52.0/65536.0,1,-nbitq), 
to_sfixed(-3935.0/65536.0,1,-nbitq), 
to_sfixed(9912.0/65536.0,1,-nbitq), 
to_sfixed(-2491.0/65536.0,1,-nbitq), 
to_sfixed(6740.0/65536.0,1,-nbitq), 
to_sfixed(-4665.0/65536.0,1,-nbitq), 
to_sfixed(-2962.0/65536.0,1,-nbitq), 
to_sfixed(-7715.0/65536.0,1,-nbitq), 
to_sfixed(-291.0/65536.0,1,-nbitq), 
to_sfixed(-1858.0/65536.0,1,-nbitq), 
to_sfixed(-2102.0/65536.0,1,-nbitq), 
to_sfixed(-1514.0/65536.0,1,-nbitq), 
to_sfixed(4130.0/65536.0,1,-nbitq), 
to_sfixed(1809.0/65536.0,1,-nbitq), 
to_sfixed(10638.0/65536.0,1,-nbitq), 
to_sfixed(-7290.0/65536.0,1,-nbitq), 
to_sfixed(-17155.0/65536.0,1,-nbitq), 
to_sfixed(5624.0/65536.0,1,-nbitq), 
to_sfixed(-3965.0/65536.0,1,-nbitq), 
to_sfixed(4124.0/65536.0,1,-nbitq), 
to_sfixed(4257.0/65536.0,1,-nbitq), 
to_sfixed(-257.0/65536.0,1,-nbitq), 
to_sfixed(2359.0/65536.0,1,-nbitq), 
to_sfixed(2728.0/65536.0,1,-nbitq), 
to_sfixed(-5040.0/65536.0,1,-nbitq), 
to_sfixed(1117.0/65536.0,1,-nbitq), 
to_sfixed(-11786.0/65536.0,1,-nbitq), 
to_sfixed(1498.0/65536.0,1,-nbitq), 
to_sfixed(-439.0/65536.0,1,-nbitq), 
to_sfixed(1209.0/65536.0,1,-nbitq), 
to_sfixed(6956.0/65536.0,1,-nbitq), 
to_sfixed(6765.0/65536.0,1,-nbitq), 
to_sfixed(7521.0/65536.0,1,-nbitq), 
to_sfixed(1593.0/65536.0,1,-nbitq), 
to_sfixed(-6833.0/65536.0,1,-nbitq), 
to_sfixed(-253.0/65536.0,1,-nbitq), 
to_sfixed(-9216.0/65536.0,1,-nbitq), 
to_sfixed(3825.0/65536.0,1,-nbitq), 
to_sfixed(-1276.0/65536.0,1,-nbitq), 
to_sfixed(-6472.0/65536.0,1,-nbitq), 
to_sfixed(1307.0/65536.0,1,-nbitq), 
to_sfixed(3915.0/65536.0,1,-nbitq), 
to_sfixed(-1463.0/65536.0,1,-nbitq), 
to_sfixed(-859.0/65536.0,1,-nbitq), 
to_sfixed(-1445.0/65536.0,1,-nbitq), 
to_sfixed(19427.0/65536.0,1,-nbitq), 
to_sfixed(-8277.0/65536.0,1,-nbitq), 
to_sfixed(8950.0/65536.0,1,-nbitq), 
to_sfixed(-560.0/65536.0,1,-nbitq), 
to_sfixed(-17542.0/65536.0,1,-nbitq), 
to_sfixed(-3514.0/65536.0,1,-nbitq), 
to_sfixed(4944.0/65536.0,1,-nbitq), 
to_sfixed(-1679.0/65536.0,1,-nbitq), 
to_sfixed(-1528.0/65536.0,1,-nbitq), 
to_sfixed(-3335.0/65536.0,1,-nbitq), 
to_sfixed(1485.0/65536.0,1,-nbitq), 
to_sfixed(949.0/65536.0,1,-nbitq), 
to_sfixed(-1097.0/65536.0,1,-nbitq), 
to_sfixed(-2929.0/65536.0,1,-nbitq), 
to_sfixed(-4723.0/65536.0,1,-nbitq), 
to_sfixed(-9449.0/65536.0,1,-nbitq), 
to_sfixed(-4860.0/65536.0,1,-nbitq), 
to_sfixed(-4413.0/65536.0,1,-nbitq), 
to_sfixed(-1452.0/65536.0,1,-nbitq), 
to_sfixed(-5379.0/65536.0,1,-nbitq), 
to_sfixed(-3110.0/65536.0,1,-nbitq), 
to_sfixed(-147.0/65536.0,1,-nbitq), 
to_sfixed(-1174.0/65536.0,1,-nbitq), 
to_sfixed(2501.0/65536.0,1,-nbitq), 
to_sfixed(6.0/65536.0,1,-nbitq), 
to_sfixed(1788.0/65536.0,1,-nbitq), 
to_sfixed(12149.0/65536.0,1,-nbitq), 
to_sfixed(-1372.0/65536.0,1,-nbitq), 
to_sfixed(14712.0/65536.0,1,-nbitq)  ), 
( to_sfixed(573.0/65536.0,1,-nbitq), 
to_sfixed(225.0/65536.0,1,-nbitq), 
to_sfixed(5958.0/65536.0,1,-nbitq), 
to_sfixed(-6342.0/65536.0,1,-nbitq), 
to_sfixed(771.0/65536.0,1,-nbitq), 
to_sfixed(20169.0/65536.0,1,-nbitq), 
to_sfixed(3622.0/65536.0,1,-nbitq), 
to_sfixed(514.0/65536.0,1,-nbitq), 
to_sfixed(13203.0/65536.0,1,-nbitq), 
to_sfixed(1572.0/65536.0,1,-nbitq), 
to_sfixed(8849.0/65536.0,1,-nbitq), 
to_sfixed(-1655.0/65536.0,1,-nbitq), 
to_sfixed(-536.0/65536.0,1,-nbitq), 
to_sfixed(-3244.0/65536.0,1,-nbitq), 
to_sfixed(2086.0/65536.0,1,-nbitq), 
to_sfixed(201.0/65536.0,1,-nbitq), 
to_sfixed(1488.0/65536.0,1,-nbitq), 
to_sfixed(-127.0/65536.0,1,-nbitq), 
to_sfixed(2578.0/65536.0,1,-nbitq), 
to_sfixed(-2154.0/65536.0,1,-nbitq), 
to_sfixed(6233.0/65536.0,1,-nbitq), 
to_sfixed(-18169.0/65536.0,1,-nbitq), 
to_sfixed(3710.0/65536.0,1,-nbitq), 
to_sfixed(10554.0/65536.0,1,-nbitq), 
to_sfixed(1314.0/65536.0,1,-nbitq), 
to_sfixed(5413.0/65536.0,1,-nbitq), 
to_sfixed(2878.0/65536.0,1,-nbitq), 
to_sfixed(-711.0/65536.0,1,-nbitq), 
to_sfixed(-3264.0/65536.0,1,-nbitq), 
to_sfixed(3198.0/65536.0,1,-nbitq), 
to_sfixed(-3100.0/65536.0,1,-nbitq), 
to_sfixed(-1984.0/65536.0,1,-nbitq), 
to_sfixed(-15328.0/65536.0,1,-nbitq), 
to_sfixed(3490.0/65536.0,1,-nbitq), 
to_sfixed(-2026.0/65536.0,1,-nbitq), 
to_sfixed(1374.0/65536.0,1,-nbitq), 
to_sfixed(5079.0/65536.0,1,-nbitq), 
to_sfixed(2118.0/65536.0,1,-nbitq), 
to_sfixed(1650.0/65536.0,1,-nbitq), 
to_sfixed(-3018.0/65536.0,1,-nbitq), 
to_sfixed(-13066.0/65536.0,1,-nbitq), 
to_sfixed(-97.0/65536.0,1,-nbitq), 
to_sfixed(-1939.0/65536.0,1,-nbitq), 
to_sfixed(-4567.0/65536.0,1,-nbitq), 
to_sfixed(-2067.0/65536.0,1,-nbitq), 
to_sfixed(-3709.0/65536.0,1,-nbitq), 
to_sfixed(-3539.0/65536.0,1,-nbitq), 
to_sfixed(7572.0/65536.0,1,-nbitq), 
to_sfixed(1299.0/65536.0,1,-nbitq), 
to_sfixed(477.0/65536.0,1,-nbitq), 
to_sfixed(167.0/65536.0,1,-nbitq), 
to_sfixed(6888.0/65536.0,1,-nbitq), 
to_sfixed(-3804.0/65536.0,1,-nbitq), 
to_sfixed(3365.0/65536.0,1,-nbitq), 
to_sfixed(4442.0/65536.0,1,-nbitq), 
to_sfixed(-13683.0/65536.0,1,-nbitq), 
to_sfixed(146.0/65536.0,1,-nbitq), 
to_sfixed(-458.0/65536.0,1,-nbitq), 
to_sfixed(-1032.0/65536.0,1,-nbitq), 
to_sfixed(3118.0/65536.0,1,-nbitq), 
to_sfixed(2080.0/65536.0,1,-nbitq), 
to_sfixed(1110.0/65536.0,1,-nbitq), 
to_sfixed(-1863.0/65536.0,1,-nbitq), 
to_sfixed(-1519.0/65536.0,1,-nbitq), 
to_sfixed(3050.0/65536.0,1,-nbitq), 
to_sfixed(-2758.0/65536.0,1,-nbitq), 
to_sfixed(-6741.0/65536.0,1,-nbitq), 
to_sfixed(6734.0/65536.0,1,-nbitq), 
to_sfixed(-6428.0/65536.0,1,-nbitq), 
to_sfixed(-6056.0/65536.0,1,-nbitq), 
to_sfixed(-6939.0/65536.0,1,-nbitq), 
to_sfixed(2373.0/65536.0,1,-nbitq), 
to_sfixed(15817.0/65536.0,1,-nbitq), 
to_sfixed(-500.0/65536.0,1,-nbitq), 
to_sfixed(1816.0/65536.0,1,-nbitq), 
to_sfixed(2894.0/65536.0,1,-nbitq), 
to_sfixed(-1603.0/65536.0,1,-nbitq), 
to_sfixed(8961.0/65536.0,1,-nbitq), 
to_sfixed(-676.0/65536.0,1,-nbitq), 
to_sfixed(9358.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2003.0/65536.0,1,-nbitq), 
to_sfixed(5271.0/65536.0,1,-nbitq), 
to_sfixed(-5728.0/65536.0,1,-nbitq), 
to_sfixed(-641.0/65536.0,1,-nbitq), 
to_sfixed(-7595.0/65536.0,1,-nbitq), 
to_sfixed(8440.0/65536.0,1,-nbitq), 
to_sfixed(4175.0/65536.0,1,-nbitq), 
to_sfixed(1448.0/65536.0,1,-nbitq), 
to_sfixed(16423.0/65536.0,1,-nbitq), 
to_sfixed(209.0/65536.0,1,-nbitq), 
to_sfixed(8068.0/65536.0,1,-nbitq), 
to_sfixed(5825.0/65536.0,1,-nbitq), 
to_sfixed(1143.0/65536.0,1,-nbitq), 
to_sfixed(-850.0/65536.0,1,-nbitq), 
to_sfixed(-1220.0/65536.0,1,-nbitq), 
to_sfixed(-1543.0/65536.0,1,-nbitq), 
to_sfixed(2316.0/65536.0,1,-nbitq), 
to_sfixed(-1095.0/65536.0,1,-nbitq), 
to_sfixed(-6144.0/65536.0,1,-nbitq), 
to_sfixed(-2204.0/65536.0,1,-nbitq), 
to_sfixed(14665.0/65536.0,1,-nbitq), 
to_sfixed(-15816.0/65536.0,1,-nbitq), 
to_sfixed(9185.0/65536.0,1,-nbitq), 
to_sfixed(12480.0/65536.0,1,-nbitq), 
to_sfixed(-4001.0/65536.0,1,-nbitq), 
to_sfixed(4376.0/65536.0,1,-nbitq), 
to_sfixed(4085.0/65536.0,1,-nbitq), 
to_sfixed(493.0/65536.0,1,-nbitq), 
to_sfixed(-7200.0/65536.0,1,-nbitq), 
to_sfixed(772.0/65536.0,1,-nbitq), 
to_sfixed(-1766.0/65536.0,1,-nbitq), 
to_sfixed(-5963.0/65536.0,1,-nbitq), 
to_sfixed(-5728.0/65536.0,1,-nbitq), 
to_sfixed(2614.0/65536.0,1,-nbitq), 
to_sfixed(1617.0/65536.0,1,-nbitq), 
to_sfixed(-2661.0/65536.0,1,-nbitq), 
to_sfixed(8336.0/65536.0,1,-nbitq), 
to_sfixed(-4236.0/65536.0,1,-nbitq), 
to_sfixed(4431.0/65536.0,1,-nbitq), 
to_sfixed(933.0/65536.0,1,-nbitq), 
to_sfixed(-7937.0/65536.0,1,-nbitq), 
to_sfixed(2761.0/65536.0,1,-nbitq), 
to_sfixed(5486.0/65536.0,1,-nbitq), 
to_sfixed(-4530.0/65536.0,1,-nbitq), 
to_sfixed(-2067.0/65536.0,1,-nbitq), 
to_sfixed(-11034.0/65536.0,1,-nbitq), 
to_sfixed(-2000.0/65536.0,1,-nbitq), 
to_sfixed(7902.0/65536.0,1,-nbitq), 
to_sfixed(-371.0/65536.0,1,-nbitq), 
to_sfixed(-1308.0/65536.0,1,-nbitq), 
to_sfixed(3003.0/65536.0,1,-nbitq), 
to_sfixed(-5294.0/65536.0,1,-nbitq), 
to_sfixed(-1350.0/65536.0,1,-nbitq), 
to_sfixed(200.0/65536.0,1,-nbitq), 
to_sfixed(6144.0/65536.0,1,-nbitq), 
to_sfixed(-4660.0/65536.0,1,-nbitq), 
to_sfixed(1068.0/65536.0,1,-nbitq), 
to_sfixed(404.0/65536.0,1,-nbitq), 
to_sfixed(2335.0/65536.0,1,-nbitq), 
to_sfixed(-4476.0/65536.0,1,-nbitq), 
to_sfixed(2346.0/65536.0,1,-nbitq), 
to_sfixed(1234.0/65536.0,1,-nbitq), 
to_sfixed(1695.0/65536.0,1,-nbitq), 
to_sfixed(-2272.0/65536.0,1,-nbitq), 
to_sfixed(4449.0/65536.0,1,-nbitq), 
to_sfixed(-3103.0/65536.0,1,-nbitq), 
to_sfixed(-2450.0/65536.0,1,-nbitq), 
to_sfixed(2820.0/65536.0,1,-nbitq), 
to_sfixed(-5724.0/65536.0,1,-nbitq), 
to_sfixed(-5908.0/65536.0,1,-nbitq), 
to_sfixed(-6279.0/65536.0,1,-nbitq), 
to_sfixed(5847.0/65536.0,1,-nbitq), 
to_sfixed(17070.0/65536.0,1,-nbitq), 
to_sfixed(1860.0/65536.0,1,-nbitq), 
to_sfixed(-1887.0/65536.0,1,-nbitq), 
to_sfixed(1165.0/65536.0,1,-nbitq), 
to_sfixed(-2222.0/65536.0,1,-nbitq), 
to_sfixed(493.0/65536.0,1,-nbitq), 
to_sfixed(-795.0/65536.0,1,-nbitq), 
to_sfixed(6818.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2599.0/65536.0,1,-nbitq), 
to_sfixed(215.0/65536.0,1,-nbitq), 
to_sfixed(1351.0/65536.0,1,-nbitq), 
to_sfixed(-1852.0/65536.0,1,-nbitq), 
to_sfixed(7188.0/65536.0,1,-nbitq), 
to_sfixed(6087.0/65536.0,1,-nbitq), 
to_sfixed(1545.0/65536.0,1,-nbitq), 
to_sfixed(2718.0/65536.0,1,-nbitq), 
to_sfixed(11270.0/65536.0,1,-nbitq), 
to_sfixed(1488.0/65536.0,1,-nbitq), 
to_sfixed(2126.0/65536.0,1,-nbitq), 
to_sfixed(3632.0/65536.0,1,-nbitq), 
to_sfixed(1589.0/65536.0,1,-nbitq), 
to_sfixed(9325.0/65536.0,1,-nbitq), 
to_sfixed(2970.0/65536.0,1,-nbitq), 
to_sfixed(-2668.0/65536.0,1,-nbitq), 
to_sfixed(-2851.0/65536.0,1,-nbitq), 
to_sfixed(-1569.0/65536.0,1,-nbitq), 
to_sfixed(-3260.0/65536.0,1,-nbitq), 
to_sfixed(216.0/65536.0,1,-nbitq), 
to_sfixed(11517.0/65536.0,1,-nbitq), 
to_sfixed(-5400.0/65536.0,1,-nbitq), 
to_sfixed(2199.0/65536.0,1,-nbitq), 
to_sfixed(9123.0/65536.0,1,-nbitq), 
to_sfixed(-1496.0/65536.0,1,-nbitq), 
to_sfixed(520.0/65536.0,1,-nbitq), 
to_sfixed(3854.0/65536.0,1,-nbitq), 
to_sfixed(-515.0/65536.0,1,-nbitq), 
to_sfixed(-6472.0/65536.0,1,-nbitq), 
to_sfixed(-1443.0/65536.0,1,-nbitq), 
to_sfixed(-2853.0/65536.0,1,-nbitq), 
to_sfixed(-6126.0/65536.0,1,-nbitq), 
to_sfixed(-5050.0/65536.0,1,-nbitq), 
to_sfixed(2579.0/65536.0,1,-nbitq), 
to_sfixed(-1406.0/65536.0,1,-nbitq), 
to_sfixed(-1783.0/65536.0,1,-nbitq), 
to_sfixed(8104.0/65536.0,1,-nbitq), 
to_sfixed(-1709.0/65536.0,1,-nbitq), 
to_sfixed(5744.0/65536.0,1,-nbitq), 
to_sfixed(-627.0/65536.0,1,-nbitq), 
to_sfixed(-2029.0/65536.0,1,-nbitq), 
to_sfixed(1201.0/65536.0,1,-nbitq), 
to_sfixed(9955.0/65536.0,1,-nbitq), 
to_sfixed(944.0/65536.0,1,-nbitq), 
to_sfixed(1020.0/65536.0,1,-nbitq), 
to_sfixed(-12210.0/65536.0,1,-nbitq), 
to_sfixed(-593.0/65536.0,1,-nbitq), 
to_sfixed(794.0/65536.0,1,-nbitq), 
to_sfixed(-1897.0/65536.0,1,-nbitq), 
to_sfixed(-1793.0/65536.0,1,-nbitq), 
to_sfixed(-1539.0/65536.0,1,-nbitq), 
to_sfixed(-5933.0/65536.0,1,-nbitq), 
to_sfixed(-2250.0/65536.0,1,-nbitq), 
to_sfixed(2865.0/65536.0,1,-nbitq), 
to_sfixed(5558.0/65536.0,1,-nbitq), 
to_sfixed(-3394.0/65536.0,1,-nbitq), 
to_sfixed(1179.0/65536.0,1,-nbitq), 
to_sfixed(-3817.0/65536.0,1,-nbitq), 
to_sfixed(409.0/65536.0,1,-nbitq), 
to_sfixed(-4626.0/65536.0,1,-nbitq), 
to_sfixed(-1086.0/65536.0,1,-nbitq), 
to_sfixed(969.0/65536.0,1,-nbitq), 
to_sfixed(-39.0/65536.0,1,-nbitq), 
to_sfixed(-3028.0/65536.0,1,-nbitq), 
to_sfixed(409.0/65536.0,1,-nbitq), 
to_sfixed(-1260.0/65536.0,1,-nbitq), 
to_sfixed(547.0/65536.0,1,-nbitq), 
to_sfixed(7603.0/65536.0,1,-nbitq), 
to_sfixed(-6180.0/65536.0,1,-nbitq), 
to_sfixed(-2074.0/65536.0,1,-nbitq), 
to_sfixed(-2063.0/65536.0,1,-nbitq), 
to_sfixed(7930.0/65536.0,1,-nbitq), 
to_sfixed(7259.0/65536.0,1,-nbitq), 
to_sfixed(-2989.0/65536.0,1,-nbitq), 
to_sfixed(762.0/65536.0,1,-nbitq), 
to_sfixed(3676.0/65536.0,1,-nbitq), 
to_sfixed(-6074.0/65536.0,1,-nbitq), 
to_sfixed(-10814.0/65536.0,1,-nbitq), 
to_sfixed(2320.0/65536.0,1,-nbitq), 
to_sfixed(954.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2323.0/65536.0,1,-nbitq), 
to_sfixed(641.0/65536.0,1,-nbitq), 
to_sfixed(3747.0/65536.0,1,-nbitq), 
to_sfixed(-4325.0/65536.0,1,-nbitq), 
to_sfixed(15583.0/65536.0,1,-nbitq), 
to_sfixed(6998.0/65536.0,1,-nbitq), 
to_sfixed(-1314.0/65536.0,1,-nbitq), 
to_sfixed(3794.0/65536.0,1,-nbitq), 
to_sfixed(3485.0/65536.0,1,-nbitq), 
to_sfixed(-2086.0/65536.0,1,-nbitq), 
to_sfixed(5172.0/65536.0,1,-nbitq), 
to_sfixed(-567.0/65536.0,1,-nbitq), 
to_sfixed(-3339.0/65536.0,1,-nbitq), 
to_sfixed(12838.0/65536.0,1,-nbitq), 
to_sfixed(4017.0/65536.0,1,-nbitq), 
to_sfixed(2907.0/65536.0,1,-nbitq), 
to_sfixed(2314.0/65536.0,1,-nbitq), 
to_sfixed(-4004.0/65536.0,1,-nbitq), 
to_sfixed(3594.0/65536.0,1,-nbitq), 
to_sfixed(-1636.0/65536.0,1,-nbitq), 
to_sfixed(8190.0/65536.0,1,-nbitq), 
to_sfixed(-11231.0/65536.0,1,-nbitq), 
to_sfixed(-2595.0/65536.0,1,-nbitq), 
to_sfixed(9896.0/65536.0,1,-nbitq), 
to_sfixed(-2232.0/65536.0,1,-nbitq), 
to_sfixed(1939.0/65536.0,1,-nbitq), 
to_sfixed(6559.0/65536.0,1,-nbitq), 
to_sfixed(3813.0/65536.0,1,-nbitq), 
to_sfixed(-6669.0/65536.0,1,-nbitq), 
to_sfixed(-1549.0/65536.0,1,-nbitq), 
to_sfixed(-2074.0/65536.0,1,-nbitq), 
to_sfixed(-2118.0/65536.0,1,-nbitq), 
to_sfixed(361.0/65536.0,1,-nbitq), 
to_sfixed(8016.0/65536.0,1,-nbitq), 
to_sfixed(-1729.0/65536.0,1,-nbitq), 
to_sfixed(-2514.0/65536.0,1,-nbitq), 
to_sfixed(9243.0/65536.0,1,-nbitq), 
to_sfixed(1307.0/65536.0,1,-nbitq), 
to_sfixed(8997.0/65536.0,1,-nbitq), 
to_sfixed(-3180.0/65536.0,1,-nbitq), 
to_sfixed(749.0/65536.0,1,-nbitq), 
to_sfixed(-1898.0/65536.0,1,-nbitq), 
to_sfixed(10820.0/65536.0,1,-nbitq), 
to_sfixed(-1960.0/65536.0,1,-nbitq), 
to_sfixed(257.0/65536.0,1,-nbitq), 
to_sfixed(-3313.0/65536.0,1,-nbitq), 
to_sfixed(-2420.0/65536.0,1,-nbitq), 
to_sfixed(-2171.0/65536.0,1,-nbitq), 
to_sfixed(-2111.0/65536.0,1,-nbitq), 
to_sfixed(-2732.0/65536.0,1,-nbitq), 
to_sfixed(406.0/65536.0,1,-nbitq), 
to_sfixed(910.0/65536.0,1,-nbitq), 
to_sfixed(-4187.0/65536.0,1,-nbitq), 
to_sfixed(-2462.0/65536.0,1,-nbitq), 
to_sfixed(-273.0/65536.0,1,-nbitq), 
to_sfixed(5927.0/65536.0,1,-nbitq), 
to_sfixed(-524.0/65536.0,1,-nbitq), 
to_sfixed(-13.0/65536.0,1,-nbitq), 
to_sfixed(-3038.0/65536.0,1,-nbitq), 
to_sfixed(-9860.0/65536.0,1,-nbitq), 
to_sfixed(2592.0/65536.0,1,-nbitq), 
to_sfixed(-1915.0/65536.0,1,-nbitq), 
to_sfixed(935.0/65536.0,1,-nbitq), 
to_sfixed(1663.0/65536.0,1,-nbitq), 
to_sfixed(1214.0/65536.0,1,-nbitq), 
to_sfixed(-3162.0/65536.0,1,-nbitq), 
to_sfixed(-3512.0/65536.0,1,-nbitq), 
to_sfixed(8020.0/65536.0,1,-nbitq), 
to_sfixed(-4406.0/65536.0,1,-nbitq), 
to_sfixed(-7181.0/65536.0,1,-nbitq), 
to_sfixed(7339.0/65536.0,1,-nbitq), 
to_sfixed(4297.0/65536.0,1,-nbitq), 
to_sfixed(4412.0/65536.0,1,-nbitq), 
to_sfixed(2432.0/65536.0,1,-nbitq), 
to_sfixed(-1990.0/65536.0,1,-nbitq), 
to_sfixed(4400.0/65536.0,1,-nbitq), 
to_sfixed(-257.0/65536.0,1,-nbitq), 
to_sfixed(-18316.0/65536.0,1,-nbitq), 
to_sfixed(-924.0/65536.0,1,-nbitq), 
to_sfixed(-4060.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1613.0/65536.0,1,-nbitq), 
to_sfixed(897.0/65536.0,1,-nbitq), 
to_sfixed(2878.0/65536.0,1,-nbitq), 
to_sfixed(-5134.0/65536.0,1,-nbitq), 
to_sfixed(9279.0/65536.0,1,-nbitq), 
to_sfixed(5339.0/65536.0,1,-nbitq), 
to_sfixed(-3921.0/65536.0,1,-nbitq), 
to_sfixed(5093.0/65536.0,1,-nbitq), 
to_sfixed(676.0/65536.0,1,-nbitq), 
to_sfixed(2212.0/65536.0,1,-nbitq), 
to_sfixed(3659.0/65536.0,1,-nbitq), 
to_sfixed(-1416.0/65536.0,1,-nbitq), 
to_sfixed(-2695.0/65536.0,1,-nbitq), 
to_sfixed(7730.0/65536.0,1,-nbitq), 
to_sfixed(1892.0/65536.0,1,-nbitq), 
to_sfixed(802.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(-6340.0/65536.0,1,-nbitq), 
to_sfixed(3757.0/65536.0,1,-nbitq), 
to_sfixed(1511.0/65536.0,1,-nbitq), 
to_sfixed(4993.0/65536.0,1,-nbitq), 
to_sfixed(-8695.0/65536.0,1,-nbitq), 
to_sfixed(1365.0/65536.0,1,-nbitq), 
to_sfixed(8179.0/65536.0,1,-nbitq), 
to_sfixed(529.0/65536.0,1,-nbitq), 
to_sfixed(9088.0/65536.0,1,-nbitq), 
to_sfixed(-505.0/65536.0,1,-nbitq), 
to_sfixed(1747.0/65536.0,1,-nbitq), 
to_sfixed(-660.0/65536.0,1,-nbitq), 
to_sfixed(-4549.0/65536.0,1,-nbitq), 
to_sfixed(-1944.0/65536.0,1,-nbitq), 
to_sfixed(-416.0/65536.0,1,-nbitq), 
to_sfixed(1519.0/65536.0,1,-nbitq), 
to_sfixed(4201.0/65536.0,1,-nbitq), 
to_sfixed(-2129.0/65536.0,1,-nbitq), 
to_sfixed(-2836.0/65536.0,1,-nbitq), 
to_sfixed(2271.0/65536.0,1,-nbitq), 
to_sfixed(-3152.0/65536.0,1,-nbitq), 
to_sfixed(8501.0/65536.0,1,-nbitq), 
to_sfixed(1065.0/65536.0,1,-nbitq), 
to_sfixed(1854.0/65536.0,1,-nbitq), 
to_sfixed(2329.0/65536.0,1,-nbitq), 
to_sfixed(10523.0/65536.0,1,-nbitq), 
to_sfixed(-1068.0/65536.0,1,-nbitq), 
to_sfixed(2312.0/65536.0,1,-nbitq), 
to_sfixed(2941.0/65536.0,1,-nbitq), 
to_sfixed(-3668.0/65536.0,1,-nbitq), 
to_sfixed(-9092.0/65536.0,1,-nbitq), 
to_sfixed(-800.0/65536.0,1,-nbitq), 
to_sfixed(-158.0/65536.0,1,-nbitq), 
to_sfixed(1666.0/65536.0,1,-nbitq), 
to_sfixed(2252.0/65536.0,1,-nbitq), 
to_sfixed(2973.0/65536.0,1,-nbitq), 
to_sfixed(-3004.0/65536.0,1,-nbitq), 
to_sfixed(-1139.0/65536.0,1,-nbitq), 
to_sfixed(5624.0/65536.0,1,-nbitq), 
to_sfixed(1353.0/65536.0,1,-nbitq), 
to_sfixed(-305.0/65536.0,1,-nbitq), 
to_sfixed(-1755.0/65536.0,1,-nbitq), 
to_sfixed(550.0/65536.0,1,-nbitq), 
to_sfixed(2825.0/65536.0,1,-nbitq), 
to_sfixed(-1898.0/65536.0,1,-nbitq), 
to_sfixed(670.0/65536.0,1,-nbitq), 
to_sfixed(-181.0/65536.0,1,-nbitq), 
to_sfixed(3912.0/65536.0,1,-nbitq), 
to_sfixed(-2809.0/65536.0,1,-nbitq), 
to_sfixed(-2456.0/65536.0,1,-nbitq), 
to_sfixed(1551.0/65536.0,1,-nbitq), 
to_sfixed(-2084.0/65536.0,1,-nbitq), 
to_sfixed(-8904.0/65536.0,1,-nbitq), 
to_sfixed(5095.0/65536.0,1,-nbitq), 
to_sfixed(3224.0/65536.0,1,-nbitq), 
to_sfixed(8032.0/65536.0,1,-nbitq), 
to_sfixed(-1973.0/65536.0,1,-nbitq), 
to_sfixed(1454.0/65536.0,1,-nbitq), 
to_sfixed(429.0/65536.0,1,-nbitq), 
to_sfixed(1592.0/65536.0,1,-nbitq), 
to_sfixed(-12117.0/65536.0,1,-nbitq), 
to_sfixed(-2784.0/65536.0,1,-nbitq), 
to_sfixed(-6506.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2315.0/65536.0,1,-nbitq), 
to_sfixed(3979.0/65536.0,1,-nbitq), 
to_sfixed(-1106.0/65536.0,1,-nbitq), 
to_sfixed(-5002.0/65536.0,1,-nbitq), 
to_sfixed(-361.0/65536.0,1,-nbitq), 
to_sfixed(2658.0/65536.0,1,-nbitq), 
to_sfixed(-94.0/65536.0,1,-nbitq), 
to_sfixed(7602.0/65536.0,1,-nbitq), 
to_sfixed(-5675.0/65536.0,1,-nbitq), 
to_sfixed(-2408.0/65536.0,1,-nbitq), 
to_sfixed(470.0/65536.0,1,-nbitq), 
to_sfixed(5390.0/65536.0,1,-nbitq), 
to_sfixed(-2674.0/65536.0,1,-nbitq), 
to_sfixed(-693.0/65536.0,1,-nbitq), 
to_sfixed(1544.0/65536.0,1,-nbitq), 
to_sfixed(1171.0/65536.0,1,-nbitq), 
to_sfixed(-2002.0/65536.0,1,-nbitq), 
to_sfixed(1669.0/65536.0,1,-nbitq), 
to_sfixed(-1456.0/65536.0,1,-nbitq), 
to_sfixed(733.0/65536.0,1,-nbitq), 
to_sfixed(4922.0/65536.0,1,-nbitq), 
to_sfixed(-3974.0/65536.0,1,-nbitq), 
to_sfixed(383.0/65536.0,1,-nbitq), 
to_sfixed(4877.0/65536.0,1,-nbitq), 
to_sfixed(-1660.0/65536.0,1,-nbitq), 
to_sfixed(6488.0/65536.0,1,-nbitq), 
to_sfixed(4748.0/65536.0,1,-nbitq), 
to_sfixed(-863.0/65536.0,1,-nbitq), 
to_sfixed(208.0/65536.0,1,-nbitq), 
to_sfixed(-4781.0/65536.0,1,-nbitq), 
to_sfixed(-1224.0/65536.0,1,-nbitq), 
to_sfixed(-2366.0/65536.0,1,-nbitq), 
to_sfixed(8596.0/65536.0,1,-nbitq), 
to_sfixed(2102.0/65536.0,1,-nbitq), 
to_sfixed(-1730.0/65536.0,1,-nbitq), 
to_sfixed(-337.0/65536.0,1,-nbitq), 
to_sfixed(1017.0/65536.0,1,-nbitq), 
to_sfixed(-3837.0/65536.0,1,-nbitq), 
to_sfixed(4161.0/65536.0,1,-nbitq), 
to_sfixed(-180.0/65536.0,1,-nbitq), 
to_sfixed(3072.0/65536.0,1,-nbitq), 
to_sfixed(-81.0/65536.0,1,-nbitq), 
to_sfixed(6350.0/65536.0,1,-nbitq), 
to_sfixed(534.0/65536.0,1,-nbitq), 
to_sfixed(1072.0/65536.0,1,-nbitq), 
to_sfixed(668.0/65536.0,1,-nbitq), 
to_sfixed(1100.0/65536.0,1,-nbitq), 
to_sfixed(-7773.0/65536.0,1,-nbitq), 
to_sfixed(-1505.0/65536.0,1,-nbitq), 
to_sfixed(1155.0/65536.0,1,-nbitq), 
to_sfixed(190.0/65536.0,1,-nbitq), 
to_sfixed(2609.0/65536.0,1,-nbitq), 
to_sfixed(5784.0/65536.0,1,-nbitq), 
to_sfixed(-349.0/65536.0,1,-nbitq), 
to_sfixed(2665.0/65536.0,1,-nbitq), 
to_sfixed(690.0/65536.0,1,-nbitq), 
to_sfixed(-38.0/65536.0,1,-nbitq), 
to_sfixed(2143.0/65536.0,1,-nbitq), 
to_sfixed(-1880.0/65536.0,1,-nbitq), 
to_sfixed(2037.0/65536.0,1,-nbitq), 
to_sfixed(-373.0/65536.0,1,-nbitq), 
to_sfixed(1722.0/65536.0,1,-nbitq), 
to_sfixed(-2200.0/65536.0,1,-nbitq), 
to_sfixed(188.0/65536.0,1,-nbitq), 
to_sfixed(-111.0/65536.0,1,-nbitq), 
to_sfixed(267.0/65536.0,1,-nbitq), 
to_sfixed(-2383.0/65536.0,1,-nbitq), 
to_sfixed(804.0/65536.0,1,-nbitq), 
to_sfixed(-5218.0/65536.0,1,-nbitq), 
to_sfixed(-5016.0/65536.0,1,-nbitq), 
to_sfixed(6013.0/65536.0,1,-nbitq), 
to_sfixed(-351.0/65536.0,1,-nbitq), 
to_sfixed(145.0/65536.0,1,-nbitq), 
to_sfixed(-2446.0/65536.0,1,-nbitq), 
to_sfixed(-1134.0/65536.0,1,-nbitq), 
to_sfixed(4546.0/65536.0,1,-nbitq), 
to_sfixed(4339.0/65536.0,1,-nbitq), 
to_sfixed(1388.0/65536.0,1,-nbitq), 
to_sfixed(-15.0/65536.0,1,-nbitq), 
to_sfixed(-9211.0/65536.0,1,-nbitq)  ), 
( to_sfixed(7460.0/65536.0,1,-nbitq), 
to_sfixed(132.0/65536.0,1,-nbitq), 
to_sfixed(612.0/65536.0,1,-nbitq), 
to_sfixed(-2687.0/65536.0,1,-nbitq), 
to_sfixed(-5538.0/65536.0,1,-nbitq), 
to_sfixed(7079.0/65536.0,1,-nbitq), 
to_sfixed(-1937.0/65536.0,1,-nbitq), 
to_sfixed(6814.0/65536.0,1,-nbitq), 
to_sfixed(-4182.0/65536.0,1,-nbitq), 
to_sfixed(-2639.0/65536.0,1,-nbitq), 
to_sfixed(-2472.0/65536.0,1,-nbitq), 
to_sfixed(7246.0/65536.0,1,-nbitq), 
to_sfixed(30.0/65536.0,1,-nbitq), 
to_sfixed(256.0/65536.0,1,-nbitq), 
to_sfixed(-1646.0/65536.0,1,-nbitq), 
to_sfixed(2844.0/65536.0,1,-nbitq), 
to_sfixed(1248.0/65536.0,1,-nbitq), 
to_sfixed(-1260.0/65536.0,1,-nbitq), 
to_sfixed(-2039.0/65536.0,1,-nbitq), 
to_sfixed(39.0/65536.0,1,-nbitq), 
to_sfixed(4046.0/65536.0,1,-nbitq), 
to_sfixed(-1453.0/65536.0,1,-nbitq), 
to_sfixed(-7355.0/65536.0,1,-nbitq), 
to_sfixed(-561.0/65536.0,1,-nbitq), 
to_sfixed(-443.0/65536.0,1,-nbitq), 
to_sfixed(2928.0/65536.0,1,-nbitq), 
to_sfixed(2435.0/65536.0,1,-nbitq), 
to_sfixed(598.0/65536.0,1,-nbitq), 
to_sfixed(2203.0/65536.0,1,-nbitq), 
to_sfixed(120.0/65536.0,1,-nbitq), 
to_sfixed(-2330.0/65536.0,1,-nbitq), 
to_sfixed(-3701.0/65536.0,1,-nbitq), 
to_sfixed(9836.0/65536.0,1,-nbitq), 
to_sfixed(190.0/65536.0,1,-nbitq), 
to_sfixed(627.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(2448.0/65536.0,1,-nbitq), 
to_sfixed(855.0/65536.0,1,-nbitq), 
to_sfixed(1950.0/65536.0,1,-nbitq), 
to_sfixed(869.0/65536.0,1,-nbitq), 
to_sfixed(5086.0/65536.0,1,-nbitq), 
to_sfixed(-536.0/65536.0,1,-nbitq), 
to_sfixed(10337.0/65536.0,1,-nbitq), 
to_sfixed(1281.0/65536.0,1,-nbitq), 
to_sfixed(-2359.0/65536.0,1,-nbitq), 
to_sfixed(-5969.0/65536.0,1,-nbitq), 
to_sfixed(-1743.0/65536.0,1,-nbitq), 
to_sfixed(-3256.0/65536.0,1,-nbitq), 
to_sfixed(-2152.0/65536.0,1,-nbitq), 
to_sfixed(4154.0/65536.0,1,-nbitq), 
to_sfixed(1401.0/65536.0,1,-nbitq), 
to_sfixed(118.0/65536.0,1,-nbitq), 
to_sfixed(12751.0/65536.0,1,-nbitq), 
to_sfixed(-5821.0/65536.0,1,-nbitq), 
to_sfixed(1585.0/65536.0,1,-nbitq), 
to_sfixed(3670.0/65536.0,1,-nbitq), 
to_sfixed(-1646.0/65536.0,1,-nbitq), 
to_sfixed(-798.0/65536.0,1,-nbitq), 
to_sfixed(-2030.0/65536.0,1,-nbitq), 
to_sfixed(5020.0/65536.0,1,-nbitq), 
to_sfixed(2191.0/65536.0,1,-nbitq), 
to_sfixed(2098.0/65536.0,1,-nbitq), 
to_sfixed(-2608.0/65536.0,1,-nbitq), 
to_sfixed(-1487.0/65536.0,1,-nbitq), 
to_sfixed(-3356.0/65536.0,1,-nbitq), 
to_sfixed(1810.0/65536.0,1,-nbitq), 
to_sfixed(4680.0/65536.0,1,-nbitq), 
to_sfixed(1325.0/65536.0,1,-nbitq), 
to_sfixed(-9545.0/65536.0,1,-nbitq), 
to_sfixed(-8824.0/65536.0,1,-nbitq), 
to_sfixed(10243.0/65536.0,1,-nbitq), 
to_sfixed(-995.0/65536.0,1,-nbitq), 
to_sfixed(2089.0/65536.0,1,-nbitq), 
to_sfixed(-1741.0/65536.0,1,-nbitq), 
to_sfixed(-2565.0/65536.0,1,-nbitq), 
to_sfixed(1993.0/65536.0,1,-nbitq), 
to_sfixed(1513.0/65536.0,1,-nbitq), 
to_sfixed(1161.0/65536.0,1,-nbitq), 
to_sfixed(64.0/65536.0,1,-nbitq), 
to_sfixed(-9853.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5410.0/65536.0,1,-nbitq), 
to_sfixed(-1564.0/65536.0,1,-nbitq), 
to_sfixed(-238.0/65536.0,1,-nbitq), 
to_sfixed(-252.0/65536.0,1,-nbitq), 
to_sfixed(-456.0/65536.0,1,-nbitq), 
to_sfixed(4434.0/65536.0,1,-nbitq), 
to_sfixed(994.0/65536.0,1,-nbitq), 
to_sfixed(1039.0/65536.0,1,-nbitq), 
to_sfixed(-2434.0/65536.0,1,-nbitq), 
to_sfixed(-1434.0/65536.0,1,-nbitq), 
to_sfixed(3169.0/65536.0,1,-nbitq), 
to_sfixed(2344.0/65536.0,1,-nbitq), 
to_sfixed(-467.0/65536.0,1,-nbitq), 
to_sfixed(-927.0/65536.0,1,-nbitq), 
to_sfixed(242.0/65536.0,1,-nbitq), 
to_sfixed(-362.0/65536.0,1,-nbitq), 
to_sfixed(2395.0/65536.0,1,-nbitq), 
to_sfixed(1629.0/65536.0,1,-nbitq), 
to_sfixed(-2509.0/65536.0,1,-nbitq), 
to_sfixed(-394.0/65536.0,1,-nbitq), 
to_sfixed(1170.0/65536.0,1,-nbitq), 
to_sfixed(-1505.0/65536.0,1,-nbitq), 
to_sfixed(-7304.0/65536.0,1,-nbitq), 
to_sfixed(4739.0/65536.0,1,-nbitq), 
to_sfixed(-2238.0/65536.0,1,-nbitq), 
to_sfixed(1874.0/65536.0,1,-nbitq), 
to_sfixed(1105.0/65536.0,1,-nbitq), 
to_sfixed(-3594.0/65536.0,1,-nbitq), 
to_sfixed(4113.0/65536.0,1,-nbitq), 
to_sfixed(2224.0/65536.0,1,-nbitq), 
to_sfixed(-3103.0/65536.0,1,-nbitq), 
to_sfixed(-679.0/65536.0,1,-nbitq), 
to_sfixed(8490.0/65536.0,1,-nbitq), 
to_sfixed(1355.0/65536.0,1,-nbitq), 
to_sfixed(-2014.0/65536.0,1,-nbitq), 
to_sfixed(-2276.0/65536.0,1,-nbitq), 
to_sfixed(879.0/65536.0,1,-nbitq), 
to_sfixed(2539.0/65536.0,1,-nbitq), 
to_sfixed(-2088.0/65536.0,1,-nbitq), 
to_sfixed(-351.0/65536.0,1,-nbitq), 
to_sfixed(1177.0/65536.0,1,-nbitq), 
to_sfixed(-2994.0/65536.0,1,-nbitq), 
to_sfixed(7828.0/65536.0,1,-nbitq), 
to_sfixed(687.0/65536.0,1,-nbitq), 
to_sfixed(1234.0/65536.0,1,-nbitq), 
to_sfixed(-4718.0/65536.0,1,-nbitq), 
to_sfixed(311.0/65536.0,1,-nbitq), 
to_sfixed(-2447.0/65536.0,1,-nbitq), 
to_sfixed(-1373.0/65536.0,1,-nbitq), 
to_sfixed(-37.0/65536.0,1,-nbitq), 
to_sfixed(3056.0/65536.0,1,-nbitq), 
to_sfixed(978.0/65536.0,1,-nbitq), 
to_sfixed(9100.0/65536.0,1,-nbitq), 
to_sfixed(-2758.0/65536.0,1,-nbitq), 
to_sfixed(3036.0/65536.0,1,-nbitq), 
to_sfixed(4312.0/65536.0,1,-nbitq), 
to_sfixed(-2243.0/65536.0,1,-nbitq), 
to_sfixed(3356.0/65536.0,1,-nbitq), 
to_sfixed(798.0/65536.0,1,-nbitq), 
to_sfixed(4249.0/65536.0,1,-nbitq), 
to_sfixed(316.0/65536.0,1,-nbitq), 
to_sfixed(-2940.0/65536.0,1,-nbitq), 
to_sfixed(260.0/65536.0,1,-nbitq), 
to_sfixed(-1061.0/65536.0,1,-nbitq), 
to_sfixed(988.0/65536.0,1,-nbitq), 
to_sfixed(658.0/65536.0,1,-nbitq), 
to_sfixed(817.0/65536.0,1,-nbitq), 
to_sfixed(1617.0/65536.0,1,-nbitq), 
to_sfixed(-7412.0/65536.0,1,-nbitq), 
to_sfixed(-9212.0/65536.0,1,-nbitq), 
to_sfixed(5919.0/65536.0,1,-nbitq), 
to_sfixed(2748.0/65536.0,1,-nbitq), 
to_sfixed(2626.0/65536.0,1,-nbitq), 
to_sfixed(702.0/65536.0,1,-nbitq), 
to_sfixed(-2461.0/65536.0,1,-nbitq), 
to_sfixed(2512.0/65536.0,1,-nbitq), 
to_sfixed(1022.0/65536.0,1,-nbitq), 
to_sfixed(1105.0/65536.0,1,-nbitq), 
to_sfixed(-40.0/65536.0,1,-nbitq), 
to_sfixed(-8730.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2256.0/65536.0,1,-nbitq), 
to_sfixed(-1993.0/65536.0,1,-nbitq), 
to_sfixed(-2575.0/65536.0,1,-nbitq), 
to_sfixed(-263.0/65536.0,1,-nbitq), 
to_sfixed(-5039.0/65536.0,1,-nbitq), 
to_sfixed(2202.0/65536.0,1,-nbitq), 
to_sfixed(-2129.0/65536.0,1,-nbitq), 
to_sfixed(2337.0/65536.0,1,-nbitq), 
to_sfixed(-210.0/65536.0,1,-nbitq), 
to_sfixed(-117.0/65536.0,1,-nbitq), 
to_sfixed(4349.0/65536.0,1,-nbitq), 
to_sfixed(1285.0/65536.0,1,-nbitq), 
to_sfixed(-2936.0/65536.0,1,-nbitq), 
to_sfixed(4287.0/65536.0,1,-nbitq), 
to_sfixed(-3632.0/65536.0,1,-nbitq), 
to_sfixed(814.0/65536.0,1,-nbitq), 
to_sfixed(1172.0/65536.0,1,-nbitq), 
to_sfixed(-4711.0/65536.0,1,-nbitq), 
to_sfixed(91.0/65536.0,1,-nbitq), 
to_sfixed(1981.0/65536.0,1,-nbitq), 
to_sfixed(98.0/65536.0,1,-nbitq), 
to_sfixed(2766.0/65536.0,1,-nbitq), 
to_sfixed(-1392.0/65536.0,1,-nbitq), 
to_sfixed(5984.0/65536.0,1,-nbitq), 
to_sfixed(3127.0/65536.0,1,-nbitq), 
to_sfixed(2242.0/65536.0,1,-nbitq), 
to_sfixed(3834.0/65536.0,1,-nbitq), 
to_sfixed(2192.0/65536.0,1,-nbitq), 
to_sfixed(-1502.0/65536.0,1,-nbitq), 
to_sfixed(2591.0/65536.0,1,-nbitq), 
to_sfixed(-772.0/65536.0,1,-nbitq), 
to_sfixed(-1033.0/65536.0,1,-nbitq), 
to_sfixed(3661.0/65536.0,1,-nbitq), 
to_sfixed(6960.0/65536.0,1,-nbitq), 
to_sfixed(-2613.0/65536.0,1,-nbitq), 
to_sfixed(1555.0/65536.0,1,-nbitq), 
to_sfixed(2853.0/65536.0,1,-nbitq), 
to_sfixed(5507.0/65536.0,1,-nbitq), 
to_sfixed(2011.0/65536.0,1,-nbitq), 
to_sfixed(2450.0/65536.0,1,-nbitq), 
to_sfixed(-590.0/65536.0,1,-nbitq), 
to_sfixed(1028.0/65536.0,1,-nbitq), 
to_sfixed(8606.0/65536.0,1,-nbitq), 
to_sfixed(-687.0/65536.0,1,-nbitq), 
to_sfixed(2297.0/65536.0,1,-nbitq), 
to_sfixed(-5257.0/65536.0,1,-nbitq), 
to_sfixed(-2352.0/65536.0,1,-nbitq), 
to_sfixed(-1280.0/65536.0,1,-nbitq), 
to_sfixed(1430.0/65536.0,1,-nbitq), 
to_sfixed(1934.0/65536.0,1,-nbitq), 
to_sfixed(-1289.0/65536.0,1,-nbitq), 
to_sfixed(-1894.0/65536.0,1,-nbitq), 
to_sfixed(7423.0/65536.0,1,-nbitq), 
to_sfixed(-475.0/65536.0,1,-nbitq), 
to_sfixed(5315.0/65536.0,1,-nbitq), 
to_sfixed(-781.0/65536.0,1,-nbitq), 
to_sfixed(2169.0/65536.0,1,-nbitq), 
to_sfixed(3668.0/65536.0,1,-nbitq), 
to_sfixed(2559.0/65536.0,1,-nbitq), 
to_sfixed(267.0/65536.0,1,-nbitq), 
to_sfixed(-2607.0/65536.0,1,-nbitq), 
to_sfixed(-1712.0/65536.0,1,-nbitq), 
to_sfixed(136.0/65536.0,1,-nbitq), 
to_sfixed(2198.0/65536.0,1,-nbitq), 
to_sfixed(-2713.0/65536.0,1,-nbitq), 
to_sfixed(-99.0/65536.0,1,-nbitq), 
to_sfixed(1815.0/65536.0,1,-nbitq), 
to_sfixed(901.0/65536.0,1,-nbitq), 
to_sfixed(-4395.0/65536.0,1,-nbitq), 
to_sfixed(-8347.0/65536.0,1,-nbitq), 
to_sfixed(2730.0/65536.0,1,-nbitq), 
to_sfixed(-2000.0/65536.0,1,-nbitq), 
to_sfixed(1636.0/65536.0,1,-nbitq), 
to_sfixed(1517.0/65536.0,1,-nbitq), 
to_sfixed(1865.0/65536.0,1,-nbitq), 
to_sfixed(1081.0/65536.0,1,-nbitq), 
to_sfixed(1687.0/65536.0,1,-nbitq), 
to_sfixed(3280.0/65536.0,1,-nbitq), 
to_sfixed(1458.0/65536.0,1,-nbitq), 
to_sfixed(-4997.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-818.0/65536.0,1,-nbitq), 
to_sfixed(-3839.0/65536.0,1,-nbitq), 
to_sfixed(-681.0/65536.0,1,-nbitq), 
to_sfixed(-1749.0/65536.0,1,-nbitq), 
to_sfixed(-4665.0/65536.0,1,-nbitq), 
to_sfixed(1432.0/65536.0,1,-nbitq), 
to_sfixed(1791.0/65536.0,1,-nbitq), 
to_sfixed(-1833.0/65536.0,1,-nbitq), 
to_sfixed(-3080.0/65536.0,1,-nbitq), 
to_sfixed(436.0/65536.0,1,-nbitq), 
to_sfixed(1480.0/65536.0,1,-nbitq), 
to_sfixed(-1498.0/65536.0,1,-nbitq), 
to_sfixed(38.0/65536.0,1,-nbitq), 
to_sfixed(-164.0/65536.0,1,-nbitq), 
to_sfixed(99.0/65536.0,1,-nbitq), 
to_sfixed(682.0/65536.0,1,-nbitq), 
to_sfixed(-1357.0/65536.0,1,-nbitq), 
to_sfixed(-5683.0/65536.0,1,-nbitq), 
to_sfixed(-3021.0/65536.0,1,-nbitq), 
to_sfixed(3130.0/65536.0,1,-nbitq), 
to_sfixed(2461.0/65536.0,1,-nbitq), 
to_sfixed(342.0/65536.0,1,-nbitq), 
to_sfixed(-3400.0/65536.0,1,-nbitq), 
to_sfixed(6628.0/65536.0,1,-nbitq), 
to_sfixed(522.0/65536.0,1,-nbitq), 
to_sfixed(1811.0/65536.0,1,-nbitq), 
to_sfixed(1189.0/65536.0,1,-nbitq), 
to_sfixed(2586.0/65536.0,1,-nbitq), 
to_sfixed(290.0/65536.0,1,-nbitq), 
to_sfixed(4096.0/65536.0,1,-nbitq), 
to_sfixed(-1441.0/65536.0,1,-nbitq), 
to_sfixed(2337.0/65536.0,1,-nbitq), 
to_sfixed(3791.0/65536.0,1,-nbitq), 
to_sfixed(1232.0/65536.0,1,-nbitq), 
to_sfixed(-1147.0/65536.0,1,-nbitq), 
to_sfixed(-570.0/65536.0,1,-nbitq), 
to_sfixed(1065.0/65536.0,1,-nbitq), 
to_sfixed(-616.0/65536.0,1,-nbitq), 
to_sfixed(-306.0/65536.0,1,-nbitq), 
to_sfixed(2792.0/65536.0,1,-nbitq), 
to_sfixed(-1977.0/65536.0,1,-nbitq), 
to_sfixed(-611.0/65536.0,1,-nbitq), 
to_sfixed(1874.0/65536.0,1,-nbitq), 
to_sfixed(4604.0/65536.0,1,-nbitq), 
to_sfixed(3322.0/65536.0,1,-nbitq), 
to_sfixed(-131.0/65536.0,1,-nbitq), 
to_sfixed(-2766.0/65536.0,1,-nbitq), 
to_sfixed(1778.0/65536.0,1,-nbitq), 
to_sfixed(2560.0/65536.0,1,-nbitq), 
to_sfixed(-434.0/65536.0,1,-nbitq), 
to_sfixed(-1310.0/65536.0,1,-nbitq), 
to_sfixed(-2126.0/65536.0,1,-nbitq), 
to_sfixed(5251.0/65536.0,1,-nbitq), 
to_sfixed(1173.0/65536.0,1,-nbitq), 
to_sfixed(1566.0/65536.0,1,-nbitq), 
to_sfixed(3665.0/65536.0,1,-nbitq), 
to_sfixed(-399.0/65536.0,1,-nbitq), 
to_sfixed(-995.0/65536.0,1,-nbitq), 
to_sfixed(2281.0/65536.0,1,-nbitq), 
to_sfixed(4053.0/65536.0,1,-nbitq), 
to_sfixed(-320.0/65536.0,1,-nbitq), 
to_sfixed(-126.0/65536.0,1,-nbitq), 
to_sfixed(-908.0/65536.0,1,-nbitq), 
to_sfixed(-1456.0/65536.0,1,-nbitq), 
to_sfixed(-2664.0/65536.0,1,-nbitq), 
to_sfixed(39.0/65536.0,1,-nbitq), 
to_sfixed(236.0/65536.0,1,-nbitq), 
to_sfixed(-1090.0/65536.0,1,-nbitq), 
to_sfixed(-4590.0/65536.0,1,-nbitq), 
to_sfixed(-2288.0/65536.0,1,-nbitq), 
to_sfixed(1303.0/65536.0,1,-nbitq), 
to_sfixed(1902.0/65536.0,1,-nbitq), 
to_sfixed(-1126.0/65536.0,1,-nbitq), 
to_sfixed(1081.0/65536.0,1,-nbitq), 
to_sfixed(2516.0/65536.0,1,-nbitq), 
to_sfixed(-1155.0/65536.0,1,-nbitq), 
to_sfixed(2476.0/65536.0,1,-nbitq), 
to_sfixed(1198.0/65536.0,1,-nbitq), 
to_sfixed(-1603.0/65536.0,1,-nbitq), 
to_sfixed(-4460.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2461.0/65536.0,1,-nbitq), 
to_sfixed(-2670.0/65536.0,1,-nbitq), 
to_sfixed(870.0/65536.0,1,-nbitq), 
to_sfixed(2052.0/65536.0,1,-nbitq), 
to_sfixed(-1980.0/65536.0,1,-nbitq), 
to_sfixed(-997.0/65536.0,1,-nbitq), 
to_sfixed(818.0/65536.0,1,-nbitq), 
to_sfixed(1947.0/65536.0,1,-nbitq), 
to_sfixed(-3353.0/65536.0,1,-nbitq), 
to_sfixed(-494.0/65536.0,1,-nbitq), 
to_sfixed(1315.0/65536.0,1,-nbitq), 
to_sfixed(926.0/65536.0,1,-nbitq), 
to_sfixed(-78.0/65536.0,1,-nbitq), 
to_sfixed(2291.0/65536.0,1,-nbitq), 
to_sfixed(445.0/65536.0,1,-nbitq), 
to_sfixed(2604.0/65536.0,1,-nbitq), 
to_sfixed(512.0/65536.0,1,-nbitq), 
to_sfixed(-2408.0/65536.0,1,-nbitq), 
to_sfixed(242.0/65536.0,1,-nbitq), 
to_sfixed(1781.0/65536.0,1,-nbitq), 
to_sfixed(-1231.0/65536.0,1,-nbitq), 
to_sfixed(-1253.0/65536.0,1,-nbitq), 
to_sfixed(1625.0/65536.0,1,-nbitq), 
to_sfixed(4393.0/65536.0,1,-nbitq), 
to_sfixed(193.0/65536.0,1,-nbitq), 
to_sfixed(3247.0/65536.0,1,-nbitq), 
to_sfixed(-4836.0/65536.0,1,-nbitq), 
to_sfixed(-194.0/65536.0,1,-nbitq), 
to_sfixed(-1690.0/65536.0,1,-nbitq), 
to_sfixed(863.0/65536.0,1,-nbitq), 
to_sfixed(-1678.0/65536.0,1,-nbitq), 
to_sfixed(2671.0/65536.0,1,-nbitq), 
to_sfixed(1182.0/65536.0,1,-nbitq), 
to_sfixed(-288.0/65536.0,1,-nbitq), 
to_sfixed(-364.0/65536.0,1,-nbitq), 
to_sfixed(2299.0/65536.0,1,-nbitq), 
to_sfixed(-1150.0/65536.0,1,-nbitq), 
to_sfixed(1364.0/65536.0,1,-nbitq), 
to_sfixed(-2610.0/65536.0,1,-nbitq), 
to_sfixed(2677.0/65536.0,1,-nbitq), 
to_sfixed(-3137.0/65536.0,1,-nbitq), 
to_sfixed(-1331.0/65536.0,1,-nbitq), 
to_sfixed(-2270.0/65536.0,1,-nbitq), 
to_sfixed(3558.0/65536.0,1,-nbitq), 
to_sfixed(-1177.0/65536.0,1,-nbitq), 
to_sfixed(4449.0/65536.0,1,-nbitq), 
to_sfixed(-2666.0/65536.0,1,-nbitq), 
to_sfixed(543.0/65536.0,1,-nbitq), 
to_sfixed(-231.0/65536.0,1,-nbitq), 
to_sfixed(4484.0/65536.0,1,-nbitq), 
to_sfixed(-336.0/65536.0,1,-nbitq), 
to_sfixed(-1392.0/65536.0,1,-nbitq), 
to_sfixed(1261.0/65536.0,1,-nbitq), 
to_sfixed(-3446.0/65536.0,1,-nbitq), 
to_sfixed(1825.0/65536.0,1,-nbitq), 
to_sfixed(-137.0/65536.0,1,-nbitq), 
to_sfixed(2052.0/65536.0,1,-nbitq), 
to_sfixed(-1129.0/65536.0,1,-nbitq), 
to_sfixed(2502.0/65536.0,1,-nbitq), 
to_sfixed(2735.0/65536.0,1,-nbitq), 
to_sfixed(386.0/65536.0,1,-nbitq), 
to_sfixed(-720.0/65536.0,1,-nbitq), 
to_sfixed(118.0/65536.0,1,-nbitq), 
to_sfixed(-40.0/65536.0,1,-nbitq), 
to_sfixed(1107.0/65536.0,1,-nbitq), 
to_sfixed(147.0/65536.0,1,-nbitq), 
to_sfixed(-2907.0/65536.0,1,-nbitq), 
to_sfixed(1552.0/65536.0,1,-nbitq), 
to_sfixed(349.0/65536.0,1,-nbitq), 
to_sfixed(-2236.0/65536.0,1,-nbitq), 
to_sfixed(2986.0/65536.0,1,-nbitq), 
to_sfixed(1135.0/65536.0,1,-nbitq), 
to_sfixed(3325.0/65536.0,1,-nbitq), 
to_sfixed(-3026.0/65536.0,1,-nbitq), 
to_sfixed(-107.0/65536.0,1,-nbitq), 
to_sfixed(860.0/65536.0,1,-nbitq), 
to_sfixed(-2698.0/65536.0,1,-nbitq), 
to_sfixed(-277.0/65536.0,1,-nbitq), 
to_sfixed(2881.0/65536.0,1,-nbitq), 
to_sfixed(-467.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-360.0/65536.0,1,-nbitq), 
to_sfixed(-2262.0/65536.0,1,-nbitq), 
to_sfixed(1805.0/65536.0,1,-nbitq), 
to_sfixed(-2492.0/65536.0,1,-nbitq), 
to_sfixed(-1850.0/65536.0,1,-nbitq), 
to_sfixed(-1370.0/65536.0,1,-nbitq), 
to_sfixed(2382.0/65536.0,1,-nbitq), 
to_sfixed(399.0/65536.0,1,-nbitq), 
to_sfixed(305.0/65536.0,1,-nbitq), 
to_sfixed(-757.0/65536.0,1,-nbitq), 
to_sfixed(2052.0/65536.0,1,-nbitq), 
to_sfixed(-1736.0/65536.0,1,-nbitq), 
to_sfixed(-545.0/65536.0,1,-nbitq), 
to_sfixed(-30.0/65536.0,1,-nbitq), 
to_sfixed(236.0/65536.0,1,-nbitq), 
to_sfixed(2000.0/65536.0,1,-nbitq), 
to_sfixed(2872.0/65536.0,1,-nbitq), 
to_sfixed(3543.0/65536.0,1,-nbitq), 
to_sfixed(-639.0/65536.0,1,-nbitq), 
to_sfixed(-677.0/65536.0,1,-nbitq), 
to_sfixed(-674.0/65536.0,1,-nbitq), 
to_sfixed(2232.0/65536.0,1,-nbitq), 
to_sfixed(511.0/65536.0,1,-nbitq), 
to_sfixed(3674.0/65536.0,1,-nbitq), 
to_sfixed(3384.0/65536.0,1,-nbitq), 
to_sfixed(-54.0/65536.0,1,-nbitq), 
to_sfixed(2191.0/65536.0,1,-nbitq), 
to_sfixed(874.0/65536.0,1,-nbitq), 
to_sfixed(667.0/65536.0,1,-nbitq), 
to_sfixed(-128.0/65536.0,1,-nbitq), 
to_sfixed(1005.0/65536.0,1,-nbitq), 
to_sfixed(-621.0/65536.0,1,-nbitq), 
to_sfixed(690.0/65536.0,1,-nbitq), 
to_sfixed(-1561.0/65536.0,1,-nbitq), 
to_sfixed(-480.0/65536.0,1,-nbitq), 
to_sfixed(1070.0/65536.0,1,-nbitq), 
to_sfixed(654.0/65536.0,1,-nbitq), 
to_sfixed(-2926.0/65536.0,1,-nbitq), 
to_sfixed(878.0/65536.0,1,-nbitq), 
to_sfixed(-1629.0/65536.0,1,-nbitq), 
to_sfixed(-3055.0/65536.0,1,-nbitq), 
to_sfixed(-3099.0/65536.0,1,-nbitq), 
to_sfixed(-1019.0/65536.0,1,-nbitq), 
to_sfixed(200.0/65536.0,1,-nbitq), 
to_sfixed(2686.0/65536.0,1,-nbitq), 
to_sfixed(3187.0/65536.0,1,-nbitq), 
to_sfixed(-1328.0/65536.0,1,-nbitq), 
to_sfixed(-435.0/65536.0,1,-nbitq), 
to_sfixed(852.0/65536.0,1,-nbitq), 
to_sfixed(-897.0/65536.0,1,-nbitq), 
to_sfixed(991.0/65536.0,1,-nbitq), 
to_sfixed(-2881.0/65536.0,1,-nbitq), 
to_sfixed(-1505.0/65536.0,1,-nbitq), 
to_sfixed(-712.0/65536.0,1,-nbitq), 
to_sfixed(1205.0/65536.0,1,-nbitq), 
to_sfixed(-321.0/65536.0,1,-nbitq), 
to_sfixed(954.0/65536.0,1,-nbitq), 
to_sfixed(1520.0/65536.0,1,-nbitq), 
to_sfixed(721.0/65536.0,1,-nbitq), 
to_sfixed(4742.0/65536.0,1,-nbitq), 
to_sfixed(-1961.0/65536.0,1,-nbitq), 
to_sfixed(-801.0/65536.0,1,-nbitq), 
to_sfixed(606.0/65536.0,1,-nbitq), 
to_sfixed(-2901.0/65536.0,1,-nbitq), 
to_sfixed(1974.0/65536.0,1,-nbitq), 
to_sfixed(-1628.0/65536.0,1,-nbitq), 
to_sfixed(478.0/65536.0,1,-nbitq), 
to_sfixed(-500.0/65536.0,1,-nbitq), 
to_sfixed(2401.0/65536.0,1,-nbitq), 
to_sfixed(-757.0/65536.0,1,-nbitq), 
to_sfixed(-1021.0/65536.0,1,-nbitq), 
to_sfixed(981.0/65536.0,1,-nbitq), 
to_sfixed(3729.0/65536.0,1,-nbitq), 
to_sfixed(-2827.0/65536.0,1,-nbitq), 
to_sfixed(2017.0/65536.0,1,-nbitq), 
to_sfixed(3950.0/65536.0,1,-nbitq), 
to_sfixed(1957.0/65536.0,1,-nbitq), 
to_sfixed(3350.0/65536.0,1,-nbitq), 
to_sfixed(-815.0/65536.0,1,-nbitq), 
to_sfixed(-10.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1607.0/65536.0,1,-nbitq), 
to_sfixed(292.0/65536.0,1,-nbitq), 
to_sfixed(-1040.0/65536.0,1,-nbitq), 
to_sfixed(2930.0/65536.0,1,-nbitq), 
to_sfixed(-1372.0/65536.0,1,-nbitq), 
to_sfixed(-388.0/65536.0,1,-nbitq), 
to_sfixed(-3177.0/65536.0,1,-nbitq), 
to_sfixed(-748.0/65536.0,1,-nbitq), 
to_sfixed(-1752.0/65536.0,1,-nbitq), 
to_sfixed(-1013.0/65536.0,1,-nbitq), 
to_sfixed(-3163.0/65536.0,1,-nbitq), 
to_sfixed(2913.0/65536.0,1,-nbitq), 
to_sfixed(-1994.0/65536.0,1,-nbitq), 
to_sfixed(-3577.0/65536.0,1,-nbitq), 
to_sfixed(2306.0/65536.0,1,-nbitq), 
to_sfixed(-626.0/65536.0,1,-nbitq), 
to_sfixed(2682.0/65536.0,1,-nbitq), 
to_sfixed(1472.0/65536.0,1,-nbitq), 
to_sfixed(2934.0/65536.0,1,-nbitq), 
to_sfixed(3236.0/65536.0,1,-nbitq), 
to_sfixed(-742.0/65536.0,1,-nbitq), 
to_sfixed(-607.0/65536.0,1,-nbitq), 
to_sfixed(2352.0/65536.0,1,-nbitq), 
to_sfixed(3469.0/65536.0,1,-nbitq), 
to_sfixed(-734.0/65536.0,1,-nbitq), 
to_sfixed(3454.0/65536.0,1,-nbitq), 
to_sfixed(960.0/65536.0,1,-nbitq), 
to_sfixed(280.0/65536.0,1,-nbitq), 
to_sfixed(1185.0/65536.0,1,-nbitq), 
to_sfixed(-1638.0/65536.0,1,-nbitq), 
to_sfixed(89.0/65536.0,1,-nbitq), 
to_sfixed(-2627.0/65536.0,1,-nbitq), 
to_sfixed(2338.0/65536.0,1,-nbitq), 
to_sfixed(-2027.0/65536.0,1,-nbitq), 
to_sfixed(2403.0/65536.0,1,-nbitq), 
to_sfixed(930.0/65536.0,1,-nbitq), 
to_sfixed(-965.0/65536.0,1,-nbitq), 
to_sfixed(-3510.0/65536.0,1,-nbitq), 
to_sfixed(1440.0/65536.0,1,-nbitq), 
to_sfixed(-1303.0/65536.0,1,-nbitq), 
to_sfixed(-2079.0/65536.0,1,-nbitq), 
to_sfixed(293.0/65536.0,1,-nbitq), 
to_sfixed(776.0/65536.0,1,-nbitq), 
to_sfixed(-184.0/65536.0,1,-nbitq), 
to_sfixed(-977.0/65536.0,1,-nbitq), 
to_sfixed(2794.0/65536.0,1,-nbitq), 
to_sfixed(-243.0/65536.0,1,-nbitq), 
to_sfixed(3410.0/65536.0,1,-nbitq), 
to_sfixed(1893.0/65536.0,1,-nbitq), 
to_sfixed(3309.0/65536.0,1,-nbitq), 
to_sfixed(1606.0/65536.0,1,-nbitq), 
to_sfixed(890.0/65536.0,1,-nbitq), 
to_sfixed(1638.0/65536.0,1,-nbitq), 
to_sfixed(1345.0/65536.0,1,-nbitq), 
to_sfixed(-70.0/65536.0,1,-nbitq), 
to_sfixed(2235.0/65536.0,1,-nbitq), 
to_sfixed(3012.0/65536.0,1,-nbitq), 
to_sfixed(916.0/65536.0,1,-nbitq), 
to_sfixed(-707.0/65536.0,1,-nbitq), 
to_sfixed(1376.0/65536.0,1,-nbitq), 
to_sfixed(-1396.0/65536.0,1,-nbitq), 
to_sfixed(2177.0/65536.0,1,-nbitq), 
to_sfixed(295.0/65536.0,1,-nbitq), 
to_sfixed(1749.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(3232.0/65536.0,1,-nbitq), 
to_sfixed(76.0/65536.0,1,-nbitq), 
to_sfixed(1603.0/65536.0,1,-nbitq), 
to_sfixed(-1294.0/65536.0,1,-nbitq), 
to_sfixed(3504.0/65536.0,1,-nbitq), 
to_sfixed(2405.0/65536.0,1,-nbitq), 
to_sfixed(-2309.0/65536.0,1,-nbitq), 
to_sfixed(-1048.0/65536.0,1,-nbitq), 
to_sfixed(702.0/65536.0,1,-nbitq), 
to_sfixed(1518.0/65536.0,1,-nbitq), 
to_sfixed(675.0/65536.0,1,-nbitq), 
to_sfixed(-1125.0/65536.0,1,-nbitq), 
to_sfixed(4443.0/65536.0,1,-nbitq), 
to_sfixed(-403.0/65536.0,1,-nbitq), 
to_sfixed(3818.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1620.0/65536.0,1,-nbitq), 
to_sfixed(2541.0/65536.0,1,-nbitq), 
to_sfixed(2991.0/65536.0,1,-nbitq), 
to_sfixed(239.0/65536.0,1,-nbitq), 
to_sfixed(-2355.0/65536.0,1,-nbitq), 
to_sfixed(-6037.0/65536.0,1,-nbitq), 
to_sfixed(239.0/65536.0,1,-nbitq), 
to_sfixed(1403.0/65536.0,1,-nbitq), 
to_sfixed(2960.0/65536.0,1,-nbitq), 
to_sfixed(840.0/65536.0,1,-nbitq), 
to_sfixed(-1193.0/65536.0,1,-nbitq), 
to_sfixed(-1228.0/65536.0,1,-nbitq), 
to_sfixed(2010.0/65536.0,1,-nbitq), 
to_sfixed(1067.0/65536.0,1,-nbitq), 
to_sfixed(555.0/65536.0,1,-nbitq), 
to_sfixed(613.0/65536.0,1,-nbitq), 
to_sfixed(-93.0/65536.0,1,-nbitq), 
to_sfixed(3270.0/65536.0,1,-nbitq), 
to_sfixed(2289.0/65536.0,1,-nbitq), 
to_sfixed(-801.0/65536.0,1,-nbitq), 
to_sfixed(837.0/65536.0,1,-nbitq), 
to_sfixed(-2652.0/65536.0,1,-nbitq), 
to_sfixed(805.0/65536.0,1,-nbitq), 
to_sfixed(2189.0/65536.0,1,-nbitq), 
to_sfixed(-373.0/65536.0,1,-nbitq), 
to_sfixed(2147.0/65536.0,1,-nbitq), 
to_sfixed(147.0/65536.0,1,-nbitq), 
to_sfixed(2662.0/65536.0,1,-nbitq), 
to_sfixed(-4330.0/65536.0,1,-nbitq), 
to_sfixed(-3627.0/65536.0,1,-nbitq), 
to_sfixed(-2137.0/65536.0,1,-nbitq), 
to_sfixed(871.0/65536.0,1,-nbitq), 
to_sfixed(-1365.0/65536.0,1,-nbitq), 
to_sfixed(-2149.0/65536.0,1,-nbitq), 
to_sfixed(-304.0/65536.0,1,-nbitq), 
to_sfixed(401.0/65536.0,1,-nbitq), 
to_sfixed(977.0/65536.0,1,-nbitq), 
to_sfixed(-250.0/65536.0,1,-nbitq), 
to_sfixed(-2748.0/65536.0,1,-nbitq), 
to_sfixed(-429.0/65536.0,1,-nbitq), 
to_sfixed(831.0/65536.0,1,-nbitq), 
to_sfixed(1955.0/65536.0,1,-nbitq), 
to_sfixed(-1776.0/65536.0,1,-nbitq), 
to_sfixed(1671.0/65536.0,1,-nbitq), 
to_sfixed(-415.0/65536.0,1,-nbitq), 
to_sfixed(2182.0/65536.0,1,-nbitq), 
to_sfixed(1291.0/65536.0,1,-nbitq), 
to_sfixed(2140.0/65536.0,1,-nbitq), 
to_sfixed(1418.0/65536.0,1,-nbitq), 
to_sfixed(3301.0/65536.0,1,-nbitq), 
to_sfixed(-1229.0/65536.0,1,-nbitq), 
to_sfixed(-228.0/65536.0,1,-nbitq), 
to_sfixed(-1507.0/65536.0,1,-nbitq), 
to_sfixed(1708.0/65536.0,1,-nbitq), 
to_sfixed(1595.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(-422.0/65536.0,1,-nbitq), 
to_sfixed(1703.0/65536.0,1,-nbitq), 
to_sfixed(1841.0/65536.0,1,-nbitq), 
to_sfixed(3916.0/65536.0,1,-nbitq), 
to_sfixed(557.0/65536.0,1,-nbitq), 
to_sfixed(-1091.0/65536.0,1,-nbitq), 
to_sfixed(2821.0/65536.0,1,-nbitq), 
to_sfixed(-2996.0/65536.0,1,-nbitq), 
to_sfixed(-1797.0/65536.0,1,-nbitq), 
to_sfixed(1215.0/65536.0,1,-nbitq), 
to_sfixed(213.0/65536.0,1,-nbitq), 
to_sfixed(-3054.0/65536.0,1,-nbitq), 
to_sfixed(-1768.0/65536.0,1,-nbitq), 
to_sfixed(-2301.0/65536.0,1,-nbitq), 
to_sfixed(-185.0/65536.0,1,-nbitq), 
to_sfixed(2888.0/65536.0,1,-nbitq), 
to_sfixed(521.0/65536.0,1,-nbitq), 
to_sfixed(-133.0/65536.0,1,-nbitq), 
to_sfixed(1342.0/65536.0,1,-nbitq), 
to_sfixed(567.0/65536.0,1,-nbitq), 
to_sfixed(-965.0/65536.0,1,-nbitq), 
to_sfixed(-104.0/65536.0,1,-nbitq), 
to_sfixed(849.0/65536.0,1,-nbitq), 
to_sfixed(398.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-227.0/65536.0,1,-nbitq), 
to_sfixed(-1181.0/65536.0,1,-nbitq), 
to_sfixed(193.0/65536.0,1,-nbitq), 
to_sfixed(2672.0/65536.0,1,-nbitq), 
to_sfixed(-866.0/65536.0,1,-nbitq), 
to_sfixed(-1147.0/65536.0,1,-nbitq), 
to_sfixed(-266.0/65536.0,1,-nbitq), 
to_sfixed(422.0/65536.0,1,-nbitq), 
to_sfixed(-1761.0/65536.0,1,-nbitq), 
to_sfixed(-2045.0/65536.0,1,-nbitq), 
to_sfixed(-2135.0/65536.0,1,-nbitq), 
to_sfixed(-382.0/65536.0,1,-nbitq), 
to_sfixed(-215.0/65536.0,1,-nbitq), 
to_sfixed(1138.0/65536.0,1,-nbitq), 
to_sfixed(-1305.0/65536.0,1,-nbitq), 
to_sfixed(-695.0/65536.0,1,-nbitq), 
to_sfixed(30.0/65536.0,1,-nbitq), 
to_sfixed(2256.0/65536.0,1,-nbitq), 
to_sfixed(478.0/65536.0,1,-nbitq), 
to_sfixed(-2007.0/65536.0,1,-nbitq), 
to_sfixed(1616.0/65536.0,1,-nbitq), 
to_sfixed(243.0/65536.0,1,-nbitq), 
to_sfixed(-828.0/65536.0,1,-nbitq), 
to_sfixed(-660.0/65536.0,1,-nbitq), 
to_sfixed(-70.0/65536.0,1,-nbitq), 
to_sfixed(2561.0/65536.0,1,-nbitq), 
to_sfixed(657.0/65536.0,1,-nbitq), 
to_sfixed(119.0/65536.0,1,-nbitq), 
to_sfixed(-1158.0/65536.0,1,-nbitq), 
to_sfixed(526.0/65536.0,1,-nbitq), 
to_sfixed(-2716.0/65536.0,1,-nbitq), 
to_sfixed(-1906.0/65536.0,1,-nbitq), 
to_sfixed(-690.0/65536.0,1,-nbitq), 
to_sfixed(1157.0/65536.0,1,-nbitq), 
to_sfixed(1995.0/65536.0,1,-nbitq), 
to_sfixed(1838.0/65536.0,1,-nbitq), 
to_sfixed(-575.0/65536.0,1,-nbitq), 
to_sfixed(-3558.0/65536.0,1,-nbitq), 
to_sfixed(-4612.0/65536.0,1,-nbitq), 
to_sfixed(-909.0/65536.0,1,-nbitq), 
to_sfixed(-1331.0/65536.0,1,-nbitq), 
to_sfixed(1780.0/65536.0,1,-nbitq), 
to_sfixed(-1643.0/65536.0,1,-nbitq), 
to_sfixed(-1864.0/65536.0,1,-nbitq), 
to_sfixed(769.0/65536.0,1,-nbitq), 
to_sfixed(5422.0/65536.0,1,-nbitq), 
to_sfixed(-569.0/65536.0,1,-nbitq), 
to_sfixed(1572.0/65536.0,1,-nbitq), 
to_sfixed(651.0/65536.0,1,-nbitq), 
to_sfixed(1292.0/65536.0,1,-nbitq), 
to_sfixed(-1964.0/65536.0,1,-nbitq), 
to_sfixed(1544.0/65536.0,1,-nbitq), 
to_sfixed(-1395.0/65536.0,1,-nbitq), 
to_sfixed(-2767.0/65536.0,1,-nbitq), 
to_sfixed(201.0/65536.0,1,-nbitq), 
to_sfixed(-1382.0/65536.0,1,-nbitq), 
to_sfixed(1234.0/65536.0,1,-nbitq), 
to_sfixed(-1352.0/65536.0,1,-nbitq), 
to_sfixed(-22.0/65536.0,1,-nbitq), 
to_sfixed(2235.0/65536.0,1,-nbitq), 
to_sfixed(-1157.0/65536.0,1,-nbitq), 
to_sfixed(2464.0/65536.0,1,-nbitq), 
to_sfixed(1443.0/65536.0,1,-nbitq), 
to_sfixed(1720.0/65536.0,1,-nbitq), 
to_sfixed(-999.0/65536.0,1,-nbitq), 
to_sfixed(3663.0/65536.0,1,-nbitq), 
to_sfixed(413.0/65536.0,1,-nbitq), 
to_sfixed(-1307.0/65536.0,1,-nbitq), 
to_sfixed(2239.0/65536.0,1,-nbitq), 
to_sfixed(1963.0/65536.0,1,-nbitq), 
to_sfixed(204.0/65536.0,1,-nbitq), 
to_sfixed(1373.0/65536.0,1,-nbitq), 
to_sfixed(-479.0/65536.0,1,-nbitq), 
to_sfixed(740.0/65536.0,1,-nbitq), 
to_sfixed(-1994.0/65536.0,1,-nbitq), 
to_sfixed(2275.0/65536.0,1,-nbitq), 
to_sfixed(3055.0/65536.0,1,-nbitq), 
to_sfixed(5244.0/65536.0,1,-nbitq), 
to_sfixed(1508.0/65536.0,1,-nbitq), 
to_sfixed(3199.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-534.0/65536.0,1,-nbitq), 
to_sfixed(-1701.0/65536.0,1,-nbitq), 
to_sfixed(3253.0/65536.0,1,-nbitq), 
to_sfixed(4121.0/65536.0,1,-nbitq), 
to_sfixed(-825.0/65536.0,1,-nbitq), 
to_sfixed(-1565.0/65536.0,1,-nbitq), 
to_sfixed(-2696.0/65536.0,1,-nbitq), 
to_sfixed(1164.0/65536.0,1,-nbitq), 
to_sfixed(-1253.0/65536.0,1,-nbitq), 
to_sfixed(3104.0/65536.0,1,-nbitq), 
to_sfixed(2951.0/65536.0,1,-nbitq), 
to_sfixed(1992.0/65536.0,1,-nbitq), 
to_sfixed(-584.0/65536.0,1,-nbitq), 
to_sfixed(2361.0/65536.0,1,-nbitq), 
to_sfixed(-203.0/65536.0,1,-nbitq), 
to_sfixed(-1856.0/65536.0,1,-nbitq), 
to_sfixed(2391.0/65536.0,1,-nbitq), 
to_sfixed(802.0/65536.0,1,-nbitq), 
to_sfixed(-1875.0/65536.0,1,-nbitq), 
to_sfixed(515.0/65536.0,1,-nbitq), 
to_sfixed(2855.0/65536.0,1,-nbitq), 
to_sfixed(213.0/65536.0,1,-nbitq), 
to_sfixed(-4001.0/65536.0,1,-nbitq), 
to_sfixed(3567.0/65536.0,1,-nbitq), 
to_sfixed(-1681.0/65536.0,1,-nbitq), 
to_sfixed(4500.0/65536.0,1,-nbitq), 
to_sfixed(775.0/65536.0,1,-nbitq), 
to_sfixed(2089.0/65536.0,1,-nbitq), 
to_sfixed(549.0/65536.0,1,-nbitq), 
to_sfixed(-2859.0/65536.0,1,-nbitq), 
to_sfixed(823.0/65536.0,1,-nbitq), 
to_sfixed(3458.0/65536.0,1,-nbitq), 
to_sfixed(1013.0/65536.0,1,-nbitq), 
to_sfixed(5692.0/65536.0,1,-nbitq), 
to_sfixed(1318.0/65536.0,1,-nbitq), 
to_sfixed(-1766.0/65536.0,1,-nbitq), 
to_sfixed(-3385.0/65536.0,1,-nbitq), 
to_sfixed(-2215.0/65536.0,1,-nbitq), 
to_sfixed(-4944.0/65536.0,1,-nbitq), 
to_sfixed(-1300.0/65536.0,1,-nbitq), 
to_sfixed(-4462.0/65536.0,1,-nbitq), 
to_sfixed(-890.0/65536.0,1,-nbitq), 
to_sfixed(32.0/65536.0,1,-nbitq), 
to_sfixed(939.0/65536.0,1,-nbitq), 
to_sfixed(-877.0/65536.0,1,-nbitq), 
to_sfixed(2083.0/65536.0,1,-nbitq), 
to_sfixed(335.0/65536.0,1,-nbitq), 
to_sfixed(2528.0/65536.0,1,-nbitq), 
to_sfixed(1442.0/65536.0,1,-nbitq), 
to_sfixed(4155.0/65536.0,1,-nbitq), 
to_sfixed(-658.0/65536.0,1,-nbitq), 
to_sfixed(-2053.0/65536.0,1,-nbitq), 
to_sfixed(2060.0/65536.0,1,-nbitq), 
to_sfixed(-2488.0/65536.0,1,-nbitq), 
to_sfixed(-426.0/65536.0,1,-nbitq), 
to_sfixed(663.0/65536.0,1,-nbitq), 
to_sfixed(-984.0/65536.0,1,-nbitq), 
to_sfixed(2798.0/65536.0,1,-nbitq), 
to_sfixed(2660.0/65536.0,1,-nbitq), 
to_sfixed(2368.0/65536.0,1,-nbitq), 
to_sfixed(1368.0/65536.0,1,-nbitq), 
to_sfixed(-1525.0/65536.0,1,-nbitq), 
to_sfixed(3065.0/65536.0,1,-nbitq), 
to_sfixed(2213.0/65536.0,1,-nbitq), 
to_sfixed(-3505.0/65536.0,1,-nbitq), 
to_sfixed(3168.0/65536.0,1,-nbitq), 
to_sfixed(-2752.0/65536.0,1,-nbitq), 
to_sfixed(440.0/65536.0,1,-nbitq), 
to_sfixed(-120.0/65536.0,1,-nbitq), 
to_sfixed(2449.0/65536.0,1,-nbitq), 
to_sfixed(862.0/65536.0,1,-nbitq), 
to_sfixed(-325.0/65536.0,1,-nbitq), 
to_sfixed(1807.0/65536.0,1,-nbitq), 
to_sfixed(1411.0/65536.0,1,-nbitq), 
to_sfixed(-1875.0/65536.0,1,-nbitq), 
to_sfixed(6838.0/65536.0,1,-nbitq), 
to_sfixed(-3688.0/65536.0,1,-nbitq), 
to_sfixed(2003.0/65536.0,1,-nbitq), 
to_sfixed(2037.0/65536.0,1,-nbitq), 
to_sfixed(2597.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-904.0/65536.0,1,-nbitq), 
to_sfixed(2238.0/65536.0,1,-nbitq), 
to_sfixed(-1204.0/65536.0,1,-nbitq), 
to_sfixed(3999.0/65536.0,1,-nbitq), 
to_sfixed(2132.0/65536.0,1,-nbitq), 
to_sfixed(-8.0/65536.0,1,-nbitq), 
to_sfixed(-657.0/65536.0,1,-nbitq), 
to_sfixed(94.0/65536.0,1,-nbitq), 
to_sfixed(920.0/65536.0,1,-nbitq), 
to_sfixed(143.0/65536.0,1,-nbitq), 
to_sfixed(1922.0/65536.0,1,-nbitq), 
to_sfixed(4537.0/65536.0,1,-nbitq), 
to_sfixed(288.0/65536.0,1,-nbitq), 
to_sfixed(-411.0/65536.0,1,-nbitq), 
to_sfixed(4621.0/65536.0,1,-nbitq), 
to_sfixed(2298.0/65536.0,1,-nbitq), 
to_sfixed(-1294.0/65536.0,1,-nbitq), 
to_sfixed(-3131.0/65536.0,1,-nbitq), 
to_sfixed(2428.0/65536.0,1,-nbitq), 
to_sfixed(-2513.0/65536.0,1,-nbitq), 
to_sfixed(3017.0/65536.0,1,-nbitq), 
to_sfixed(-526.0/65536.0,1,-nbitq), 
to_sfixed(-5847.0/65536.0,1,-nbitq), 
to_sfixed(-3869.0/65536.0,1,-nbitq), 
to_sfixed(-490.0/65536.0,1,-nbitq), 
to_sfixed(2552.0/65536.0,1,-nbitq), 
to_sfixed(1148.0/65536.0,1,-nbitq), 
to_sfixed(218.0/65536.0,1,-nbitq), 
to_sfixed(4018.0/65536.0,1,-nbitq), 
to_sfixed(3370.0/65536.0,1,-nbitq), 
to_sfixed(-2195.0/65536.0,1,-nbitq), 
to_sfixed(1633.0/65536.0,1,-nbitq), 
to_sfixed(845.0/65536.0,1,-nbitq), 
to_sfixed(1812.0/65536.0,1,-nbitq), 
to_sfixed(33.0/65536.0,1,-nbitq), 
to_sfixed(-2640.0/65536.0,1,-nbitq), 
to_sfixed(-3009.0/65536.0,1,-nbitq), 
to_sfixed(3229.0/65536.0,1,-nbitq), 
to_sfixed(-1519.0/65536.0,1,-nbitq), 
to_sfixed(3232.0/65536.0,1,-nbitq), 
to_sfixed(-8394.0/65536.0,1,-nbitq), 
to_sfixed(-2473.0/65536.0,1,-nbitq), 
to_sfixed(8072.0/65536.0,1,-nbitq), 
to_sfixed(2355.0/65536.0,1,-nbitq), 
to_sfixed(-782.0/65536.0,1,-nbitq), 
to_sfixed(7218.0/65536.0,1,-nbitq), 
to_sfixed(559.0/65536.0,1,-nbitq), 
to_sfixed(-3805.0/65536.0,1,-nbitq), 
to_sfixed(-875.0/65536.0,1,-nbitq), 
to_sfixed(263.0/65536.0,1,-nbitq), 
to_sfixed(2240.0/65536.0,1,-nbitq), 
to_sfixed(-3673.0/65536.0,1,-nbitq), 
to_sfixed(2556.0/65536.0,1,-nbitq), 
to_sfixed(-1582.0/65536.0,1,-nbitq), 
to_sfixed(-2679.0/65536.0,1,-nbitq), 
to_sfixed(2082.0/65536.0,1,-nbitq), 
to_sfixed(-2260.0/65536.0,1,-nbitq), 
to_sfixed(2415.0/65536.0,1,-nbitq), 
to_sfixed(1639.0/65536.0,1,-nbitq), 
to_sfixed(1256.0/65536.0,1,-nbitq), 
to_sfixed(532.0/65536.0,1,-nbitq), 
to_sfixed(1499.0/65536.0,1,-nbitq), 
to_sfixed(-1855.0/65536.0,1,-nbitq), 
to_sfixed(-3105.0/65536.0,1,-nbitq), 
to_sfixed(-3752.0/65536.0,1,-nbitq), 
to_sfixed(2015.0/65536.0,1,-nbitq), 
to_sfixed(-24.0/65536.0,1,-nbitq), 
to_sfixed(1129.0/65536.0,1,-nbitq), 
to_sfixed(-691.0/65536.0,1,-nbitq), 
to_sfixed(-659.0/65536.0,1,-nbitq), 
to_sfixed(384.0/65536.0,1,-nbitq), 
to_sfixed(2237.0/65536.0,1,-nbitq), 
to_sfixed(-148.0/65536.0,1,-nbitq), 
to_sfixed(2503.0/65536.0,1,-nbitq), 
to_sfixed(97.0/65536.0,1,-nbitq), 
to_sfixed(7541.0/65536.0,1,-nbitq), 
to_sfixed(-2547.0/65536.0,1,-nbitq), 
to_sfixed(5549.0/65536.0,1,-nbitq), 
to_sfixed(146.0/65536.0,1,-nbitq), 
to_sfixed(21.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-717.0/65536.0,1,-nbitq), 
to_sfixed(-652.0/65536.0,1,-nbitq), 
to_sfixed(946.0/65536.0,1,-nbitq), 
to_sfixed(6555.0/65536.0,1,-nbitq), 
to_sfixed(743.0/65536.0,1,-nbitq), 
to_sfixed(414.0/65536.0,1,-nbitq), 
to_sfixed(-744.0/65536.0,1,-nbitq), 
to_sfixed(1397.0/65536.0,1,-nbitq), 
to_sfixed(2037.0/65536.0,1,-nbitq), 
to_sfixed(-1217.0/65536.0,1,-nbitq), 
to_sfixed(-1031.0/65536.0,1,-nbitq), 
to_sfixed(18216.0/65536.0,1,-nbitq), 
to_sfixed(751.0/65536.0,1,-nbitq), 
to_sfixed(1981.0/65536.0,1,-nbitq), 
to_sfixed(5260.0/65536.0,1,-nbitq), 
to_sfixed(-1190.0/65536.0,1,-nbitq), 
to_sfixed(828.0/65536.0,1,-nbitq), 
to_sfixed(-6307.0/65536.0,1,-nbitq), 
to_sfixed(5365.0/65536.0,1,-nbitq), 
to_sfixed(211.0/65536.0,1,-nbitq), 
to_sfixed(5225.0/65536.0,1,-nbitq), 
to_sfixed(2139.0/65536.0,1,-nbitq), 
to_sfixed(-3201.0/65536.0,1,-nbitq), 
to_sfixed(-7382.0/65536.0,1,-nbitq), 
to_sfixed(-4878.0/65536.0,1,-nbitq), 
to_sfixed(3231.0/65536.0,1,-nbitq), 
to_sfixed(2898.0/65536.0,1,-nbitq), 
to_sfixed(-2144.0/65536.0,1,-nbitq), 
to_sfixed(3792.0/65536.0,1,-nbitq), 
to_sfixed(1775.0/65536.0,1,-nbitq), 
to_sfixed(-1166.0/65536.0,1,-nbitq), 
to_sfixed(2656.0/65536.0,1,-nbitq), 
to_sfixed(2223.0/65536.0,1,-nbitq), 
to_sfixed(-534.0/65536.0,1,-nbitq), 
to_sfixed(-1925.0/65536.0,1,-nbitq), 
to_sfixed(-1999.0/65536.0,1,-nbitq), 
to_sfixed(-5452.0/65536.0,1,-nbitq), 
to_sfixed(3007.0/65536.0,1,-nbitq), 
to_sfixed(-2104.0/65536.0,1,-nbitq), 
to_sfixed(-2273.0/65536.0,1,-nbitq), 
to_sfixed(-11602.0/65536.0,1,-nbitq), 
to_sfixed(-197.0/65536.0,1,-nbitq), 
to_sfixed(11746.0/65536.0,1,-nbitq), 
to_sfixed(1085.0/65536.0,1,-nbitq), 
to_sfixed(-1703.0/65536.0,1,-nbitq), 
to_sfixed(3695.0/65536.0,1,-nbitq), 
to_sfixed(-589.0/65536.0,1,-nbitq), 
to_sfixed(-2039.0/65536.0,1,-nbitq), 
to_sfixed(2650.0/65536.0,1,-nbitq), 
to_sfixed(5504.0/65536.0,1,-nbitq), 
to_sfixed(3082.0/65536.0,1,-nbitq), 
to_sfixed(-3175.0/65536.0,1,-nbitq), 
to_sfixed(2342.0/65536.0,1,-nbitq), 
to_sfixed(3471.0/65536.0,1,-nbitq), 
to_sfixed(-1644.0/65536.0,1,-nbitq), 
to_sfixed(6187.0/65536.0,1,-nbitq), 
to_sfixed(-359.0/65536.0,1,-nbitq), 
to_sfixed(776.0/65536.0,1,-nbitq), 
to_sfixed(-2040.0/65536.0,1,-nbitq), 
to_sfixed(-2983.0/65536.0,1,-nbitq), 
to_sfixed(-2697.0/65536.0,1,-nbitq), 
to_sfixed(481.0/65536.0,1,-nbitq), 
to_sfixed(-125.0/65536.0,1,-nbitq), 
to_sfixed(430.0/65536.0,1,-nbitq), 
to_sfixed(-93.0/65536.0,1,-nbitq), 
to_sfixed(2043.0/65536.0,1,-nbitq), 
to_sfixed(-1135.0/65536.0,1,-nbitq), 
to_sfixed(-5592.0/65536.0,1,-nbitq), 
to_sfixed(-7125.0/65536.0,1,-nbitq), 
to_sfixed(215.0/65536.0,1,-nbitq), 
to_sfixed(2424.0/65536.0,1,-nbitq), 
to_sfixed(-1449.0/65536.0,1,-nbitq), 
to_sfixed(-4082.0/65536.0,1,-nbitq), 
to_sfixed(-654.0/65536.0,1,-nbitq), 
to_sfixed(-1234.0/65536.0,1,-nbitq), 
to_sfixed(769.0/65536.0,1,-nbitq), 
to_sfixed(1384.0/65536.0,1,-nbitq), 
to_sfixed(4482.0/65536.0,1,-nbitq), 
to_sfixed(935.0/65536.0,1,-nbitq), 
to_sfixed(-1668.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2147.0/65536.0,1,-nbitq), 
to_sfixed(-2971.0/65536.0,1,-nbitq), 
to_sfixed(5731.0/65536.0,1,-nbitq), 
to_sfixed(2295.0/65536.0,1,-nbitq), 
to_sfixed(-1407.0/65536.0,1,-nbitq), 
to_sfixed(-698.0/65536.0,1,-nbitq), 
to_sfixed(-1392.0/65536.0,1,-nbitq), 
to_sfixed(-1562.0/65536.0,1,-nbitq), 
to_sfixed(-2482.0/65536.0,1,-nbitq), 
to_sfixed(970.0/65536.0,1,-nbitq), 
to_sfixed(5050.0/65536.0,1,-nbitq), 
to_sfixed(18467.0/65536.0,1,-nbitq), 
to_sfixed(-2499.0/65536.0,1,-nbitq), 
to_sfixed(-170.0/65536.0,1,-nbitq), 
to_sfixed(3820.0/65536.0,1,-nbitq), 
to_sfixed(2912.0/65536.0,1,-nbitq), 
to_sfixed(-2504.0/65536.0,1,-nbitq), 
to_sfixed(-8524.0/65536.0,1,-nbitq), 
to_sfixed(3991.0/65536.0,1,-nbitq), 
to_sfixed(-1605.0/65536.0,1,-nbitq), 
to_sfixed(7305.0/65536.0,1,-nbitq), 
to_sfixed(431.0/65536.0,1,-nbitq), 
to_sfixed(-450.0/65536.0,1,-nbitq), 
to_sfixed(-4329.0/65536.0,1,-nbitq), 
to_sfixed(-1412.0/65536.0,1,-nbitq), 
to_sfixed(2453.0/65536.0,1,-nbitq), 
to_sfixed(-2481.0/65536.0,1,-nbitq), 
to_sfixed(2021.0/65536.0,1,-nbitq), 
to_sfixed(1940.0/65536.0,1,-nbitq), 
to_sfixed(6080.0/65536.0,1,-nbitq), 
to_sfixed(1738.0/65536.0,1,-nbitq), 
to_sfixed(2442.0/65536.0,1,-nbitq), 
to_sfixed(4822.0/65536.0,1,-nbitq), 
to_sfixed(-136.0/65536.0,1,-nbitq), 
to_sfixed(-1251.0/65536.0,1,-nbitq), 
to_sfixed(1625.0/65536.0,1,-nbitq), 
to_sfixed(-6904.0/65536.0,1,-nbitq), 
to_sfixed(-1383.0/65536.0,1,-nbitq), 
to_sfixed(3889.0/65536.0,1,-nbitq), 
to_sfixed(-5091.0/65536.0,1,-nbitq), 
to_sfixed(-14035.0/65536.0,1,-nbitq), 
to_sfixed(410.0/65536.0,1,-nbitq), 
to_sfixed(10448.0/65536.0,1,-nbitq), 
to_sfixed(-2216.0/65536.0,1,-nbitq), 
to_sfixed(3276.0/65536.0,1,-nbitq), 
to_sfixed(-3829.0/65536.0,1,-nbitq), 
to_sfixed(-445.0/65536.0,1,-nbitq), 
to_sfixed(-1936.0/65536.0,1,-nbitq), 
to_sfixed(3902.0/65536.0,1,-nbitq), 
to_sfixed(-514.0/65536.0,1,-nbitq), 
to_sfixed(-2002.0/65536.0,1,-nbitq), 
to_sfixed(-4374.0/65536.0,1,-nbitq), 
to_sfixed(1822.0/65536.0,1,-nbitq), 
to_sfixed(2644.0/65536.0,1,-nbitq), 
to_sfixed(-3225.0/65536.0,1,-nbitq), 
to_sfixed(4052.0/65536.0,1,-nbitq), 
to_sfixed(1649.0/65536.0,1,-nbitq), 
to_sfixed(338.0/65536.0,1,-nbitq), 
to_sfixed(-87.0/65536.0,1,-nbitq), 
to_sfixed(-3367.0/65536.0,1,-nbitq), 
to_sfixed(-1277.0/65536.0,1,-nbitq), 
to_sfixed(-326.0/65536.0,1,-nbitq), 
to_sfixed(-808.0/65536.0,1,-nbitq), 
to_sfixed(-3284.0/65536.0,1,-nbitq), 
to_sfixed(-1650.0/65536.0,1,-nbitq), 
to_sfixed(3359.0/65536.0,1,-nbitq), 
to_sfixed(-4843.0/65536.0,1,-nbitq), 
to_sfixed(-9098.0/65536.0,1,-nbitq), 
to_sfixed(-7069.0/65536.0,1,-nbitq), 
to_sfixed(-7426.0/65536.0,1,-nbitq), 
to_sfixed(2315.0/65536.0,1,-nbitq), 
to_sfixed(-4292.0/65536.0,1,-nbitq), 
to_sfixed(-4892.0/65536.0,1,-nbitq), 
to_sfixed(574.0/65536.0,1,-nbitq), 
to_sfixed(-2493.0/65536.0,1,-nbitq), 
to_sfixed(1276.0/65536.0,1,-nbitq), 
to_sfixed(2377.0/65536.0,1,-nbitq), 
to_sfixed(718.0/65536.0,1,-nbitq), 
to_sfixed(-1789.0/65536.0,1,-nbitq), 
to_sfixed(-2362.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3524.0/65536.0,1,-nbitq), 
to_sfixed(-373.0/65536.0,1,-nbitq), 
to_sfixed(3546.0/65536.0,1,-nbitq), 
to_sfixed(2922.0/65536.0,1,-nbitq), 
to_sfixed(-6079.0/65536.0,1,-nbitq), 
to_sfixed(3008.0/65536.0,1,-nbitq), 
to_sfixed(4088.0/65536.0,1,-nbitq), 
to_sfixed(5675.0/65536.0,1,-nbitq), 
to_sfixed(3267.0/65536.0,1,-nbitq), 
to_sfixed(-932.0/65536.0,1,-nbitq), 
to_sfixed(7489.0/65536.0,1,-nbitq), 
to_sfixed(11578.0/65536.0,1,-nbitq), 
to_sfixed(-1744.0/65536.0,1,-nbitq), 
to_sfixed(-2664.0/65536.0,1,-nbitq), 
to_sfixed(-1111.0/65536.0,1,-nbitq), 
to_sfixed(2260.0/65536.0,1,-nbitq), 
to_sfixed(-1017.0/65536.0,1,-nbitq), 
to_sfixed(-2396.0/65536.0,1,-nbitq), 
to_sfixed(-1310.0/65536.0,1,-nbitq), 
to_sfixed(-1448.0/65536.0,1,-nbitq), 
to_sfixed(6416.0/65536.0,1,-nbitq), 
to_sfixed(-2361.0/65536.0,1,-nbitq), 
to_sfixed(-1543.0/65536.0,1,-nbitq), 
to_sfixed(587.0/65536.0,1,-nbitq), 
to_sfixed(2490.0/65536.0,1,-nbitq), 
to_sfixed(2359.0/65536.0,1,-nbitq), 
to_sfixed(-6032.0/65536.0,1,-nbitq), 
to_sfixed(-327.0/65536.0,1,-nbitq), 
to_sfixed(519.0/65536.0,1,-nbitq), 
to_sfixed(7002.0/65536.0,1,-nbitq), 
to_sfixed(217.0/65536.0,1,-nbitq), 
to_sfixed(4455.0/65536.0,1,-nbitq), 
to_sfixed(7046.0/65536.0,1,-nbitq), 
to_sfixed(1149.0/65536.0,1,-nbitq), 
to_sfixed(-2877.0/65536.0,1,-nbitq), 
to_sfixed(-1013.0/65536.0,1,-nbitq), 
to_sfixed(-9736.0/65536.0,1,-nbitq), 
to_sfixed(2165.0/65536.0,1,-nbitq), 
to_sfixed(2648.0/65536.0,1,-nbitq), 
to_sfixed(-4928.0/65536.0,1,-nbitq), 
to_sfixed(-16097.0/65536.0,1,-nbitq), 
to_sfixed(-1914.0/65536.0,1,-nbitq), 
to_sfixed(12357.0/65536.0,1,-nbitq), 
to_sfixed(-2631.0/65536.0,1,-nbitq), 
to_sfixed(-1376.0/65536.0,1,-nbitq), 
to_sfixed(-11140.0/65536.0,1,-nbitq), 
to_sfixed(172.0/65536.0,1,-nbitq), 
to_sfixed(1258.0/65536.0,1,-nbitq), 
to_sfixed(-461.0/65536.0,1,-nbitq), 
to_sfixed(734.0/65536.0,1,-nbitq), 
to_sfixed(1527.0/65536.0,1,-nbitq), 
to_sfixed(-60.0/65536.0,1,-nbitq), 
to_sfixed(262.0/65536.0,1,-nbitq), 
to_sfixed(6040.0/65536.0,1,-nbitq), 
to_sfixed(-4432.0/65536.0,1,-nbitq), 
to_sfixed(2719.0/65536.0,1,-nbitq), 
to_sfixed(-1340.0/65536.0,1,-nbitq), 
to_sfixed(-133.0/65536.0,1,-nbitq), 
to_sfixed(933.0/65536.0,1,-nbitq), 
to_sfixed(923.0/65536.0,1,-nbitq), 
to_sfixed(329.0/65536.0,1,-nbitq), 
to_sfixed(-1642.0/65536.0,1,-nbitq), 
to_sfixed(-1444.0/65536.0,1,-nbitq), 
to_sfixed(581.0/65536.0,1,-nbitq), 
to_sfixed(-279.0/65536.0,1,-nbitq), 
to_sfixed(3837.0/65536.0,1,-nbitq), 
to_sfixed(-2179.0/65536.0,1,-nbitq), 
to_sfixed(-6444.0/65536.0,1,-nbitq), 
to_sfixed(-42.0/65536.0,1,-nbitq), 
to_sfixed(6001.0/65536.0,1,-nbitq), 
to_sfixed(878.0/65536.0,1,-nbitq), 
to_sfixed(2550.0/65536.0,1,-nbitq), 
to_sfixed(-1854.0/65536.0,1,-nbitq), 
to_sfixed(-3217.0/65536.0,1,-nbitq), 
to_sfixed(537.0/65536.0,1,-nbitq), 
to_sfixed(-443.0/65536.0,1,-nbitq), 
to_sfixed(-1398.0/65536.0,1,-nbitq), 
to_sfixed(957.0/65536.0,1,-nbitq), 
to_sfixed(355.0/65536.0,1,-nbitq), 
to_sfixed(2759.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3067.0/65536.0,1,-nbitq), 
to_sfixed(513.0/65536.0,1,-nbitq), 
to_sfixed(6605.0/65536.0,1,-nbitq), 
to_sfixed(3168.0/65536.0,1,-nbitq), 
to_sfixed(3026.0/65536.0,1,-nbitq), 
to_sfixed(-3272.0/65536.0,1,-nbitq), 
to_sfixed(3387.0/65536.0,1,-nbitq), 
to_sfixed(-2284.0/65536.0,1,-nbitq), 
to_sfixed(1492.0/65536.0,1,-nbitq), 
to_sfixed(665.0/65536.0,1,-nbitq), 
to_sfixed(5862.0/65536.0,1,-nbitq), 
to_sfixed(310.0/65536.0,1,-nbitq), 
to_sfixed(1147.0/65536.0,1,-nbitq), 
to_sfixed(5449.0/65536.0,1,-nbitq), 
to_sfixed(4290.0/65536.0,1,-nbitq), 
to_sfixed(-878.0/65536.0,1,-nbitq), 
to_sfixed(1742.0/65536.0,1,-nbitq), 
to_sfixed(4458.0/65536.0,1,-nbitq), 
to_sfixed(4202.0/65536.0,1,-nbitq), 
to_sfixed(-2214.0/65536.0,1,-nbitq), 
to_sfixed(2275.0/65536.0,1,-nbitq), 
to_sfixed(-801.0/65536.0,1,-nbitq), 
to_sfixed(3221.0/65536.0,1,-nbitq), 
to_sfixed(-4353.0/65536.0,1,-nbitq), 
to_sfixed(1010.0/65536.0,1,-nbitq), 
to_sfixed(-103.0/65536.0,1,-nbitq), 
to_sfixed(-3934.0/65536.0,1,-nbitq), 
to_sfixed(-2041.0/65536.0,1,-nbitq), 
to_sfixed(-908.0/65536.0,1,-nbitq), 
to_sfixed(3476.0/65536.0,1,-nbitq), 
to_sfixed(-2720.0/65536.0,1,-nbitq), 
to_sfixed(5868.0/65536.0,1,-nbitq), 
to_sfixed(6899.0/65536.0,1,-nbitq), 
to_sfixed(3396.0/65536.0,1,-nbitq), 
to_sfixed(-832.0/65536.0,1,-nbitq), 
to_sfixed(2702.0/65536.0,1,-nbitq), 
to_sfixed(3293.0/65536.0,1,-nbitq), 
to_sfixed(-986.0/65536.0,1,-nbitq), 
to_sfixed(-1501.0/65536.0,1,-nbitq), 
to_sfixed(-877.0/65536.0,1,-nbitq), 
to_sfixed(-6785.0/65536.0,1,-nbitq), 
to_sfixed(1176.0/65536.0,1,-nbitq), 
to_sfixed(7396.0/65536.0,1,-nbitq), 
to_sfixed(-1808.0/65536.0,1,-nbitq), 
to_sfixed(-782.0/65536.0,1,-nbitq), 
to_sfixed(-16794.0/65536.0,1,-nbitq), 
to_sfixed(1638.0/65536.0,1,-nbitq), 
to_sfixed(1528.0/65536.0,1,-nbitq), 
to_sfixed(3328.0/65536.0,1,-nbitq), 
to_sfixed(2260.0/65536.0,1,-nbitq), 
to_sfixed(-380.0/65536.0,1,-nbitq), 
to_sfixed(-2311.0/65536.0,1,-nbitq), 
to_sfixed(1600.0/65536.0,1,-nbitq), 
to_sfixed(8316.0/65536.0,1,-nbitq), 
to_sfixed(-5527.0/65536.0,1,-nbitq), 
to_sfixed(6541.0/65536.0,1,-nbitq), 
to_sfixed(1364.0/65536.0,1,-nbitq), 
to_sfixed(3059.0/65536.0,1,-nbitq), 
to_sfixed(-2698.0/65536.0,1,-nbitq), 
to_sfixed(2360.0/65536.0,1,-nbitq), 
to_sfixed(1114.0/65536.0,1,-nbitq), 
to_sfixed(1262.0/65536.0,1,-nbitq), 
to_sfixed(1238.0/65536.0,1,-nbitq), 
to_sfixed(781.0/65536.0,1,-nbitq), 
to_sfixed(-4334.0/65536.0,1,-nbitq), 
to_sfixed(10820.0/65536.0,1,-nbitq), 
to_sfixed(-1403.0/65536.0,1,-nbitq), 
to_sfixed(-6993.0/65536.0,1,-nbitq), 
to_sfixed(3276.0/65536.0,1,-nbitq), 
to_sfixed(463.0/65536.0,1,-nbitq), 
to_sfixed(-1840.0/65536.0,1,-nbitq), 
to_sfixed(5041.0/65536.0,1,-nbitq), 
to_sfixed(-2544.0/65536.0,1,-nbitq), 
to_sfixed(2140.0/65536.0,1,-nbitq), 
to_sfixed(-2207.0/65536.0,1,-nbitq), 
to_sfixed(6426.0/65536.0,1,-nbitq), 
to_sfixed(3794.0/65536.0,1,-nbitq), 
to_sfixed(802.0/65536.0,1,-nbitq), 
to_sfixed(-2215.0/65536.0,1,-nbitq), 
to_sfixed(-564.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1445.0/65536.0,1,-nbitq), 
to_sfixed(-1097.0/65536.0,1,-nbitq), 
to_sfixed(6705.0/65536.0,1,-nbitq), 
to_sfixed(2181.0/65536.0,1,-nbitq), 
to_sfixed(-2691.0/65536.0,1,-nbitq), 
to_sfixed(-4020.0/65536.0,1,-nbitq), 
to_sfixed(19.0/65536.0,1,-nbitq), 
to_sfixed(-1540.0/65536.0,1,-nbitq), 
to_sfixed(-129.0/65536.0,1,-nbitq), 
to_sfixed(-487.0/65536.0,1,-nbitq), 
to_sfixed(7293.0/65536.0,1,-nbitq), 
to_sfixed(4797.0/65536.0,1,-nbitq), 
to_sfixed(4817.0/65536.0,1,-nbitq), 
to_sfixed(1677.0/65536.0,1,-nbitq), 
to_sfixed(8527.0/65536.0,1,-nbitq), 
to_sfixed(-1614.0/65536.0,1,-nbitq), 
to_sfixed(-645.0/65536.0,1,-nbitq), 
to_sfixed(371.0/65536.0,1,-nbitq), 
to_sfixed(8214.0/65536.0,1,-nbitq), 
to_sfixed(-1805.0/65536.0,1,-nbitq), 
to_sfixed(5590.0/65536.0,1,-nbitq), 
to_sfixed(-5454.0/65536.0,1,-nbitq), 
to_sfixed(4255.0/65536.0,1,-nbitq), 
to_sfixed(302.0/65536.0,1,-nbitq), 
to_sfixed(226.0/65536.0,1,-nbitq), 
to_sfixed(-5213.0/65536.0,1,-nbitq), 
to_sfixed(-1383.0/65536.0,1,-nbitq), 
to_sfixed(-786.0/65536.0,1,-nbitq), 
to_sfixed(-2293.0/65536.0,1,-nbitq), 
to_sfixed(6248.0/65536.0,1,-nbitq), 
to_sfixed(486.0/65536.0,1,-nbitq), 
to_sfixed(8664.0/65536.0,1,-nbitq), 
to_sfixed(3741.0/65536.0,1,-nbitq), 
to_sfixed(4122.0/65536.0,1,-nbitq), 
to_sfixed(-2242.0/65536.0,1,-nbitq), 
to_sfixed(1960.0/65536.0,1,-nbitq), 
to_sfixed(11597.0/65536.0,1,-nbitq), 
to_sfixed(-7117.0/65536.0,1,-nbitq), 
to_sfixed(-3607.0/65536.0,1,-nbitq), 
to_sfixed(2620.0/65536.0,1,-nbitq), 
to_sfixed(-2115.0/65536.0,1,-nbitq), 
to_sfixed(-336.0/65536.0,1,-nbitq), 
to_sfixed(9053.0/65536.0,1,-nbitq), 
to_sfixed(-4782.0/65536.0,1,-nbitq), 
to_sfixed(1862.0/65536.0,1,-nbitq), 
to_sfixed(-20155.0/65536.0,1,-nbitq), 
to_sfixed(-3719.0/65536.0,1,-nbitq), 
to_sfixed(-1242.0/65536.0,1,-nbitq), 
to_sfixed(2715.0/65536.0,1,-nbitq), 
to_sfixed(3337.0/65536.0,1,-nbitq), 
to_sfixed(1384.0/65536.0,1,-nbitq), 
to_sfixed(-1826.0/65536.0,1,-nbitq), 
to_sfixed(1925.0/65536.0,1,-nbitq), 
to_sfixed(5489.0/65536.0,1,-nbitq), 
to_sfixed(-1883.0/65536.0,1,-nbitq), 
to_sfixed(4393.0/65536.0,1,-nbitq), 
to_sfixed(999.0/65536.0,1,-nbitq), 
to_sfixed(1598.0/65536.0,1,-nbitq), 
to_sfixed(1249.0/65536.0,1,-nbitq), 
to_sfixed(-3372.0/65536.0,1,-nbitq), 
to_sfixed(2068.0/65536.0,1,-nbitq), 
to_sfixed(-1228.0/65536.0,1,-nbitq), 
to_sfixed(-1525.0/65536.0,1,-nbitq), 
to_sfixed(-945.0/65536.0,1,-nbitq), 
to_sfixed(-1555.0/65536.0,1,-nbitq), 
to_sfixed(7888.0/65536.0,1,-nbitq), 
to_sfixed(-4815.0/65536.0,1,-nbitq), 
to_sfixed(-10431.0/65536.0,1,-nbitq), 
to_sfixed(-784.0/65536.0,1,-nbitq), 
to_sfixed(4693.0/65536.0,1,-nbitq), 
to_sfixed(-4456.0/65536.0,1,-nbitq), 
to_sfixed(11096.0/65536.0,1,-nbitq), 
to_sfixed(-5288.0/65536.0,1,-nbitq), 
to_sfixed(-864.0/65536.0,1,-nbitq), 
to_sfixed(-801.0/65536.0,1,-nbitq), 
to_sfixed(5602.0/65536.0,1,-nbitq), 
to_sfixed(-1220.0/65536.0,1,-nbitq), 
to_sfixed(-3727.0/65536.0,1,-nbitq), 
to_sfixed(-1572.0/65536.0,1,-nbitq), 
to_sfixed(-3918.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1939.0/65536.0,1,-nbitq), 
to_sfixed(-1127.0/65536.0,1,-nbitq), 
to_sfixed(-8972.0/65536.0,1,-nbitq), 
to_sfixed(5026.0/65536.0,1,-nbitq), 
to_sfixed(3608.0/65536.0,1,-nbitq), 
to_sfixed(-7303.0/65536.0,1,-nbitq), 
to_sfixed(1027.0/65536.0,1,-nbitq), 
to_sfixed(846.0/65536.0,1,-nbitq), 
to_sfixed(-1997.0/65536.0,1,-nbitq), 
to_sfixed(1946.0/65536.0,1,-nbitq), 
to_sfixed(6849.0/65536.0,1,-nbitq), 
to_sfixed(6958.0/65536.0,1,-nbitq), 
to_sfixed(4882.0/65536.0,1,-nbitq), 
to_sfixed(-5586.0/65536.0,1,-nbitq), 
to_sfixed(154.0/65536.0,1,-nbitq), 
to_sfixed(-1836.0/65536.0,1,-nbitq), 
to_sfixed(2183.0/65536.0,1,-nbitq), 
to_sfixed(1592.0/65536.0,1,-nbitq), 
to_sfixed(48.0/65536.0,1,-nbitq), 
to_sfixed(2283.0/65536.0,1,-nbitq), 
to_sfixed(-413.0/65536.0,1,-nbitq), 
to_sfixed(-9537.0/65536.0,1,-nbitq), 
to_sfixed(7550.0/65536.0,1,-nbitq), 
to_sfixed(-1705.0/65536.0,1,-nbitq), 
to_sfixed(962.0/65536.0,1,-nbitq), 
to_sfixed(-3353.0/65536.0,1,-nbitq), 
to_sfixed(-5462.0/65536.0,1,-nbitq), 
to_sfixed(-3478.0/65536.0,1,-nbitq), 
to_sfixed(-13846.0/65536.0,1,-nbitq), 
to_sfixed(9125.0/65536.0,1,-nbitq), 
to_sfixed(3733.0/65536.0,1,-nbitq), 
to_sfixed(10536.0/65536.0,1,-nbitq), 
to_sfixed(2107.0/65536.0,1,-nbitq), 
to_sfixed(9821.0/65536.0,1,-nbitq), 
to_sfixed(-1898.0/65536.0,1,-nbitq), 
to_sfixed(1939.0/65536.0,1,-nbitq), 
to_sfixed(11857.0/65536.0,1,-nbitq), 
to_sfixed(-15366.0/65536.0,1,-nbitq), 
to_sfixed(-10848.0/65536.0,1,-nbitq), 
to_sfixed(1670.0/65536.0,1,-nbitq), 
to_sfixed(-2206.0/65536.0,1,-nbitq), 
to_sfixed(-645.0/65536.0,1,-nbitq), 
to_sfixed(4622.0/65536.0,1,-nbitq), 
to_sfixed(-10890.0/65536.0,1,-nbitq), 
to_sfixed(523.0/65536.0,1,-nbitq), 
to_sfixed(-17324.0/65536.0,1,-nbitq), 
to_sfixed(-3517.0/65536.0,1,-nbitq), 
to_sfixed(4265.0/65536.0,1,-nbitq), 
to_sfixed(-632.0/65536.0,1,-nbitq), 
to_sfixed(-552.0/65536.0,1,-nbitq), 
to_sfixed(-1075.0/65536.0,1,-nbitq), 
to_sfixed(-5167.0/65536.0,1,-nbitq), 
to_sfixed(2065.0/65536.0,1,-nbitq), 
to_sfixed(-1992.0/65536.0,1,-nbitq), 
to_sfixed(-5133.0/65536.0,1,-nbitq), 
to_sfixed(4558.0/65536.0,1,-nbitq), 
to_sfixed(1588.0/65536.0,1,-nbitq), 
to_sfixed(-2522.0/65536.0,1,-nbitq), 
to_sfixed(-2343.0/65536.0,1,-nbitq), 
to_sfixed(-1061.0/65536.0,1,-nbitq), 
to_sfixed(1367.0/65536.0,1,-nbitq), 
to_sfixed(-2737.0/65536.0,1,-nbitq), 
to_sfixed(936.0/65536.0,1,-nbitq), 
to_sfixed(-1932.0/65536.0,1,-nbitq), 
to_sfixed(-5344.0/65536.0,1,-nbitq), 
to_sfixed(7211.0/65536.0,1,-nbitq), 
to_sfixed(-2649.0/65536.0,1,-nbitq), 
to_sfixed(-11231.0/65536.0,1,-nbitq), 
to_sfixed(-6894.0/65536.0,1,-nbitq), 
to_sfixed(1657.0/65536.0,1,-nbitq), 
to_sfixed(736.0/65536.0,1,-nbitq), 
to_sfixed(10360.0/65536.0,1,-nbitq), 
to_sfixed(-3461.0/65536.0,1,-nbitq), 
to_sfixed(-2217.0/65536.0,1,-nbitq), 
to_sfixed(-2412.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(-4101.0/65536.0,1,-nbitq), 
to_sfixed(-20712.0/65536.0,1,-nbitq), 
to_sfixed(2094.0/65536.0,1,-nbitq), 
to_sfixed(-10092.0/65536.0,1,-nbitq)  ), 
( to_sfixed(851.0/65536.0,1,-nbitq), 
to_sfixed(1239.0/65536.0,1,-nbitq), 
to_sfixed(-16887.0/65536.0,1,-nbitq), 
to_sfixed(2099.0/65536.0,1,-nbitq), 
to_sfixed(17072.0/65536.0,1,-nbitq), 
to_sfixed(-4738.0/65536.0,1,-nbitq), 
to_sfixed(3318.0/65536.0,1,-nbitq), 
to_sfixed(-213.0/65536.0,1,-nbitq), 
to_sfixed(-3185.0/65536.0,1,-nbitq), 
to_sfixed(-2799.0/65536.0,1,-nbitq), 
to_sfixed(10682.0/65536.0,1,-nbitq), 
to_sfixed(1635.0/65536.0,1,-nbitq), 
to_sfixed(4291.0/65536.0,1,-nbitq), 
to_sfixed(-2713.0/65536.0,1,-nbitq), 
to_sfixed(-318.0/65536.0,1,-nbitq), 
to_sfixed(-1540.0/65536.0,1,-nbitq), 
to_sfixed(-150.0/65536.0,1,-nbitq), 
to_sfixed(8663.0/65536.0,1,-nbitq), 
to_sfixed(564.0/65536.0,1,-nbitq), 
to_sfixed(-1228.0/65536.0,1,-nbitq), 
to_sfixed(6785.0/65536.0,1,-nbitq), 
to_sfixed(338.0/65536.0,1,-nbitq), 
to_sfixed(15287.0/65536.0,1,-nbitq), 
to_sfixed(-4848.0/65536.0,1,-nbitq), 
to_sfixed(4491.0/65536.0,1,-nbitq), 
to_sfixed(-6527.0/65536.0,1,-nbitq), 
to_sfixed(-5036.0/65536.0,1,-nbitq), 
to_sfixed(-3439.0/65536.0,1,-nbitq), 
to_sfixed(-2949.0/65536.0,1,-nbitq), 
to_sfixed(6210.0/65536.0,1,-nbitq), 
to_sfixed(2209.0/65536.0,1,-nbitq), 
to_sfixed(5635.0/65536.0,1,-nbitq), 
to_sfixed(5755.0/65536.0,1,-nbitq), 
to_sfixed(5601.0/65536.0,1,-nbitq), 
to_sfixed(986.0/65536.0,1,-nbitq), 
to_sfixed(-3164.0/65536.0,1,-nbitq), 
to_sfixed(15928.0/65536.0,1,-nbitq), 
to_sfixed(-10608.0/65536.0,1,-nbitq), 
to_sfixed(-12307.0/65536.0,1,-nbitq), 
to_sfixed(2384.0/65536.0,1,-nbitq), 
to_sfixed(-9128.0/65536.0,1,-nbitq), 
to_sfixed(-1698.0/65536.0,1,-nbitq), 
to_sfixed(-3487.0/65536.0,1,-nbitq), 
to_sfixed(-12040.0/65536.0,1,-nbitq), 
to_sfixed(-2720.0/65536.0,1,-nbitq), 
to_sfixed(1094.0/65536.0,1,-nbitq), 
to_sfixed(-3716.0/65536.0,1,-nbitq), 
to_sfixed(-3149.0/65536.0,1,-nbitq), 
to_sfixed(-2488.0/65536.0,1,-nbitq), 
to_sfixed(-316.0/65536.0,1,-nbitq), 
to_sfixed(-2052.0/65536.0,1,-nbitq), 
to_sfixed(-7472.0/65536.0,1,-nbitq), 
to_sfixed(242.0/65536.0,1,-nbitq), 
to_sfixed(-7141.0/65536.0,1,-nbitq), 
to_sfixed(-7267.0/65536.0,1,-nbitq), 
to_sfixed(7774.0/65536.0,1,-nbitq), 
to_sfixed(-2925.0/65536.0,1,-nbitq), 
to_sfixed(3816.0/65536.0,1,-nbitq), 
to_sfixed(-2978.0/65536.0,1,-nbitq), 
to_sfixed(-3463.0/65536.0,1,-nbitq), 
to_sfixed(3818.0/65536.0,1,-nbitq), 
to_sfixed(1324.0/65536.0,1,-nbitq), 
to_sfixed(1692.0/65536.0,1,-nbitq), 
to_sfixed(-2809.0/65536.0,1,-nbitq), 
to_sfixed(-12926.0/65536.0,1,-nbitq), 
to_sfixed(2991.0/65536.0,1,-nbitq), 
to_sfixed(114.0/65536.0,1,-nbitq), 
to_sfixed(-6896.0/65536.0,1,-nbitq), 
to_sfixed(-6274.0/65536.0,1,-nbitq), 
to_sfixed(690.0/65536.0,1,-nbitq), 
to_sfixed(-979.0/65536.0,1,-nbitq), 
to_sfixed(8390.0/65536.0,1,-nbitq), 
to_sfixed(-6133.0/65536.0,1,-nbitq), 
to_sfixed(2900.0/65536.0,1,-nbitq), 
to_sfixed(-1890.0/65536.0,1,-nbitq), 
to_sfixed(-8193.0/65536.0,1,-nbitq), 
to_sfixed(-4815.0/65536.0,1,-nbitq), 
to_sfixed(-7731.0/65536.0,1,-nbitq), 
to_sfixed(266.0/65536.0,1,-nbitq), 
to_sfixed(-6502.0/65536.0,1,-nbitq)  ), 
( to_sfixed(7219.0/65536.0,1,-nbitq), 
to_sfixed(-4953.0/65536.0,1,-nbitq), 
to_sfixed(-16974.0/65536.0,1,-nbitq), 
to_sfixed(2926.0/65536.0,1,-nbitq), 
to_sfixed(14220.0/65536.0,1,-nbitq), 
to_sfixed(-6225.0/65536.0,1,-nbitq), 
to_sfixed(5362.0/65536.0,1,-nbitq), 
to_sfixed(4255.0/65536.0,1,-nbitq), 
to_sfixed(-1881.0/65536.0,1,-nbitq), 
to_sfixed(1041.0/65536.0,1,-nbitq), 
to_sfixed(9053.0/65536.0,1,-nbitq), 
to_sfixed(5057.0/65536.0,1,-nbitq), 
to_sfixed(377.0/65536.0,1,-nbitq), 
to_sfixed(-627.0/65536.0,1,-nbitq), 
to_sfixed(-4242.0/65536.0,1,-nbitq), 
to_sfixed(-238.0/65536.0,1,-nbitq), 
to_sfixed(-1315.0/65536.0,1,-nbitq), 
to_sfixed(3102.0/65536.0,1,-nbitq), 
to_sfixed(-1087.0/65536.0,1,-nbitq), 
to_sfixed(-1053.0/65536.0,1,-nbitq), 
to_sfixed(7053.0/65536.0,1,-nbitq), 
to_sfixed(1722.0/65536.0,1,-nbitq), 
to_sfixed(15693.0/65536.0,1,-nbitq), 
to_sfixed(-149.0/65536.0,1,-nbitq), 
to_sfixed(357.0/65536.0,1,-nbitq), 
to_sfixed(-3090.0/65536.0,1,-nbitq), 
to_sfixed(-4735.0/65536.0,1,-nbitq), 
to_sfixed(-1362.0/65536.0,1,-nbitq), 
to_sfixed(8650.0/65536.0,1,-nbitq), 
to_sfixed(975.0/65536.0,1,-nbitq), 
to_sfixed(4093.0/65536.0,1,-nbitq), 
to_sfixed(-386.0/65536.0,1,-nbitq), 
to_sfixed(4880.0/65536.0,1,-nbitq), 
to_sfixed(3336.0/65536.0,1,-nbitq), 
to_sfixed(-2274.0/65536.0,1,-nbitq), 
to_sfixed(-407.0/65536.0,1,-nbitq), 
to_sfixed(13329.0/65536.0,1,-nbitq), 
to_sfixed(-3938.0/65536.0,1,-nbitq), 
to_sfixed(-13831.0/65536.0,1,-nbitq), 
to_sfixed(-2643.0/65536.0,1,-nbitq), 
to_sfixed(-6308.0/65536.0,1,-nbitq), 
to_sfixed(-2094.0/65536.0,1,-nbitq), 
to_sfixed(-10359.0/65536.0,1,-nbitq), 
to_sfixed(-11481.0/65536.0,1,-nbitq), 
to_sfixed(1528.0/65536.0,1,-nbitq), 
to_sfixed(11809.0/65536.0,1,-nbitq), 
to_sfixed(-116.0/65536.0,1,-nbitq), 
to_sfixed(4390.0/65536.0,1,-nbitq), 
to_sfixed(1669.0/65536.0,1,-nbitq), 
to_sfixed(-5019.0/65536.0,1,-nbitq), 
to_sfixed(-2580.0/65536.0,1,-nbitq), 
to_sfixed(-8823.0/65536.0,1,-nbitq), 
to_sfixed(-1917.0/65536.0,1,-nbitq), 
to_sfixed(-689.0/65536.0,1,-nbitq), 
to_sfixed(-6540.0/65536.0,1,-nbitq), 
to_sfixed(-1038.0/65536.0,1,-nbitq), 
to_sfixed(-2163.0/65536.0,1,-nbitq), 
to_sfixed(96.0/65536.0,1,-nbitq), 
to_sfixed(-2617.0/65536.0,1,-nbitq), 
to_sfixed(-4802.0/65536.0,1,-nbitq), 
to_sfixed(8348.0/65536.0,1,-nbitq), 
to_sfixed(1414.0/65536.0,1,-nbitq), 
to_sfixed(-1393.0/65536.0,1,-nbitq), 
to_sfixed(-532.0/65536.0,1,-nbitq), 
to_sfixed(-12168.0/65536.0,1,-nbitq), 
to_sfixed(-11580.0/65536.0,1,-nbitq), 
to_sfixed(-446.0/65536.0,1,-nbitq), 
to_sfixed(-4509.0/65536.0,1,-nbitq), 
to_sfixed(-11158.0/65536.0,1,-nbitq), 
to_sfixed(2276.0/65536.0,1,-nbitq), 
to_sfixed(1895.0/65536.0,1,-nbitq), 
to_sfixed(-4163.0/65536.0,1,-nbitq), 
to_sfixed(-3243.0/65536.0,1,-nbitq), 
to_sfixed(2117.0/65536.0,1,-nbitq), 
to_sfixed(-2498.0/65536.0,1,-nbitq), 
to_sfixed(-7341.0/65536.0,1,-nbitq), 
to_sfixed(-1913.0/65536.0,1,-nbitq), 
to_sfixed(-1091.0/65536.0,1,-nbitq), 
to_sfixed(56.0/65536.0,1,-nbitq), 
to_sfixed(-2626.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4506.0/65536.0,1,-nbitq), 
to_sfixed(-3115.0/65536.0,1,-nbitq), 
to_sfixed(-13167.0/65536.0,1,-nbitq), 
to_sfixed(-2031.0/65536.0,1,-nbitq), 
to_sfixed(-9335.0/65536.0,1,-nbitq), 
to_sfixed(-15041.0/65536.0,1,-nbitq), 
to_sfixed(4156.0/65536.0,1,-nbitq), 
to_sfixed(-29.0/65536.0,1,-nbitq), 
to_sfixed(-2866.0/65536.0,1,-nbitq), 
to_sfixed(1126.0/65536.0,1,-nbitq), 
to_sfixed(3384.0/65536.0,1,-nbitq), 
to_sfixed(4498.0/65536.0,1,-nbitq), 
to_sfixed(-1381.0/65536.0,1,-nbitq), 
to_sfixed(1440.0/65536.0,1,-nbitq), 
to_sfixed(-10418.0/65536.0,1,-nbitq), 
to_sfixed(-1320.0/65536.0,1,-nbitq), 
to_sfixed(-2750.0/65536.0,1,-nbitq), 
to_sfixed(-2873.0/65536.0,1,-nbitq), 
to_sfixed(-2051.0/65536.0,1,-nbitq), 
to_sfixed(1763.0/65536.0,1,-nbitq), 
to_sfixed(5955.0/65536.0,1,-nbitq), 
to_sfixed(4636.0/65536.0,1,-nbitq), 
to_sfixed(19359.0/65536.0,1,-nbitq), 
to_sfixed(3604.0/65536.0,1,-nbitq), 
to_sfixed(104.0/65536.0,1,-nbitq), 
to_sfixed(-718.0/65536.0,1,-nbitq), 
to_sfixed(-7692.0/65536.0,1,-nbitq), 
to_sfixed(784.0/65536.0,1,-nbitq), 
to_sfixed(3118.0/65536.0,1,-nbitq), 
to_sfixed(1627.0/65536.0,1,-nbitq), 
to_sfixed(2621.0/65536.0,1,-nbitq), 
to_sfixed(7373.0/65536.0,1,-nbitq), 
to_sfixed(7651.0/65536.0,1,-nbitq), 
to_sfixed(-2253.0/65536.0,1,-nbitq), 
to_sfixed(-240.0/65536.0,1,-nbitq), 
to_sfixed(-179.0/65536.0,1,-nbitq), 
to_sfixed(650.0/65536.0,1,-nbitq), 
to_sfixed(-2891.0/65536.0,1,-nbitq), 
to_sfixed(-3221.0/65536.0,1,-nbitq), 
to_sfixed(-5617.0/65536.0,1,-nbitq), 
to_sfixed(-3789.0/65536.0,1,-nbitq), 
to_sfixed(674.0/65536.0,1,-nbitq), 
to_sfixed(-11510.0/65536.0,1,-nbitq), 
to_sfixed(-8384.0/65536.0,1,-nbitq), 
to_sfixed(1501.0/65536.0,1,-nbitq), 
to_sfixed(7919.0/65536.0,1,-nbitq), 
to_sfixed(-3078.0/65536.0,1,-nbitq), 
to_sfixed(5310.0/65536.0,1,-nbitq), 
to_sfixed(-1008.0/65536.0,1,-nbitq), 
to_sfixed(-140.0/65536.0,1,-nbitq), 
to_sfixed(-1223.0/65536.0,1,-nbitq), 
to_sfixed(-1805.0/65536.0,1,-nbitq), 
to_sfixed(1250.0/65536.0,1,-nbitq), 
to_sfixed(-5519.0/65536.0,1,-nbitq), 
to_sfixed(-3814.0/65536.0,1,-nbitq), 
to_sfixed(-267.0/65536.0,1,-nbitq), 
to_sfixed(-1474.0/65536.0,1,-nbitq), 
to_sfixed(-1976.0/65536.0,1,-nbitq), 
to_sfixed(1143.0/65536.0,1,-nbitq), 
to_sfixed(-5610.0/65536.0,1,-nbitq), 
to_sfixed(2753.0/65536.0,1,-nbitq), 
to_sfixed(1710.0/65536.0,1,-nbitq), 
to_sfixed(1717.0/65536.0,1,-nbitq), 
to_sfixed(-1690.0/65536.0,1,-nbitq), 
to_sfixed(-1466.0/65536.0,1,-nbitq), 
to_sfixed(-8276.0/65536.0,1,-nbitq), 
to_sfixed(-4100.0/65536.0,1,-nbitq), 
to_sfixed(-1643.0/65536.0,1,-nbitq), 
to_sfixed(-7475.0/65536.0,1,-nbitq), 
to_sfixed(-11019.0/65536.0,1,-nbitq), 
to_sfixed(1192.0/65536.0,1,-nbitq), 
to_sfixed(384.0/65536.0,1,-nbitq), 
to_sfixed(-12706.0/65536.0,1,-nbitq), 
to_sfixed(2158.0/65536.0,1,-nbitq), 
to_sfixed(-933.0/65536.0,1,-nbitq), 
to_sfixed(-3953.0/65536.0,1,-nbitq), 
to_sfixed(4203.0/65536.0,1,-nbitq), 
to_sfixed(3595.0/65536.0,1,-nbitq), 
to_sfixed(-7.0/65536.0,1,-nbitq), 
to_sfixed(3831.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2835.0/65536.0,1,-nbitq), 
to_sfixed(2437.0/65536.0,1,-nbitq), 
to_sfixed(-2618.0/65536.0,1,-nbitq), 
to_sfixed(-7391.0/65536.0,1,-nbitq), 
to_sfixed(-7817.0/65536.0,1,-nbitq), 
to_sfixed(-5986.0/65536.0,1,-nbitq), 
to_sfixed(517.0/65536.0,1,-nbitq), 
to_sfixed(-6906.0/65536.0,1,-nbitq), 
to_sfixed(1828.0/65536.0,1,-nbitq), 
to_sfixed(1172.0/65536.0,1,-nbitq), 
to_sfixed(2609.0/65536.0,1,-nbitq), 
to_sfixed(-3726.0/65536.0,1,-nbitq), 
to_sfixed(-1332.0/65536.0,1,-nbitq), 
to_sfixed(-8939.0/65536.0,1,-nbitq), 
to_sfixed(-3187.0/65536.0,1,-nbitq), 
to_sfixed(1337.0/65536.0,1,-nbitq), 
to_sfixed(-2967.0/65536.0,1,-nbitq), 
to_sfixed(-851.0/65536.0,1,-nbitq), 
to_sfixed(3051.0/65536.0,1,-nbitq), 
to_sfixed(1844.0/65536.0,1,-nbitq), 
to_sfixed(14698.0/65536.0,1,-nbitq), 
to_sfixed(-1097.0/65536.0,1,-nbitq), 
to_sfixed(-4951.0/65536.0,1,-nbitq), 
to_sfixed(437.0/65536.0,1,-nbitq), 
to_sfixed(-5810.0/65536.0,1,-nbitq), 
to_sfixed(-830.0/65536.0,1,-nbitq), 
to_sfixed(766.0/65536.0,1,-nbitq), 
to_sfixed(1688.0/65536.0,1,-nbitq), 
to_sfixed(4014.0/65536.0,1,-nbitq), 
to_sfixed(-2402.0/65536.0,1,-nbitq), 
to_sfixed(-118.0/65536.0,1,-nbitq), 
to_sfixed(7386.0/65536.0,1,-nbitq), 
to_sfixed(-5007.0/65536.0,1,-nbitq), 
to_sfixed(930.0/65536.0,1,-nbitq), 
to_sfixed(245.0/65536.0,1,-nbitq), 
to_sfixed(530.0/65536.0,1,-nbitq), 
to_sfixed(1164.0/65536.0,1,-nbitq), 
to_sfixed(-822.0/65536.0,1,-nbitq), 
to_sfixed(14282.0/65536.0,1,-nbitq), 
to_sfixed(-3017.0/65536.0,1,-nbitq), 
to_sfixed(-4117.0/65536.0,1,-nbitq), 
to_sfixed(-2604.0/65536.0,1,-nbitq), 
to_sfixed(-12489.0/65536.0,1,-nbitq), 
to_sfixed(-583.0/65536.0,1,-nbitq), 
to_sfixed(-1325.0/65536.0,1,-nbitq), 
to_sfixed(7640.0/65536.0,1,-nbitq), 
to_sfixed(-1668.0/65536.0,1,-nbitq), 
to_sfixed(6538.0/65536.0,1,-nbitq), 
to_sfixed(1601.0/65536.0,1,-nbitq), 
to_sfixed(-941.0/65536.0,1,-nbitq), 
to_sfixed(-1149.0/65536.0,1,-nbitq), 
to_sfixed(4664.0/65536.0,1,-nbitq), 
to_sfixed(595.0/65536.0,1,-nbitq), 
to_sfixed(1760.0/65536.0,1,-nbitq), 
to_sfixed(-3654.0/65536.0,1,-nbitq), 
to_sfixed(-1836.0/65536.0,1,-nbitq), 
to_sfixed(-1802.0/65536.0,1,-nbitq), 
to_sfixed(30.0/65536.0,1,-nbitq), 
to_sfixed(-3053.0/65536.0,1,-nbitq), 
to_sfixed(633.0/65536.0,1,-nbitq), 
to_sfixed(-6166.0/65536.0,1,-nbitq), 
to_sfixed(554.0/65536.0,1,-nbitq), 
to_sfixed(1255.0/65536.0,1,-nbitq), 
to_sfixed(-1510.0/65536.0,1,-nbitq), 
to_sfixed(-1499.0/65536.0,1,-nbitq), 
to_sfixed(-7732.0/65536.0,1,-nbitq), 
to_sfixed(-12644.0/65536.0,1,-nbitq), 
to_sfixed(1235.0/65536.0,1,-nbitq), 
to_sfixed(-6376.0/65536.0,1,-nbitq), 
to_sfixed(-6163.0/65536.0,1,-nbitq), 
to_sfixed(-2783.0/65536.0,1,-nbitq), 
to_sfixed(3425.0/65536.0,1,-nbitq), 
to_sfixed(-6266.0/65536.0,1,-nbitq), 
to_sfixed(1607.0/65536.0,1,-nbitq), 
to_sfixed(-854.0/65536.0,1,-nbitq), 
to_sfixed(-5952.0/65536.0,1,-nbitq), 
to_sfixed(2854.0/65536.0,1,-nbitq), 
to_sfixed(6822.0/65536.0,1,-nbitq), 
to_sfixed(1972.0/65536.0,1,-nbitq), 
to_sfixed(8422.0/65536.0,1,-nbitq)  ), 
( to_sfixed(792.0/65536.0,1,-nbitq), 
to_sfixed(7858.0/65536.0,1,-nbitq), 
to_sfixed(11614.0/65536.0,1,-nbitq), 
to_sfixed(-9507.0/65536.0,1,-nbitq), 
to_sfixed(-2227.0/65536.0,1,-nbitq), 
to_sfixed(5951.0/65536.0,1,-nbitq), 
to_sfixed(4215.0/65536.0,1,-nbitq), 
to_sfixed(-6385.0/65536.0,1,-nbitq), 
to_sfixed(11524.0/65536.0,1,-nbitq), 
to_sfixed(-2257.0/65536.0,1,-nbitq), 
to_sfixed(4846.0/65536.0,1,-nbitq), 
to_sfixed(-8558.0/65536.0,1,-nbitq), 
to_sfixed(1991.0/65536.0,1,-nbitq), 
to_sfixed(-3142.0/65536.0,1,-nbitq), 
to_sfixed(1765.0/65536.0,1,-nbitq), 
to_sfixed(-613.0/65536.0,1,-nbitq), 
to_sfixed(2048.0/65536.0,1,-nbitq), 
to_sfixed(-501.0/65536.0,1,-nbitq), 
to_sfixed(4627.0/65536.0,1,-nbitq), 
to_sfixed(2975.0/65536.0,1,-nbitq), 
to_sfixed(13735.0/65536.0,1,-nbitq), 
to_sfixed(1424.0/65536.0,1,-nbitq), 
to_sfixed(-13319.0/65536.0,1,-nbitq), 
to_sfixed(3057.0/65536.0,1,-nbitq), 
to_sfixed(-3710.0/65536.0,1,-nbitq), 
to_sfixed(-2802.0/65536.0,1,-nbitq), 
to_sfixed(-1937.0/65536.0,1,-nbitq), 
to_sfixed(2818.0/65536.0,1,-nbitq), 
to_sfixed(-363.0/65536.0,1,-nbitq), 
to_sfixed(-2244.0/65536.0,1,-nbitq), 
to_sfixed(156.0/65536.0,1,-nbitq), 
to_sfixed(-4544.0/65536.0,1,-nbitq), 
to_sfixed(-7020.0/65536.0,1,-nbitq), 
to_sfixed(-2828.0/65536.0,1,-nbitq), 
to_sfixed(-775.0/65536.0,1,-nbitq), 
to_sfixed(3245.0/65536.0,1,-nbitq), 
to_sfixed(4264.0/65536.0,1,-nbitq), 
to_sfixed(3380.0/65536.0,1,-nbitq), 
to_sfixed(13804.0/65536.0,1,-nbitq), 
to_sfixed(455.0/65536.0,1,-nbitq), 
to_sfixed(-14189.0/65536.0,1,-nbitq), 
to_sfixed(-895.0/65536.0,1,-nbitq), 
to_sfixed(-12981.0/65536.0,1,-nbitq), 
to_sfixed(-2088.0/65536.0,1,-nbitq), 
to_sfixed(-2194.0/65536.0,1,-nbitq), 
to_sfixed(-400.0/65536.0,1,-nbitq), 
to_sfixed(-658.0/65536.0,1,-nbitq), 
to_sfixed(3402.0/65536.0,1,-nbitq), 
to_sfixed(792.0/65536.0,1,-nbitq), 
to_sfixed(2394.0/65536.0,1,-nbitq), 
to_sfixed(-1725.0/65536.0,1,-nbitq), 
to_sfixed(15212.0/65536.0,1,-nbitq), 
to_sfixed(-4165.0/65536.0,1,-nbitq), 
to_sfixed(12647.0/65536.0,1,-nbitq), 
to_sfixed(-4739.0/65536.0,1,-nbitq), 
to_sfixed(-12984.0/65536.0,1,-nbitq), 
to_sfixed(966.0/65536.0,1,-nbitq), 
to_sfixed(4386.0/65536.0,1,-nbitq), 
to_sfixed(-2820.0/65536.0,1,-nbitq), 
to_sfixed(3141.0/65536.0,1,-nbitq), 
to_sfixed(-3036.0/65536.0,1,-nbitq), 
to_sfixed(1759.0/65536.0,1,-nbitq), 
to_sfixed(2700.0/65536.0,1,-nbitq), 
to_sfixed(1259.0/65536.0,1,-nbitq), 
to_sfixed(1165.0/65536.0,1,-nbitq), 
to_sfixed(-5349.0/65536.0,1,-nbitq), 
to_sfixed(-8953.0/65536.0,1,-nbitq), 
to_sfixed(4251.0/65536.0,1,-nbitq), 
to_sfixed(-4651.0/65536.0,1,-nbitq), 
to_sfixed(-584.0/65536.0,1,-nbitq), 
to_sfixed(-1910.0/65536.0,1,-nbitq), 
to_sfixed(5692.0/65536.0,1,-nbitq), 
to_sfixed(2574.0/65536.0,1,-nbitq), 
to_sfixed(-2286.0/65536.0,1,-nbitq), 
to_sfixed(587.0/65536.0,1,-nbitq), 
to_sfixed(-7377.0/65536.0,1,-nbitq), 
to_sfixed(-3179.0/65536.0,1,-nbitq), 
to_sfixed(11458.0/65536.0,1,-nbitq), 
to_sfixed(-1570.0/65536.0,1,-nbitq), 
to_sfixed(8131.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2895.0/65536.0,1,-nbitq), 
to_sfixed(1646.0/65536.0,1,-nbitq), 
to_sfixed(6824.0/65536.0,1,-nbitq), 
to_sfixed(-5426.0/65536.0,1,-nbitq), 
to_sfixed(-4440.0/65536.0,1,-nbitq), 
to_sfixed(17011.0/65536.0,1,-nbitq), 
to_sfixed(253.0/65536.0,1,-nbitq), 
to_sfixed(-2063.0/65536.0,1,-nbitq), 
to_sfixed(16627.0/65536.0,1,-nbitq), 
to_sfixed(-212.0/65536.0,1,-nbitq), 
to_sfixed(7383.0/65536.0,1,-nbitq), 
to_sfixed(-6560.0/65536.0,1,-nbitq), 
to_sfixed(-2747.0/65536.0,1,-nbitq), 
to_sfixed(-1996.0/65536.0,1,-nbitq), 
to_sfixed(1107.0/65536.0,1,-nbitq), 
to_sfixed(-1218.0/65536.0,1,-nbitq), 
to_sfixed(-2080.0/65536.0,1,-nbitq), 
to_sfixed(347.0/65536.0,1,-nbitq), 
to_sfixed(-1987.0/65536.0,1,-nbitq), 
to_sfixed(348.0/65536.0,1,-nbitq), 
to_sfixed(9981.0/65536.0,1,-nbitq), 
to_sfixed(-7068.0/65536.0,1,-nbitq), 
to_sfixed(3532.0/65536.0,1,-nbitq), 
to_sfixed(5705.0/65536.0,1,-nbitq), 
to_sfixed(-314.0/65536.0,1,-nbitq), 
to_sfixed(-458.0/65536.0,1,-nbitq), 
to_sfixed(310.0/65536.0,1,-nbitq), 
to_sfixed(-411.0/65536.0,1,-nbitq), 
to_sfixed(100.0/65536.0,1,-nbitq), 
to_sfixed(2002.0/65536.0,1,-nbitq), 
to_sfixed(1985.0/65536.0,1,-nbitq), 
to_sfixed(-4265.0/65536.0,1,-nbitq), 
to_sfixed(-10820.0/65536.0,1,-nbitq), 
to_sfixed(1880.0/65536.0,1,-nbitq), 
to_sfixed(595.0/65536.0,1,-nbitq), 
to_sfixed(-96.0/65536.0,1,-nbitq), 
to_sfixed(6565.0/65536.0,1,-nbitq), 
to_sfixed(1671.0/65536.0,1,-nbitq), 
to_sfixed(4274.0/65536.0,1,-nbitq), 
to_sfixed(-2303.0/65536.0,1,-nbitq), 
to_sfixed(-12909.0/65536.0,1,-nbitq), 
to_sfixed(-67.0/65536.0,1,-nbitq), 
to_sfixed(-10905.0/65536.0,1,-nbitq), 
to_sfixed(-5966.0/65536.0,1,-nbitq), 
to_sfixed(1245.0/65536.0,1,-nbitq), 
to_sfixed(-5972.0/65536.0,1,-nbitq), 
to_sfixed(-6294.0/65536.0,1,-nbitq), 
to_sfixed(6413.0/65536.0,1,-nbitq), 
to_sfixed(-2100.0/65536.0,1,-nbitq), 
to_sfixed(2563.0/65536.0,1,-nbitq), 
to_sfixed(2031.0/65536.0,1,-nbitq), 
to_sfixed(11455.0/65536.0,1,-nbitq), 
to_sfixed(-2777.0/65536.0,1,-nbitq), 
to_sfixed(5672.0/65536.0,1,-nbitq), 
to_sfixed(2093.0/65536.0,1,-nbitq), 
to_sfixed(-5486.0/65536.0,1,-nbitq), 
to_sfixed(739.0/65536.0,1,-nbitq), 
to_sfixed(-1541.0/65536.0,1,-nbitq), 
to_sfixed(-2460.0/65536.0,1,-nbitq), 
to_sfixed(1870.0/65536.0,1,-nbitq), 
to_sfixed(-1965.0/65536.0,1,-nbitq), 
to_sfixed(733.0/65536.0,1,-nbitq), 
to_sfixed(-966.0/65536.0,1,-nbitq), 
to_sfixed(-2905.0/65536.0,1,-nbitq), 
to_sfixed(4230.0/65536.0,1,-nbitq), 
to_sfixed(-5689.0/65536.0,1,-nbitq), 
to_sfixed(-7553.0/65536.0,1,-nbitq), 
to_sfixed(7440.0/65536.0,1,-nbitq), 
to_sfixed(-2929.0/65536.0,1,-nbitq), 
to_sfixed(-2806.0/65536.0,1,-nbitq), 
to_sfixed(-4746.0/65536.0,1,-nbitq), 
to_sfixed(6735.0/65536.0,1,-nbitq), 
to_sfixed(12369.0/65536.0,1,-nbitq), 
to_sfixed(-2527.0/65536.0,1,-nbitq), 
to_sfixed(1950.0/65536.0,1,-nbitq), 
to_sfixed(2013.0/65536.0,1,-nbitq), 
to_sfixed(2995.0/65536.0,1,-nbitq), 
to_sfixed(11304.0/65536.0,1,-nbitq), 
to_sfixed(1621.0/65536.0,1,-nbitq), 
to_sfixed(6018.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1170.0/65536.0,1,-nbitq), 
to_sfixed(2094.0/65536.0,1,-nbitq), 
to_sfixed(4255.0/65536.0,1,-nbitq), 
to_sfixed(1684.0/65536.0,1,-nbitq), 
to_sfixed(-4414.0/65536.0,1,-nbitq), 
to_sfixed(10812.0/65536.0,1,-nbitq), 
to_sfixed(522.0/65536.0,1,-nbitq), 
to_sfixed(-1581.0/65536.0,1,-nbitq), 
to_sfixed(11177.0/65536.0,1,-nbitq), 
to_sfixed(-530.0/65536.0,1,-nbitq), 
to_sfixed(1183.0/65536.0,1,-nbitq), 
to_sfixed(820.0/65536.0,1,-nbitq), 
to_sfixed(-883.0/65536.0,1,-nbitq), 
to_sfixed(-1962.0/65536.0,1,-nbitq), 
to_sfixed(1347.0/65536.0,1,-nbitq), 
to_sfixed(255.0/65536.0,1,-nbitq), 
to_sfixed(-900.0/65536.0,1,-nbitq), 
to_sfixed(-2363.0/65536.0,1,-nbitq), 
to_sfixed(-4849.0/65536.0,1,-nbitq), 
to_sfixed(-161.0/65536.0,1,-nbitq), 
to_sfixed(11853.0/65536.0,1,-nbitq), 
to_sfixed(-12775.0/65536.0,1,-nbitq), 
to_sfixed(10448.0/65536.0,1,-nbitq), 
to_sfixed(5819.0/65536.0,1,-nbitq), 
to_sfixed(-1954.0/65536.0,1,-nbitq), 
to_sfixed(5507.0/65536.0,1,-nbitq), 
to_sfixed(737.0/65536.0,1,-nbitq), 
to_sfixed(2771.0/65536.0,1,-nbitq), 
to_sfixed(-3906.0/65536.0,1,-nbitq), 
to_sfixed(114.0/65536.0,1,-nbitq), 
to_sfixed(-1052.0/65536.0,1,-nbitq), 
to_sfixed(-2064.0/65536.0,1,-nbitq), 
to_sfixed(-6923.0/65536.0,1,-nbitq), 
to_sfixed(5341.0/65536.0,1,-nbitq), 
to_sfixed(1193.0/65536.0,1,-nbitq), 
to_sfixed(-3032.0/65536.0,1,-nbitq), 
to_sfixed(4403.0/65536.0,1,-nbitq), 
to_sfixed(-2401.0/65536.0,1,-nbitq), 
to_sfixed(2277.0/65536.0,1,-nbitq), 
to_sfixed(-2192.0/65536.0,1,-nbitq), 
to_sfixed(-6524.0/65536.0,1,-nbitq), 
to_sfixed(2681.0/65536.0,1,-nbitq), 
to_sfixed(4121.0/65536.0,1,-nbitq), 
to_sfixed(-7481.0/65536.0,1,-nbitq), 
to_sfixed(912.0/65536.0,1,-nbitq), 
to_sfixed(-6503.0/65536.0,1,-nbitq), 
to_sfixed(-6222.0/65536.0,1,-nbitq), 
to_sfixed(3153.0/65536.0,1,-nbitq), 
to_sfixed(-3002.0/65536.0,1,-nbitq), 
to_sfixed(2531.0/65536.0,1,-nbitq), 
to_sfixed(21.0/65536.0,1,-nbitq), 
to_sfixed(912.0/65536.0,1,-nbitq), 
to_sfixed(-875.0/65536.0,1,-nbitq), 
to_sfixed(9726.0/65536.0,1,-nbitq), 
to_sfixed(90.0/65536.0,1,-nbitq), 
to_sfixed(-259.0/65536.0,1,-nbitq), 
to_sfixed(1654.0/65536.0,1,-nbitq), 
to_sfixed(-3708.0/65536.0,1,-nbitq), 
to_sfixed(-1426.0/65536.0,1,-nbitq), 
to_sfixed(-3409.0/65536.0,1,-nbitq), 
to_sfixed(6184.0/65536.0,1,-nbitq), 
to_sfixed(1388.0/65536.0,1,-nbitq), 
to_sfixed(360.0/65536.0,1,-nbitq), 
to_sfixed(2056.0/65536.0,1,-nbitq), 
to_sfixed(43.0/65536.0,1,-nbitq), 
to_sfixed(-139.0/65536.0,1,-nbitq), 
to_sfixed(-3706.0/65536.0,1,-nbitq), 
to_sfixed(1490.0/65536.0,1,-nbitq), 
to_sfixed(-2430.0/65536.0,1,-nbitq), 
to_sfixed(-1633.0/65536.0,1,-nbitq), 
to_sfixed(-5783.0/65536.0,1,-nbitq), 
to_sfixed(7583.0/65536.0,1,-nbitq), 
to_sfixed(10384.0/65536.0,1,-nbitq), 
to_sfixed(-1132.0/65536.0,1,-nbitq), 
to_sfixed(137.0/65536.0,1,-nbitq), 
to_sfixed(4910.0/65536.0,1,-nbitq), 
to_sfixed(3561.0/65536.0,1,-nbitq), 
to_sfixed(114.0/65536.0,1,-nbitq), 
to_sfixed(-184.0/65536.0,1,-nbitq), 
to_sfixed(2786.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3338.0/65536.0,1,-nbitq), 
to_sfixed(2210.0/65536.0,1,-nbitq), 
to_sfixed(-726.0/65536.0,1,-nbitq), 
to_sfixed(-4712.0/65536.0,1,-nbitq), 
to_sfixed(14327.0/65536.0,1,-nbitq), 
to_sfixed(12439.0/65536.0,1,-nbitq), 
to_sfixed(1444.0/65536.0,1,-nbitq), 
to_sfixed(598.0/65536.0,1,-nbitq), 
to_sfixed(6277.0/65536.0,1,-nbitq), 
to_sfixed(-219.0/65536.0,1,-nbitq), 
to_sfixed(2068.0/65536.0,1,-nbitq), 
to_sfixed(1248.0/65536.0,1,-nbitq), 
to_sfixed(75.0/65536.0,1,-nbitq), 
to_sfixed(3103.0/65536.0,1,-nbitq), 
to_sfixed(1084.0/65536.0,1,-nbitq), 
to_sfixed(629.0/65536.0,1,-nbitq), 
to_sfixed(-2398.0/65536.0,1,-nbitq), 
to_sfixed(-4436.0/65536.0,1,-nbitq), 
to_sfixed(-2983.0/65536.0,1,-nbitq), 
to_sfixed(1294.0/65536.0,1,-nbitq), 
to_sfixed(12665.0/65536.0,1,-nbitq), 
to_sfixed(-7078.0/65536.0,1,-nbitq), 
to_sfixed(2665.0/65536.0,1,-nbitq), 
to_sfixed(7541.0/65536.0,1,-nbitq), 
to_sfixed(3357.0/65536.0,1,-nbitq), 
to_sfixed(3582.0/65536.0,1,-nbitq), 
to_sfixed(1130.0/65536.0,1,-nbitq), 
to_sfixed(2778.0/65536.0,1,-nbitq), 
to_sfixed(-406.0/65536.0,1,-nbitq), 
to_sfixed(-4093.0/65536.0,1,-nbitq), 
to_sfixed(-5240.0/65536.0,1,-nbitq), 
to_sfixed(-2187.0/65536.0,1,-nbitq), 
to_sfixed(-856.0/65536.0,1,-nbitq), 
to_sfixed(6239.0/65536.0,1,-nbitq), 
to_sfixed(1372.0/65536.0,1,-nbitq), 
to_sfixed(737.0/65536.0,1,-nbitq), 
to_sfixed(9154.0/65536.0,1,-nbitq), 
to_sfixed(1664.0/65536.0,1,-nbitq), 
to_sfixed(2927.0/65536.0,1,-nbitq), 
to_sfixed(-330.0/65536.0,1,-nbitq), 
to_sfixed(-4576.0/65536.0,1,-nbitq), 
to_sfixed(-3067.0/65536.0,1,-nbitq), 
to_sfixed(15022.0/65536.0,1,-nbitq), 
to_sfixed(-2313.0/65536.0,1,-nbitq), 
to_sfixed(-1276.0/65536.0,1,-nbitq), 
to_sfixed(-8677.0/65536.0,1,-nbitq), 
to_sfixed(-3618.0/65536.0,1,-nbitq), 
to_sfixed(986.0/65536.0,1,-nbitq), 
to_sfixed(-2070.0/65536.0,1,-nbitq), 
to_sfixed(-2770.0/65536.0,1,-nbitq), 
to_sfixed(-2186.0/65536.0,1,-nbitq), 
to_sfixed(-7647.0/65536.0,1,-nbitq), 
to_sfixed(-3705.0/65536.0,1,-nbitq), 
to_sfixed(-972.0/65536.0,1,-nbitq), 
to_sfixed(4879.0/65536.0,1,-nbitq), 
to_sfixed(3631.0/65536.0,1,-nbitq), 
to_sfixed(2965.0/65536.0,1,-nbitq), 
to_sfixed(-1964.0/65536.0,1,-nbitq), 
to_sfixed(-991.0/65536.0,1,-nbitq), 
to_sfixed(-9138.0/65536.0,1,-nbitq), 
to_sfixed(4459.0/65536.0,1,-nbitq), 
to_sfixed(-600.0/65536.0,1,-nbitq), 
to_sfixed(314.0/65536.0,1,-nbitq), 
to_sfixed(492.0/65536.0,1,-nbitq), 
to_sfixed(4984.0/65536.0,1,-nbitq), 
to_sfixed(-1848.0/65536.0,1,-nbitq), 
to_sfixed(-4959.0/65536.0,1,-nbitq), 
to_sfixed(4964.0/65536.0,1,-nbitq), 
to_sfixed(-10766.0/65536.0,1,-nbitq), 
to_sfixed(-4167.0/65536.0,1,-nbitq), 
to_sfixed(-1755.0/65536.0,1,-nbitq), 
to_sfixed(9987.0/65536.0,1,-nbitq), 
to_sfixed(-190.0/65536.0,1,-nbitq), 
to_sfixed(1303.0/65536.0,1,-nbitq), 
to_sfixed(-1386.0/65536.0,1,-nbitq), 
to_sfixed(4918.0/65536.0,1,-nbitq), 
to_sfixed(8043.0/65536.0,1,-nbitq), 
to_sfixed(-11196.0/65536.0,1,-nbitq), 
to_sfixed(1873.0/65536.0,1,-nbitq), 
to_sfixed(-957.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4585.0/65536.0,1,-nbitq), 
to_sfixed(1358.0/65536.0,1,-nbitq), 
to_sfixed(-1036.0/65536.0,1,-nbitq), 
to_sfixed(-6543.0/65536.0,1,-nbitq), 
to_sfixed(11025.0/65536.0,1,-nbitq), 
to_sfixed(6182.0/65536.0,1,-nbitq), 
to_sfixed(245.0/65536.0,1,-nbitq), 
to_sfixed(5367.0/65536.0,1,-nbitq), 
to_sfixed(1901.0/65536.0,1,-nbitq), 
to_sfixed(-482.0/65536.0,1,-nbitq), 
to_sfixed(5591.0/65536.0,1,-nbitq), 
to_sfixed(-1546.0/65536.0,1,-nbitq), 
to_sfixed(439.0/65536.0,1,-nbitq), 
to_sfixed(11032.0/65536.0,1,-nbitq), 
to_sfixed(2253.0/65536.0,1,-nbitq), 
to_sfixed(-1283.0/65536.0,1,-nbitq), 
to_sfixed(943.0/65536.0,1,-nbitq), 
to_sfixed(-4215.0/65536.0,1,-nbitq), 
to_sfixed(-2960.0/65536.0,1,-nbitq), 
to_sfixed(-1181.0/65536.0,1,-nbitq), 
to_sfixed(6738.0/65536.0,1,-nbitq), 
to_sfixed(-6952.0/65536.0,1,-nbitq), 
to_sfixed(1692.0/65536.0,1,-nbitq), 
to_sfixed(9402.0/65536.0,1,-nbitq), 
to_sfixed(-1383.0/65536.0,1,-nbitq), 
to_sfixed(3659.0/65536.0,1,-nbitq), 
to_sfixed(540.0/65536.0,1,-nbitq), 
to_sfixed(4316.0/65536.0,1,-nbitq), 
to_sfixed(-5703.0/65536.0,1,-nbitq), 
to_sfixed(-1582.0/65536.0,1,-nbitq), 
to_sfixed(-5679.0/65536.0,1,-nbitq), 
to_sfixed(-4144.0/65536.0,1,-nbitq), 
to_sfixed(-1529.0/65536.0,1,-nbitq), 
to_sfixed(8943.0/65536.0,1,-nbitq), 
to_sfixed(-2044.0/65536.0,1,-nbitq), 
to_sfixed(-2451.0/65536.0,1,-nbitq), 
to_sfixed(11138.0/65536.0,1,-nbitq), 
to_sfixed(3280.0/65536.0,1,-nbitq), 
to_sfixed(12607.0/65536.0,1,-nbitq), 
to_sfixed(-1623.0/65536.0,1,-nbitq), 
to_sfixed(3165.0/65536.0,1,-nbitq), 
to_sfixed(737.0/65536.0,1,-nbitq), 
to_sfixed(4552.0/65536.0,1,-nbitq), 
to_sfixed(-349.0/65536.0,1,-nbitq), 
to_sfixed(-1600.0/65536.0,1,-nbitq), 
to_sfixed(-3362.0/65536.0,1,-nbitq), 
to_sfixed(-522.0/65536.0,1,-nbitq), 
to_sfixed(-1538.0/65536.0,1,-nbitq), 
to_sfixed(17.0/65536.0,1,-nbitq), 
to_sfixed(-1435.0/65536.0,1,-nbitq), 
to_sfixed(-2380.0/65536.0,1,-nbitq), 
to_sfixed(-7882.0/65536.0,1,-nbitq), 
to_sfixed(-8026.0/65536.0,1,-nbitq), 
to_sfixed(4426.0/65536.0,1,-nbitq), 
to_sfixed(5107.0/65536.0,1,-nbitq), 
to_sfixed(-4856.0/65536.0,1,-nbitq), 
to_sfixed(-918.0/65536.0,1,-nbitq), 
to_sfixed(-2609.0/65536.0,1,-nbitq), 
to_sfixed(-1519.0/65536.0,1,-nbitq), 
to_sfixed(-6025.0/65536.0,1,-nbitq), 
to_sfixed(4702.0/65536.0,1,-nbitq), 
to_sfixed(-2544.0/65536.0,1,-nbitq), 
to_sfixed(1332.0/65536.0,1,-nbitq), 
to_sfixed(-1891.0/65536.0,1,-nbitq), 
to_sfixed(576.0/65536.0,1,-nbitq), 
to_sfixed(-4782.0/65536.0,1,-nbitq), 
to_sfixed(-2743.0/65536.0,1,-nbitq), 
to_sfixed(3684.0/65536.0,1,-nbitq), 
to_sfixed(-3588.0/65536.0,1,-nbitq), 
to_sfixed(-1544.0/65536.0,1,-nbitq), 
to_sfixed(1058.0/65536.0,1,-nbitq), 
to_sfixed(8909.0/65536.0,1,-nbitq), 
to_sfixed(543.0/65536.0,1,-nbitq), 
to_sfixed(42.0/65536.0,1,-nbitq), 
to_sfixed(1962.0/65536.0,1,-nbitq), 
to_sfixed(2198.0/65536.0,1,-nbitq), 
to_sfixed(5460.0/65536.0,1,-nbitq), 
to_sfixed(-13510.0/65536.0,1,-nbitq), 
to_sfixed(-1659.0/65536.0,1,-nbitq), 
to_sfixed(-5834.0/65536.0,1,-nbitq)  ), 
( to_sfixed(962.0/65536.0,1,-nbitq), 
to_sfixed(379.0/65536.0,1,-nbitq), 
to_sfixed(3446.0/65536.0,1,-nbitq), 
to_sfixed(-3636.0/65536.0,1,-nbitq), 
to_sfixed(2885.0/65536.0,1,-nbitq), 
to_sfixed(5244.0/65536.0,1,-nbitq), 
to_sfixed(-982.0/65536.0,1,-nbitq), 
to_sfixed(5510.0/65536.0,1,-nbitq), 
to_sfixed(125.0/65536.0,1,-nbitq), 
to_sfixed(-65.0/65536.0,1,-nbitq), 
to_sfixed(-1726.0/65536.0,1,-nbitq), 
to_sfixed(3886.0/65536.0,1,-nbitq), 
to_sfixed(1454.0/65536.0,1,-nbitq), 
to_sfixed(12997.0/65536.0,1,-nbitq), 
to_sfixed(-2565.0/65536.0,1,-nbitq), 
to_sfixed(-1303.0/65536.0,1,-nbitq), 
to_sfixed(329.0/65536.0,1,-nbitq), 
to_sfixed(-5172.0/65536.0,1,-nbitq), 
to_sfixed(-28.0/65536.0,1,-nbitq), 
to_sfixed(3087.0/65536.0,1,-nbitq), 
to_sfixed(7374.0/65536.0,1,-nbitq), 
to_sfixed(-265.0/65536.0,1,-nbitq), 
to_sfixed(913.0/65536.0,1,-nbitq), 
to_sfixed(13050.0/65536.0,1,-nbitq), 
to_sfixed(-290.0/65536.0,1,-nbitq), 
to_sfixed(5888.0/65536.0,1,-nbitq), 
to_sfixed(1404.0/65536.0,1,-nbitq), 
to_sfixed(-570.0/65536.0,1,-nbitq), 
to_sfixed(-1699.0/65536.0,1,-nbitq), 
to_sfixed(-6576.0/65536.0,1,-nbitq), 
to_sfixed(-4608.0/65536.0,1,-nbitq), 
to_sfixed(2186.0/65536.0,1,-nbitq), 
to_sfixed(2179.0/65536.0,1,-nbitq), 
to_sfixed(3979.0/65536.0,1,-nbitq), 
to_sfixed(-1762.0/65536.0,1,-nbitq), 
to_sfixed(-4224.0/65536.0,1,-nbitq), 
to_sfixed(3451.0/65536.0,1,-nbitq), 
to_sfixed(2647.0/65536.0,1,-nbitq), 
to_sfixed(8867.0/65536.0,1,-nbitq), 
to_sfixed(-65.0/65536.0,1,-nbitq), 
to_sfixed(3752.0/65536.0,1,-nbitq), 
to_sfixed(-1532.0/65536.0,1,-nbitq), 
to_sfixed(5562.0/65536.0,1,-nbitq), 
to_sfixed(-948.0/65536.0,1,-nbitq), 
to_sfixed(3035.0/65536.0,1,-nbitq), 
to_sfixed(-1665.0/65536.0,1,-nbitq), 
to_sfixed(-2299.0/65536.0,1,-nbitq), 
to_sfixed(-9009.0/65536.0,1,-nbitq), 
to_sfixed(311.0/65536.0,1,-nbitq), 
to_sfixed(-426.0/65536.0,1,-nbitq), 
to_sfixed(-218.0/65536.0,1,-nbitq), 
to_sfixed(-2748.0/65536.0,1,-nbitq), 
to_sfixed(-7799.0/65536.0,1,-nbitq), 
to_sfixed(-2375.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(4191.0/65536.0,1,-nbitq), 
to_sfixed(1368.0/65536.0,1,-nbitq), 
to_sfixed(168.0/65536.0,1,-nbitq), 
to_sfixed(2447.0/65536.0,1,-nbitq), 
to_sfixed(-1598.0/65536.0,1,-nbitq), 
to_sfixed(1532.0/65536.0,1,-nbitq), 
to_sfixed(-2484.0/65536.0,1,-nbitq), 
to_sfixed(2953.0/65536.0,1,-nbitq), 
to_sfixed(608.0/65536.0,1,-nbitq), 
to_sfixed(329.0/65536.0,1,-nbitq), 
to_sfixed(-3556.0/65536.0,1,-nbitq), 
to_sfixed(-766.0/65536.0,1,-nbitq), 
to_sfixed(1062.0/65536.0,1,-nbitq), 
to_sfixed(-4338.0/65536.0,1,-nbitq), 
to_sfixed(-4987.0/65536.0,1,-nbitq), 
to_sfixed(3783.0/65536.0,1,-nbitq), 
to_sfixed(2291.0/65536.0,1,-nbitq), 
to_sfixed(2910.0/65536.0,1,-nbitq), 
to_sfixed(-43.0/65536.0,1,-nbitq), 
to_sfixed(642.0/65536.0,1,-nbitq), 
to_sfixed(-2230.0/65536.0,1,-nbitq), 
to_sfixed(-590.0/65536.0,1,-nbitq), 
to_sfixed(-10264.0/65536.0,1,-nbitq), 
to_sfixed(120.0/65536.0,1,-nbitq), 
to_sfixed(-4247.0/65536.0,1,-nbitq)  ), 
( to_sfixed(167.0/65536.0,1,-nbitq), 
to_sfixed(3628.0/65536.0,1,-nbitq), 
to_sfixed(-477.0/65536.0,1,-nbitq), 
to_sfixed(-512.0/65536.0,1,-nbitq), 
to_sfixed(-1933.0/65536.0,1,-nbitq), 
to_sfixed(607.0/65536.0,1,-nbitq), 
to_sfixed(-2338.0/65536.0,1,-nbitq), 
to_sfixed(7177.0/65536.0,1,-nbitq), 
to_sfixed(787.0/65536.0,1,-nbitq), 
to_sfixed(-2148.0/65536.0,1,-nbitq), 
to_sfixed(-1728.0/65536.0,1,-nbitq), 
to_sfixed(5560.0/65536.0,1,-nbitq), 
to_sfixed(1003.0/65536.0,1,-nbitq), 
to_sfixed(5984.0/65536.0,1,-nbitq), 
to_sfixed(-4201.0/65536.0,1,-nbitq), 
to_sfixed(1582.0/65536.0,1,-nbitq), 
to_sfixed(1770.0/65536.0,1,-nbitq), 
to_sfixed(-104.0/65536.0,1,-nbitq), 
to_sfixed(-228.0/65536.0,1,-nbitq), 
to_sfixed(-2539.0/65536.0,1,-nbitq), 
to_sfixed(3806.0/65536.0,1,-nbitq), 
to_sfixed(2358.0/65536.0,1,-nbitq), 
to_sfixed(-762.0/65536.0,1,-nbitq), 
to_sfixed(1145.0/65536.0,1,-nbitq), 
to_sfixed(-980.0/65536.0,1,-nbitq), 
to_sfixed(559.0/65536.0,1,-nbitq), 
to_sfixed(1220.0/65536.0,1,-nbitq), 
to_sfixed(1270.0/65536.0,1,-nbitq), 
to_sfixed(-3280.0/65536.0,1,-nbitq), 
to_sfixed(157.0/65536.0,1,-nbitq), 
to_sfixed(-5837.0/65536.0,1,-nbitq), 
to_sfixed(-3437.0/65536.0,1,-nbitq), 
to_sfixed(5599.0/65536.0,1,-nbitq), 
to_sfixed(5774.0/65536.0,1,-nbitq), 
to_sfixed(-1665.0/65536.0,1,-nbitq), 
to_sfixed(-793.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(-1208.0/65536.0,1,-nbitq), 
to_sfixed(5553.0/65536.0,1,-nbitq), 
to_sfixed(634.0/65536.0,1,-nbitq), 
to_sfixed(5291.0/65536.0,1,-nbitq), 
to_sfixed(1872.0/65536.0,1,-nbitq), 
to_sfixed(8540.0/65536.0,1,-nbitq), 
to_sfixed(-1966.0/65536.0,1,-nbitq), 
to_sfixed(2289.0/65536.0,1,-nbitq), 
to_sfixed(-893.0/65536.0,1,-nbitq), 
to_sfixed(90.0/65536.0,1,-nbitq), 
to_sfixed(-3759.0/65536.0,1,-nbitq), 
to_sfixed(727.0/65536.0,1,-nbitq), 
to_sfixed(1753.0/65536.0,1,-nbitq), 
to_sfixed(2687.0/65536.0,1,-nbitq), 
to_sfixed(985.0/65536.0,1,-nbitq), 
to_sfixed(-873.0/65536.0,1,-nbitq), 
to_sfixed(-7507.0/65536.0,1,-nbitq), 
to_sfixed(-484.0/65536.0,1,-nbitq), 
to_sfixed(5157.0/65536.0,1,-nbitq), 
to_sfixed(-2571.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(-1805.0/65536.0,1,-nbitq), 
to_sfixed(-4165.0/65536.0,1,-nbitq), 
to_sfixed(-3404.0/65536.0,1,-nbitq), 
to_sfixed(655.0/65536.0,1,-nbitq), 
to_sfixed(1938.0/65536.0,1,-nbitq), 
to_sfixed(-3182.0/65536.0,1,-nbitq), 
to_sfixed(-3146.0/65536.0,1,-nbitq), 
to_sfixed(-6485.0/65536.0,1,-nbitq), 
to_sfixed(-377.0/65536.0,1,-nbitq), 
to_sfixed(-229.0/65536.0,1,-nbitq), 
to_sfixed(-4725.0/65536.0,1,-nbitq), 
to_sfixed(-8126.0/65536.0,1,-nbitq), 
to_sfixed(6414.0/65536.0,1,-nbitq), 
to_sfixed(1778.0/65536.0,1,-nbitq), 
to_sfixed(-80.0/65536.0,1,-nbitq), 
to_sfixed(1191.0/65536.0,1,-nbitq), 
to_sfixed(2325.0/65536.0,1,-nbitq), 
to_sfixed(4510.0/65536.0,1,-nbitq), 
to_sfixed(6312.0/65536.0,1,-nbitq), 
to_sfixed(-2037.0/65536.0,1,-nbitq), 
to_sfixed(2321.0/65536.0,1,-nbitq), 
to_sfixed(-6896.0/65536.0,1,-nbitq)  ), 
( to_sfixed(6533.0/65536.0,1,-nbitq), 
to_sfixed(2267.0/65536.0,1,-nbitq), 
to_sfixed(-192.0/65536.0,1,-nbitq), 
to_sfixed(1246.0/65536.0,1,-nbitq), 
to_sfixed(-7013.0/65536.0,1,-nbitq), 
to_sfixed(723.0/65536.0,1,-nbitq), 
to_sfixed(765.0/65536.0,1,-nbitq), 
to_sfixed(1941.0/65536.0,1,-nbitq), 
to_sfixed(-2878.0/65536.0,1,-nbitq), 
to_sfixed(-2439.0/65536.0,1,-nbitq), 
to_sfixed(-615.0/65536.0,1,-nbitq), 
to_sfixed(6244.0/65536.0,1,-nbitq), 
to_sfixed(1898.0/65536.0,1,-nbitq), 
to_sfixed(-1010.0/65536.0,1,-nbitq), 
to_sfixed(-2632.0/65536.0,1,-nbitq), 
to_sfixed(-2638.0/65536.0,1,-nbitq), 
to_sfixed(2410.0/65536.0,1,-nbitq), 
to_sfixed(-1970.0/65536.0,1,-nbitq), 
to_sfixed(-5332.0/65536.0,1,-nbitq), 
to_sfixed(3441.0/65536.0,1,-nbitq), 
to_sfixed(1116.0/65536.0,1,-nbitq), 
to_sfixed(2493.0/65536.0,1,-nbitq), 
to_sfixed(-6432.0/65536.0,1,-nbitq), 
to_sfixed(-1065.0/65536.0,1,-nbitq), 
to_sfixed(1991.0/65536.0,1,-nbitq), 
to_sfixed(-2974.0/65536.0,1,-nbitq), 
to_sfixed(2419.0/65536.0,1,-nbitq), 
to_sfixed(1347.0/65536.0,1,-nbitq), 
to_sfixed(-219.0/65536.0,1,-nbitq), 
to_sfixed(1278.0/65536.0,1,-nbitq), 
to_sfixed(-4182.0/65536.0,1,-nbitq), 
to_sfixed(-1068.0/65536.0,1,-nbitq), 
to_sfixed(7257.0/65536.0,1,-nbitq), 
to_sfixed(8506.0/65536.0,1,-nbitq), 
to_sfixed(-735.0/65536.0,1,-nbitq), 
to_sfixed(1424.0/65536.0,1,-nbitq), 
to_sfixed(-1439.0/65536.0,1,-nbitq), 
to_sfixed(3400.0/65536.0,1,-nbitq), 
to_sfixed(6546.0/65536.0,1,-nbitq), 
to_sfixed(-1353.0/65536.0,1,-nbitq), 
to_sfixed(6076.0/65536.0,1,-nbitq), 
to_sfixed(-2902.0/65536.0,1,-nbitq), 
to_sfixed(8185.0/65536.0,1,-nbitq), 
to_sfixed(-5501.0/65536.0,1,-nbitq), 
to_sfixed(-1502.0/65536.0,1,-nbitq), 
to_sfixed(-8973.0/65536.0,1,-nbitq), 
to_sfixed(-3216.0/65536.0,1,-nbitq), 
to_sfixed(-2634.0/65536.0,1,-nbitq), 
to_sfixed(-457.0/65536.0,1,-nbitq), 
to_sfixed(-755.0/65536.0,1,-nbitq), 
to_sfixed(2269.0/65536.0,1,-nbitq), 
to_sfixed(-2942.0/65536.0,1,-nbitq), 
to_sfixed(6097.0/65536.0,1,-nbitq), 
to_sfixed(-4741.0/65536.0,1,-nbitq), 
to_sfixed(486.0/65536.0,1,-nbitq), 
to_sfixed(555.0/65536.0,1,-nbitq), 
to_sfixed(-2958.0/65536.0,1,-nbitq), 
to_sfixed(2143.0/65536.0,1,-nbitq), 
to_sfixed(-506.0/65536.0,1,-nbitq), 
to_sfixed(918.0/65536.0,1,-nbitq), 
to_sfixed(-1679.0/65536.0,1,-nbitq), 
to_sfixed(-2265.0/65536.0,1,-nbitq), 
to_sfixed(3127.0/65536.0,1,-nbitq), 
to_sfixed(1135.0/65536.0,1,-nbitq), 
to_sfixed(-6156.0/65536.0,1,-nbitq), 
to_sfixed(-69.0/65536.0,1,-nbitq), 
to_sfixed(-1944.0/65536.0,1,-nbitq), 
to_sfixed(77.0/65536.0,1,-nbitq), 
to_sfixed(-9851.0/65536.0,1,-nbitq), 
to_sfixed(-7786.0/65536.0,1,-nbitq), 
to_sfixed(6405.0/65536.0,1,-nbitq), 
to_sfixed(-205.0/65536.0,1,-nbitq), 
to_sfixed(572.0/65536.0,1,-nbitq), 
to_sfixed(-1358.0/65536.0,1,-nbitq), 
to_sfixed(-1116.0/65536.0,1,-nbitq), 
to_sfixed(1689.0/65536.0,1,-nbitq), 
to_sfixed(-1866.0/65536.0,1,-nbitq), 
to_sfixed(-2479.0/65536.0,1,-nbitq), 
to_sfixed(582.0/65536.0,1,-nbitq), 
to_sfixed(-13563.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4552.0/65536.0,1,-nbitq), 
to_sfixed(2667.0/65536.0,1,-nbitq), 
to_sfixed(-2050.0/65536.0,1,-nbitq), 
to_sfixed(-98.0/65536.0,1,-nbitq), 
to_sfixed(-1939.0/65536.0,1,-nbitq), 
to_sfixed(3954.0/65536.0,1,-nbitq), 
to_sfixed(2220.0/65536.0,1,-nbitq), 
to_sfixed(-1720.0/65536.0,1,-nbitq), 
to_sfixed(-1952.0/65536.0,1,-nbitq), 
to_sfixed(31.0/65536.0,1,-nbitq), 
to_sfixed(677.0/65536.0,1,-nbitq), 
to_sfixed(2181.0/65536.0,1,-nbitq), 
to_sfixed(195.0/65536.0,1,-nbitq), 
to_sfixed(3338.0/65536.0,1,-nbitq), 
to_sfixed(-1362.0/65536.0,1,-nbitq), 
to_sfixed(-166.0/65536.0,1,-nbitq), 
to_sfixed(144.0/65536.0,1,-nbitq), 
to_sfixed(-844.0/65536.0,1,-nbitq), 
to_sfixed(79.0/65536.0,1,-nbitq), 
to_sfixed(-940.0/65536.0,1,-nbitq), 
to_sfixed(3306.0/65536.0,1,-nbitq), 
to_sfixed(1138.0/65536.0,1,-nbitq), 
to_sfixed(-4684.0/65536.0,1,-nbitq), 
to_sfixed(7230.0/65536.0,1,-nbitq), 
to_sfixed(2518.0/65536.0,1,-nbitq), 
to_sfixed(5941.0/65536.0,1,-nbitq), 
to_sfixed(3931.0/65536.0,1,-nbitq), 
to_sfixed(-1771.0/65536.0,1,-nbitq), 
to_sfixed(1201.0/65536.0,1,-nbitq), 
to_sfixed(1235.0/65536.0,1,-nbitq), 
to_sfixed(-3949.0/65536.0,1,-nbitq), 
to_sfixed(2325.0/65536.0,1,-nbitq), 
to_sfixed(8439.0/65536.0,1,-nbitq), 
to_sfixed(3967.0/65536.0,1,-nbitq), 
to_sfixed(-1818.0/65536.0,1,-nbitq), 
to_sfixed(-628.0/65536.0,1,-nbitq), 
to_sfixed(556.0/65536.0,1,-nbitq), 
to_sfixed(1724.0/65536.0,1,-nbitq), 
to_sfixed(-846.0/65536.0,1,-nbitq), 
to_sfixed(2606.0/65536.0,1,-nbitq), 
to_sfixed(3189.0/65536.0,1,-nbitq), 
to_sfixed(461.0/65536.0,1,-nbitq), 
to_sfixed(3726.0/65536.0,1,-nbitq), 
to_sfixed(-2563.0/65536.0,1,-nbitq), 
to_sfixed(948.0/65536.0,1,-nbitq), 
to_sfixed(-3450.0/65536.0,1,-nbitq), 
to_sfixed(-1056.0/65536.0,1,-nbitq), 
to_sfixed(-3497.0/65536.0,1,-nbitq), 
to_sfixed(-1085.0/65536.0,1,-nbitq), 
to_sfixed(1067.0/65536.0,1,-nbitq), 
to_sfixed(1018.0/65536.0,1,-nbitq), 
to_sfixed(-842.0/65536.0,1,-nbitq), 
to_sfixed(8978.0/65536.0,1,-nbitq), 
to_sfixed(-6605.0/65536.0,1,-nbitq), 
to_sfixed(6728.0/65536.0,1,-nbitq), 
to_sfixed(147.0/65536.0,1,-nbitq), 
to_sfixed(2748.0/65536.0,1,-nbitq), 
to_sfixed(-1399.0/65536.0,1,-nbitq), 
to_sfixed(-1449.0/65536.0,1,-nbitq), 
to_sfixed(169.0/65536.0,1,-nbitq), 
to_sfixed(-1296.0/65536.0,1,-nbitq), 
to_sfixed(-265.0/65536.0,1,-nbitq), 
to_sfixed(2050.0/65536.0,1,-nbitq), 
to_sfixed(134.0/65536.0,1,-nbitq), 
to_sfixed(-1137.0/65536.0,1,-nbitq), 
to_sfixed(3148.0/65536.0,1,-nbitq), 
to_sfixed(-3199.0/65536.0,1,-nbitq), 
to_sfixed(-167.0/65536.0,1,-nbitq), 
to_sfixed(-6853.0/65536.0,1,-nbitq), 
to_sfixed(-7615.0/65536.0,1,-nbitq), 
to_sfixed(5972.0/65536.0,1,-nbitq), 
to_sfixed(578.0/65536.0,1,-nbitq), 
to_sfixed(1548.0/65536.0,1,-nbitq), 
to_sfixed(-2501.0/65536.0,1,-nbitq), 
to_sfixed(2293.0/65536.0,1,-nbitq), 
to_sfixed(1717.0/65536.0,1,-nbitq), 
to_sfixed(-1305.0/65536.0,1,-nbitq), 
to_sfixed(-2416.0/65536.0,1,-nbitq), 
to_sfixed(-2109.0/65536.0,1,-nbitq), 
to_sfixed(-5751.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-299.0/65536.0,1,-nbitq), 
to_sfixed(-1637.0/65536.0,1,-nbitq), 
to_sfixed(2020.0/65536.0,1,-nbitq), 
to_sfixed(-2844.0/65536.0,1,-nbitq), 
to_sfixed(-642.0/65536.0,1,-nbitq), 
to_sfixed(1221.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(-2360.0/65536.0,1,-nbitq), 
to_sfixed(-556.0/65536.0,1,-nbitq), 
to_sfixed(1771.0/65536.0,1,-nbitq), 
to_sfixed(-131.0/65536.0,1,-nbitq), 
to_sfixed(-2613.0/65536.0,1,-nbitq), 
to_sfixed(-2349.0/65536.0,1,-nbitq), 
to_sfixed(1403.0/65536.0,1,-nbitq), 
to_sfixed(-3676.0/65536.0,1,-nbitq), 
to_sfixed(2177.0/65536.0,1,-nbitq), 
to_sfixed(-2783.0/65536.0,1,-nbitq), 
to_sfixed(-2407.0/65536.0,1,-nbitq), 
to_sfixed(112.0/65536.0,1,-nbitq), 
to_sfixed(1600.0/65536.0,1,-nbitq), 
to_sfixed(-190.0/65536.0,1,-nbitq), 
to_sfixed(962.0/65536.0,1,-nbitq), 
to_sfixed(-771.0/65536.0,1,-nbitq), 
to_sfixed(3487.0/65536.0,1,-nbitq), 
to_sfixed(3219.0/65536.0,1,-nbitq), 
to_sfixed(2871.0/65536.0,1,-nbitq), 
to_sfixed(4452.0/65536.0,1,-nbitq), 
to_sfixed(2576.0/65536.0,1,-nbitq), 
to_sfixed(1256.0/65536.0,1,-nbitq), 
to_sfixed(674.0/65536.0,1,-nbitq), 
to_sfixed(-2674.0/65536.0,1,-nbitq), 
to_sfixed(4393.0/65536.0,1,-nbitq), 
to_sfixed(4878.0/65536.0,1,-nbitq), 
to_sfixed(1878.0/65536.0,1,-nbitq), 
to_sfixed(1005.0/65536.0,1,-nbitq), 
to_sfixed(-1420.0/65536.0,1,-nbitq), 
to_sfixed(3703.0/65536.0,1,-nbitq), 
to_sfixed(240.0/65536.0,1,-nbitq), 
to_sfixed(-1865.0/65536.0,1,-nbitq), 
to_sfixed(3678.0/65536.0,1,-nbitq), 
to_sfixed(3222.0/65536.0,1,-nbitq), 
to_sfixed(1929.0/65536.0,1,-nbitq), 
to_sfixed(4036.0/65536.0,1,-nbitq), 
to_sfixed(1548.0/65536.0,1,-nbitq), 
to_sfixed(2213.0/65536.0,1,-nbitq), 
to_sfixed(-1268.0/65536.0,1,-nbitq), 
to_sfixed(-2132.0/65536.0,1,-nbitq), 
to_sfixed(-4600.0/65536.0,1,-nbitq), 
to_sfixed(-463.0/65536.0,1,-nbitq), 
to_sfixed(4446.0/65536.0,1,-nbitq), 
to_sfixed(-782.0/65536.0,1,-nbitq), 
to_sfixed(-2620.0/65536.0,1,-nbitq), 
to_sfixed(9458.0/65536.0,1,-nbitq), 
to_sfixed(-5788.0/65536.0,1,-nbitq), 
to_sfixed(6886.0/65536.0,1,-nbitq), 
to_sfixed(4429.0/65536.0,1,-nbitq), 
to_sfixed(903.0/65536.0,1,-nbitq), 
to_sfixed(-1745.0/65536.0,1,-nbitq), 
to_sfixed(3033.0/65536.0,1,-nbitq), 
to_sfixed(3859.0/65536.0,1,-nbitq), 
to_sfixed(846.0/65536.0,1,-nbitq), 
to_sfixed(-232.0/65536.0,1,-nbitq), 
to_sfixed(413.0/65536.0,1,-nbitq), 
to_sfixed(-2017.0/65536.0,1,-nbitq), 
to_sfixed(-828.0/65536.0,1,-nbitq), 
to_sfixed(-2110.0/65536.0,1,-nbitq), 
to_sfixed(86.0/65536.0,1,-nbitq), 
to_sfixed(-2398.0/65536.0,1,-nbitq), 
to_sfixed(-6768.0/65536.0,1,-nbitq), 
to_sfixed(-6439.0/65536.0,1,-nbitq), 
to_sfixed(5850.0/65536.0,1,-nbitq), 
to_sfixed(-2027.0/65536.0,1,-nbitq), 
to_sfixed(-161.0/65536.0,1,-nbitq), 
to_sfixed(1489.0/65536.0,1,-nbitq), 
to_sfixed(908.0/65536.0,1,-nbitq), 
to_sfixed(1746.0/65536.0,1,-nbitq), 
to_sfixed(-1593.0/65536.0,1,-nbitq), 
to_sfixed(-722.0/65536.0,1,-nbitq), 
to_sfixed(1580.0/65536.0,1,-nbitq), 
to_sfixed(-2660.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2190.0/65536.0,1,-nbitq), 
to_sfixed(-3890.0/65536.0,1,-nbitq), 
to_sfixed(3198.0/65536.0,1,-nbitq), 
to_sfixed(-1807.0/65536.0,1,-nbitq), 
to_sfixed(-2269.0/65536.0,1,-nbitq), 
to_sfixed(-725.0/65536.0,1,-nbitq), 
to_sfixed(-886.0/65536.0,1,-nbitq), 
to_sfixed(2230.0/65536.0,1,-nbitq), 
to_sfixed(520.0/65536.0,1,-nbitq), 
to_sfixed(1037.0/65536.0,1,-nbitq), 
to_sfixed(526.0/65536.0,1,-nbitq), 
to_sfixed(-833.0/65536.0,1,-nbitq), 
to_sfixed(-2453.0/65536.0,1,-nbitq), 
to_sfixed(-3529.0/65536.0,1,-nbitq), 
to_sfixed(-3082.0/65536.0,1,-nbitq), 
to_sfixed(2198.0/65536.0,1,-nbitq), 
to_sfixed(-1406.0/65536.0,1,-nbitq), 
to_sfixed(-5141.0/65536.0,1,-nbitq), 
to_sfixed(-2989.0/65536.0,1,-nbitq), 
to_sfixed(1967.0/65536.0,1,-nbitq), 
to_sfixed(-905.0/65536.0,1,-nbitq), 
to_sfixed(250.0/65536.0,1,-nbitq), 
to_sfixed(-3425.0/65536.0,1,-nbitq), 
to_sfixed(5198.0/65536.0,1,-nbitq), 
to_sfixed(3742.0/65536.0,1,-nbitq), 
to_sfixed(700.0/65536.0,1,-nbitq), 
to_sfixed(3178.0/65536.0,1,-nbitq), 
to_sfixed(-1445.0/65536.0,1,-nbitq), 
to_sfixed(2658.0/65536.0,1,-nbitq), 
to_sfixed(2995.0/65536.0,1,-nbitq), 
to_sfixed(2320.0/65536.0,1,-nbitq), 
to_sfixed(965.0/65536.0,1,-nbitq), 
to_sfixed(4293.0/65536.0,1,-nbitq), 
to_sfixed(742.0/65536.0,1,-nbitq), 
to_sfixed(-2715.0/65536.0,1,-nbitq), 
to_sfixed(770.0/65536.0,1,-nbitq), 
to_sfixed(-1172.0/65536.0,1,-nbitq), 
to_sfixed(-3816.0/65536.0,1,-nbitq), 
to_sfixed(-317.0/65536.0,1,-nbitq), 
to_sfixed(384.0/65536.0,1,-nbitq), 
to_sfixed(-489.0/65536.0,1,-nbitq), 
to_sfixed(1650.0/65536.0,1,-nbitq), 
to_sfixed(2936.0/65536.0,1,-nbitq), 
to_sfixed(1992.0/65536.0,1,-nbitq), 
to_sfixed(-984.0/65536.0,1,-nbitq), 
to_sfixed(3738.0/65536.0,1,-nbitq), 
to_sfixed(651.0/65536.0,1,-nbitq), 
to_sfixed(-3701.0/65536.0,1,-nbitq), 
to_sfixed(1423.0/65536.0,1,-nbitq), 
to_sfixed(509.0/65536.0,1,-nbitq), 
to_sfixed(-393.0/65536.0,1,-nbitq), 
to_sfixed(-594.0/65536.0,1,-nbitq), 
to_sfixed(7720.0/65536.0,1,-nbitq), 
to_sfixed(-2287.0/65536.0,1,-nbitq), 
to_sfixed(6159.0/65536.0,1,-nbitq), 
to_sfixed(816.0/65536.0,1,-nbitq), 
to_sfixed(2493.0/65536.0,1,-nbitq), 
to_sfixed(-3765.0/65536.0,1,-nbitq), 
to_sfixed(1862.0/65536.0,1,-nbitq), 
to_sfixed(5232.0/65536.0,1,-nbitq), 
to_sfixed(845.0/65536.0,1,-nbitq), 
to_sfixed(2156.0/65536.0,1,-nbitq), 
to_sfixed(-690.0/65536.0,1,-nbitq), 
to_sfixed(1846.0/65536.0,1,-nbitq), 
to_sfixed(585.0/65536.0,1,-nbitq), 
to_sfixed(3972.0/65536.0,1,-nbitq), 
to_sfixed(-1818.0/65536.0,1,-nbitq), 
to_sfixed(-3009.0/65536.0,1,-nbitq), 
to_sfixed(-1772.0/65536.0,1,-nbitq), 
to_sfixed(-2433.0/65536.0,1,-nbitq), 
to_sfixed(1417.0/65536.0,1,-nbitq), 
to_sfixed(-495.0/65536.0,1,-nbitq), 
to_sfixed(1825.0/65536.0,1,-nbitq), 
to_sfixed(-3215.0/65536.0,1,-nbitq), 
to_sfixed(-2573.0/65536.0,1,-nbitq), 
to_sfixed(1627.0/65536.0,1,-nbitq), 
to_sfixed(-2583.0/65536.0,1,-nbitq), 
to_sfixed(1323.0/65536.0,1,-nbitq), 
to_sfixed(-1591.0/65536.0,1,-nbitq), 
to_sfixed(2218.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-541.0/65536.0,1,-nbitq), 
to_sfixed(-3400.0/65536.0,1,-nbitq), 
to_sfixed(-978.0/65536.0,1,-nbitq), 
to_sfixed(-1461.0/65536.0,1,-nbitq), 
to_sfixed(-2692.0/65536.0,1,-nbitq), 
to_sfixed(-1970.0/65536.0,1,-nbitq), 
to_sfixed(1519.0/65536.0,1,-nbitq), 
to_sfixed(-1651.0/65536.0,1,-nbitq), 
to_sfixed(-2763.0/65536.0,1,-nbitq), 
to_sfixed(-1642.0/65536.0,1,-nbitq), 
to_sfixed(-3774.0/65536.0,1,-nbitq), 
to_sfixed(1269.0/65536.0,1,-nbitq), 
to_sfixed(2735.0/65536.0,1,-nbitq), 
to_sfixed(-2354.0/65536.0,1,-nbitq), 
to_sfixed(-3215.0/65536.0,1,-nbitq), 
to_sfixed(-643.0/65536.0,1,-nbitq), 
to_sfixed(1015.0/65536.0,1,-nbitq), 
to_sfixed(-2801.0/65536.0,1,-nbitq), 
to_sfixed(-1796.0/65536.0,1,-nbitq), 
to_sfixed(-1336.0/65536.0,1,-nbitq), 
to_sfixed(-3127.0/65536.0,1,-nbitq), 
to_sfixed(506.0/65536.0,1,-nbitq), 
to_sfixed(-1325.0/65536.0,1,-nbitq), 
to_sfixed(2005.0/65536.0,1,-nbitq), 
to_sfixed(1661.0/65536.0,1,-nbitq), 
to_sfixed(-682.0/65536.0,1,-nbitq), 
to_sfixed(81.0/65536.0,1,-nbitq), 
to_sfixed(-251.0/65536.0,1,-nbitq), 
to_sfixed(525.0/65536.0,1,-nbitq), 
to_sfixed(-2434.0/65536.0,1,-nbitq), 
to_sfixed(2135.0/65536.0,1,-nbitq), 
to_sfixed(-2023.0/65536.0,1,-nbitq), 
to_sfixed(1870.0/65536.0,1,-nbitq), 
to_sfixed(-2462.0/65536.0,1,-nbitq), 
to_sfixed(-2657.0/65536.0,1,-nbitq), 
to_sfixed(-822.0/65536.0,1,-nbitq), 
to_sfixed(-987.0/65536.0,1,-nbitq), 
to_sfixed(-1451.0/65536.0,1,-nbitq), 
to_sfixed(-2586.0/65536.0,1,-nbitq), 
to_sfixed(-2705.0/65536.0,1,-nbitq), 
to_sfixed(1541.0/65536.0,1,-nbitq), 
to_sfixed(330.0/65536.0,1,-nbitq), 
to_sfixed(1190.0/65536.0,1,-nbitq), 
to_sfixed(1150.0/65536.0,1,-nbitq), 
to_sfixed(3160.0/65536.0,1,-nbitq), 
to_sfixed(914.0/65536.0,1,-nbitq), 
to_sfixed(-3347.0/65536.0,1,-nbitq), 
to_sfixed(1991.0/65536.0,1,-nbitq), 
to_sfixed(-365.0/65536.0,1,-nbitq), 
to_sfixed(-23.0/65536.0,1,-nbitq), 
to_sfixed(3340.0/65536.0,1,-nbitq), 
to_sfixed(-4250.0/65536.0,1,-nbitq), 
to_sfixed(803.0/65536.0,1,-nbitq), 
to_sfixed(1348.0/65536.0,1,-nbitq), 
to_sfixed(-103.0/65536.0,1,-nbitq), 
to_sfixed(2807.0/65536.0,1,-nbitq), 
to_sfixed(1078.0/65536.0,1,-nbitq), 
to_sfixed(2177.0/65536.0,1,-nbitq), 
to_sfixed(-824.0/65536.0,1,-nbitq), 
to_sfixed(3827.0/65536.0,1,-nbitq), 
to_sfixed(-2255.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(-1617.0/65536.0,1,-nbitq), 
to_sfixed(709.0/65536.0,1,-nbitq), 
to_sfixed(-1298.0/65536.0,1,-nbitq), 
to_sfixed(64.0/65536.0,1,-nbitq), 
to_sfixed(1629.0/65536.0,1,-nbitq), 
to_sfixed(-1532.0/65536.0,1,-nbitq), 
to_sfixed(-4308.0/65536.0,1,-nbitq), 
to_sfixed(1648.0/65536.0,1,-nbitq), 
to_sfixed(1422.0/65536.0,1,-nbitq), 
to_sfixed(-2915.0/65536.0,1,-nbitq), 
to_sfixed(2752.0/65536.0,1,-nbitq), 
to_sfixed(1465.0/65536.0,1,-nbitq), 
to_sfixed(2336.0/65536.0,1,-nbitq), 
to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(-2321.0/65536.0,1,-nbitq), 
to_sfixed(1313.0/65536.0,1,-nbitq), 
to_sfixed(408.0/65536.0,1,-nbitq), 
to_sfixed(-973.0/65536.0,1,-nbitq)  ), 
( to_sfixed(689.0/65536.0,1,-nbitq), 
to_sfixed(893.0/65536.0,1,-nbitq), 
to_sfixed(591.0/65536.0,1,-nbitq), 
to_sfixed(1140.0/65536.0,1,-nbitq), 
to_sfixed(1784.0/65536.0,1,-nbitq), 
to_sfixed(-4097.0/65536.0,1,-nbitq), 
to_sfixed(-1321.0/65536.0,1,-nbitq), 
to_sfixed(-59.0/65536.0,1,-nbitq), 
to_sfixed(-1966.0/65536.0,1,-nbitq), 
to_sfixed(-804.0/65536.0,1,-nbitq), 
to_sfixed(1555.0/65536.0,1,-nbitq), 
to_sfixed(2907.0/65536.0,1,-nbitq), 
to_sfixed(1259.0/65536.0,1,-nbitq), 
to_sfixed(-4156.0/65536.0,1,-nbitq), 
to_sfixed(-954.0/65536.0,1,-nbitq), 
to_sfixed(1432.0/65536.0,1,-nbitq), 
to_sfixed(1585.0/65536.0,1,-nbitq), 
to_sfixed(2385.0/65536.0,1,-nbitq), 
to_sfixed(2059.0/65536.0,1,-nbitq), 
to_sfixed(1360.0/65536.0,1,-nbitq), 
to_sfixed(296.0/65536.0,1,-nbitq), 
to_sfixed(1544.0/65536.0,1,-nbitq), 
to_sfixed(-3022.0/65536.0,1,-nbitq), 
to_sfixed(-86.0/65536.0,1,-nbitq), 
to_sfixed(-361.0/65536.0,1,-nbitq), 
to_sfixed(63.0/65536.0,1,-nbitq), 
to_sfixed(-3567.0/65536.0,1,-nbitq), 
to_sfixed(100.0/65536.0,1,-nbitq), 
to_sfixed(-2633.0/65536.0,1,-nbitq), 
to_sfixed(-1432.0/65536.0,1,-nbitq), 
to_sfixed(-1243.0/65536.0,1,-nbitq), 
to_sfixed(1011.0/65536.0,1,-nbitq), 
to_sfixed(-2490.0/65536.0,1,-nbitq), 
to_sfixed(-4104.0/65536.0,1,-nbitq), 
to_sfixed(-1374.0/65536.0,1,-nbitq), 
to_sfixed(-1206.0/65536.0,1,-nbitq), 
to_sfixed(-3535.0/65536.0,1,-nbitq), 
to_sfixed(-2477.0/65536.0,1,-nbitq), 
to_sfixed(-2464.0/65536.0,1,-nbitq), 
to_sfixed(2903.0/65536.0,1,-nbitq), 
to_sfixed(-1399.0/65536.0,1,-nbitq), 
to_sfixed(1103.0/65536.0,1,-nbitq), 
to_sfixed(-3569.0/65536.0,1,-nbitq), 
to_sfixed(-947.0/65536.0,1,-nbitq), 
to_sfixed(881.0/65536.0,1,-nbitq), 
to_sfixed(3624.0/65536.0,1,-nbitq), 
to_sfixed(-944.0/65536.0,1,-nbitq), 
to_sfixed(1194.0/65536.0,1,-nbitq), 
to_sfixed(2957.0/65536.0,1,-nbitq), 
to_sfixed(2634.0/65536.0,1,-nbitq), 
to_sfixed(-331.0/65536.0,1,-nbitq), 
to_sfixed(-1705.0/65536.0,1,-nbitq), 
to_sfixed(-806.0/65536.0,1,-nbitq), 
to_sfixed(1515.0/65536.0,1,-nbitq), 
to_sfixed(-908.0/65536.0,1,-nbitq), 
to_sfixed(2592.0/65536.0,1,-nbitq), 
to_sfixed(274.0/65536.0,1,-nbitq), 
to_sfixed(-1123.0/65536.0,1,-nbitq), 
to_sfixed(-2907.0/65536.0,1,-nbitq), 
to_sfixed(5331.0/65536.0,1,-nbitq), 
to_sfixed(1375.0/65536.0,1,-nbitq), 
to_sfixed(2379.0/65536.0,1,-nbitq), 
to_sfixed(-1028.0/65536.0,1,-nbitq), 
to_sfixed(-1238.0/65536.0,1,-nbitq), 
to_sfixed(-1155.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(-2057.0/65536.0,1,-nbitq), 
to_sfixed(-2850.0/65536.0,1,-nbitq), 
to_sfixed(2101.0/65536.0,1,-nbitq), 
to_sfixed(2543.0/65536.0,1,-nbitq), 
to_sfixed(178.0/65536.0,1,-nbitq), 
to_sfixed(1775.0/65536.0,1,-nbitq), 
to_sfixed(684.0/65536.0,1,-nbitq), 
to_sfixed(1094.0/65536.0,1,-nbitq), 
to_sfixed(2193.0/65536.0,1,-nbitq), 
to_sfixed(1318.0/65536.0,1,-nbitq), 
to_sfixed(41.0/65536.0,1,-nbitq), 
to_sfixed(3754.0/65536.0,1,-nbitq), 
to_sfixed(1943.0/65536.0,1,-nbitq), 
to_sfixed(2660.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1153.0/65536.0,1,-nbitq), 
to_sfixed(-1471.0/65536.0,1,-nbitq), 
to_sfixed(-1979.0/65536.0,1,-nbitq), 
to_sfixed(1640.0/65536.0,1,-nbitq), 
to_sfixed(1444.0/65536.0,1,-nbitq), 
to_sfixed(-439.0/65536.0,1,-nbitq), 
to_sfixed(-334.0/65536.0,1,-nbitq), 
to_sfixed(-1705.0/65536.0,1,-nbitq), 
to_sfixed(-1984.0/65536.0,1,-nbitq), 
to_sfixed(411.0/65536.0,1,-nbitq), 
to_sfixed(-1851.0/65536.0,1,-nbitq), 
to_sfixed(-1499.0/65536.0,1,-nbitq), 
to_sfixed(3216.0/65536.0,1,-nbitq), 
to_sfixed(582.0/65536.0,1,-nbitq), 
to_sfixed(1518.0/65536.0,1,-nbitq), 
to_sfixed(-360.0/65536.0,1,-nbitq), 
to_sfixed(-2891.0/65536.0,1,-nbitq), 
to_sfixed(-1363.0/65536.0,1,-nbitq), 
to_sfixed(-1531.0/65536.0,1,-nbitq), 
to_sfixed(-1622.0/65536.0,1,-nbitq), 
to_sfixed(-313.0/65536.0,1,-nbitq), 
to_sfixed(-1392.0/65536.0,1,-nbitq), 
to_sfixed(1531.0/65536.0,1,-nbitq), 
to_sfixed(-162.0/65536.0,1,-nbitq), 
to_sfixed(407.0/65536.0,1,-nbitq), 
to_sfixed(-483.0/65536.0,1,-nbitq), 
to_sfixed(901.0/65536.0,1,-nbitq), 
to_sfixed(2730.0/65536.0,1,-nbitq), 
to_sfixed(-1948.0/65536.0,1,-nbitq), 
to_sfixed(-1521.0/65536.0,1,-nbitq), 
to_sfixed(2499.0/65536.0,1,-nbitq), 
to_sfixed(-1663.0/65536.0,1,-nbitq), 
to_sfixed(1026.0/65536.0,1,-nbitq), 
to_sfixed(-1128.0/65536.0,1,-nbitq), 
to_sfixed(-1714.0/65536.0,1,-nbitq), 
to_sfixed(-788.0/65536.0,1,-nbitq), 
to_sfixed(-2188.0/65536.0,1,-nbitq), 
to_sfixed(1322.0/65536.0,1,-nbitq), 
to_sfixed(-2074.0/65536.0,1,-nbitq), 
to_sfixed(2305.0/65536.0,1,-nbitq), 
to_sfixed(-3374.0/65536.0,1,-nbitq), 
to_sfixed(691.0/65536.0,1,-nbitq), 
to_sfixed(-1793.0/65536.0,1,-nbitq), 
to_sfixed(-1725.0/65536.0,1,-nbitq), 
to_sfixed(1326.0/65536.0,1,-nbitq), 
to_sfixed(212.0/65536.0,1,-nbitq), 
to_sfixed(802.0/65536.0,1,-nbitq), 
to_sfixed(653.0/65536.0,1,-nbitq), 
to_sfixed(3524.0/65536.0,1,-nbitq), 
to_sfixed(-915.0/65536.0,1,-nbitq), 
to_sfixed(182.0/65536.0,1,-nbitq), 
to_sfixed(-3258.0/65536.0,1,-nbitq), 
to_sfixed(3162.0/65536.0,1,-nbitq), 
to_sfixed(-1164.0/65536.0,1,-nbitq), 
to_sfixed(-1201.0/65536.0,1,-nbitq), 
to_sfixed(692.0/65536.0,1,-nbitq), 
to_sfixed(-2463.0/65536.0,1,-nbitq), 
to_sfixed(2344.0/65536.0,1,-nbitq), 
to_sfixed(-1537.0/65536.0,1,-nbitq), 
to_sfixed(3162.0/65536.0,1,-nbitq), 
to_sfixed(170.0/65536.0,1,-nbitq), 
to_sfixed(87.0/65536.0,1,-nbitq), 
to_sfixed(-1629.0/65536.0,1,-nbitq), 
to_sfixed(-455.0/65536.0,1,-nbitq), 
to_sfixed(976.0/65536.0,1,-nbitq), 
to_sfixed(-1333.0/65536.0,1,-nbitq), 
to_sfixed(-1673.0/65536.0,1,-nbitq), 
to_sfixed(-1230.0/65536.0,1,-nbitq), 
to_sfixed(1165.0/65536.0,1,-nbitq), 
to_sfixed(684.0/65536.0,1,-nbitq), 
to_sfixed(2836.0/65536.0,1,-nbitq), 
to_sfixed(408.0/65536.0,1,-nbitq), 
to_sfixed(-1755.0/65536.0,1,-nbitq), 
to_sfixed(2233.0/65536.0,1,-nbitq), 
to_sfixed(-2554.0/65536.0,1,-nbitq), 
to_sfixed(818.0/65536.0,1,-nbitq), 
to_sfixed(-3073.0/65536.0,1,-nbitq), 
to_sfixed(3692.0/65536.0,1,-nbitq), 
to_sfixed(2578.0/65536.0,1,-nbitq), 
to_sfixed(2834.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-612.0/65536.0,1,-nbitq), 
to_sfixed(-2546.0/65536.0,1,-nbitq), 
to_sfixed(-1823.0/65536.0,1,-nbitq), 
to_sfixed(-1187.0/65536.0,1,-nbitq), 
to_sfixed(-295.0/65536.0,1,-nbitq), 
to_sfixed(-1075.0/65536.0,1,-nbitq), 
to_sfixed(-278.0/65536.0,1,-nbitq), 
to_sfixed(-1366.0/65536.0,1,-nbitq), 
to_sfixed(277.0/65536.0,1,-nbitq), 
to_sfixed(-1498.0/65536.0,1,-nbitq), 
to_sfixed(-3186.0/65536.0,1,-nbitq), 
to_sfixed(-2549.0/65536.0,1,-nbitq), 
to_sfixed(469.0/65536.0,1,-nbitq), 
to_sfixed(-886.0/65536.0,1,-nbitq), 
to_sfixed(1317.0/65536.0,1,-nbitq), 
to_sfixed(2157.0/65536.0,1,-nbitq), 
to_sfixed(-1489.0/65536.0,1,-nbitq), 
to_sfixed(1907.0/65536.0,1,-nbitq), 
to_sfixed(-1402.0/65536.0,1,-nbitq), 
to_sfixed(2035.0/65536.0,1,-nbitq), 
to_sfixed(-4163.0/65536.0,1,-nbitq), 
to_sfixed(-457.0/65536.0,1,-nbitq), 
to_sfixed(-1510.0/65536.0,1,-nbitq), 
to_sfixed(3750.0/65536.0,1,-nbitq), 
to_sfixed(2223.0/65536.0,1,-nbitq), 
to_sfixed(-3259.0/65536.0,1,-nbitq), 
to_sfixed(-1560.0/65536.0,1,-nbitq), 
to_sfixed(1282.0/65536.0,1,-nbitq), 
to_sfixed(-5223.0/65536.0,1,-nbitq), 
to_sfixed(-1360.0/65536.0,1,-nbitq), 
to_sfixed(-2310.0/65536.0,1,-nbitq), 
to_sfixed(-180.0/65536.0,1,-nbitq), 
to_sfixed(-433.0/65536.0,1,-nbitq), 
to_sfixed(-2930.0/65536.0,1,-nbitq), 
to_sfixed(2492.0/65536.0,1,-nbitq), 
to_sfixed(-1494.0/65536.0,1,-nbitq), 
to_sfixed(2079.0/65536.0,1,-nbitq), 
to_sfixed(-3463.0/65536.0,1,-nbitq), 
to_sfixed(-3658.0/65536.0,1,-nbitq), 
to_sfixed(-486.0/65536.0,1,-nbitq), 
to_sfixed(-2057.0/65536.0,1,-nbitq), 
to_sfixed(-2569.0/65536.0,1,-nbitq), 
to_sfixed(-2480.0/65536.0,1,-nbitq), 
to_sfixed(3614.0/65536.0,1,-nbitq), 
to_sfixed(1382.0/65536.0,1,-nbitq), 
to_sfixed(4186.0/65536.0,1,-nbitq), 
to_sfixed(-201.0/65536.0,1,-nbitq), 
to_sfixed(-1133.0/65536.0,1,-nbitq), 
to_sfixed(29.0/65536.0,1,-nbitq), 
to_sfixed(-596.0/65536.0,1,-nbitq), 
to_sfixed(-1744.0/65536.0,1,-nbitq), 
to_sfixed(-2077.0/65536.0,1,-nbitq), 
to_sfixed(2061.0/65536.0,1,-nbitq), 
to_sfixed(1179.0/65536.0,1,-nbitq), 
to_sfixed(834.0/65536.0,1,-nbitq), 
to_sfixed(-675.0/65536.0,1,-nbitq), 
to_sfixed(1667.0/65536.0,1,-nbitq), 
to_sfixed(208.0/65536.0,1,-nbitq), 
to_sfixed(210.0/65536.0,1,-nbitq), 
to_sfixed(887.0/65536.0,1,-nbitq), 
to_sfixed(-2266.0/65536.0,1,-nbitq), 
to_sfixed(-957.0/65536.0,1,-nbitq), 
to_sfixed(-2261.0/65536.0,1,-nbitq), 
to_sfixed(2208.0/65536.0,1,-nbitq), 
to_sfixed(1564.0/65536.0,1,-nbitq), 
to_sfixed(-1522.0/65536.0,1,-nbitq), 
to_sfixed(-494.0/65536.0,1,-nbitq), 
to_sfixed(-1599.0/65536.0,1,-nbitq), 
to_sfixed(608.0/65536.0,1,-nbitq), 
to_sfixed(-91.0/65536.0,1,-nbitq), 
to_sfixed(3112.0/65536.0,1,-nbitq), 
to_sfixed(-1173.0/65536.0,1,-nbitq), 
to_sfixed(3522.0/65536.0,1,-nbitq), 
to_sfixed(1283.0/65536.0,1,-nbitq), 
to_sfixed(49.0/65536.0,1,-nbitq), 
to_sfixed(-103.0/65536.0,1,-nbitq), 
to_sfixed(1659.0/65536.0,1,-nbitq), 
to_sfixed(5282.0/65536.0,1,-nbitq), 
to_sfixed(-1794.0/65536.0,1,-nbitq), 
to_sfixed(2742.0/65536.0,1,-nbitq)  ), 
( to_sfixed(810.0/65536.0,1,-nbitq), 
to_sfixed(-3123.0/65536.0,1,-nbitq), 
to_sfixed(-858.0/65536.0,1,-nbitq), 
to_sfixed(240.0/65536.0,1,-nbitq), 
to_sfixed(1234.0/65536.0,1,-nbitq), 
to_sfixed(-3128.0/65536.0,1,-nbitq), 
to_sfixed(-1996.0/65536.0,1,-nbitq), 
to_sfixed(-1032.0/65536.0,1,-nbitq), 
to_sfixed(2179.0/65536.0,1,-nbitq), 
to_sfixed(-38.0/65536.0,1,-nbitq), 
to_sfixed(-3632.0/65536.0,1,-nbitq), 
to_sfixed(-386.0/65536.0,1,-nbitq), 
to_sfixed(2411.0/65536.0,1,-nbitq), 
to_sfixed(-60.0/65536.0,1,-nbitq), 
to_sfixed(1386.0/65536.0,1,-nbitq), 
to_sfixed(-2633.0/65536.0,1,-nbitq), 
to_sfixed(-404.0/65536.0,1,-nbitq), 
to_sfixed(-6.0/65536.0,1,-nbitq), 
to_sfixed(3159.0/65536.0,1,-nbitq), 
to_sfixed(-22.0/65536.0,1,-nbitq), 
to_sfixed(-4230.0/65536.0,1,-nbitq), 
to_sfixed(1167.0/65536.0,1,-nbitq), 
to_sfixed(-509.0/65536.0,1,-nbitq), 
to_sfixed(53.0/65536.0,1,-nbitq), 
to_sfixed(2920.0/65536.0,1,-nbitq), 
to_sfixed(1417.0/65536.0,1,-nbitq), 
to_sfixed(287.0/65536.0,1,-nbitq), 
to_sfixed(-1614.0/65536.0,1,-nbitq), 
to_sfixed(-1257.0/65536.0,1,-nbitq), 
to_sfixed(155.0/65536.0,1,-nbitq), 
to_sfixed(-2343.0/65536.0,1,-nbitq), 
to_sfixed(3230.0/65536.0,1,-nbitq), 
to_sfixed(-3973.0/65536.0,1,-nbitq), 
to_sfixed(-2961.0/65536.0,1,-nbitq), 
to_sfixed(-1640.0/65536.0,1,-nbitq), 
to_sfixed(-1237.0/65536.0,1,-nbitq), 
to_sfixed(-480.0/65536.0,1,-nbitq), 
to_sfixed(-1897.0/65536.0,1,-nbitq), 
to_sfixed(1024.0/65536.0,1,-nbitq), 
to_sfixed(-273.0/65536.0,1,-nbitq), 
to_sfixed(-287.0/65536.0,1,-nbitq), 
to_sfixed(1547.0/65536.0,1,-nbitq), 
to_sfixed(-4864.0/65536.0,1,-nbitq), 
to_sfixed(-1445.0/65536.0,1,-nbitq), 
to_sfixed(-2293.0/65536.0,1,-nbitq), 
to_sfixed(1669.0/65536.0,1,-nbitq), 
to_sfixed(877.0/65536.0,1,-nbitq), 
to_sfixed(2449.0/65536.0,1,-nbitq), 
to_sfixed(-87.0/65536.0,1,-nbitq), 
to_sfixed(1874.0/65536.0,1,-nbitq), 
to_sfixed(-933.0/65536.0,1,-nbitq), 
to_sfixed(-106.0/65536.0,1,-nbitq), 
to_sfixed(2209.0/65536.0,1,-nbitq), 
to_sfixed(-3277.0/65536.0,1,-nbitq), 
to_sfixed(-1076.0/65536.0,1,-nbitq), 
to_sfixed(-2168.0/65536.0,1,-nbitq), 
to_sfixed(-203.0/65536.0,1,-nbitq), 
to_sfixed(3190.0/65536.0,1,-nbitq), 
to_sfixed(-2546.0/65536.0,1,-nbitq), 
to_sfixed(4563.0/65536.0,1,-nbitq), 
to_sfixed(-348.0/65536.0,1,-nbitq), 
to_sfixed(-283.0/65536.0,1,-nbitq), 
to_sfixed(-59.0/65536.0,1,-nbitq), 
to_sfixed(-166.0/65536.0,1,-nbitq), 
to_sfixed(-789.0/65536.0,1,-nbitq), 
to_sfixed(2562.0/65536.0,1,-nbitq), 
to_sfixed(2576.0/65536.0,1,-nbitq), 
to_sfixed(-831.0/65536.0,1,-nbitq), 
to_sfixed(1169.0/65536.0,1,-nbitq), 
to_sfixed(-1616.0/65536.0,1,-nbitq), 
to_sfixed(1227.0/65536.0,1,-nbitq), 
to_sfixed(4184.0/65536.0,1,-nbitq), 
to_sfixed(3149.0/65536.0,1,-nbitq), 
to_sfixed(-3211.0/65536.0,1,-nbitq), 
to_sfixed(627.0/65536.0,1,-nbitq), 
to_sfixed(-1250.0/65536.0,1,-nbitq), 
to_sfixed(-590.0/65536.0,1,-nbitq), 
to_sfixed(4609.0/65536.0,1,-nbitq), 
to_sfixed(-2977.0/65536.0,1,-nbitq), 
to_sfixed(2804.0/65536.0,1,-nbitq)  ), 
( to_sfixed(739.0/65536.0,1,-nbitq), 
to_sfixed(-3531.0/65536.0,1,-nbitq), 
to_sfixed(-569.0/65536.0,1,-nbitq), 
to_sfixed(-1179.0/65536.0,1,-nbitq), 
to_sfixed(351.0/65536.0,1,-nbitq), 
to_sfixed(-391.0/65536.0,1,-nbitq), 
to_sfixed(770.0/65536.0,1,-nbitq), 
to_sfixed(-196.0/65536.0,1,-nbitq), 
to_sfixed(422.0/65536.0,1,-nbitq), 
to_sfixed(681.0/65536.0,1,-nbitq), 
to_sfixed(-3668.0/65536.0,1,-nbitq), 
to_sfixed(-3196.0/65536.0,1,-nbitq), 
to_sfixed(1772.0/65536.0,1,-nbitq), 
to_sfixed(-3105.0/65536.0,1,-nbitq), 
to_sfixed(-2371.0/65536.0,1,-nbitq), 
to_sfixed(304.0/65536.0,1,-nbitq), 
to_sfixed(-666.0/65536.0,1,-nbitq), 
to_sfixed(2942.0/65536.0,1,-nbitq), 
to_sfixed(1091.0/65536.0,1,-nbitq), 
to_sfixed(3247.0/65536.0,1,-nbitq), 
to_sfixed(-2020.0/65536.0,1,-nbitq), 
to_sfixed(-699.0/65536.0,1,-nbitq), 
to_sfixed(301.0/65536.0,1,-nbitq), 
to_sfixed(4674.0/65536.0,1,-nbitq), 
to_sfixed(4395.0/65536.0,1,-nbitq), 
to_sfixed(2215.0/65536.0,1,-nbitq), 
to_sfixed(-2321.0/65536.0,1,-nbitq), 
to_sfixed(-1537.0/65536.0,1,-nbitq), 
to_sfixed(-3146.0/65536.0,1,-nbitq), 
to_sfixed(-938.0/65536.0,1,-nbitq), 
to_sfixed(710.0/65536.0,1,-nbitq), 
to_sfixed(-179.0/65536.0,1,-nbitq), 
to_sfixed(447.0/65536.0,1,-nbitq), 
to_sfixed(2651.0/65536.0,1,-nbitq), 
to_sfixed(-2777.0/65536.0,1,-nbitq), 
to_sfixed(-1363.0/65536.0,1,-nbitq), 
to_sfixed(1386.0/65536.0,1,-nbitq), 
to_sfixed(-2388.0/65536.0,1,-nbitq), 
to_sfixed(-2790.0/65536.0,1,-nbitq), 
to_sfixed(582.0/65536.0,1,-nbitq), 
to_sfixed(-2573.0/65536.0,1,-nbitq), 
to_sfixed(-1134.0/65536.0,1,-nbitq), 
to_sfixed(-2122.0/65536.0,1,-nbitq), 
to_sfixed(2790.0/65536.0,1,-nbitq), 
to_sfixed(932.0/65536.0,1,-nbitq), 
to_sfixed(3896.0/65536.0,1,-nbitq), 
to_sfixed(-1181.0/65536.0,1,-nbitq), 
to_sfixed(724.0/65536.0,1,-nbitq), 
to_sfixed(180.0/65536.0,1,-nbitq), 
to_sfixed(1168.0/65536.0,1,-nbitq), 
to_sfixed(-124.0/65536.0,1,-nbitq), 
to_sfixed(-132.0/65536.0,1,-nbitq), 
to_sfixed(2018.0/65536.0,1,-nbitq), 
to_sfixed(1334.0/65536.0,1,-nbitq), 
to_sfixed(1866.0/65536.0,1,-nbitq), 
to_sfixed(4503.0/65536.0,1,-nbitq), 
to_sfixed(-2083.0/65536.0,1,-nbitq), 
to_sfixed(-1754.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(4961.0/65536.0,1,-nbitq), 
to_sfixed(1424.0/65536.0,1,-nbitq), 
to_sfixed(-1954.0/65536.0,1,-nbitq), 
to_sfixed(479.0/65536.0,1,-nbitq), 
to_sfixed(308.0/65536.0,1,-nbitq), 
to_sfixed(3054.0/65536.0,1,-nbitq), 
to_sfixed(6126.0/65536.0,1,-nbitq), 
to_sfixed(-2097.0/65536.0,1,-nbitq), 
to_sfixed(-1962.0/65536.0,1,-nbitq), 
to_sfixed(-818.0/65536.0,1,-nbitq), 
to_sfixed(-2164.0/65536.0,1,-nbitq), 
to_sfixed(-2753.0/65536.0,1,-nbitq), 
to_sfixed(987.0/65536.0,1,-nbitq), 
to_sfixed(-796.0/65536.0,1,-nbitq), 
to_sfixed(-3049.0/65536.0,1,-nbitq), 
to_sfixed(659.0/65536.0,1,-nbitq), 
to_sfixed(-167.0/65536.0,1,-nbitq), 
to_sfixed(96.0/65536.0,1,-nbitq), 
to_sfixed(-223.0/65536.0,1,-nbitq), 
to_sfixed(2609.0/65536.0,1,-nbitq), 
to_sfixed(677.0/65536.0,1,-nbitq)  ), 
( to_sfixed(416.0/65536.0,1,-nbitq), 
to_sfixed(-3622.0/65536.0,1,-nbitq), 
to_sfixed(1288.0/65536.0,1,-nbitq), 
to_sfixed(1050.0/65536.0,1,-nbitq), 
to_sfixed(-468.0/65536.0,1,-nbitq), 
to_sfixed(-2246.0/65536.0,1,-nbitq), 
to_sfixed(-3789.0/65536.0,1,-nbitq), 
to_sfixed(2314.0/65536.0,1,-nbitq), 
to_sfixed(1456.0/65536.0,1,-nbitq), 
to_sfixed(1438.0/65536.0,1,-nbitq), 
to_sfixed(1792.0/65536.0,1,-nbitq), 
to_sfixed(3511.0/65536.0,1,-nbitq), 
to_sfixed(-955.0/65536.0,1,-nbitq), 
to_sfixed(3183.0/65536.0,1,-nbitq), 
to_sfixed(2548.0/65536.0,1,-nbitq), 
to_sfixed(3088.0/65536.0,1,-nbitq), 
to_sfixed(-551.0/65536.0,1,-nbitq), 
to_sfixed(1898.0/65536.0,1,-nbitq), 
to_sfixed(2553.0/65536.0,1,-nbitq), 
to_sfixed(-1908.0/65536.0,1,-nbitq), 
to_sfixed(-770.0/65536.0,1,-nbitq), 
to_sfixed(1016.0/65536.0,1,-nbitq), 
to_sfixed(-1960.0/65536.0,1,-nbitq), 
to_sfixed(1277.0/65536.0,1,-nbitq), 
to_sfixed(1407.0/65536.0,1,-nbitq), 
to_sfixed(3983.0/65536.0,1,-nbitq), 
to_sfixed(-395.0/65536.0,1,-nbitq), 
to_sfixed(-2465.0/65536.0,1,-nbitq), 
to_sfixed(-5943.0/65536.0,1,-nbitq), 
to_sfixed(-2994.0/65536.0,1,-nbitq), 
to_sfixed(-3168.0/65536.0,1,-nbitq), 
to_sfixed(2084.0/65536.0,1,-nbitq), 
to_sfixed(-413.0/65536.0,1,-nbitq), 
to_sfixed(6303.0/65536.0,1,-nbitq), 
to_sfixed(1962.0/65536.0,1,-nbitq), 
to_sfixed(2622.0/65536.0,1,-nbitq), 
to_sfixed(840.0/65536.0,1,-nbitq), 
to_sfixed(-2169.0/65536.0,1,-nbitq), 
to_sfixed(1665.0/65536.0,1,-nbitq), 
to_sfixed(-864.0/65536.0,1,-nbitq), 
to_sfixed(-7175.0/65536.0,1,-nbitq), 
to_sfixed(1601.0/65536.0,1,-nbitq), 
to_sfixed(5092.0/65536.0,1,-nbitq), 
to_sfixed(174.0/65536.0,1,-nbitq), 
to_sfixed(-2612.0/65536.0,1,-nbitq), 
to_sfixed(2716.0/65536.0,1,-nbitq), 
to_sfixed(2642.0/65536.0,1,-nbitq), 
to_sfixed(-2546.0/65536.0,1,-nbitq), 
to_sfixed(-355.0/65536.0,1,-nbitq), 
to_sfixed(4413.0/65536.0,1,-nbitq), 
to_sfixed(-1674.0/65536.0,1,-nbitq), 
to_sfixed(-1631.0/65536.0,1,-nbitq), 
to_sfixed(1513.0/65536.0,1,-nbitq), 
to_sfixed(186.0/65536.0,1,-nbitq), 
to_sfixed(-2940.0/65536.0,1,-nbitq), 
to_sfixed(1446.0/65536.0,1,-nbitq), 
to_sfixed(1129.0/65536.0,1,-nbitq), 
to_sfixed(2849.0/65536.0,1,-nbitq), 
to_sfixed(25.0/65536.0,1,-nbitq), 
to_sfixed(1718.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(-1386.0/65536.0,1,-nbitq), 
to_sfixed(-1625.0/65536.0,1,-nbitq), 
to_sfixed(-1606.0/65536.0,1,-nbitq), 
to_sfixed(924.0/65536.0,1,-nbitq), 
to_sfixed(1584.0/65536.0,1,-nbitq), 
to_sfixed(-215.0/65536.0,1,-nbitq), 
to_sfixed(218.0/65536.0,1,-nbitq), 
to_sfixed(-45.0/65536.0,1,-nbitq), 
to_sfixed(-1185.0/65536.0,1,-nbitq), 
to_sfixed(748.0/65536.0,1,-nbitq), 
to_sfixed(1092.0/65536.0,1,-nbitq), 
to_sfixed(1963.0/65536.0,1,-nbitq), 
to_sfixed(-268.0/65536.0,1,-nbitq), 
to_sfixed(-1648.0/65536.0,1,-nbitq), 
to_sfixed(-470.0/65536.0,1,-nbitq), 
to_sfixed(-835.0/65536.0,1,-nbitq), 
to_sfixed(2944.0/65536.0,1,-nbitq), 
to_sfixed(60.0/65536.0,1,-nbitq), 
to_sfixed(-1713.0/65536.0,1,-nbitq)  ), 
( to_sfixed(682.0/65536.0,1,-nbitq), 
to_sfixed(1904.0/65536.0,1,-nbitq), 
to_sfixed(7615.0/65536.0,1,-nbitq), 
to_sfixed(496.0/65536.0,1,-nbitq), 
to_sfixed(2951.0/65536.0,1,-nbitq), 
to_sfixed(396.0/65536.0,1,-nbitq), 
to_sfixed(-1576.0/65536.0,1,-nbitq), 
to_sfixed(582.0/65536.0,1,-nbitq), 
to_sfixed(3507.0/65536.0,1,-nbitq), 
to_sfixed(1818.0/65536.0,1,-nbitq), 
to_sfixed(-1705.0/65536.0,1,-nbitq), 
to_sfixed(13044.0/65536.0,1,-nbitq), 
to_sfixed(631.0/65536.0,1,-nbitq), 
to_sfixed(3867.0/65536.0,1,-nbitq), 
to_sfixed(2690.0/65536.0,1,-nbitq), 
to_sfixed(666.0/65536.0,1,-nbitq), 
to_sfixed(761.0/65536.0,1,-nbitq), 
to_sfixed(-4754.0/65536.0,1,-nbitq), 
to_sfixed(1311.0/65536.0,1,-nbitq), 
to_sfixed(2517.0/65536.0,1,-nbitq), 
to_sfixed(-670.0/65536.0,1,-nbitq), 
to_sfixed(2281.0/65536.0,1,-nbitq), 
to_sfixed(1812.0/65536.0,1,-nbitq), 
to_sfixed(-252.0/65536.0,1,-nbitq), 
to_sfixed(-4390.0/65536.0,1,-nbitq), 
to_sfixed(4898.0/65536.0,1,-nbitq), 
to_sfixed(-3330.0/65536.0,1,-nbitq), 
to_sfixed(1946.0/65536.0,1,-nbitq), 
to_sfixed(-3567.0/65536.0,1,-nbitq), 
to_sfixed(5737.0/65536.0,1,-nbitq), 
to_sfixed(-1314.0/65536.0,1,-nbitq), 
to_sfixed(6132.0/65536.0,1,-nbitq), 
to_sfixed(2244.0/65536.0,1,-nbitq), 
to_sfixed(7715.0/65536.0,1,-nbitq), 
to_sfixed(-1638.0/65536.0,1,-nbitq), 
to_sfixed(-1801.0/65536.0,1,-nbitq), 
to_sfixed(-5220.0/65536.0,1,-nbitq), 
to_sfixed(730.0/65536.0,1,-nbitq), 
to_sfixed(-1749.0/65536.0,1,-nbitq), 
to_sfixed(-1471.0/65536.0,1,-nbitq), 
to_sfixed(-10003.0/65536.0,1,-nbitq), 
to_sfixed(-1060.0/65536.0,1,-nbitq), 
to_sfixed(9997.0/65536.0,1,-nbitq), 
to_sfixed(2186.0/65536.0,1,-nbitq), 
to_sfixed(258.0/65536.0,1,-nbitq), 
to_sfixed(1576.0/65536.0,1,-nbitq), 
to_sfixed(2936.0/65536.0,1,-nbitq), 
to_sfixed(-2726.0/65536.0,1,-nbitq), 
to_sfixed(1401.0/65536.0,1,-nbitq), 
to_sfixed(2385.0/65536.0,1,-nbitq), 
to_sfixed(1526.0/65536.0,1,-nbitq), 
to_sfixed(-4956.0/65536.0,1,-nbitq), 
to_sfixed(1279.0/65536.0,1,-nbitq), 
to_sfixed(9206.0/65536.0,1,-nbitq), 
to_sfixed(-4908.0/65536.0,1,-nbitq), 
to_sfixed(3126.0/65536.0,1,-nbitq), 
to_sfixed(-766.0/65536.0,1,-nbitq), 
to_sfixed(-468.0/65536.0,1,-nbitq), 
to_sfixed(-2401.0/65536.0,1,-nbitq), 
to_sfixed(-2187.0/65536.0,1,-nbitq), 
to_sfixed(2735.0/65536.0,1,-nbitq), 
to_sfixed(-1408.0/65536.0,1,-nbitq), 
to_sfixed(-2556.0/65536.0,1,-nbitq), 
to_sfixed(-1255.0/65536.0,1,-nbitq), 
to_sfixed(3064.0/65536.0,1,-nbitq), 
to_sfixed(307.0/65536.0,1,-nbitq), 
to_sfixed(-5050.0/65536.0,1,-nbitq), 
to_sfixed(-2655.0/65536.0,1,-nbitq), 
to_sfixed(-2806.0/65536.0,1,-nbitq), 
to_sfixed(-1373.0/65536.0,1,-nbitq), 
to_sfixed(709.0/65536.0,1,-nbitq), 
to_sfixed(-1153.0/65536.0,1,-nbitq), 
to_sfixed(1505.0/65536.0,1,-nbitq), 
to_sfixed(-694.0/65536.0,1,-nbitq), 
to_sfixed(-2728.0/65536.0,1,-nbitq), 
to_sfixed(2205.0/65536.0,1,-nbitq), 
to_sfixed(2370.0/65536.0,1,-nbitq), 
to_sfixed(-953.0/65536.0,1,-nbitq), 
to_sfixed(-2533.0/65536.0,1,-nbitq), 
to_sfixed(-2418.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1261.0/65536.0,1,-nbitq), 
to_sfixed(-1870.0/65536.0,1,-nbitq), 
to_sfixed(9579.0/65536.0,1,-nbitq), 
to_sfixed(-376.0/65536.0,1,-nbitq), 
to_sfixed(-2754.0/65536.0,1,-nbitq), 
to_sfixed(795.0/65536.0,1,-nbitq), 
to_sfixed(2347.0/65536.0,1,-nbitq), 
to_sfixed(2519.0/65536.0,1,-nbitq), 
to_sfixed(531.0/65536.0,1,-nbitq), 
to_sfixed(-1405.0/65536.0,1,-nbitq), 
to_sfixed(-1043.0/65536.0,1,-nbitq), 
to_sfixed(12144.0/65536.0,1,-nbitq), 
to_sfixed(-1236.0/65536.0,1,-nbitq), 
to_sfixed(5643.0/65536.0,1,-nbitq), 
to_sfixed(-3429.0/65536.0,1,-nbitq), 
to_sfixed(398.0/65536.0,1,-nbitq), 
to_sfixed(-1217.0/65536.0,1,-nbitq), 
to_sfixed(-7353.0/65536.0,1,-nbitq), 
to_sfixed(5411.0/65536.0,1,-nbitq), 
to_sfixed(-146.0/65536.0,1,-nbitq), 
to_sfixed(-335.0/65536.0,1,-nbitq), 
to_sfixed(2037.0/65536.0,1,-nbitq), 
to_sfixed(-1403.0/65536.0,1,-nbitq), 
to_sfixed(-3640.0/65536.0,1,-nbitq), 
to_sfixed(-1750.0/65536.0,1,-nbitq), 
to_sfixed(5790.0/65536.0,1,-nbitq), 
to_sfixed(-2549.0/65536.0,1,-nbitq), 
to_sfixed(-2458.0/65536.0,1,-nbitq), 
to_sfixed(-4269.0/65536.0,1,-nbitq), 
to_sfixed(7638.0/65536.0,1,-nbitq), 
to_sfixed(2060.0/65536.0,1,-nbitq), 
to_sfixed(7171.0/65536.0,1,-nbitq), 
to_sfixed(2125.0/65536.0,1,-nbitq), 
to_sfixed(2153.0/65536.0,1,-nbitq), 
to_sfixed(-2261.0/65536.0,1,-nbitq), 
to_sfixed(1358.0/65536.0,1,-nbitq), 
to_sfixed(-5314.0/65536.0,1,-nbitq), 
to_sfixed(297.0/65536.0,1,-nbitq), 
to_sfixed(3069.0/65536.0,1,-nbitq), 
to_sfixed(-2600.0/65536.0,1,-nbitq), 
to_sfixed(-10322.0/65536.0,1,-nbitq), 
to_sfixed(1709.0/65536.0,1,-nbitq), 
to_sfixed(11184.0/65536.0,1,-nbitq), 
to_sfixed(-4176.0/65536.0,1,-nbitq), 
to_sfixed(2072.0/65536.0,1,-nbitq), 
to_sfixed(-1022.0/65536.0,1,-nbitq), 
to_sfixed(-1948.0/65536.0,1,-nbitq), 
to_sfixed(-3597.0/65536.0,1,-nbitq), 
to_sfixed(2453.0/65536.0,1,-nbitq), 
to_sfixed(1206.0/65536.0,1,-nbitq), 
to_sfixed(605.0/65536.0,1,-nbitq), 
to_sfixed(-8114.0/65536.0,1,-nbitq), 
to_sfixed(1318.0/65536.0,1,-nbitq), 
to_sfixed(9272.0/65536.0,1,-nbitq), 
to_sfixed(-4476.0/65536.0,1,-nbitq), 
to_sfixed(1014.0/65536.0,1,-nbitq), 
to_sfixed(-1804.0/65536.0,1,-nbitq), 
to_sfixed(3968.0/65536.0,1,-nbitq), 
to_sfixed(-1587.0/65536.0,1,-nbitq), 
to_sfixed(791.0/65536.0,1,-nbitq), 
to_sfixed(1566.0/65536.0,1,-nbitq), 
to_sfixed(-2749.0/65536.0,1,-nbitq), 
to_sfixed(2380.0/65536.0,1,-nbitq), 
to_sfixed(753.0/65536.0,1,-nbitq), 
to_sfixed(1466.0/65536.0,1,-nbitq), 
to_sfixed(-1434.0/65536.0,1,-nbitq), 
to_sfixed(-1751.0/65536.0,1,-nbitq), 
to_sfixed(-4103.0/65536.0,1,-nbitq), 
to_sfixed(-218.0/65536.0,1,-nbitq), 
to_sfixed(-4885.0/65536.0,1,-nbitq), 
to_sfixed(865.0/65536.0,1,-nbitq), 
to_sfixed(5536.0/65536.0,1,-nbitq), 
to_sfixed(-3405.0/65536.0,1,-nbitq), 
to_sfixed(-2181.0/65536.0,1,-nbitq), 
to_sfixed(-326.0/65536.0,1,-nbitq), 
to_sfixed(-2447.0/65536.0,1,-nbitq), 
to_sfixed(5492.0/65536.0,1,-nbitq), 
to_sfixed(-306.0/65536.0,1,-nbitq), 
to_sfixed(827.0/65536.0,1,-nbitq), 
to_sfixed(-336.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-493.0/65536.0,1,-nbitq), 
to_sfixed(-3412.0/65536.0,1,-nbitq), 
to_sfixed(9507.0/65536.0,1,-nbitq), 
to_sfixed(-897.0/65536.0,1,-nbitq), 
to_sfixed(-477.0/65536.0,1,-nbitq), 
to_sfixed(-2256.0/65536.0,1,-nbitq), 
to_sfixed(-712.0/65536.0,1,-nbitq), 
to_sfixed(2352.0/65536.0,1,-nbitq), 
to_sfixed(1345.0/65536.0,1,-nbitq), 
to_sfixed(2589.0/65536.0,1,-nbitq), 
to_sfixed(696.0/65536.0,1,-nbitq), 
to_sfixed(7334.0/65536.0,1,-nbitq), 
to_sfixed(323.0/65536.0,1,-nbitq), 
to_sfixed(4257.0/65536.0,1,-nbitq), 
to_sfixed(55.0/65536.0,1,-nbitq), 
to_sfixed(-1239.0/65536.0,1,-nbitq), 
to_sfixed(-2754.0/65536.0,1,-nbitq), 
to_sfixed(-6759.0/65536.0,1,-nbitq), 
to_sfixed(6400.0/65536.0,1,-nbitq), 
to_sfixed(-1123.0/65536.0,1,-nbitq), 
to_sfixed(-2041.0/65536.0,1,-nbitq), 
to_sfixed(-756.0/65536.0,1,-nbitq), 
to_sfixed(2781.0/65536.0,1,-nbitq), 
to_sfixed(585.0/65536.0,1,-nbitq), 
to_sfixed(1427.0/65536.0,1,-nbitq), 
to_sfixed(3616.0/65536.0,1,-nbitq), 
to_sfixed(-6237.0/65536.0,1,-nbitq), 
to_sfixed(-832.0/65536.0,1,-nbitq), 
to_sfixed(-1676.0/65536.0,1,-nbitq), 
to_sfixed(3786.0/65536.0,1,-nbitq), 
to_sfixed(-1433.0/65536.0,1,-nbitq), 
to_sfixed(6179.0/65536.0,1,-nbitq), 
to_sfixed(965.0/65536.0,1,-nbitq), 
to_sfixed(4736.0/65536.0,1,-nbitq), 
to_sfixed(-287.0/65536.0,1,-nbitq), 
to_sfixed(-1793.0/65536.0,1,-nbitq), 
to_sfixed(-6410.0/65536.0,1,-nbitq), 
to_sfixed(4497.0/65536.0,1,-nbitq), 
to_sfixed(2115.0/65536.0,1,-nbitq), 
to_sfixed(-3118.0/65536.0,1,-nbitq), 
to_sfixed(-8410.0/65536.0,1,-nbitq), 
to_sfixed(1475.0/65536.0,1,-nbitq), 
to_sfixed(10500.0/65536.0,1,-nbitq), 
to_sfixed(-4303.0/65536.0,1,-nbitq), 
to_sfixed(115.0/65536.0,1,-nbitq), 
to_sfixed(-8062.0/65536.0,1,-nbitq), 
to_sfixed(340.0/65536.0,1,-nbitq), 
to_sfixed(2277.0/65536.0,1,-nbitq), 
to_sfixed(-996.0/65536.0,1,-nbitq), 
to_sfixed(677.0/65536.0,1,-nbitq), 
to_sfixed(-2688.0/65536.0,1,-nbitq), 
to_sfixed(-3550.0/65536.0,1,-nbitq), 
to_sfixed(2438.0/65536.0,1,-nbitq), 
to_sfixed(2274.0/65536.0,1,-nbitq), 
to_sfixed(-5927.0/65536.0,1,-nbitq), 
to_sfixed(3422.0/65536.0,1,-nbitq), 
to_sfixed(861.0/65536.0,1,-nbitq), 
to_sfixed(840.0/65536.0,1,-nbitq), 
to_sfixed(-2792.0/65536.0,1,-nbitq), 
to_sfixed(1214.0/65536.0,1,-nbitq), 
to_sfixed(4027.0/65536.0,1,-nbitq), 
to_sfixed(-1667.0/65536.0,1,-nbitq), 
to_sfixed(-1806.0/65536.0,1,-nbitq), 
to_sfixed(1228.0/65536.0,1,-nbitq), 
to_sfixed(3344.0/65536.0,1,-nbitq), 
to_sfixed(7200.0/65536.0,1,-nbitq), 
to_sfixed(-5673.0/65536.0,1,-nbitq), 
to_sfixed(-2975.0/65536.0,1,-nbitq), 
to_sfixed(-2755.0/65536.0,1,-nbitq), 
to_sfixed(-5709.0/65536.0,1,-nbitq), 
to_sfixed(-1579.0/65536.0,1,-nbitq), 
to_sfixed(3014.0/65536.0,1,-nbitq), 
to_sfixed(-3744.0/65536.0,1,-nbitq), 
to_sfixed(648.0/65536.0,1,-nbitq), 
to_sfixed(1293.0/65536.0,1,-nbitq), 
to_sfixed(-2968.0/65536.0,1,-nbitq), 
to_sfixed(4134.0/65536.0,1,-nbitq), 
to_sfixed(2663.0/65536.0,1,-nbitq), 
to_sfixed(2954.0/65536.0,1,-nbitq), 
to_sfixed(4353.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2846.0/65536.0,1,-nbitq), 
to_sfixed(-1787.0/65536.0,1,-nbitq), 
to_sfixed(8354.0/65536.0,1,-nbitq), 
to_sfixed(-4515.0/65536.0,1,-nbitq), 
to_sfixed(-5243.0/65536.0,1,-nbitq), 
to_sfixed(-5053.0/65536.0,1,-nbitq), 
to_sfixed(2612.0/65536.0,1,-nbitq), 
to_sfixed(-1365.0/65536.0,1,-nbitq), 
to_sfixed(1782.0/65536.0,1,-nbitq), 
to_sfixed(2357.0/65536.0,1,-nbitq), 
to_sfixed(3954.0/65536.0,1,-nbitq), 
to_sfixed(-2981.0/65536.0,1,-nbitq), 
to_sfixed(-340.0/65536.0,1,-nbitq), 
to_sfixed(1826.0/65536.0,1,-nbitq), 
to_sfixed(337.0/65536.0,1,-nbitq), 
to_sfixed(-2771.0/65536.0,1,-nbitq), 
to_sfixed(-243.0/65536.0,1,-nbitq), 
to_sfixed(-272.0/65536.0,1,-nbitq), 
to_sfixed(635.0/65536.0,1,-nbitq), 
to_sfixed(2001.0/65536.0,1,-nbitq), 
to_sfixed(1996.0/65536.0,1,-nbitq), 
to_sfixed(725.0/65536.0,1,-nbitq), 
to_sfixed(694.0/65536.0,1,-nbitq), 
to_sfixed(-2317.0/65536.0,1,-nbitq), 
to_sfixed(2893.0/65536.0,1,-nbitq), 
to_sfixed(-936.0/65536.0,1,-nbitq), 
to_sfixed(-6826.0/65536.0,1,-nbitq), 
to_sfixed(1249.0/65536.0,1,-nbitq), 
to_sfixed(-7189.0/65536.0,1,-nbitq), 
to_sfixed(-389.0/65536.0,1,-nbitq), 
to_sfixed(-474.0/65536.0,1,-nbitq), 
to_sfixed(7983.0/65536.0,1,-nbitq), 
to_sfixed(1145.0/65536.0,1,-nbitq), 
to_sfixed(7366.0/65536.0,1,-nbitq), 
to_sfixed(-2958.0/65536.0,1,-nbitq), 
to_sfixed(3259.0/65536.0,1,-nbitq), 
to_sfixed(3865.0/65536.0,1,-nbitq), 
to_sfixed(969.0/65536.0,1,-nbitq), 
to_sfixed(-423.0/65536.0,1,-nbitq), 
to_sfixed(3879.0/65536.0,1,-nbitq), 
to_sfixed(-6313.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(10019.0/65536.0,1,-nbitq), 
to_sfixed(-3697.0/65536.0,1,-nbitq), 
to_sfixed(2958.0/65536.0,1,-nbitq), 
to_sfixed(-16912.0/65536.0,1,-nbitq), 
to_sfixed(3173.0/65536.0,1,-nbitq), 
to_sfixed(1989.0/65536.0,1,-nbitq), 
to_sfixed(1281.0/65536.0,1,-nbitq), 
to_sfixed(2267.0/65536.0,1,-nbitq), 
to_sfixed(-1130.0/65536.0,1,-nbitq), 
to_sfixed(-5695.0/65536.0,1,-nbitq), 
to_sfixed(-2548.0/65536.0,1,-nbitq), 
to_sfixed(-2187.0/65536.0,1,-nbitq), 
to_sfixed(-3890.0/65536.0,1,-nbitq), 
to_sfixed(4144.0/65536.0,1,-nbitq), 
to_sfixed(-1106.0/65536.0,1,-nbitq), 
to_sfixed(484.0/65536.0,1,-nbitq), 
to_sfixed(-3377.0/65536.0,1,-nbitq), 
to_sfixed(-3755.0/65536.0,1,-nbitq), 
to_sfixed(2253.0/65536.0,1,-nbitq), 
to_sfixed(-732.0/65536.0,1,-nbitq), 
to_sfixed(153.0/65536.0,1,-nbitq), 
to_sfixed(-2664.0/65536.0,1,-nbitq), 
to_sfixed(387.0/65536.0,1,-nbitq), 
to_sfixed(4780.0/65536.0,1,-nbitq), 
to_sfixed(-5198.0/65536.0,1,-nbitq), 
to_sfixed(-6317.0/65536.0,1,-nbitq), 
to_sfixed(-108.0/65536.0,1,-nbitq), 
to_sfixed(-2178.0/65536.0,1,-nbitq), 
to_sfixed(-1468.0/65536.0,1,-nbitq), 
to_sfixed(7528.0/65536.0,1,-nbitq), 
to_sfixed(-1943.0/65536.0,1,-nbitq), 
to_sfixed(-2562.0/65536.0,1,-nbitq), 
to_sfixed(1312.0/65536.0,1,-nbitq), 
to_sfixed(3274.0/65536.0,1,-nbitq), 
to_sfixed(4925.0/65536.0,1,-nbitq), 
to_sfixed(-963.0/65536.0,1,-nbitq), 
to_sfixed(638.0/65536.0,1,-nbitq), 
to_sfixed(-2445.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4301.0/65536.0,1,-nbitq), 
to_sfixed(-132.0/65536.0,1,-nbitq), 
to_sfixed(3468.0/65536.0,1,-nbitq), 
to_sfixed(-2288.0/65536.0,1,-nbitq), 
to_sfixed(-354.0/65536.0,1,-nbitq), 
to_sfixed(-7236.0/65536.0,1,-nbitq), 
to_sfixed(4274.0/65536.0,1,-nbitq), 
to_sfixed(-885.0/65536.0,1,-nbitq), 
to_sfixed(-2592.0/65536.0,1,-nbitq), 
to_sfixed(-2700.0/65536.0,1,-nbitq), 
to_sfixed(7034.0/65536.0,1,-nbitq), 
to_sfixed(11706.0/65536.0,1,-nbitq), 
to_sfixed(-927.0/65536.0,1,-nbitq), 
to_sfixed(1576.0/65536.0,1,-nbitq), 
to_sfixed(3273.0/65536.0,1,-nbitq), 
to_sfixed(1217.0/65536.0,1,-nbitq), 
to_sfixed(647.0/65536.0,1,-nbitq), 
to_sfixed(-3216.0/65536.0,1,-nbitq), 
to_sfixed(3248.0/65536.0,1,-nbitq), 
to_sfixed(218.0/65536.0,1,-nbitq), 
to_sfixed(-1041.0/65536.0,1,-nbitq), 
to_sfixed(-427.0/65536.0,1,-nbitq), 
to_sfixed(583.0/65536.0,1,-nbitq), 
to_sfixed(2269.0/65536.0,1,-nbitq), 
to_sfixed(-1466.0/65536.0,1,-nbitq), 
to_sfixed(167.0/65536.0,1,-nbitq), 
to_sfixed(-7328.0/65536.0,1,-nbitq), 
to_sfixed(1521.0/65536.0,1,-nbitq), 
to_sfixed(-9928.0/65536.0,1,-nbitq), 
to_sfixed(4689.0/65536.0,1,-nbitq), 
to_sfixed(-590.0/65536.0,1,-nbitq), 
to_sfixed(8670.0/65536.0,1,-nbitq), 
to_sfixed(295.0/65536.0,1,-nbitq), 
to_sfixed(5361.0/65536.0,1,-nbitq), 
to_sfixed(-208.0/65536.0,1,-nbitq), 
to_sfixed(3239.0/65536.0,1,-nbitq), 
to_sfixed(6464.0/65536.0,1,-nbitq), 
to_sfixed(-8239.0/65536.0,1,-nbitq), 
to_sfixed(-7847.0/65536.0,1,-nbitq), 
to_sfixed(-553.0/65536.0,1,-nbitq), 
to_sfixed(-2269.0/65536.0,1,-nbitq), 
to_sfixed(1147.0/65536.0,1,-nbitq), 
to_sfixed(9768.0/65536.0,1,-nbitq), 
to_sfixed(-3506.0/65536.0,1,-nbitq), 
to_sfixed(2366.0/65536.0,1,-nbitq), 
to_sfixed(-17322.0/65536.0,1,-nbitq), 
to_sfixed(-2521.0/65536.0,1,-nbitq), 
to_sfixed(1771.0/65536.0,1,-nbitq), 
to_sfixed(-2461.0/65536.0,1,-nbitq), 
to_sfixed(1671.0/65536.0,1,-nbitq), 
to_sfixed(1360.0/65536.0,1,-nbitq), 
to_sfixed(-4601.0/65536.0,1,-nbitq), 
to_sfixed(3965.0/65536.0,1,-nbitq), 
to_sfixed(851.0/65536.0,1,-nbitq), 
to_sfixed(-3090.0/65536.0,1,-nbitq), 
to_sfixed(7936.0/65536.0,1,-nbitq), 
to_sfixed(-1282.0/65536.0,1,-nbitq), 
to_sfixed(-1741.0/65536.0,1,-nbitq), 
to_sfixed(-1851.0/65536.0,1,-nbitq), 
to_sfixed(-1565.0/65536.0,1,-nbitq), 
to_sfixed(5197.0/65536.0,1,-nbitq), 
to_sfixed(-1723.0/65536.0,1,-nbitq), 
to_sfixed(-2577.0/65536.0,1,-nbitq), 
to_sfixed(645.0/65536.0,1,-nbitq), 
to_sfixed(1961.0/65536.0,1,-nbitq), 
to_sfixed(2571.0/65536.0,1,-nbitq), 
to_sfixed(-3573.0/65536.0,1,-nbitq), 
to_sfixed(-6198.0/65536.0,1,-nbitq), 
to_sfixed(-2959.0/65536.0,1,-nbitq), 
to_sfixed(4084.0/65536.0,1,-nbitq), 
to_sfixed(216.0/65536.0,1,-nbitq), 
to_sfixed(5678.0/65536.0,1,-nbitq), 
to_sfixed(-2804.0/65536.0,1,-nbitq), 
to_sfixed(2601.0/65536.0,1,-nbitq), 
to_sfixed(2580.0/65536.0,1,-nbitq), 
to_sfixed(4307.0/65536.0,1,-nbitq), 
to_sfixed(-419.0/65536.0,1,-nbitq), 
to_sfixed(-6681.0/65536.0,1,-nbitq), 
to_sfixed(4.0/65536.0,1,-nbitq), 
to_sfixed(-4409.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-485.0/65536.0,1,-nbitq), 
to_sfixed(-1168.0/65536.0,1,-nbitq), 
to_sfixed(-5135.0/65536.0,1,-nbitq), 
to_sfixed(164.0/65536.0,1,-nbitq), 
to_sfixed(4746.0/65536.0,1,-nbitq), 
to_sfixed(-2062.0/65536.0,1,-nbitq), 
to_sfixed(2095.0/65536.0,1,-nbitq), 
to_sfixed(-4144.0/65536.0,1,-nbitq), 
to_sfixed(-6313.0/65536.0,1,-nbitq), 
to_sfixed(-1177.0/65536.0,1,-nbitq), 
to_sfixed(5510.0/65536.0,1,-nbitq), 
to_sfixed(11476.0/65536.0,1,-nbitq), 
to_sfixed(2757.0/65536.0,1,-nbitq), 
to_sfixed(-1055.0/65536.0,1,-nbitq), 
to_sfixed(8674.0/65536.0,1,-nbitq), 
to_sfixed(-2743.0/65536.0,1,-nbitq), 
to_sfixed(-2236.0/65536.0,1,-nbitq), 
to_sfixed(2339.0/65536.0,1,-nbitq), 
to_sfixed(6818.0/65536.0,1,-nbitq), 
to_sfixed(693.0/65536.0,1,-nbitq), 
to_sfixed(-2792.0/65536.0,1,-nbitq), 
to_sfixed(-5519.0/65536.0,1,-nbitq), 
to_sfixed(7341.0/65536.0,1,-nbitq), 
to_sfixed(-761.0/65536.0,1,-nbitq), 
to_sfixed(-1047.0/65536.0,1,-nbitq), 
to_sfixed(1036.0/65536.0,1,-nbitq), 
to_sfixed(-6097.0/65536.0,1,-nbitq), 
to_sfixed(2081.0/65536.0,1,-nbitq), 
to_sfixed(-18995.0/65536.0,1,-nbitq), 
to_sfixed(8654.0/65536.0,1,-nbitq), 
to_sfixed(777.0/65536.0,1,-nbitq), 
to_sfixed(10424.0/65536.0,1,-nbitq), 
to_sfixed(3093.0/65536.0,1,-nbitq), 
to_sfixed(-1815.0/65536.0,1,-nbitq), 
to_sfixed(-1317.0/65536.0,1,-nbitq), 
to_sfixed(343.0/65536.0,1,-nbitq), 
to_sfixed(8953.0/65536.0,1,-nbitq), 
to_sfixed(-10712.0/65536.0,1,-nbitq), 
to_sfixed(-6263.0/65536.0,1,-nbitq), 
to_sfixed(2150.0/65536.0,1,-nbitq), 
to_sfixed(-3671.0/65536.0,1,-nbitq), 
to_sfixed(2669.0/65536.0,1,-nbitq), 
to_sfixed(4060.0/65536.0,1,-nbitq), 
to_sfixed(-6898.0/65536.0,1,-nbitq), 
to_sfixed(-1198.0/65536.0,1,-nbitq), 
to_sfixed(-6014.0/65536.0,1,-nbitq), 
to_sfixed(178.0/65536.0,1,-nbitq), 
to_sfixed(-3336.0/65536.0,1,-nbitq), 
to_sfixed(-41.0/65536.0,1,-nbitq), 
to_sfixed(-2296.0/65536.0,1,-nbitq), 
to_sfixed(2271.0/65536.0,1,-nbitq), 
to_sfixed(-7255.0/65536.0,1,-nbitq), 
to_sfixed(3965.0/65536.0,1,-nbitq), 
to_sfixed(-4781.0/65536.0,1,-nbitq), 
to_sfixed(-8063.0/65536.0,1,-nbitq), 
to_sfixed(4912.0/65536.0,1,-nbitq), 
to_sfixed(1660.0/65536.0,1,-nbitq), 
to_sfixed(1982.0/65536.0,1,-nbitq), 
to_sfixed(-808.0/65536.0,1,-nbitq), 
to_sfixed(-3580.0/65536.0,1,-nbitq), 
to_sfixed(3815.0/65536.0,1,-nbitq), 
to_sfixed(2244.0/65536.0,1,-nbitq), 
to_sfixed(2380.0/65536.0,1,-nbitq), 
to_sfixed(1568.0/65536.0,1,-nbitq), 
to_sfixed(-4874.0/65536.0,1,-nbitq), 
to_sfixed(5556.0/65536.0,1,-nbitq), 
to_sfixed(-5612.0/65536.0,1,-nbitq), 
to_sfixed(-3555.0/65536.0,1,-nbitq), 
to_sfixed(-944.0/65536.0,1,-nbitq), 
to_sfixed(-1322.0/65536.0,1,-nbitq), 
to_sfixed(-230.0/65536.0,1,-nbitq), 
to_sfixed(2981.0/65536.0,1,-nbitq), 
to_sfixed(-5772.0/65536.0,1,-nbitq), 
to_sfixed(-2935.0/65536.0,1,-nbitq), 
to_sfixed(1891.0/65536.0,1,-nbitq), 
to_sfixed(-2805.0/65536.0,1,-nbitq), 
to_sfixed(-785.0/65536.0,1,-nbitq), 
to_sfixed(-17663.0/65536.0,1,-nbitq), 
to_sfixed(-320.0/65536.0,1,-nbitq), 
to_sfixed(-5612.0/65536.0,1,-nbitq)  ), 
( to_sfixed(80.0/65536.0,1,-nbitq), 
to_sfixed(-3817.0/65536.0,1,-nbitq), 
to_sfixed(-12696.0/65536.0,1,-nbitq), 
to_sfixed(-2176.0/65536.0,1,-nbitq), 
to_sfixed(16590.0/65536.0,1,-nbitq), 
to_sfixed(-8327.0/65536.0,1,-nbitq), 
to_sfixed(5676.0/65536.0,1,-nbitq), 
to_sfixed(-8084.0/65536.0,1,-nbitq), 
to_sfixed(-4040.0/65536.0,1,-nbitq), 
to_sfixed(-2632.0/65536.0,1,-nbitq), 
to_sfixed(6522.0/65536.0,1,-nbitq), 
to_sfixed(-1128.0/65536.0,1,-nbitq), 
to_sfixed(2907.0/65536.0,1,-nbitq), 
to_sfixed(2251.0/65536.0,1,-nbitq), 
to_sfixed(2779.0/65536.0,1,-nbitq), 
to_sfixed(835.0/65536.0,1,-nbitq), 
to_sfixed(-1196.0/65536.0,1,-nbitq), 
to_sfixed(9492.0/65536.0,1,-nbitq), 
to_sfixed(7329.0/65536.0,1,-nbitq), 
to_sfixed(1883.0/65536.0,1,-nbitq), 
to_sfixed(-260.0/65536.0,1,-nbitq), 
to_sfixed(1251.0/65536.0,1,-nbitq), 
to_sfixed(14362.0/65536.0,1,-nbitq), 
to_sfixed(-5306.0/65536.0,1,-nbitq), 
to_sfixed(562.0/65536.0,1,-nbitq), 
to_sfixed(-6420.0/65536.0,1,-nbitq), 
to_sfixed(-7347.0/65536.0,1,-nbitq), 
to_sfixed(1013.0/65536.0,1,-nbitq), 
to_sfixed(-13965.0/65536.0,1,-nbitq), 
to_sfixed(4951.0/65536.0,1,-nbitq), 
to_sfixed(2925.0/65536.0,1,-nbitq), 
to_sfixed(4289.0/65536.0,1,-nbitq), 
to_sfixed(1706.0/65536.0,1,-nbitq), 
to_sfixed(175.0/65536.0,1,-nbitq), 
to_sfixed(-109.0/65536.0,1,-nbitq), 
to_sfixed(-908.0/65536.0,1,-nbitq), 
to_sfixed(12358.0/65536.0,1,-nbitq), 
to_sfixed(-9896.0/65536.0,1,-nbitq), 
to_sfixed(-3492.0/65536.0,1,-nbitq), 
to_sfixed(-305.0/65536.0,1,-nbitq), 
to_sfixed(-9157.0/65536.0,1,-nbitq), 
to_sfixed(-1612.0/65536.0,1,-nbitq), 
to_sfixed(-5508.0/65536.0,1,-nbitq), 
to_sfixed(-5299.0/65536.0,1,-nbitq), 
to_sfixed(2252.0/65536.0,1,-nbitq), 
to_sfixed(410.0/65536.0,1,-nbitq), 
to_sfixed(-3265.0/65536.0,1,-nbitq), 
to_sfixed(-2401.0/65536.0,1,-nbitq), 
to_sfixed(707.0/65536.0,1,-nbitq), 
to_sfixed(-4813.0/65536.0,1,-nbitq), 
to_sfixed(183.0/65536.0,1,-nbitq), 
to_sfixed(-7382.0/65536.0,1,-nbitq), 
to_sfixed(1416.0/65536.0,1,-nbitq), 
to_sfixed(-1713.0/65536.0,1,-nbitq), 
to_sfixed(-4324.0/65536.0,1,-nbitq), 
to_sfixed(2441.0/65536.0,1,-nbitq), 
to_sfixed(88.0/65536.0,1,-nbitq), 
to_sfixed(280.0/65536.0,1,-nbitq), 
to_sfixed(-123.0/65536.0,1,-nbitq), 
to_sfixed(-9051.0/65536.0,1,-nbitq), 
to_sfixed(6603.0/65536.0,1,-nbitq), 
to_sfixed(2733.0/65536.0,1,-nbitq), 
to_sfixed(-2151.0/65536.0,1,-nbitq), 
to_sfixed(1247.0/65536.0,1,-nbitq), 
to_sfixed(-5807.0/65536.0,1,-nbitq), 
to_sfixed(-4289.0/65536.0,1,-nbitq), 
to_sfixed(811.0/65536.0,1,-nbitq), 
to_sfixed(-1805.0/65536.0,1,-nbitq), 
to_sfixed(-3174.0/65536.0,1,-nbitq), 
to_sfixed(8265.0/65536.0,1,-nbitq), 
to_sfixed(501.0/65536.0,1,-nbitq), 
to_sfixed(2242.0/65536.0,1,-nbitq), 
to_sfixed(-290.0/65536.0,1,-nbitq), 
to_sfixed(-1393.0/65536.0,1,-nbitq), 
to_sfixed(2449.0/65536.0,1,-nbitq), 
to_sfixed(-6435.0/65536.0,1,-nbitq), 
to_sfixed(-1563.0/65536.0,1,-nbitq), 
to_sfixed(-10069.0/65536.0,1,-nbitq), 
to_sfixed(972.0/65536.0,1,-nbitq), 
to_sfixed(-7839.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3933.0/65536.0,1,-nbitq), 
to_sfixed(-1671.0/65536.0,1,-nbitq), 
to_sfixed(-13857.0/65536.0,1,-nbitq), 
to_sfixed(1310.0/65536.0,1,-nbitq), 
to_sfixed(9376.0/65536.0,1,-nbitq), 
to_sfixed(-8599.0/65536.0,1,-nbitq), 
to_sfixed(1036.0/65536.0,1,-nbitq), 
to_sfixed(-2164.0/65536.0,1,-nbitq), 
to_sfixed(-4102.0/65536.0,1,-nbitq), 
to_sfixed(1228.0/65536.0,1,-nbitq), 
to_sfixed(8212.0/65536.0,1,-nbitq), 
to_sfixed(2649.0/65536.0,1,-nbitq), 
to_sfixed(3772.0/65536.0,1,-nbitq), 
to_sfixed(2909.0/65536.0,1,-nbitq), 
to_sfixed(-4158.0/65536.0,1,-nbitq), 
to_sfixed(50.0/65536.0,1,-nbitq), 
to_sfixed(-2872.0/65536.0,1,-nbitq), 
to_sfixed(1703.0/65536.0,1,-nbitq), 
to_sfixed(85.0/65536.0,1,-nbitq), 
to_sfixed(642.0/65536.0,1,-nbitq), 
to_sfixed(-1891.0/65536.0,1,-nbitq), 
to_sfixed(-2742.0/65536.0,1,-nbitq), 
to_sfixed(17729.0/65536.0,1,-nbitq), 
to_sfixed(-1429.0/65536.0,1,-nbitq), 
to_sfixed(1237.0/65536.0,1,-nbitq), 
to_sfixed(150.0/65536.0,1,-nbitq), 
to_sfixed(-8296.0/65536.0,1,-nbitq), 
to_sfixed(-2027.0/65536.0,1,-nbitq), 
to_sfixed(259.0/65536.0,1,-nbitq), 
to_sfixed(4774.0/65536.0,1,-nbitq), 
to_sfixed(772.0/65536.0,1,-nbitq), 
to_sfixed(3637.0/65536.0,1,-nbitq), 
to_sfixed(-87.0/65536.0,1,-nbitq), 
to_sfixed(-4915.0/65536.0,1,-nbitq), 
to_sfixed(2854.0/65536.0,1,-nbitq), 
to_sfixed(1828.0/65536.0,1,-nbitq), 
to_sfixed(12216.0/65536.0,1,-nbitq), 
to_sfixed(-6447.0/65536.0,1,-nbitq), 
to_sfixed(-7630.0/65536.0,1,-nbitq), 
to_sfixed(6.0/65536.0,1,-nbitq), 
to_sfixed(-6599.0/65536.0,1,-nbitq), 
to_sfixed(-884.0/65536.0,1,-nbitq), 
to_sfixed(-767.0/65536.0,1,-nbitq), 
to_sfixed(-7925.0/65536.0,1,-nbitq), 
to_sfixed(-1247.0/65536.0,1,-nbitq), 
to_sfixed(3364.0/65536.0,1,-nbitq), 
to_sfixed(224.0/65536.0,1,-nbitq), 
to_sfixed(3644.0/65536.0,1,-nbitq), 
to_sfixed(-59.0/65536.0,1,-nbitq), 
to_sfixed(21.0/65536.0,1,-nbitq), 
to_sfixed(-1253.0/65536.0,1,-nbitq), 
to_sfixed(-11035.0/65536.0,1,-nbitq), 
to_sfixed(-1698.0/65536.0,1,-nbitq), 
to_sfixed(-4119.0/65536.0,1,-nbitq), 
to_sfixed(-7004.0/65536.0,1,-nbitq), 
to_sfixed(-1544.0/65536.0,1,-nbitq), 
to_sfixed(-3307.0/65536.0,1,-nbitq), 
to_sfixed(-4216.0/65536.0,1,-nbitq), 
to_sfixed(609.0/65536.0,1,-nbitq), 
to_sfixed(-7252.0/65536.0,1,-nbitq), 
to_sfixed(10657.0/65536.0,1,-nbitq), 
to_sfixed(1455.0/65536.0,1,-nbitq), 
to_sfixed(2089.0/65536.0,1,-nbitq), 
to_sfixed(-849.0/65536.0,1,-nbitq), 
to_sfixed(-7385.0/65536.0,1,-nbitq), 
to_sfixed(-10528.0/65536.0,1,-nbitq), 
to_sfixed(-1974.0/65536.0,1,-nbitq), 
to_sfixed(7225.0/65536.0,1,-nbitq), 
to_sfixed(-717.0/65536.0,1,-nbitq), 
to_sfixed(1808.0/65536.0,1,-nbitq), 
to_sfixed(3416.0/65536.0,1,-nbitq), 
to_sfixed(-1931.0/65536.0,1,-nbitq), 
to_sfixed(-1069.0/65536.0,1,-nbitq), 
to_sfixed(-1644.0/65536.0,1,-nbitq), 
to_sfixed(1488.0/65536.0,1,-nbitq), 
to_sfixed(-7678.0/65536.0,1,-nbitq), 
to_sfixed(-2777.0/65536.0,1,-nbitq), 
to_sfixed(917.0/65536.0,1,-nbitq), 
to_sfixed(1647.0/65536.0,1,-nbitq), 
to_sfixed(-3277.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2383.0/65536.0,1,-nbitq), 
to_sfixed(-1425.0/65536.0,1,-nbitq), 
to_sfixed(-13879.0/65536.0,1,-nbitq), 
to_sfixed(-6632.0/65536.0,1,-nbitq), 
to_sfixed(-4745.0/65536.0,1,-nbitq), 
to_sfixed(-14063.0/65536.0,1,-nbitq), 
to_sfixed(3909.0/65536.0,1,-nbitq), 
to_sfixed(6050.0/65536.0,1,-nbitq), 
to_sfixed(2296.0/65536.0,1,-nbitq), 
to_sfixed(2127.0/65536.0,1,-nbitq), 
to_sfixed(5293.0/65536.0,1,-nbitq), 
to_sfixed(-4664.0/65536.0,1,-nbitq), 
to_sfixed(-845.0/65536.0,1,-nbitq), 
to_sfixed(-179.0/65536.0,1,-nbitq), 
to_sfixed(-7542.0/65536.0,1,-nbitq), 
to_sfixed(2416.0/65536.0,1,-nbitq), 
to_sfixed(1428.0/65536.0,1,-nbitq), 
to_sfixed(-5323.0/65536.0,1,-nbitq), 
to_sfixed(1380.0/65536.0,1,-nbitq), 
to_sfixed(-1200.0/65536.0,1,-nbitq), 
to_sfixed(-3553.0/65536.0,1,-nbitq), 
to_sfixed(340.0/65536.0,1,-nbitq), 
to_sfixed(11556.0/65536.0,1,-nbitq), 
to_sfixed(1354.0/65536.0,1,-nbitq), 
to_sfixed(-4991.0/65536.0,1,-nbitq), 
to_sfixed(1319.0/65536.0,1,-nbitq), 
to_sfixed(-10126.0/65536.0,1,-nbitq), 
to_sfixed(-2099.0/65536.0,1,-nbitq), 
to_sfixed(1528.0/65536.0,1,-nbitq), 
to_sfixed(2470.0/65536.0,1,-nbitq), 
to_sfixed(1942.0/65536.0,1,-nbitq), 
to_sfixed(10016.0/65536.0,1,-nbitq), 
to_sfixed(-2557.0/65536.0,1,-nbitq), 
to_sfixed(-7394.0/65536.0,1,-nbitq), 
to_sfixed(1932.0/65536.0,1,-nbitq), 
to_sfixed(-588.0/65536.0,1,-nbitq), 
to_sfixed(4432.0/65536.0,1,-nbitq), 
to_sfixed(-4436.0/65536.0,1,-nbitq), 
to_sfixed(-5479.0/65536.0,1,-nbitq), 
to_sfixed(-2307.0/65536.0,1,-nbitq), 
to_sfixed(-6012.0/65536.0,1,-nbitq), 
to_sfixed(-608.0/65536.0,1,-nbitq), 
to_sfixed(-2252.0/65536.0,1,-nbitq), 
to_sfixed(-1954.0/65536.0,1,-nbitq), 
to_sfixed(1473.0/65536.0,1,-nbitq), 
to_sfixed(-564.0/65536.0,1,-nbitq), 
to_sfixed(536.0/65536.0,1,-nbitq), 
to_sfixed(7900.0/65536.0,1,-nbitq), 
to_sfixed(-2157.0/65536.0,1,-nbitq), 
to_sfixed(-3253.0/65536.0,1,-nbitq), 
to_sfixed(2489.0/65536.0,1,-nbitq), 
to_sfixed(-13733.0/65536.0,1,-nbitq), 
to_sfixed(138.0/65536.0,1,-nbitq), 
to_sfixed(940.0/65536.0,1,-nbitq), 
to_sfixed(-4293.0/65536.0,1,-nbitq), 
to_sfixed(-2561.0/65536.0,1,-nbitq), 
to_sfixed(2115.0/65536.0,1,-nbitq), 
to_sfixed(567.0/65536.0,1,-nbitq), 
to_sfixed(-3624.0/65536.0,1,-nbitq), 
to_sfixed(85.0/65536.0,1,-nbitq), 
to_sfixed(6359.0/65536.0,1,-nbitq), 
to_sfixed(2509.0/65536.0,1,-nbitq), 
to_sfixed(-146.0/65536.0,1,-nbitq), 
to_sfixed(-583.0/65536.0,1,-nbitq), 
to_sfixed(1189.0/65536.0,1,-nbitq), 
to_sfixed(-6248.0/65536.0,1,-nbitq), 
to_sfixed(-6373.0/65536.0,1,-nbitq), 
to_sfixed(9120.0/65536.0,1,-nbitq), 
to_sfixed(344.0/65536.0,1,-nbitq), 
to_sfixed(-2901.0/65536.0,1,-nbitq), 
to_sfixed(-1747.0/65536.0,1,-nbitq), 
to_sfixed(2710.0/65536.0,1,-nbitq), 
to_sfixed(-6861.0/65536.0,1,-nbitq), 
to_sfixed(-2526.0/65536.0,1,-nbitq), 
to_sfixed(-1858.0/65536.0,1,-nbitq), 
to_sfixed(-4267.0/65536.0,1,-nbitq), 
to_sfixed(1785.0/65536.0,1,-nbitq), 
to_sfixed(5171.0/65536.0,1,-nbitq), 
to_sfixed(1483.0/65536.0,1,-nbitq), 
to_sfixed(-432.0/65536.0,1,-nbitq)  ), 
( to_sfixed(284.0/65536.0,1,-nbitq), 
to_sfixed(5470.0/65536.0,1,-nbitq), 
to_sfixed(225.0/65536.0,1,-nbitq), 
to_sfixed(-7818.0/65536.0,1,-nbitq), 
to_sfixed(-1252.0/65536.0,1,-nbitq), 
to_sfixed(-2225.0/65536.0,1,-nbitq), 
to_sfixed(-1263.0/65536.0,1,-nbitq), 
to_sfixed(1353.0/65536.0,1,-nbitq), 
to_sfixed(8094.0/65536.0,1,-nbitq), 
to_sfixed(-2628.0/65536.0,1,-nbitq), 
to_sfixed(-1202.0/65536.0,1,-nbitq), 
to_sfixed(-5165.0/65536.0,1,-nbitq), 
to_sfixed(380.0/65536.0,1,-nbitq), 
to_sfixed(445.0/65536.0,1,-nbitq), 
to_sfixed(-5637.0/65536.0,1,-nbitq), 
to_sfixed(1141.0/65536.0,1,-nbitq), 
to_sfixed(1081.0/65536.0,1,-nbitq), 
to_sfixed(-4634.0/65536.0,1,-nbitq), 
to_sfixed(5171.0/65536.0,1,-nbitq), 
to_sfixed(-2221.0/65536.0,1,-nbitq), 
to_sfixed(1978.0/65536.0,1,-nbitq), 
to_sfixed(-1010.0/65536.0,1,-nbitq), 
to_sfixed(-1336.0/65536.0,1,-nbitq), 
to_sfixed(-2597.0/65536.0,1,-nbitq), 
to_sfixed(-5585.0/65536.0,1,-nbitq), 
to_sfixed(2574.0/65536.0,1,-nbitq), 
to_sfixed(-3990.0/65536.0,1,-nbitq), 
to_sfixed(3899.0/65536.0,1,-nbitq), 
to_sfixed(4894.0/65536.0,1,-nbitq), 
to_sfixed(-3244.0/65536.0,1,-nbitq), 
to_sfixed(-391.0/65536.0,1,-nbitq), 
to_sfixed(-386.0/65536.0,1,-nbitq), 
to_sfixed(-3687.0/65536.0,1,-nbitq), 
to_sfixed(-2255.0/65536.0,1,-nbitq), 
to_sfixed(-511.0/65536.0,1,-nbitq), 
to_sfixed(3577.0/65536.0,1,-nbitq), 
to_sfixed(1068.0/65536.0,1,-nbitq), 
to_sfixed(-4810.0/65536.0,1,-nbitq), 
to_sfixed(10634.0/65536.0,1,-nbitq), 
to_sfixed(-1795.0/65536.0,1,-nbitq), 
to_sfixed(-8799.0/65536.0,1,-nbitq), 
to_sfixed(1411.0/65536.0,1,-nbitq), 
to_sfixed(-2379.0/65536.0,1,-nbitq), 
to_sfixed(-33.0/65536.0,1,-nbitq), 
to_sfixed(82.0/65536.0,1,-nbitq), 
to_sfixed(6031.0/65536.0,1,-nbitq), 
to_sfixed(-3349.0/65536.0,1,-nbitq), 
to_sfixed(6747.0/65536.0,1,-nbitq), 
to_sfixed(2952.0/65536.0,1,-nbitq), 
to_sfixed(19.0/65536.0,1,-nbitq), 
to_sfixed(1422.0/65536.0,1,-nbitq), 
to_sfixed(-12391.0/65536.0,1,-nbitq), 
to_sfixed(-2435.0/65536.0,1,-nbitq), 
to_sfixed(9277.0/65536.0,1,-nbitq), 
to_sfixed(-1194.0/65536.0,1,-nbitq), 
to_sfixed(-2997.0/65536.0,1,-nbitq), 
to_sfixed(-3376.0/65536.0,1,-nbitq), 
to_sfixed(291.0/65536.0,1,-nbitq), 
to_sfixed(-1807.0/65536.0,1,-nbitq), 
to_sfixed(908.0/65536.0,1,-nbitq), 
to_sfixed(-924.0/65536.0,1,-nbitq), 
to_sfixed(-1516.0/65536.0,1,-nbitq), 
to_sfixed(2207.0/65536.0,1,-nbitq), 
to_sfixed(-504.0/65536.0,1,-nbitq), 
to_sfixed(2781.0/65536.0,1,-nbitq), 
to_sfixed(-9858.0/65536.0,1,-nbitq), 
to_sfixed(-8993.0/65536.0,1,-nbitq), 
to_sfixed(6245.0/65536.0,1,-nbitq), 
to_sfixed(-117.0/65536.0,1,-nbitq), 
to_sfixed(493.0/65536.0,1,-nbitq), 
to_sfixed(-1860.0/65536.0,1,-nbitq), 
to_sfixed(10993.0/65536.0,1,-nbitq), 
to_sfixed(-10037.0/65536.0,1,-nbitq), 
to_sfixed(2537.0/65536.0,1,-nbitq), 
to_sfixed(65.0/65536.0,1,-nbitq), 
to_sfixed(-3074.0/65536.0,1,-nbitq), 
to_sfixed(2127.0/65536.0,1,-nbitq), 
to_sfixed(3576.0/65536.0,1,-nbitq), 
to_sfixed(1200.0/65536.0,1,-nbitq), 
to_sfixed(7279.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-36.0/65536.0,1,-nbitq), 
to_sfixed(5735.0/65536.0,1,-nbitq), 
to_sfixed(4592.0/65536.0,1,-nbitq), 
to_sfixed(-8683.0/65536.0,1,-nbitq), 
to_sfixed(838.0/65536.0,1,-nbitq), 
to_sfixed(7070.0/65536.0,1,-nbitq), 
to_sfixed(2009.0/65536.0,1,-nbitq), 
to_sfixed(-1171.0/65536.0,1,-nbitq), 
to_sfixed(11939.0/65536.0,1,-nbitq), 
to_sfixed(-3035.0/65536.0,1,-nbitq), 
to_sfixed(2250.0/65536.0,1,-nbitq), 
to_sfixed(-9702.0/65536.0,1,-nbitq), 
to_sfixed(83.0/65536.0,1,-nbitq), 
to_sfixed(-2632.0/65536.0,1,-nbitq), 
to_sfixed(237.0/65536.0,1,-nbitq), 
to_sfixed(2355.0/65536.0,1,-nbitq), 
to_sfixed(2738.0/65536.0,1,-nbitq), 
to_sfixed(-3832.0/65536.0,1,-nbitq), 
to_sfixed(2621.0/65536.0,1,-nbitq), 
to_sfixed(-1971.0/65536.0,1,-nbitq), 
to_sfixed(1551.0/65536.0,1,-nbitq), 
to_sfixed(288.0/65536.0,1,-nbitq), 
to_sfixed(-14378.0/65536.0,1,-nbitq), 
to_sfixed(4800.0/65536.0,1,-nbitq), 
to_sfixed(1020.0/65536.0,1,-nbitq), 
to_sfixed(1860.0/65536.0,1,-nbitq), 
to_sfixed(-1747.0/65536.0,1,-nbitq), 
to_sfixed(-1126.0/65536.0,1,-nbitq), 
to_sfixed(2055.0/65536.0,1,-nbitq), 
to_sfixed(-2014.0/65536.0,1,-nbitq), 
to_sfixed(-2572.0/65536.0,1,-nbitq), 
to_sfixed(-7775.0/65536.0,1,-nbitq), 
to_sfixed(-8654.0/65536.0,1,-nbitq), 
to_sfixed(1498.0/65536.0,1,-nbitq), 
to_sfixed(-2391.0/65536.0,1,-nbitq), 
to_sfixed(2933.0/65536.0,1,-nbitq), 
to_sfixed(3490.0/65536.0,1,-nbitq), 
to_sfixed(562.0/65536.0,1,-nbitq), 
to_sfixed(14732.0/65536.0,1,-nbitq), 
to_sfixed(-317.0/65536.0,1,-nbitq), 
to_sfixed(-7720.0/65536.0,1,-nbitq), 
to_sfixed(-2193.0/65536.0,1,-nbitq), 
to_sfixed(-9074.0/65536.0,1,-nbitq), 
to_sfixed(-1420.0/65536.0,1,-nbitq), 
to_sfixed(-1228.0/65536.0,1,-nbitq), 
to_sfixed(3943.0/65536.0,1,-nbitq), 
to_sfixed(-1342.0/65536.0,1,-nbitq), 
to_sfixed(1927.0/65536.0,1,-nbitq), 
to_sfixed(-2095.0/65536.0,1,-nbitq), 
to_sfixed(541.0/65536.0,1,-nbitq), 
to_sfixed(36.0/65536.0,1,-nbitq), 
to_sfixed(590.0/65536.0,1,-nbitq), 
to_sfixed(-3415.0/65536.0,1,-nbitq), 
to_sfixed(588.0/65536.0,1,-nbitq), 
to_sfixed(-4842.0/65536.0,1,-nbitq), 
to_sfixed(-4104.0/65536.0,1,-nbitq), 
to_sfixed(-2596.0/65536.0,1,-nbitq), 
to_sfixed(2118.0/65536.0,1,-nbitq), 
to_sfixed(-586.0/65536.0,1,-nbitq), 
to_sfixed(874.0/65536.0,1,-nbitq), 
to_sfixed(-973.0/65536.0,1,-nbitq), 
to_sfixed(504.0/65536.0,1,-nbitq), 
to_sfixed(848.0/65536.0,1,-nbitq), 
to_sfixed(-858.0/65536.0,1,-nbitq), 
to_sfixed(4477.0/65536.0,1,-nbitq), 
to_sfixed(-7763.0/65536.0,1,-nbitq), 
to_sfixed(-9604.0/65536.0,1,-nbitq), 
to_sfixed(3507.0/65536.0,1,-nbitq), 
to_sfixed(5424.0/65536.0,1,-nbitq), 
to_sfixed(-1125.0/65536.0,1,-nbitq), 
to_sfixed(-30.0/65536.0,1,-nbitq), 
to_sfixed(5962.0/65536.0,1,-nbitq), 
to_sfixed(-6490.0/65536.0,1,-nbitq), 
to_sfixed(737.0/65536.0,1,-nbitq), 
to_sfixed(-2140.0/65536.0,1,-nbitq), 
to_sfixed(-2686.0/65536.0,1,-nbitq), 
to_sfixed(5302.0/65536.0,1,-nbitq), 
to_sfixed(8813.0/65536.0,1,-nbitq), 
to_sfixed(-2194.0/65536.0,1,-nbitq), 
to_sfixed(4534.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2407.0/65536.0,1,-nbitq), 
to_sfixed(2481.0/65536.0,1,-nbitq), 
to_sfixed(1844.0/65536.0,1,-nbitq), 
to_sfixed(-4700.0/65536.0,1,-nbitq), 
to_sfixed(-1945.0/65536.0,1,-nbitq), 
to_sfixed(14455.0/65536.0,1,-nbitq), 
to_sfixed(-2017.0/65536.0,1,-nbitq), 
to_sfixed(329.0/65536.0,1,-nbitq), 
to_sfixed(11563.0/65536.0,1,-nbitq), 
to_sfixed(-3112.0/65536.0,1,-nbitq), 
to_sfixed(3130.0/65536.0,1,-nbitq), 
to_sfixed(-6457.0/65536.0,1,-nbitq), 
to_sfixed(-215.0/65536.0,1,-nbitq), 
to_sfixed(-2776.0/65536.0,1,-nbitq), 
to_sfixed(1853.0/65536.0,1,-nbitq), 
to_sfixed(1058.0/65536.0,1,-nbitq), 
to_sfixed(469.0/65536.0,1,-nbitq), 
to_sfixed(-3144.0/65536.0,1,-nbitq), 
to_sfixed(221.0/65536.0,1,-nbitq), 
to_sfixed(2582.0/65536.0,1,-nbitq), 
to_sfixed(2208.0/65536.0,1,-nbitq), 
to_sfixed(-6485.0/65536.0,1,-nbitq), 
to_sfixed(-262.0/65536.0,1,-nbitq), 
to_sfixed(6148.0/65536.0,1,-nbitq), 
to_sfixed(415.0/65536.0,1,-nbitq), 
to_sfixed(930.0/65536.0,1,-nbitq), 
to_sfixed(1810.0/65536.0,1,-nbitq), 
to_sfixed(-1370.0/65536.0,1,-nbitq), 
to_sfixed(-523.0/65536.0,1,-nbitq), 
to_sfixed(886.0/65536.0,1,-nbitq), 
to_sfixed(-356.0/65536.0,1,-nbitq), 
to_sfixed(-6961.0/65536.0,1,-nbitq), 
to_sfixed(-6811.0/65536.0,1,-nbitq), 
to_sfixed(2751.0/65536.0,1,-nbitq), 
to_sfixed(-1854.0/65536.0,1,-nbitq), 
to_sfixed(3399.0/65536.0,1,-nbitq), 
to_sfixed(2301.0/65536.0,1,-nbitq), 
to_sfixed(5203.0/65536.0,1,-nbitq), 
to_sfixed(7558.0/65536.0,1,-nbitq), 
to_sfixed(-2038.0/65536.0,1,-nbitq), 
to_sfixed(-8477.0/65536.0,1,-nbitq), 
to_sfixed(-2894.0/65536.0,1,-nbitq), 
to_sfixed(-15677.0/65536.0,1,-nbitq), 
to_sfixed(-2414.0/65536.0,1,-nbitq), 
to_sfixed(-1736.0/65536.0,1,-nbitq), 
to_sfixed(-5371.0/65536.0,1,-nbitq), 
to_sfixed(-650.0/65536.0,1,-nbitq), 
to_sfixed(4065.0/65536.0,1,-nbitq), 
to_sfixed(-1325.0/65536.0,1,-nbitq), 
to_sfixed(1713.0/65536.0,1,-nbitq), 
to_sfixed(-2126.0/65536.0,1,-nbitq), 
to_sfixed(6263.0/65536.0,1,-nbitq), 
to_sfixed(2754.0/65536.0,1,-nbitq), 
to_sfixed(7302.0/65536.0,1,-nbitq), 
to_sfixed(-3278.0/65536.0,1,-nbitq), 
to_sfixed(-1887.0/65536.0,1,-nbitq), 
to_sfixed(-2851.0/65536.0,1,-nbitq), 
to_sfixed(539.0/65536.0,1,-nbitq), 
to_sfixed(-1856.0/65536.0,1,-nbitq), 
to_sfixed(2544.0/65536.0,1,-nbitq), 
to_sfixed(4799.0/65536.0,1,-nbitq), 
to_sfixed(-2086.0/65536.0,1,-nbitq), 
to_sfixed(2341.0/65536.0,1,-nbitq), 
to_sfixed(1827.0/65536.0,1,-nbitq), 
to_sfixed(2109.0/65536.0,1,-nbitq), 
to_sfixed(-8736.0/65536.0,1,-nbitq), 
to_sfixed(-13704.0/65536.0,1,-nbitq), 
to_sfixed(5442.0/65536.0,1,-nbitq), 
to_sfixed(4431.0/65536.0,1,-nbitq), 
to_sfixed(870.0/65536.0,1,-nbitq), 
to_sfixed(-2019.0/65536.0,1,-nbitq), 
to_sfixed(1551.0/65536.0,1,-nbitq), 
to_sfixed(6344.0/65536.0,1,-nbitq), 
to_sfixed(-2940.0/65536.0,1,-nbitq), 
to_sfixed(2821.0/65536.0,1,-nbitq), 
to_sfixed(282.0/65536.0,1,-nbitq), 
to_sfixed(4412.0/65536.0,1,-nbitq), 
to_sfixed(2846.0/65536.0,1,-nbitq), 
to_sfixed(1797.0/65536.0,1,-nbitq), 
to_sfixed(3876.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2276.0/65536.0,1,-nbitq), 
to_sfixed(-2684.0/65536.0,1,-nbitq), 
to_sfixed(3487.0/65536.0,1,-nbitq), 
to_sfixed(-54.0/65536.0,1,-nbitq), 
to_sfixed(-731.0/65536.0,1,-nbitq), 
to_sfixed(13202.0/65536.0,1,-nbitq), 
to_sfixed(2157.0/65536.0,1,-nbitq), 
to_sfixed(2375.0/65536.0,1,-nbitq), 
to_sfixed(8318.0/65536.0,1,-nbitq), 
to_sfixed(1251.0/65536.0,1,-nbitq), 
to_sfixed(3442.0/65536.0,1,-nbitq), 
to_sfixed(-1017.0/65536.0,1,-nbitq), 
to_sfixed(-255.0/65536.0,1,-nbitq), 
to_sfixed(-468.0/65536.0,1,-nbitq), 
to_sfixed(-216.0/65536.0,1,-nbitq), 
to_sfixed(968.0/65536.0,1,-nbitq), 
to_sfixed(-2782.0/65536.0,1,-nbitq), 
to_sfixed(-6713.0/65536.0,1,-nbitq), 
to_sfixed(-1627.0/65536.0,1,-nbitq), 
to_sfixed(-862.0/65536.0,1,-nbitq), 
to_sfixed(7582.0/65536.0,1,-nbitq), 
to_sfixed(-1985.0/65536.0,1,-nbitq), 
to_sfixed(4521.0/65536.0,1,-nbitq), 
to_sfixed(4815.0/65536.0,1,-nbitq), 
to_sfixed(-191.0/65536.0,1,-nbitq), 
to_sfixed(4380.0/65536.0,1,-nbitq), 
to_sfixed(202.0/65536.0,1,-nbitq), 
to_sfixed(-1819.0/65536.0,1,-nbitq), 
to_sfixed(4258.0/65536.0,1,-nbitq), 
to_sfixed(-1124.0/65536.0,1,-nbitq), 
to_sfixed(978.0/65536.0,1,-nbitq), 
to_sfixed(-4520.0/65536.0,1,-nbitq), 
to_sfixed(-7984.0/65536.0,1,-nbitq), 
to_sfixed(5536.0/65536.0,1,-nbitq), 
to_sfixed(705.0/65536.0,1,-nbitq), 
to_sfixed(4036.0/65536.0,1,-nbitq), 
to_sfixed(2501.0/65536.0,1,-nbitq), 
to_sfixed(-4814.0/65536.0,1,-nbitq), 
to_sfixed(-1016.0/65536.0,1,-nbitq), 
to_sfixed(-3569.0/65536.0,1,-nbitq), 
to_sfixed(-5666.0/65536.0,1,-nbitq), 
to_sfixed(1690.0/65536.0,1,-nbitq), 
to_sfixed(-7762.0/65536.0,1,-nbitq), 
to_sfixed(-6999.0/65536.0,1,-nbitq), 
to_sfixed(-1560.0/65536.0,1,-nbitq), 
to_sfixed(-6005.0/65536.0,1,-nbitq), 
to_sfixed(-670.0/65536.0,1,-nbitq), 
to_sfixed(163.0/65536.0,1,-nbitq), 
to_sfixed(-924.0/65536.0,1,-nbitq), 
to_sfixed(1976.0/65536.0,1,-nbitq), 
to_sfixed(208.0/65536.0,1,-nbitq), 
to_sfixed(-596.0/65536.0,1,-nbitq), 
to_sfixed(-2012.0/65536.0,1,-nbitq), 
to_sfixed(7384.0/65536.0,1,-nbitq), 
to_sfixed(151.0/65536.0,1,-nbitq), 
to_sfixed(-3098.0/65536.0,1,-nbitq), 
to_sfixed(1588.0/65536.0,1,-nbitq), 
to_sfixed(-4771.0/65536.0,1,-nbitq), 
to_sfixed(-2872.0/65536.0,1,-nbitq), 
to_sfixed(-172.0/65536.0,1,-nbitq), 
to_sfixed(3818.0/65536.0,1,-nbitq), 
to_sfixed(-1503.0/65536.0,1,-nbitq), 
to_sfixed(2042.0/65536.0,1,-nbitq), 
to_sfixed(530.0/65536.0,1,-nbitq), 
to_sfixed(-5134.0/65536.0,1,-nbitq), 
to_sfixed(-4277.0/65536.0,1,-nbitq), 
to_sfixed(-10105.0/65536.0,1,-nbitq), 
to_sfixed(1423.0/65536.0,1,-nbitq), 
to_sfixed(-4303.0/65536.0,1,-nbitq), 
to_sfixed(-6996.0/65536.0,1,-nbitq), 
to_sfixed(-2544.0/65536.0,1,-nbitq), 
to_sfixed(5444.0/65536.0,1,-nbitq), 
to_sfixed(8843.0/65536.0,1,-nbitq), 
to_sfixed(1372.0/65536.0,1,-nbitq), 
to_sfixed(-2793.0/65536.0,1,-nbitq), 
to_sfixed(5143.0/65536.0,1,-nbitq), 
to_sfixed(4664.0/65536.0,1,-nbitq), 
to_sfixed(-3188.0/65536.0,1,-nbitq), 
to_sfixed(3004.0/65536.0,1,-nbitq), 
to_sfixed(1171.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-5222.0/65536.0,1,-nbitq), 
to_sfixed(-2924.0/65536.0,1,-nbitq), 
to_sfixed(1346.0/65536.0,1,-nbitq), 
to_sfixed(-5331.0/65536.0,1,-nbitq), 
to_sfixed(7432.0/65536.0,1,-nbitq), 
to_sfixed(14161.0/65536.0,1,-nbitq), 
to_sfixed(-1959.0/65536.0,1,-nbitq), 
to_sfixed(450.0/65536.0,1,-nbitq), 
to_sfixed(546.0/65536.0,1,-nbitq), 
to_sfixed(2280.0/65536.0,1,-nbitq), 
to_sfixed(-1948.0/65536.0,1,-nbitq), 
to_sfixed(-475.0/65536.0,1,-nbitq), 
to_sfixed(1729.0/65536.0,1,-nbitq), 
to_sfixed(4533.0/65536.0,1,-nbitq), 
to_sfixed(-1372.0/65536.0,1,-nbitq), 
to_sfixed(-125.0/65536.0,1,-nbitq), 
to_sfixed(-1873.0/65536.0,1,-nbitq), 
to_sfixed(-6970.0/65536.0,1,-nbitq), 
to_sfixed(-1550.0/65536.0,1,-nbitq), 
to_sfixed(-180.0/65536.0,1,-nbitq), 
to_sfixed(2283.0/65536.0,1,-nbitq), 
to_sfixed(-4234.0/65536.0,1,-nbitq), 
to_sfixed(7191.0/65536.0,1,-nbitq), 
to_sfixed(708.0/65536.0,1,-nbitq), 
to_sfixed(2127.0/65536.0,1,-nbitq), 
to_sfixed(6265.0/65536.0,1,-nbitq), 
to_sfixed(3997.0/65536.0,1,-nbitq), 
to_sfixed(2598.0/65536.0,1,-nbitq), 
to_sfixed(1496.0/65536.0,1,-nbitq), 
to_sfixed(3009.0/65536.0,1,-nbitq), 
to_sfixed(1560.0/65536.0,1,-nbitq), 
to_sfixed(-2662.0/65536.0,1,-nbitq), 
to_sfixed(-4743.0/65536.0,1,-nbitq), 
to_sfixed(4027.0/65536.0,1,-nbitq), 
to_sfixed(1958.0/65536.0,1,-nbitq), 
to_sfixed(1212.0/65536.0,1,-nbitq), 
to_sfixed(4890.0/65536.0,1,-nbitq), 
to_sfixed(-2342.0/65536.0,1,-nbitq), 
to_sfixed(5773.0/65536.0,1,-nbitq), 
to_sfixed(2271.0/65536.0,1,-nbitq), 
to_sfixed(3927.0/65536.0,1,-nbitq), 
to_sfixed(2185.0/65536.0,1,-nbitq), 
to_sfixed(5133.0/65536.0,1,-nbitq), 
to_sfixed(485.0/65536.0,1,-nbitq), 
to_sfixed(1529.0/65536.0,1,-nbitq), 
to_sfixed(-9322.0/65536.0,1,-nbitq), 
to_sfixed(353.0/65536.0,1,-nbitq), 
to_sfixed(-7515.0/65536.0,1,-nbitq), 
to_sfixed(1220.0/65536.0,1,-nbitq), 
to_sfixed(267.0/65536.0,1,-nbitq), 
to_sfixed(-695.0/65536.0,1,-nbitq), 
to_sfixed(-2546.0/65536.0,1,-nbitq), 
to_sfixed(-8882.0/65536.0,1,-nbitq), 
to_sfixed(-5759.0/65536.0,1,-nbitq), 
to_sfixed(2397.0/65536.0,1,-nbitq), 
to_sfixed(3120.0/65536.0,1,-nbitq), 
to_sfixed(3744.0/65536.0,1,-nbitq), 
to_sfixed(158.0/65536.0,1,-nbitq), 
to_sfixed(-2918.0/65536.0,1,-nbitq), 
to_sfixed(-3690.0/65536.0,1,-nbitq), 
to_sfixed(-4274.0/65536.0,1,-nbitq), 
to_sfixed(-549.0/65536.0,1,-nbitq), 
to_sfixed(753.0/65536.0,1,-nbitq), 
to_sfixed(1973.0/65536.0,1,-nbitq), 
to_sfixed(1459.0/65536.0,1,-nbitq), 
to_sfixed(226.0/65536.0,1,-nbitq), 
to_sfixed(-2175.0/65536.0,1,-nbitq), 
to_sfixed(8425.0/65536.0,1,-nbitq), 
to_sfixed(-8364.0/65536.0,1,-nbitq), 
to_sfixed(-8119.0/65536.0,1,-nbitq), 
to_sfixed(-3870.0/65536.0,1,-nbitq), 
to_sfixed(8337.0/65536.0,1,-nbitq), 
to_sfixed(3627.0/65536.0,1,-nbitq), 
to_sfixed(-332.0/65536.0,1,-nbitq), 
to_sfixed(2379.0/65536.0,1,-nbitq), 
to_sfixed(1730.0/65536.0,1,-nbitq), 
to_sfixed(9529.0/65536.0,1,-nbitq), 
to_sfixed(-11083.0/65536.0,1,-nbitq), 
to_sfixed(-992.0/65536.0,1,-nbitq), 
to_sfixed(-1380.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-6011.0/65536.0,1,-nbitq), 
to_sfixed(1454.0/65536.0,1,-nbitq), 
to_sfixed(-2596.0/65536.0,1,-nbitq), 
to_sfixed(-2221.0/65536.0,1,-nbitq), 
to_sfixed(2891.0/65536.0,1,-nbitq), 
to_sfixed(7164.0/65536.0,1,-nbitq), 
to_sfixed(2580.0/65536.0,1,-nbitq), 
to_sfixed(4567.0/65536.0,1,-nbitq), 
to_sfixed(1329.0/65536.0,1,-nbitq), 
to_sfixed(2363.0/65536.0,1,-nbitq), 
to_sfixed(-417.0/65536.0,1,-nbitq), 
to_sfixed(-1187.0/65536.0,1,-nbitq), 
to_sfixed(-1796.0/65536.0,1,-nbitq), 
to_sfixed(12364.0/65536.0,1,-nbitq), 
to_sfixed(-4680.0/65536.0,1,-nbitq), 
to_sfixed(556.0/65536.0,1,-nbitq), 
to_sfixed(-2782.0/65536.0,1,-nbitq), 
to_sfixed(-5129.0/65536.0,1,-nbitq), 
to_sfixed(-2105.0/65536.0,1,-nbitq), 
to_sfixed(-2692.0/65536.0,1,-nbitq), 
to_sfixed(4393.0/65536.0,1,-nbitq), 
to_sfixed(687.0/65536.0,1,-nbitq), 
to_sfixed(-611.0/65536.0,1,-nbitq), 
to_sfixed(12412.0/65536.0,1,-nbitq), 
to_sfixed(-3789.0/65536.0,1,-nbitq), 
to_sfixed(1776.0/65536.0,1,-nbitq), 
to_sfixed(2739.0/65536.0,1,-nbitq), 
to_sfixed(2403.0/65536.0,1,-nbitq), 
to_sfixed(1408.0/65536.0,1,-nbitq), 
to_sfixed(-2993.0/65536.0,1,-nbitq), 
to_sfixed(-1060.0/65536.0,1,-nbitq), 
to_sfixed(-1993.0/65536.0,1,-nbitq), 
to_sfixed(3009.0/65536.0,1,-nbitq), 
to_sfixed(5428.0/65536.0,1,-nbitq), 
to_sfixed(-665.0/65536.0,1,-nbitq), 
to_sfixed(-325.0/65536.0,1,-nbitq), 
to_sfixed(9449.0/65536.0,1,-nbitq), 
to_sfixed(4027.0/65536.0,1,-nbitq), 
to_sfixed(5455.0/65536.0,1,-nbitq), 
to_sfixed(2090.0/65536.0,1,-nbitq), 
to_sfixed(5910.0/65536.0,1,-nbitq), 
to_sfixed(-844.0/65536.0,1,-nbitq), 
to_sfixed(6914.0/65536.0,1,-nbitq), 
to_sfixed(-4274.0/65536.0,1,-nbitq), 
to_sfixed(-2691.0/65536.0,1,-nbitq), 
to_sfixed(-1806.0/65536.0,1,-nbitq), 
to_sfixed(-1873.0/65536.0,1,-nbitq), 
to_sfixed(-3808.0/65536.0,1,-nbitq), 
to_sfixed(1951.0/65536.0,1,-nbitq), 
to_sfixed(2530.0/65536.0,1,-nbitq), 
to_sfixed(362.0/65536.0,1,-nbitq), 
to_sfixed(-6177.0/65536.0,1,-nbitq), 
to_sfixed(-10731.0/65536.0,1,-nbitq), 
to_sfixed(-2017.0/65536.0,1,-nbitq), 
to_sfixed(7320.0/65536.0,1,-nbitq), 
to_sfixed(2690.0/65536.0,1,-nbitq), 
to_sfixed(1439.0/65536.0,1,-nbitq), 
to_sfixed(-570.0/65536.0,1,-nbitq), 
to_sfixed(-1731.0/65536.0,1,-nbitq), 
to_sfixed(-4315.0/65536.0,1,-nbitq), 
to_sfixed(1274.0/65536.0,1,-nbitq), 
to_sfixed(498.0/65536.0,1,-nbitq), 
to_sfixed(1999.0/65536.0,1,-nbitq), 
to_sfixed(-1991.0/65536.0,1,-nbitq), 
to_sfixed(-3887.0/65536.0,1,-nbitq), 
to_sfixed(-5084.0/65536.0,1,-nbitq), 
to_sfixed(-7914.0/65536.0,1,-nbitq), 
to_sfixed(2133.0/65536.0,1,-nbitq), 
to_sfixed(-2022.0/65536.0,1,-nbitq), 
to_sfixed(-2045.0/65536.0,1,-nbitq), 
to_sfixed(-762.0/65536.0,1,-nbitq), 
to_sfixed(4979.0/65536.0,1,-nbitq), 
to_sfixed(1190.0/65536.0,1,-nbitq), 
to_sfixed(-2854.0/65536.0,1,-nbitq), 
to_sfixed(-1155.0/65536.0,1,-nbitq), 
to_sfixed(2746.0/65536.0,1,-nbitq), 
to_sfixed(4824.0/65536.0,1,-nbitq), 
to_sfixed(-14217.0/65536.0,1,-nbitq), 
to_sfixed(276.0/65536.0,1,-nbitq), 
to_sfixed(-2003.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-517.0/65536.0,1,-nbitq), 
to_sfixed(-1123.0/65536.0,1,-nbitq), 
to_sfixed(-652.0/65536.0,1,-nbitq), 
to_sfixed(-3012.0/65536.0,1,-nbitq), 
to_sfixed(2084.0/65536.0,1,-nbitq), 
to_sfixed(4864.0/65536.0,1,-nbitq), 
to_sfixed(-243.0/65536.0,1,-nbitq), 
to_sfixed(4480.0/65536.0,1,-nbitq), 
to_sfixed(472.0/65536.0,1,-nbitq), 
to_sfixed(1837.0/65536.0,1,-nbitq), 
to_sfixed(-1240.0/65536.0,1,-nbitq), 
to_sfixed(4847.0/65536.0,1,-nbitq), 
to_sfixed(-569.0/65536.0,1,-nbitq), 
to_sfixed(9615.0/65536.0,1,-nbitq), 
to_sfixed(-2006.0/65536.0,1,-nbitq), 
to_sfixed(-1187.0/65536.0,1,-nbitq), 
to_sfixed(-2535.0/65536.0,1,-nbitq), 
to_sfixed(1430.0/65536.0,1,-nbitq), 
to_sfixed(-3964.0/65536.0,1,-nbitq), 
to_sfixed(2406.0/65536.0,1,-nbitq), 
to_sfixed(2124.0/65536.0,1,-nbitq), 
to_sfixed(2834.0/65536.0,1,-nbitq), 
to_sfixed(1936.0/65536.0,1,-nbitq), 
to_sfixed(7570.0/65536.0,1,-nbitq), 
to_sfixed(-1216.0/65536.0,1,-nbitq), 
to_sfixed(2395.0/65536.0,1,-nbitq), 
to_sfixed(3614.0/65536.0,1,-nbitq), 
to_sfixed(-1349.0/65536.0,1,-nbitq), 
to_sfixed(1805.0/65536.0,1,-nbitq), 
to_sfixed(-175.0/65536.0,1,-nbitq), 
to_sfixed(-3411.0/65536.0,1,-nbitq), 
to_sfixed(6.0/65536.0,1,-nbitq), 
to_sfixed(2514.0/65536.0,1,-nbitq), 
to_sfixed(1150.0/65536.0,1,-nbitq), 
to_sfixed(-2221.0/65536.0,1,-nbitq), 
to_sfixed(-222.0/65536.0,1,-nbitq), 
to_sfixed(6620.0/65536.0,1,-nbitq), 
to_sfixed(-3636.0/65536.0,1,-nbitq), 
to_sfixed(4804.0/65536.0,1,-nbitq), 
to_sfixed(1497.0/65536.0,1,-nbitq), 
to_sfixed(10412.0/65536.0,1,-nbitq), 
to_sfixed(-2179.0/65536.0,1,-nbitq), 
to_sfixed(5704.0/65536.0,1,-nbitq), 
to_sfixed(-3804.0/65536.0,1,-nbitq), 
to_sfixed(2062.0/65536.0,1,-nbitq), 
to_sfixed(492.0/65536.0,1,-nbitq), 
to_sfixed(2977.0/65536.0,1,-nbitq), 
to_sfixed(-1937.0/65536.0,1,-nbitq), 
to_sfixed(-2158.0/65536.0,1,-nbitq), 
to_sfixed(-1254.0/65536.0,1,-nbitq), 
to_sfixed(-1984.0/65536.0,1,-nbitq), 
to_sfixed(-3535.0/65536.0,1,-nbitq), 
to_sfixed(-7635.0/65536.0,1,-nbitq), 
to_sfixed(-2314.0/65536.0,1,-nbitq), 
to_sfixed(6407.0/65536.0,1,-nbitq), 
to_sfixed(6902.0/65536.0,1,-nbitq), 
to_sfixed(-2730.0/65536.0,1,-nbitq), 
to_sfixed(3566.0/65536.0,1,-nbitq), 
to_sfixed(-675.0/65536.0,1,-nbitq), 
to_sfixed(-1201.0/65536.0,1,-nbitq), 
to_sfixed(383.0/65536.0,1,-nbitq), 
to_sfixed(-1540.0/65536.0,1,-nbitq), 
to_sfixed(-1932.0/65536.0,1,-nbitq), 
to_sfixed(-2993.0/65536.0,1,-nbitq), 
to_sfixed(-5670.0/65536.0,1,-nbitq), 
to_sfixed(-3414.0/65536.0,1,-nbitq), 
to_sfixed(-6309.0/65536.0,1,-nbitq), 
to_sfixed(4717.0/65536.0,1,-nbitq), 
to_sfixed(-4024.0/65536.0,1,-nbitq), 
to_sfixed(-3864.0/65536.0,1,-nbitq), 
to_sfixed(1978.0/65536.0,1,-nbitq), 
to_sfixed(3184.0/65536.0,1,-nbitq), 
to_sfixed(254.0/65536.0,1,-nbitq), 
to_sfixed(-1174.0/65536.0,1,-nbitq), 
to_sfixed(659.0/65536.0,1,-nbitq), 
to_sfixed(4352.0/65536.0,1,-nbitq), 
to_sfixed(209.0/65536.0,1,-nbitq), 
to_sfixed(-10028.0/65536.0,1,-nbitq), 
to_sfixed(-53.0/65536.0,1,-nbitq), 
to_sfixed(-5550.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5185.0/65536.0,1,-nbitq), 
to_sfixed(5008.0/65536.0,1,-nbitq), 
to_sfixed(-5218.0/65536.0,1,-nbitq), 
to_sfixed(-4049.0/65536.0,1,-nbitq), 
to_sfixed(580.0/65536.0,1,-nbitq), 
to_sfixed(719.0/65536.0,1,-nbitq), 
to_sfixed(-1009.0/65536.0,1,-nbitq), 
to_sfixed(-13.0/65536.0,1,-nbitq), 
to_sfixed(-3703.0/65536.0,1,-nbitq), 
to_sfixed(-690.0/65536.0,1,-nbitq), 
to_sfixed(-3276.0/65536.0,1,-nbitq), 
to_sfixed(518.0/65536.0,1,-nbitq), 
to_sfixed(-2835.0/65536.0,1,-nbitq), 
to_sfixed(3679.0/65536.0,1,-nbitq), 
to_sfixed(-730.0/65536.0,1,-nbitq), 
to_sfixed(-1059.0/65536.0,1,-nbitq), 
to_sfixed(303.0/65536.0,1,-nbitq), 
to_sfixed(-38.0/65536.0,1,-nbitq), 
to_sfixed(-318.0/65536.0,1,-nbitq), 
to_sfixed(2687.0/65536.0,1,-nbitq), 
to_sfixed(463.0/65536.0,1,-nbitq), 
to_sfixed(2204.0/65536.0,1,-nbitq), 
to_sfixed(-1163.0/65536.0,1,-nbitq), 
to_sfixed(3918.0/65536.0,1,-nbitq), 
to_sfixed(-2394.0/65536.0,1,-nbitq), 
to_sfixed(193.0/65536.0,1,-nbitq), 
to_sfixed(1831.0/65536.0,1,-nbitq), 
to_sfixed(-2329.0/65536.0,1,-nbitq), 
to_sfixed(1025.0/65536.0,1,-nbitq), 
to_sfixed(-2834.0/65536.0,1,-nbitq), 
to_sfixed(-4007.0/65536.0,1,-nbitq), 
to_sfixed(-121.0/65536.0,1,-nbitq), 
to_sfixed(1876.0/65536.0,1,-nbitq), 
to_sfixed(-90.0/65536.0,1,-nbitq), 
to_sfixed(-1670.0/65536.0,1,-nbitq), 
to_sfixed(-376.0/65536.0,1,-nbitq), 
to_sfixed(2005.0/65536.0,1,-nbitq), 
to_sfixed(408.0/65536.0,1,-nbitq), 
to_sfixed(6786.0/65536.0,1,-nbitq), 
to_sfixed(-1506.0/65536.0,1,-nbitq), 
to_sfixed(7459.0/65536.0,1,-nbitq), 
to_sfixed(1160.0/65536.0,1,-nbitq), 
to_sfixed(6323.0/65536.0,1,-nbitq), 
to_sfixed(-3348.0/65536.0,1,-nbitq), 
to_sfixed(2229.0/65536.0,1,-nbitq), 
to_sfixed(-1612.0/65536.0,1,-nbitq), 
to_sfixed(1568.0/65536.0,1,-nbitq), 
to_sfixed(-3630.0/65536.0,1,-nbitq), 
to_sfixed(413.0/65536.0,1,-nbitq), 
to_sfixed(3026.0/65536.0,1,-nbitq), 
to_sfixed(-955.0/65536.0,1,-nbitq), 
to_sfixed(-2444.0/65536.0,1,-nbitq), 
to_sfixed(-2863.0/65536.0,1,-nbitq), 
to_sfixed(-3463.0/65536.0,1,-nbitq), 
to_sfixed(5115.0/65536.0,1,-nbitq), 
to_sfixed(-17.0/65536.0,1,-nbitq), 
to_sfixed(2060.0/65536.0,1,-nbitq), 
to_sfixed(3200.0/65536.0,1,-nbitq), 
to_sfixed(-2877.0/65536.0,1,-nbitq), 
to_sfixed(1348.0/65536.0,1,-nbitq), 
to_sfixed(-2362.0/65536.0,1,-nbitq), 
to_sfixed(-2.0/65536.0,1,-nbitq), 
to_sfixed(-818.0/65536.0,1,-nbitq), 
to_sfixed(1305.0/65536.0,1,-nbitq), 
to_sfixed(-6909.0/65536.0,1,-nbitq), 
to_sfixed(-3401.0/65536.0,1,-nbitq), 
to_sfixed(-5654.0/65536.0,1,-nbitq), 
to_sfixed(-2645.0/65536.0,1,-nbitq), 
to_sfixed(-6868.0/65536.0,1,-nbitq), 
to_sfixed(-2991.0/65536.0,1,-nbitq), 
to_sfixed(2661.0/65536.0,1,-nbitq), 
to_sfixed(2088.0/65536.0,1,-nbitq), 
to_sfixed(3232.0/65536.0,1,-nbitq), 
to_sfixed(-127.0/65536.0,1,-nbitq), 
to_sfixed(-622.0/65536.0,1,-nbitq), 
to_sfixed(2484.0/65536.0,1,-nbitq), 
to_sfixed(714.0/65536.0,1,-nbitq), 
to_sfixed(1296.0/65536.0,1,-nbitq), 
to_sfixed(-1901.0/65536.0,1,-nbitq), 
to_sfixed(-9363.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2437.0/65536.0,1,-nbitq), 
to_sfixed(3055.0/65536.0,1,-nbitq), 
to_sfixed(-2037.0/65536.0,1,-nbitq), 
to_sfixed(-1613.0/65536.0,1,-nbitq), 
to_sfixed(-2902.0/65536.0,1,-nbitq), 
to_sfixed(2460.0/65536.0,1,-nbitq), 
to_sfixed(-2174.0/65536.0,1,-nbitq), 
to_sfixed(809.0/65536.0,1,-nbitq), 
to_sfixed(-2872.0/65536.0,1,-nbitq), 
to_sfixed(2549.0/65536.0,1,-nbitq), 
to_sfixed(1986.0/65536.0,1,-nbitq), 
to_sfixed(7152.0/65536.0,1,-nbitq), 
to_sfixed(-2096.0/65536.0,1,-nbitq), 
to_sfixed(1430.0/65536.0,1,-nbitq), 
to_sfixed(-1975.0/65536.0,1,-nbitq), 
to_sfixed(-805.0/65536.0,1,-nbitq), 
to_sfixed(175.0/65536.0,1,-nbitq), 
to_sfixed(3359.0/65536.0,1,-nbitq), 
to_sfixed(-3788.0/65536.0,1,-nbitq), 
to_sfixed(1816.0/65536.0,1,-nbitq), 
to_sfixed(-1898.0/65536.0,1,-nbitq), 
to_sfixed(8472.0/65536.0,1,-nbitq), 
to_sfixed(-1349.0/65536.0,1,-nbitq), 
to_sfixed(3075.0/65536.0,1,-nbitq), 
to_sfixed(701.0/65536.0,1,-nbitq), 
to_sfixed(-223.0/65536.0,1,-nbitq), 
to_sfixed(4359.0/65536.0,1,-nbitq), 
to_sfixed(83.0/65536.0,1,-nbitq), 
to_sfixed(1682.0/65536.0,1,-nbitq), 
to_sfixed(546.0/65536.0,1,-nbitq), 
to_sfixed(-2786.0/65536.0,1,-nbitq), 
to_sfixed(-648.0/65536.0,1,-nbitq), 
to_sfixed(9017.0/65536.0,1,-nbitq), 
to_sfixed(1137.0/65536.0,1,-nbitq), 
to_sfixed(-613.0/65536.0,1,-nbitq), 
to_sfixed(1405.0/65536.0,1,-nbitq), 
to_sfixed(-1639.0/65536.0,1,-nbitq), 
to_sfixed(1844.0/65536.0,1,-nbitq), 
to_sfixed(3481.0/65536.0,1,-nbitq), 
to_sfixed(3988.0/65536.0,1,-nbitq), 
to_sfixed(2344.0/65536.0,1,-nbitq), 
to_sfixed(2798.0/65536.0,1,-nbitq), 
to_sfixed(3790.0/65536.0,1,-nbitq), 
to_sfixed(-1512.0/65536.0,1,-nbitq), 
to_sfixed(-1109.0/65536.0,1,-nbitq), 
to_sfixed(-2973.0/65536.0,1,-nbitq), 
to_sfixed(2095.0/65536.0,1,-nbitq), 
to_sfixed(-1297.0/65536.0,1,-nbitq), 
to_sfixed(-2991.0/65536.0,1,-nbitq), 
to_sfixed(-385.0/65536.0,1,-nbitq), 
to_sfixed(616.0/65536.0,1,-nbitq), 
to_sfixed(-1629.0/65536.0,1,-nbitq), 
to_sfixed(554.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(3169.0/65536.0,1,-nbitq), 
to_sfixed(-110.0/65536.0,1,-nbitq), 
to_sfixed(-2661.0/65536.0,1,-nbitq), 
to_sfixed(-343.0/65536.0,1,-nbitq), 
to_sfixed(1151.0/65536.0,1,-nbitq), 
to_sfixed(-1621.0/65536.0,1,-nbitq), 
to_sfixed(238.0/65536.0,1,-nbitq), 
to_sfixed(-452.0/65536.0,1,-nbitq), 
to_sfixed(-2629.0/65536.0,1,-nbitq), 
to_sfixed(1381.0/65536.0,1,-nbitq), 
to_sfixed(-2859.0/65536.0,1,-nbitq), 
to_sfixed(2055.0/65536.0,1,-nbitq), 
to_sfixed(-5213.0/65536.0,1,-nbitq), 
to_sfixed(-2570.0/65536.0,1,-nbitq), 
to_sfixed(-10458.0/65536.0,1,-nbitq), 
to_sfixed(-10623.0/65536.0,1,-nbitq), 
to_sfixed(4415.0/65536.0,1,-nbitq), 
to_sfixed(-1959.0/65536.0,1,-nbitq), 
to_sfixed(848.0/65536.0,1,-nbitq), 
to_sfixed(-1241.0/65536.0,1,-nbitq), 
to_sfixed(1702.0/65536.0,1,-nbitq), 
to_sfixed(1692.0/65536.0,1,-nbitq), 
to_sfixed(1412.0/65536.0,1,-nbitq), 
to_sfixed(-4335.0/65536.0,1,-nbitq), 
to_sfixed(1447.0/65536.0,1,-nbitq), 
to_sfixed(-10593.0/65536.0,1,-nbitq)  ), 
( to_sfixed(227.0/65536.0,1,-nbitq), 
to_sfixed(-1912.0/65536.0,1,-nbitq), 
to_sfixed(-1447.0/65536.0,1,-nbitq), 
to_sfixed(3370.0/65536.0,1,-nbitq), 
to_sfixed(-3668.0/65536.0,1,-nbitq), 
to_sfixed(1572.0/65536.0,1,-nbitq), 
to_sfixed(553.0/65536.0,1,-nbitq), 
to_sfixed(2893.0/65536.0,1,-nbitq), 
to_sfixed(2274.0/65536.0,1,-nbitq), 
to_sfixed(377.0/65536.0,1,-nbitq), 
to_sfixed(-1049.0/65536.0,1,-nbitq), 
to_sfixed(3159.0/65536.0,1,-nbitq), 
to_sfixed(-1052.0/65536.0,1,-nbitq), 
to_sfixed(-1507.0/65536.0,1,-nbitq), 
to_sfixed(-3468.0/65536.0,1,-nbitq), 
to_sfixed(-2656.0/65536.0,1,-nbitq), 
to_sfixed(450.0/65536.0,1,-nbitq), 
to_sfixed(-3425.0/65536.0,1,-nbitq), 
to_sfixed(187.0/65536.0,1,-nbitq), 
to_sfixed(-1357.0/65536.0,1,-nbitq), 
to_sfixed(2783.0/65536.0,1,-nbitq), 
to_sfixed(4108.0/65536.0,1,-nbitq), 
to_sfixed(-1133.0/65536.0,1,-nbitq), 
to_sfixed(4968.0/65536.0,1,-nbitq), 
to_sfixed(1610.0/65536.0,1,-nbitq), 
to_sfixed(3117.0/65536.0,1,-nbitq), 
to_sfixed(4631.0/65536.0,1,-nbitq), 
to_sfixed(-1406.0/65536.0,1,-nbitq), 
to_sfixed(-1050.0/65536.0,1,-nbitq), 
to_sfixed(1426.0/65536.0,1,-nbitq), 
to_sfixed(-613.0/65536.0,1,-nbitq), 
to_sfixed(2782.0/65536.0,1,-nbitq), 
to_sfixed(3240.0/65536.0,1,-nbitq), 
to_sfixed(-960.0/65536.0,1,-nbitq), 
to_sfixed(-2157.0/65536.0,1,-nbitq), 
to_sfixed(2112.0/65536.0,1,-nbitq), 
to_sfixed(-640.0/65536.0,1,-nbitq), 
to_sfixed(1754.0/65536.0,1,-nbitq), 
to_sfixed(3815.0/65536.0,1,-nbitq), 
to_sfixed(3044.0/65536.0,1,-nbitq), 
to_sfixed(-321.0/65536.0,1,-nbitq), 
to_sfixed(-2879.0/65536.0,1,-nbitq), 
to_sfixed(6453.0/65536.0,1,-nbitq), 
to_sfixed(-1418.0/65536.0,1,-nbitq), 
to_sfixed(-2304.0/65536.0,1,-nbitq), 
to_sfixed(-298.0/65536.0,1,-nbitq), 
to_sfixed(-2016.0/65536.0,1,-nbitq), 
to_sfixed(-2519.0/65536.0,1,-nbitq), 
to_sfixed(-2894.0/65536.0,1,-nbitq), 
to_sfixed(1916.0/65536.0,1,-nbitq), 
to_sfixed(2664.0/65536.0,1,-nbitq), 
to_sfixed(-2087.0/65536.0,1,-nbitq), 
to_sfixed(7617.0/65536.0,1,-nbitq), 
to_sfixed(-5073.0/65536.0,1,-nbitq), 
to_sfixed(3312.0/65536.0,1,-nbitq), 
to_sfixed(2000.0/65536.0,1,-nbitq), 
to_sfixed(39.0/65536.0,1,-nbitq), 
to_sfixed(2665.0/65536.0,1,-nbitq), 
to_sfixed(-422.0/65536.0,1,-nbitq), 
to_sfixed(4496.0/65536.0,1,-nbitq), 
to_sfixed(3169.0/65536.0,1,-nbitq), 
to_sfixed(-1960.0/65536.0,1,-nbitq), 
to_sfixed(2523.0/65536.0,1,-nbitq), 
to_sfixed(896.0/65536.0,1,-nbitq), 
to_sfixed(-3436.0/65536.0,1,-nbitq), 
to_sfixed(2189.0/65536.0,1,-nbitq), 
to_sfixed(-4497.0/65536.0,1,-nbitq), 
to_sfixed(-972.0/65536.0,1,-nbitq), 
to_sfixed(-6902.0/65536.0,1,-nbitq), 
to_sfixed(-5963.0/65536.0,1,-nbitq), 
to_sfixed(3473.0/65536.0,1,-nbitq), 
to_sfixed(-2468.0/65536.0,1,-nbitq), 
to_sfixed(1771.0/65536.0,1,-nbitq), 
to_sfixed(-3248.0/65536.0,1,-nbitq), 
to_sfixed(-2027.0/65536.0,1,-nbitq), 
to_sfixed(4519.0/65536.0,1,-nbitq), 
to_sfixed(1441.0/65536.0,1,-nbitq), 
to_sfixed(2493.0/65536.0,1,-nbitq), 
to_sfixed(-1955.0/65536.0,1,-nbitq), 
to_sfixed(-7570.0/65536.0,1,-nbitq)  ), 
( to_sfixed(9.0/65536.0,1,-nbitq), 
to_sfixed(-1605.0/65536.0,1,-nbitq), 
to_sfixed(1940.0/65536.0,1,-nbitq), 
to_sfixed(-359.0/65536.0,1,-nbitq), 
to_sfixed(1514.0/65536.0,1,-nbitq), 
to_sfixed(105.0/65536.0,1,-nbitq), 
to_sfixed(-42.0/65536.0,1,-nbitq), 
to_sfixed(-2875.0/65536.0,1,-nbitq), 
to_sfixed(-495.0/65536.0,1,-nbitq), 
to_sfixed(745.0/65536.0,1,-nbitq), 
to_sfixed(-1532.0/65536.0,1,-nbitq), 
to_sfixed(-2937.0/65536.0,1,-nbitq), 
to_sfixed(1572.0/65536.0,1,-nbitq), 
to_sfixed(-1013.0/65536.0,1,-nbitq), 
to_sfixed(-817.0/65536.0,1,-nbitq), 
to_sfixed(-2398.0/65536.0,1,-nbitq), 
to_sfixed(2373.0/65536.0,1,-nbitq), 
to_sfixed(-4511.0/65536.0,1,-nbitq), 
to_sfixed(-4122.0/65536.0,1,-nbitq), 
to_sfixed(2934.0/65536.0,1,-nbitq), 
to_sfixed(1882.0/65536.0,1,-nbitq), 
to_sfixed(265.0/65536.0,1,-nbitq), 
to_sfixed(-839.0/65536.0,1,-nbitq), 
to_sfixed(1792.0/65536.0,1,-nbitq), 
to_sfixed(-489.0/65536.0,1,-nbitq), 
to_sfixed(5208.0/65536.0,1,-nbitq), 
to_sfixed(1200.0/65536.0,1,-nbitq), 
to_sfixed(2159.0/65536.0,1,-nbitq), 
to_sfixed(-1627.0/65536.0,1,-nbitq), 
to_sfixed(445.0/65536.0,1,-nbitq), 
to_sfixed(4602.0/65536.0,1,-nbitq), 
to_sfixed(1229.0/65536.0,1,-nbitq), 
to_sfixed(3940.0/65536.0,1,-nbitq), 
to_sfixed(4186.0/65536.0,1,-nbitq), 
to_sfixed(-1126.0/65536.0,1,-nbitq), 
to_sfixed(2180.0/65536.0,1,-nbitq), 
to_sfixed(2743.0/65536.0,1,-nbitq), 
to_sfixed(513.0/65536.0,1,-nbitq), 
to_sfixed(832.0/65536.0,1,-nbitq), 
to_sfixed(-1014.0/65536.0,1,-nbitq), 
to_sfixed(-3619.0/65536.0,1,-nbitq), 
to_sfixed(2503.0/65536.0,1,-nbitq), 
to_sfixed(4826.0/65536.0,1,-nbitq), 
to_sfixed(-280.0/65536.0,1,-nbitq), 
to_sfixed(342.0/65536.0,1,-nbitq), 
to_sfixed(-23.0/65536.0,1,-nbitq), 
to_sfixed(243.0/65536.0,1,-nbitq), 
to_sfixed(-3254.0/65536.0,1,-nbitq), 
to_sfixed(-1327.0/65536.0,1,-nbitq), 
to_sfixed(4361.0/65536.0,1,-nbitq), 
to_sfixed(-988.0/65536.0,1,-nbitq), 
to_sfixed(-335.0/65536.0,1,-nbitq), 
to_sfixed(7909.0/65536.0,1,-nbitq), 
to_sfixed(-6112.0/65536.0,1,-nbitq), 
to_sfixed(1688.0/65536.0,1,-nbitq), 
to_sfixed(3559.0/65536.0,1,-nbitq), 
to_sfixed(2701.0/65536.0,1,-nbitq), 
to_sfixed(738.0/65536.0,1,-nbitq), 
to_sfixed(1445.0/65536.0,1,-nbitq), 
to_sfixed(-11.0/65536.0,1,-nbitq), 
to_sfixed(-1965.0/65536.0,1,-nbitq), 
to_sfixed(-3071.0/65536.0,1,-nbitq), 
to_sfixed(-1322.0/65536.0,1,-nbitq), 
to_sfixed(1739.0/65536.0,1,-nbitq), 
to_sfixed(1987.0/65536.0,1,-nbitq), 
to_sfixed(-525.0/65536.0,1,-nbitq), 
to_sfixed(-2050.0/65536.0,1,-nbitq), 
to_sfixed(-1295.0/65536.0,1,-nbitq), 
to_sfixed(-6903.0/65536.0,1,-nbitq), 
to_sfixed(-5946.0/65536.0,1,-nbitq), 
to_sfixed(5876.0/65536.0,1,-nbitq), 
to_sfixed(-4803.0/65536.0,1,-nbitq), 
to_sfixed(5843.0/65536.0,1,-nbitq), 
to_sfixed(-744.0/65536.0,1,-nbitq), 
to_sfixed(-411.0/65536.0,1,-nbitq), 
to_sfixed(2787.0/65536.0,1,-nbitq), 
to_sfixed(-571.0/65536.0,1,-nbitq), 
to_sfixed(1608.0/65536.0,1,-nbitq), 
to_sfixed(1295.0/65536.0,1,-nbitq), 
to_sfixed(-706.0/65536.0,1,-nbitq)  ), 
( to_sfixed(576.0/65536.0,1,-nbitq), 
to_sfixed(413.0/65536.0,1,-nbitq), 
to_sfixed(875.0/65536.0,1,-nbitq), 
to_sfixed(-1830.0/65536.0,1,-nbitq), 
to_sfixed(1346.0/65536.0,1,-nbitq), 
to_sfixed(-2633.0/65536.0,1,-nbitq), 
to_sfixed(-1733.0/65536.0,1,-nbitq), 
to_sfixed(2324.0/65536.0,1,-nbitq), 
to_sfixed(648.0/65536.0,1,-nbitq), 
to_sfixed(-1838.0/65536.0,1,-nbitq), 
to_sfixed(1052.0/65536.0,1,-nbitq), 
to_sfixed(3226.0/65536.0,1,-nbitq), 
to_sfixed(-1151.0/65536.0,1,-nbitq), 
to_sfixed(-1903.0/65536.0,1,-nbitq), 
to_sfixed(-565.0/65536.0,1,-nbitq), 
to_sfixed(836.0/65536.0,1,-nbitq), 
to_sfixed(-1813.0/65536.0,1,-nbitq), 
to_sfixed(244.0/65536.0,1,-nbitq), 
to_sfixed(607.0/65536.0,1,-nbitq), 
to_sfixed(-2090.0/65536.0,1,-nbitq), 
to_sfixed(-539.0/65536.0,1,-nbitq), 
to_sfixed(-1345.0/65536.0,1,-nbitq), 
to_sfixed(-3279.0/65536.0,1,-nbitq), 
to_sfixed(-50.0/65536.0,1,-nbitq), 
to_sfixed(4400.0/65536.0,1,-nbitq), 
to_sfixed(-1129.0/65536.0,1,-nbitq), 
to_sfixed(392.0/65536.0,1,-nbitq), 
to_sfixed(1821.0/65536.0,1,-nbitq), 
to_sfixed(-1655.0/65536.0,1,-nbitq), 
to_sfixed(-599.0/65536.0,1,-nbitq), 
to_sfixed(-846.0/65536.0,1,-nbitq), 
to_sfixed(1917.0/65536.0,1,-nbitq), 
to_sfixed(276.0/65536.0,1,-nbitq), 
to_sfixed(880.0/65536.0,1,-nbitq), 
to_sfixed(2473.0/65536.0,1,-nbitq), 
to_sfixed(-3011.0/65536.0,1,-nbitq), 
to_sfixed(-739.0/65536.0,1,-nbitq), 
to_sfixed(-3011.0/65536.0,1,-nbitq), 
to_sfixed(-3362.0/65536.0,1,-nbitq), 
to_sfixed(-1884.0/65536.0,1,-nbitq), 
to_sfixed(-2262.0/65536.0,1,-nbitq), 
to_sfixed(-1195.0/65536.0,1,-nbitq), 
to_sfixed(1801.0/65536.0,1,-nbitq), 
to_sfixed(3525.0/65536.0,1,-nbitq), 
to_sfixed(1158.0/65536.0,1,-nbitq), 
to_sfixed(1349.0/65536.0,1,-nbitq), 
to_sfixed(-2521.0/65536.0,1,-nbitq), 
to_sfixed(994.0/65536.0,1,-nbitq), 
to_sfixed(1641.0/65536.0,1,-nbitq), 
to_sfixed(-1000.0/65536.0,1,-nbitq), 
to_sfixed(-579.0/65536.0,1,-nbitq), 
to_sfixed(-1468.0/65536.0,1,-nbitq), 
to_sfixed(3081.0/65536.0,1,-nbitq), 
to_sfixed(-5840.0/65536.0,1,-nbitq), 
to_sfixed(861.0/65536.0,1,-nbitq), 
to_sfixed(2098.0/65536.0,1,-nbitq), 
to_sfixed(372.0/65536.0,1,-nbitq), 
to_sfixed(-417.0/65536.0,1,-nbitq), 
to_sfixed(925.0/65536.0,1,-nbitq), 
to_sfixed(3521.0/65536.0,1,-nbitq), 
to_sfixed(188.0/65536.0,1,-nbitq), 
to_sfixed(2514.0/65536.0,1,-nbitq), 
to_sfixed(2706.0/65536.0,1,-nbitq), 
to_sfixed(-1109.0/65536.0,1,-nbitq), 
to_sfixed(-1728.0/65536.0,1,-nbitq), 
to_sfixed(-285.0/65536.0,1,-nbitq), 
to_sfixed(1692.0/65536.0,1,-nbitq), 
to_sfixed(-1547.0/65536.0,1,-nbitq), 
to_sfixed(-929.0/65536.0,1,-nbitq), 
to_sfixed(1446.0/65536.0,1,-nbitq), 
to_sfixed(473.0/65536.0,1,-nbitq), 
to_sfixed(-1942.0/65536.0,1,-nbitq), 
to_sfixed(-1738.0/65536.0,1,-nbitq), 
to_sfixed(2566.0/65536.0,1,-nbitq), 
to_sfixed(1803.0/65536.0,1,-nbitq), 
to_sfixed(1616.0/65536.0,1,-nbitq), 
to_sfixed(-735.0/65536.0,1,-nbitq), 
to_sfixed(587.0/65536.0,1,-nbitq), 
to_sfixed(-3095.0/65536.0,1,-nbitq), 
to_sfixed(3029.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2852.0/65536.0,1,-nbitq), 
to_sfixed(1786.0/65536.0,1,-nbitq), 
to_sfixed(1956.0/65536.0,1,-nbitq), 
to_sfixed(249.0/65536.0,1,-nbitq), 
to_sfixed(-754.0/65536.0,1,-nbitq), 
to_sfixed(1633.0/65536.0,1,-nbitq), 
to_sfixed(-1372.0/65536.0,1,-nbitq), 
to_sfixed(2354.0/65536.0,1,-nbitq), 
to_sfixed(510.0/65536.0,1,-nbitq), 
to_sfixed(-1422.0/65536.0,1,-nbitq), 
to_sfixed(-3758.0/65536.0,1,-nbitq), 
to_sfixed(-1750.0/65536.0,1,-nbitq), 
to_sfixed(959.0/65536.0,1,-nbitq), 
to_sfixed(-1875.0/65536.0,1,-nbitq), 
to_sfixed(-1211.0/65536.0,1,-nbitq), 
to_sfixed(1594.0/65536.0,1,-nbitq), 
to_sfixed(206.0/65536.0,1,-nbitq), 
to_sfixed(3323.0/65536.0,1,-nbitq), 
to_sfixed(-329.0/65536.0,1,-nbitq), 
to_sfixed(-197.0/65536.0,1,-nbitq), 
to_sfixed(122.0/65536.0,1,-nbitq), 
to_sfixed(3639.0/65536.0,1,-nbitq), 
to_sfixed(-1636.0/65536.0,1,-nbitq), 
to_sfixed(1379.0/65536.0,1,-nbitq), 
to_sfixed(3252.0/65536.0,1,-nbitq), 
to_sfixed(2681.0/65536.0,1,-nbitq), 
to_sfixed(-2663.0/65536.0,1,-nbitq), 
to_sfixed(-1958.0/65536.0,1,-nbitq), 
to_sfixed(-646.0/65536.0,1,-nbitq), 
to_sfixed(-762.0/65536.0,1,-nbitq), 
to_sfixed(-1611.0/65536.0,1,-nbitq), 
to_sfixed(-93.0/65536.0,1,-nbitq), 
to_sfixed(894.0/65536.0,1,-nbitq), 
to_sfixed(-1764.0/65536.0,1,-nbitq), 
to_sfixed(-145.0/65536.0,1,-nbitq), 
to_sfixed(-2588.0/65536.0,1,-nbitq), 
to_sfixed(-3570.0/65536.0,1,-nbitq), 
to_sfixed(-2244.0/65536.0,1,-nbitq), 
to_sfixed(-626.0/65536.0,1,-nbitq), 
to_sfixed(487.0/65536.0,1,-nbitq), 
to_sfixed(-950.0/65536.0,1,-nbitq), 
to_sfixed(-3140.0/65536.0,1,-nbitq), 
to_sfixed(-905.0/65536.0,1,-nbitq), 
to_sfixed(1574.0/65536.0,1,-nbitq), 
to_sfixed(632.0/65536.0,1,-nbitq), 
to_sfixed(4747.0/65536.0,1,-nbitq), 
to_sfixed(1411.0/65536.0,1,-nbitq), 
to_sfixed(2110.0/65536.0,1,-nbitq), 
to_sfixed(1994.0/65536.0,1,-nbitq), 
to_sfixed(-186.0/65536.0,1,-nbitq), 
to_sfixed(2827.0/65536.0,1,-nbitq), 
to_sfixed(-910.0/65536.0,1,-nbitq), 
to_sfixed(345.0/65536.0,1,-nbitq), 
to_sfixed(761.0/65536.0,1,-nbitq), 
to_sfixed(3972.0/65536.0,1,-nbitq), 
to_sfixed(-1365.0/65536.0,1,-nbitq), 
to_sfixed(1770.0/65536.0,1,-nbitq), 
to_sfixed(-63.0/65536.0,1,-nbitq), 
to_sfixed(-818.0/65536.0,1,-nbitq), 
to_sfixed(1062.0/65536.0,1,-nbitq), 
to_sfixed(-2928.0/65536.0,1,-nbitq), 
to_sfixed(-2870.0/65536.0,1,-nbitq), 
to_sfixed(-89.0/65536.0,1,-nbitq), 
to_sfixed(2236.0/65536.0,1,-nbitq), 
to_sfixed(71.0/65536.0,1,-nbitq), 
to_sfixed(-1813.0/65536.0,1,-nbitq), 
to_sfixed(676.0/65536.0,1,-nbitq), 
to_sfixed(491.0/65536.0,1,-nbitq), 
to_sfixed(-822.0/65536.0,1,-nbitq), 
to_sfixed(430.0/65536.0,1,-nbitq), 
to_sfixed(-1954.0/65536.0,1,-nbitq), 
to_sfixed(-3026.0/65536.0,1,-nbitq), 
to_sfixed(3256.0/65536.0,1,-nbitq), 
to_sfixed(-335.0/65536.0,1,-nbitq), 
to_sfixed(438.0/65536.0,1,-nbitq), 
to_sfixed(981.0/65536.0,1,-nbitq), 
to_sfixed(-1137.0/65536.0,1,-nbitq), 
to_sfixed(3290.0/65536.0,1,-nbitq), 
to_sfixed(-2985.0/65536.0,1,-nbitq), 
to_sfixed(-1889.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1579.0/65536.0,1,-nbitq), 
to_sfixed(-902.0/65536.0,1,-nbitq), 
to_sfixed(-1725.0/65536.0,1,-nbitq), 
to_sfixed(2082.0/65536.0,1,-nbitq), 
to_sfixed(976.0/65536.0,1,-nbitq), 
to_sfixed(-2832.0/65536.0,1,-nbitq), 
to_sfixed(-637.0/65536.0,1,-nbitq), 
to_sfixed(-2069.0/65536.0,1,-nbitq), 
to_sfixed(-3438.0/65536.0,1,-nbitq), 
to_sfixed(-419.0/65536.0,1,-nbitq), 
to_sfixed(-2530.0/65536.0,1,-nbitq), 
to_sfixed(2463.0/65536.0,1,-nbitq), 
to_sfixed(-2101.0/65536.0,1,-nbitq), 
to_sfixed(637.0/65536.0,1,-nbitq), 
to_sfixed(2434.0/65536.0,1,-nbitq), 
to_sfixed(1129.0/65536.0,1,-nbitq), 
to_sfixed(1501.0/65536.0,1,-nbitq), 
to_sfixed(2882.0/65536.0,1,-nbitq), 
to_sfixed(1903.0/65536.0,1,-nbitq), 
to_sfixed(1107.0/65536.0,1,-nbitq), 
to_sfixed(-3695.0/65536.0,1,-nbitq), 
to_sfixed(524.0/65536.0,1,-nbitq), 
to_sfixed(40.0/65536.0,1,-nbitq), 
to_sfixed(1721.0/65536.0,1,-nbitq), 
to_sfixed(-95.0/65536.0,1,-nbitq), 
to_sfixed(2753.0/65536.0,1,-nbitq), 
to_sfixed(-1622.0/65536.0,1,-nbitq), 
to_sfixed(856.0/65536.0,1,-nbitq), 
to_sfixed(-1915.0/65536.0,1,-nbitq), 
to_sfixed(1922.0/65536.0,1,-nbitq), 
to_sfixed(170.0/65536.0,1,-nbitq), 
to_sfixed(193.0/65536.0,1,-nbitq), 
to_sfixed(-3106.0/65536.0,1,-nbitq), 
to_sfixed(-2252.0/65536.0,1,-nbitq), 
to_sfixed(-2167.0/65536.0,1,-nbitq), 
to_sfixed(-2796.0/65536.0,1,-nbitq), 
to_sfixed(-2617.0/65536.0,1,-nbitq), 
to_sfixed(-1685.0/65536.0,1,-nbitq), 
to_sfixed(-3538.0/65536.0,1,-nbitq), 
to_sfixed(1071.0/65536.0,1,-nbitq), 
to_sfixed(-2918.0/65536.0,1,-nbitq), 
to_sfixed(1969.0/65536.0,1,-nbitq), 
to_sfixed(-79.0/65536.0,1,-nbitq), 
to_sfixed(448.0/65536.0,1,-nbitq), 
to_sfixed(-114.0/65536.0,1,-nbitq), 
to_sfixed(5267.0/65536.0,1,-nbitq), 
to_sfixed(-1686.0/65536.0,1,-nbitq), 
to_sfixed(163.0/65536.0,1,-nbitq), 
to_sfixed(2690.0/65536.0,1,-nbitq), 
to_sfixed(-185.0/65536.0,1,-nbitq), 
to_sfixed(-338.0/65536.0,1,-nbitq), 
to_sfixed(-3104.0/65536.0,1,-nbitq), 
to_sfixed(2606.0/65536.0,1,-nbitq), 
to_sfixed(-3192.0/65536.0,1,-nbitq), 
to_sfixed(1298.0/65536.0,1,-nbitq), 
to_sfixed(347.0/65536.0,1,-nbitq), 
to_sfixed(403.0/65536.0,1,-nbitq), 
to_sfixed(-105.0/65536.0,1,-nbitq), 
to_sfixed(152.0/65536.0,1,-nbitq), 
to_sfixed(1499.0/65536.0,1,-nbitq), 
to_sfixed(-1636.0/65536.0,1,-nbitq), 
to_sfixed(-1920.0/65536.0,1,-nbitq), 
to_sfixed(-1772.0/65536.0,1,-nbitq), 
to_sfixed(598.0/65536.0,1,-nbitq), 
to_sfixed(617.0/65536.0,1,-nbitq), 
to_sfixed(-1837.0/65536.0,1,-nbitq), 
to_sfixed(2762.0/65536.0,1,-nbitq), 
to_sfixed(-2399.0/65536.0,1,-nbitq), 
to_sfixed(-1378.0/65536.0,1,-nbitq), 
to_sfixed(2682.0/65536.0,1,-nbitq), 
to_sfixed(-2570.0/65536.0,1,-nbitq), 
to_sfixed(-3646.0/65536.0,1,-nbitq), 
to_sfixed(3047.0/65536.0,1,-nbitq), 
to_sfixed(-2905.0/65536.0,1,-nbitq), 
to_sfixed(-1568.0/65536.0,1,-nbitq), 
to_sfixed(-74.0/65536.0,1,-nbitq), 
to_sfixed(-2233.0/65536.0,1,-nbitq), 
to_sfixed(1272.0/65536.0,1,-nbitq), 
to_sfixed(-2963.0/65536.0,1,-nbitq), 
to_sfixed(-30.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2580.0/65536.0,1,-nbitq), 
to_sfixed(-2498.0/65536.0,1,-nbitq), 
to_sfixed(-251.0/65536.0,1,-nbitq), 
to_sfixed(-2801.0/65536.0,1,-nbitq), 
to_sfixed(-348.0/65536.0,1,-nbitq), 
to_sfixed(849.0/65536.0,1,-nbitq), 
to_sfixed(2103.0/65536.0,1,-nbitq), 
to_sfixed(-1993.0/65536.0,1,-nbitq), 
to_sfixed(-2914.0/65536.0,1,-nbitq), 
to_sfixed(-2616.0/65536.0,1,-nbitq), 
to_sfixed(-1880.0/65536.0,1,-nbitq), 
to_sfixed(3239.0/65536.0,1,-nbitq), 
to_sfixed(2529.0/65536.0,1,-nbitq), 
to_sfixed(-1206.0/65536.0,1,-nbitq), 
to_sfixed(333.0/65536.0,1,-nbitq), 
to_sfixed(281.0/65536.0,1,-nbitq), 
to_sfixed(-60.0/65536.0,1,-nbitq), 
to_sfixed(-1559.0/65536.0,1,-nbitq), 
to_sfixed(2526.0/65536.0,1,-nbitq), 
to_sfixed(-2482.0/65536.0,1,-nbitq), 
to_sfixed(1337.0/65536.0,1,-nbitq), 
to_sfixed(-2562.0/65536.0,1,-nbitq), 
to_sfixed(-1474.0/65536.0,1,-nbitq), 
to_sfixed(-631.0/65536.0,1,-nbitq), 
to_sfixed(-2775.0/65536.0,1,-nbitq), 
to_sfixed(-1773.0/65536.0,1,-nbitq), 
to_sfixed(-2133.0/65536.0,1,-nbitq), 
to_sfixed(-1737.0/65536.0,1,-nbitq), 
to_sfixed(-3973.0/65536.0,1,-nbitq), 
to_sfixed(-2244.0/65536.0,1,-nbitq), 
to_sfixed(-2650.0/65536.0,1,-nbitq), 
to_sfixed(1271.0/65536.0,1,-nbitq), 
to_sfixed(-4737.0/65536.0,1,-nbitq), 
to_sfixed(-592.0/65536.0,1,-nbitq), 
to_sfixed(-1594.0/65536.0,1,-nbitq), 
to_sfixed(-1543.0/65536.0,1,-nbitq), 
to_sfixed(2078.0/65536.0,1,-nbitq), 
to_sfixed(-2629.0/65536.0,1,-nbitq), 
to_sfixed(-2899.0/65536.0,1,-nbitq), 
to_sfixed(2077.0/65536.0,1,-nbitq), 
to_sfixed(-2255.0/65536.0,1,-nbitq), 
to_sfixed(1426.0/65536.0,1,-nbitq), 
to_sfixed(254.0/65536.0,1,-nbitq), 
to_sfixed(-749.0/65536.0,1,-nbitq), 
to_sfixed(2373.0/65536.0,1,-nbitq), 
to_sfixed(4946.0/65536.0,1,-nbitq), 
to_sfixed(1528.0/65536.0,1,-nbitq), 
to_sfixed(-634.0/65536.0,1,-nbitq), 
to_sfixed(457.0/65536.0,1,-nbitq), 
to_sfixed(2529.0/65536.0,1,-nbitq), 
to_sfixed(1899.0/65536.0,1,-nbitq), 
to_sfixed(2565.0/65536.0,1,-nbitq), 
to_sfixed(-963.0/65536.0,1,-nbitq), 
to_sfixed(-1210.0/65536.0,1,-nbitq), 
to_sfixed(2802.0/65536.0,1,-nbitq), 
to_sfixed(915.0/65536.0,1,-nbitq), 
to_sfixed(-2538.0/65536.0,1,-nbitq), 
to_sfixed(-670.0/65536.0,1,-nbitq), 
to_sfixed(336.0/65536.0,1,-nbitq), 
to_sfixed(5179.0/65536.0,1,-nbitq), 
to_sfixed(137.0/65536.0,1,-nbitq), 
to_sfixed(2602.0/65536.0,1,-nbitq), 
to_sfixed(-479.0/65536.0,1,-nbitq), 
to_sfixed(-18.0/65536.0,1,-nbitq), 
to_sfixed(-365.0/65536.0,1,-nbitq), 
to_sfixed(-744.0/65536.0,1,-nbitq), 
to_sfixed(1464.0/65536.0,1,-nbitq), 
to_sfixed(-1769.0/65536.0,1,-nbitq), 
to_sfixed(-2236.0/65536.0,1,-nbitq), 
to_sfixed(5057.0/65536.0,1,-nbitq), 
to_sfixed(-1348.0/65536.0,1,-nbitq), 
to_sfixed(-2029.0/65536.0,1,-nbitq), 
to_sfixed(3218.0/65536.0,1,-nbitq), 
to_sfixed(-2901.0/65536.0,1,-nbitq), 
to_sfixed(-2003.0/65536.0,1,-nbitq), 
to_sfixed(-819.0/65536.0,1,-nbitq), 
to_sfixed(-3006.0/65536.0,1,-nbitq), 
to_sfixed(3177.0/65536.0,1,-nbitq), 
to_sfixed(-3036.0/65536.0,1,-nbitq), 
to_sfixed(2695.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-890.0/65536.0,1,-nbitq), 
to_sfixed(2803.0/65536.0,1,-nbitq), 
to_sfixed(705.0/65536.0,1,-nbitq), 
to_sfixed(-3411.0/65536.0,1,-nbitq), 
to_sfixed(-1903.0/65536.0,1,-nbitq), 
to_sfixed(-3286.0/65536.0,1,-nbitq), 
to_sfixed(2142.0/65536.0,1,-nbitq), 
to_sfixed(-1294.0/65536.0,1,-nbitq), 
to_sfixed(-865.0/65536.0,1,-nbitq), 
to_sfixed(247.0/65536.0,1,-nbitq), 
to_sfixed(-756.0/65536.0,1,-nbitq), 
to_sfixed(294.0/65536.0,1,-nbitq), 
to_sfixed(-101.0/65536.0,1,-nbitq), 
to_sfixed(-358.0/65536.0,1,-nbitq), 
to_sfixed(5.0/65536.0,1,-nbitq), 
to_sfixed(3169.0/65536.0,1,-nbitq), 
to_sfixed(1331.0/65536.0,1,-nbitq), 
to_sfixed(1403.0/65536.0,1,-nbitq), 
to_sfixed(1333.0/65536.0,1,-nbitq), 
to_sfixed(150.0/65536.0,1,-nbitq), 
to_sfixed(-274.0/65536.0,1,-nbitq), 
to_sfixed(-388.0/65536.0,1,-nbitq), 
to_sfixed(199.0/65536.0,1,-nbitq), 
to_sfixed(316.0/65536.0,1,-nbitq), 
to_sfixed(2635.0/65536.0,1,-nbitq), 
to_sfixed(-716.0/65536.0,1,-nbitq), 
to_sfixed(-1165.0/65536.0,1,-nbitq), 
to_sfixed(807.0/65536.0,1,-nbitq), 
to_sfixed(-4512.0/65536.0,1,-nbitq), 
to_sfixed(-680.0/65536.0,1,-nbitq), 
to_sfixed(-700.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(254.0/65536.0,1,-nbitq), 
to_sfixed(-441.0/65536.0,1,-nbitq), 
to_sfixed(-2218.0/65536.0,1,-nbitq), 
to_sfixed(-1897.0/65536.0,1,-nbitq), 
to_sfixed(-2806.0/65536.0,1,-nbitq), 
to_sfixed(1642.0/65536.0,1,-nbitq), 
to_sfixed(-3024.0/65536.0,1,-nbitq), 
to_sfixed(1189.0/65536.0,1,-nbitq), 
to_sfixed(-547.0/65536.0,1,-nbitq), 
to_sfixed(1438.0/65536.0,1,-nbitq), 
to_sfixed(69.0/65536.0,1,-nbitq), 
to_sfixed(1908.0/65536.0,1,-nbitq), 
to_sfixed(971.0/65536.0,1,-nbitq), 
to_sfixed(-240.0/65536.0,1,-nbitq), 
to_sfixed(-2016.0/65536.0,1,-nbitq), 
to_sfixed(-699.0/65536.0,1,-nbitq), 
to_sfixed(2077.0/65536.0,1,-nbitq), 
to_sfixed(3233.0/65536.0,1,-nbitq), 
to_sfixed(-520.0/65536.0,1,-nbitq), 
to_sfixed(-2829.0/65536.0,1,-nbitq), 
to_sfixed(124.0/65536.0,1,-nbitq), 
to_sfixed(-442.0/65536.0,1,-nbitq), 
to_sfixed(-1614.0/65536.0,1,-nbitq), 
to_sfixed(763.0/65536.0,1,-nbitq), 
to_sfixed(-556.0/65536.0,1,-nbitq), 
to_sfixed(-617.0/65536.0,1,-nbitq), 
to_sfixed(871.0/65536.0,1,-nbitq), 
to_sfixed(1525.0/65536.0,1,-nbitq), 
to_sfixed(1314.0/65536.0,1,-nbitq), 
to_sfixed(1331.0/65536.0,1,-nbitq), 
to_sfixed(-2706.0/65536.0,1,-nbitq), 
to_sfixed(1715.0/65536.0,1,-nbitq), 
to_sfixed(1420.0/65536.0,1,-nbitq), 
to_sfixed(-1623.0/65536.0,1,-nbitq), 
to_sfixed(1330.0/65536.0,1,-nbitq), 
to_sfixed(-2857.0/65536.0,1,-nbitq), 
to_sfixed(-355.0/65536.0,1,-nbitq), 
to_sfixed(1322.0/65536.0,1,-nbitq), 
to_sfixed(2483.0/65536.0,1,-nbitq), 
to_sfixed(1376.0/65536.0,1,-nbitq), 
to_sfixed(248.0/65536.0,1,-nbitq), 
to_sfixed(-1512.0/65536.0,1,-nbitq), 
to_sfixed(1354.0/65536.0,1,-nbitq), 
to_sfixed(428.0/65536.0,1,-nbitq), 
to_sfixed(-662.0/65536.0,1,-nbitq), 
to_sfixed(4524.0/65536.0,1,-nbitq), 
to_sfixed(2724.0/65536.0,1,-nbitq), 
to_sfixed(2494.0/65536.0,1,-nbitq)  ), 
( to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(-2781.0/65536.0,1,-nbitq), 
to_sfixed(702.0/65536.0,1,-nbitq), 
to_sfixed(-1847.0/65536.0,1,-nbitq), 
to_sfixed(173.0/65536.0,1,-nbitq), 
to_sfixed(-5284.0/65536.0,1,-nbitq), 
to_sfixed(1061.0/65536.0,1,-nbitq), 
to_sfixed(271.0/65536.0,1,-nbitq), 
to_sfixed(-2309.0/65536.0,1,-nbitq), 
to_sfixed(1628.0/65536.0,1,-nbitq), 
to_sfixed(-1683.0/65536.0,1,-nbitq), 
to_sfixed(-359.0/65536.0,1,-nbitq), 
to_sfixed(-180.0/65536.0,1,-nbitq), 
to_sfixed(1510.0/65536.0,1,-nbitq), 
to_sfixed(-528.0/65536.0,1,-nbitq), 
to_sfixed(1756.0/65536.0,1,-nbitq), 
to_sfixed(1676.0/65536.0,1,-nbitq), 
to_sfixed(-3224.0/65536.0,1,-nbitq), 
to_sfixed(1021.0/65536.0,1,-nbitq), 
to_sfixed(1229.0/65536.0,1,-nbitq), 
to_sfixed(1080.0/65536.0,1,-nbitq), 
to_sfixed(-3094.0/65536.0,1,-nbitq), 
to_sfixed(3908.0/65536.0,1,-nbitq), 
to_sfixed(1089.0/65536.0,1,-nbitq), 
to_sfixed(2151.0/65536.0,1,-nbitq), 
to_sfixed(-449.0/65536.0,1,-nbitq), 
to_sfixed(-3621.0/65536.0,1,-nbitq), 
to_sfixed(1226.0/65536.0,1,-nbitq), 
to_sfixed(-3280.0/65536.0,1,-nbitq), 
to_sfixed(-3902.0/65536.0,1,-nbitq), 
to_sfixed(3023.0/65536.0,1,-nbitq), 
to_sfixed(2710.0/65536.0,1,-nbitq), 
to_sfixed(-1524.0/65536.0,1,-nbitq), 
to_sfixed(1854.0/65536.0,1,-nbitq), 
to_sfixed(-1169.0/65536.0,1,-nbitq), 
to_sfixed(1829.0/65536.0,1,-nbitq), 
to_sfixed(379.0/65536.0,1,-nbitq), 
to_sfixed(-1941.0/65536.0,1,-nbitq), 
to_sfixed(-326.0/65536.0,1,-nbitq), 
to_sfixed(-2328.0/65536.0,1,-nbitq), 
to_sfixed(-456.0/65536.0,1,-nbitq), 
to_sfixed(-1721.0/65536.0,1,-nbitq), 
to_sfixed(-4148.0/65536.0,1,-nbitq), 
to_sfixed(2691.0/65536.0,1,-nbitq), 
to_sfixed(2892.0/65536.0,1,-nbitq), 
to_sfixed(4650.0/65536.0,1,-nbitq), 
to_sfixed(-927.0/65536.0,1,-nbitq), 
to_sfixed(411.0/65536.0,1,-nbitq), 
to_sfixed(265.0/65536.0,1,-nbitq), 
to_sfixed(2423.0/65536.0,1,-nbitq), 
to_sfixed(-1279.0/65536.0,1,-nbitq), 
to_sfixed(2515.0/65536.0,1,-nbitq), 
to_sfixed(3440.0/65536.0,1,-nbitq), 
to_sfixed(-2310.0/65536.0,1,-nbitq), 
to_sfixed(2123.0/65536.0,1,-nbitq), 
to_sfixed(-1701.0/65536.0,1,-nbitq), 
to_sfixed(597.0/65536.0,1,-nbitq), 
to_sfixed(2053.0/65536.0,1,-nbitq), 
to_sfixed(405.0/65536.0,1,-nbitq), 
to_sfixed(2140.0/65536.0,1,-nbitq), 
to_sfixed(-2355.0/65536.0,1,-nbitq), 
to_sfixed(-1144.0/65536.0,1,-nbitq), 
to_sfixed(-1555.0/65536.0,1,-nbitq), 
to_sfixed(44.0/65536.0,1,-nbitq), 
to_sfixed(4076.0/65536.0,1,-nbitq), 
to_sfixed(-1995.0/65536.0,1,-nbitq), 
to_sfixed(-2327.0/65536.0,1,-nbitq), 
to_sfixed(-1204.0/65536.0,1,-nbitq), 
to_sfixed(-1607.0/65536.0,1,-nbitq), 
to_sfixed(5259.0/65536.0,1,-nbitq), 
to_sfixed(1366.0/65536.0,1,-nbitq), 
to_sfixed(-3030.0/65536.0,1,-nbitq), 
to_sfixed(-941.0/65536.0,1,-nbitq), 
to_sfixed(1465.0/65536.0,1,-nbitq), 
to_sfixed(2152.0/65536.0,1,-nbitq), 
to_sfixed(-2341.0/65536.0,1,-nbitq), 
to_sfixed(2195.0/65536.0,1,-nbitq), 
to_sfixed(3948.0/65536.0,1,-nbitq), 
to_sfixed(-2039.0/65536.0,1,-nbitq), 
to_sfixed(304.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1506.0/65536.0,1,-nbitq), 
to_sfixed(184.0/65536.0,1,-nbitq), 
to_sfixed(-3756.0/65536.0,1,-nbitq), 
to_sfixed(-586.0/65536.0,1,-nbitq), 
to_sfixed(2048.0/65536.0,1,-nbitq), 
to_sfixed(-771.0/65536.0,1,-nbitq), 
to_sfixed(-1389.0/65536.0,1,-nbitq), 
to_sfixed(-1952.0/65536.0,1,-nbitq), 
to_sfixed(-1934.0/65536.0,1,-nbitq), 
to_sfixed(1953.0/65536.0,1,-nbitq), 
to_sfixed(1026.0/65536.0,1,-nbitq), 
to_sfixed(742.0/65536.0,1,-nbitq), 
to_sfixed(-245.0/65536.0,1,-nbitq), 
to_sfixed(1645.0/65536.0,1,-nbitq), 
to_sfixed(628.0/65536.0,1,-nbitq), 
to_sfixed(1841.0/65536.0,1,-nbitq), 
to_sfixed(-1834.0/65536.0,1,-nbitq), 
to_sfixed(-2380.0/65536.0,1,-nbitq), 
to_sfixed(-596.0/65536.0,1,-nbitq), 
to_sfixed(580.0/65536.0,1,-nbitq), 
to_sfixed(820.0/65536.0,1,-nbitq), 
to_sfixed(-1084.0/65536.0,1,-nbitq), 
to_sfixed(551.0/65536.0,1,-nbitq), 
to_sfixed(259.0/65536.0,1,-nbitq), 
to_sfixed(271.0/65536.0,1,-nbitq), 
to_sfixed(-2142.0/65536.0,1,-nbitq), 
to_sfixed(-3521.0/65536.0,1,-nbitq), 
to_sfixed(1126.0/65536.0,1,-nbitq), 
to_sfixed(-3544.0/65536.0,1,-nbitq), 
to_sfixed(-1053.0/65536.0,1,-nbitq), 
to_sfixed(-1519.0/65536.0,1,-nbitq), 
to_sfixed(-53.0/65536.0,1,-nbitq), 
to_sfixed(-1234.0/65536.0,1,-nbitq), 
to_sfixed(7009.0/65536.0,1,-nbitq), 
to_sfixed(1166.0/65536.0,1,-nbitq), 
to_sfixed(-2066.0/65536.0,1,-nbitq), 
to_sfixed(2473.0/65536.0,1,-nbitq), 
to_sfixed(2474.0/65536.0,1,-nbitq), 
to_sfixed(3900.0/65536.0,1,-nbitq), 
to_sfixed(-3297.0/65536.0,1,-nbitq), 
to_sfixed(184.0/65536.0,1,-nbitq), 
to_sfixed(2258.0/65536.0,1,-nbitq), 
to_sfixed(112.0/65536.0,1,-nbitq), 
to_sfixed(3470.0/65536.0,1,-nbitq), 
to_sfixed(497.0/65536.0,1,-nbitq), 
to_sfixed(762.0/65536.0,1,-nbitq), 
to_sfixed(-1438.0/65536.0,1,-nbitq), 
to_sfixed(-4236.0/65536.0,1,-nbitq), 
to_sfixed(3826.0/65536.0,1,-nbitq), 
to_sfixed(613.0/65536.0,1,-nbitq), 
to_sfixed(-1675.0/65536.0,1,-nbitq), 
to_sfixed(-6060.0/65536.0,1,-nbitq), 
to_sfixed(1264.0/65536.0,1,-nbitq), 
to_sfixed(-1130.0/65536.0,1,-nbitq), 
to_sfixed(-2060.0/65536.0,1,-nbitq), 
to_sfixed(1231.0/65536.0,1,-nbitq), 
to_sfixed(-1574.0/65536.0,1,-nbitq), 
to_sfixed(2565.0/65536.0,1,-nbitq), 
to_sfixed(-1760.0/65536.0,1,-nbitq), 
to_sfixed(133.0/65536.0,1,-nbitq), 
to_sfixed(-508.0/65536.0,1,-nbitq), 
to_sfixed(-3413.0/65536.0,1,-nbitq), 
to_sfixed(472.0/65536.0,1,-nbitq), 
to_sfixed(-1141.0/65536.0,1,-nbitq), 
to_sfixed(958.0/65536.0,1,-nbitq), 
to_sfixed(1959.0/65536.0,1,-nbitq), 
to_sfixed(-2485.0/65536.0,1,-nbitq), 
to_sfixed(2423.0/65536.0,1,-nbitq), 
to_sfixed(-5437.0/65536.0,1,-nbitq), 
to_sfixed(773.0/65536.0,1,-nbitq), 
to_sfixed(2430.0/65536.0,1,-nbitq), 
to_sfixed(1040.0/65536.0,1,-nbitq), 
to_sfixed(-1652.0/65536.0,1,-nbitq), 
to_sfixed(2633.0/65536.0,1,-nbitq), 
to_sfixed(-641.0/65536.0,1,-nbitq), 
to_sfixed(-1450.0/65536.0,1,-nbitq), 
to_sfixed(2851.0/65536.0,1,-nbitq), 
to_sfixed(1676.0/65536.0,1,-nbitq), 
to_sfixed(-3081.0/65536.0,1,-nbitq), 
to_sfixed(1600.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2887.0/65536.0,1,-nbitq), 
to_sfixed(49.0/65536.0,1,-nbitq), 
to_sfixed(-1720.0/65536.0,1,-nbitq), 
to_sfixed(-768.0/65536.0,1,-nbitq), 
to_sfixed(894.0/65536.0,1,-nbitq), 
to_sfixed(-828.0/65536.0,1,-nbitq), 
to_sfixed(94.0/65536.0,1,-nbitq), 
to_sfixed(715.0/65536.0,1,-nbitq), 
to_sfixed(3431.0/65536.0,1,-nbitq), 
to_sfixed(-2241.0/65536.0,1,-nbitq), 
to_sfixed(-3222.0/65536.0,1,-nbitq), 
to_sfixed(4724.0/65536.0,1,-nbitq), 
to_sfixed(-2077.0/65536.0,1,-nbitq), 
to_sfixed(2646.0/65536.0,1,-nbitq), 
to_sfixed(-2476.0/65536.0,1,-nbitq), 
to_sfixed(-857.0/65536.0,1,-nbitq), 
to_sfixed(737.0/65536.0,1,-nbitq), 
to_sfixed(-3161.0/65536.0,1,-nbitq), 
to_sfixed(-169.0/65536.0,1,-nbitq), 
to_sfixed(-686.0/65536.0,1,-nbitq), 
to_sfixed(711.0/65536.0,1,-nbitq), 
to_sfixed(-684.0/65536.0,1,-nbitq), 
to_sfixed(-922.0/65536.0,1,-nbitq), 
to_sfixed(-805.0/65536.0,1,-nbitq), 
to_sfixed(2320.0/65536.0,1,-nbitq), 
to_sfixed(7.0/65536.0,1,-nbitq), 
to_sfixed(2813.0/65536.0,1,-nbitq), 
to_sfixed(2531.0/65536.0,1,-nbitq), 
to_sfixed(-2967.0/65536.0,1,-nbitq), 
to_sfixed(-77.0/65536.0,1,-nbitq), 
to_sfixed(3860.0/65536.0,1,-nbitq), 
to_sfixed(2925.0/65536.0,1,-nbitq), 
to_sfixed(-144.0/65536.0,1,-nbitq), 
to_sfixed(10504.0/65536.0,1,-nbitq), 
to_sfixed(-539.0/65536.0,1,-nbitq), 
to_sfixed(-1168.0/65536.0,1,-nbitq), 
to_sfixed(-2778.0/65536.0,1,-nbitq), 
to_sfixed(2954.0/65536.0,1,-nbitq), 
to_sfixed(1691.0/65536.0,1,-nbitq), 
to_sfixed(-779.0/65536.0,1,-nbitq), 
to_sfixed(-8016.0/65536.0,1,-nbitq), 
to_sfixed(-1922.0/65536.0,1,-nbitq), 
to_sfixed(9568.0/65536.0,1,-nbitq), 
to_sfixed(1893.0/65536.0,1,-nbitq), 
to_sfixed(-894.0/65536.0,1,-nbitq), 
to_sfixed(1912.0/65536.0,1,-nbitq), 
to_sfixed(2714.0/65536.0,1,-nbitq), 
to_sfixed(-4227.0/65536.0,1,-nbitq), 
to_sfixed(1286.0/65536.0,1,-nbitq), 
to_sfixed(641.0/65536.0,1,-nbitq), 
to_sfixed(3127.0/65536.0,1,-nbitq), 
to_sfixed(-1831.0/65536.0,1,-nbitq), 
to_sfixed(-404.0/65536.0,1,-nbitq), 
to_sfixed(98.0/65536.0,1,-nbitq), 
to_sfixed(-1515.0/65536.0,1,-nbitq), 
to_sfixed(1756.0/65536.0,1,-nbitq), 
to_sfixed(1432.0/65536.0,1,-nbitq), 
to_sfixed(2992.0/65536.0,1,-nbitq), 
to_sfixed(-2017.0/65536.0,1,-nbitq), 
to_sfixed(2083.0/65536.0,1,-nbitq), 
to_sfixed(-2707.0/65536.0,1,-nbitq), 
to_sfixed(-2295.0/65536.0,1,-nbitq), 
to_sfixed(1850.0/65536.0,1,-nbitq), 
to_sfixed(-2772.0/65536.0,1,-nbitq), 
to_sfixed(-318.0/65536.0,1,-nbitq), 
to_sfixed(3021.0/65536.0,1,-nbitq), 
to_sfixed(-2564.0/65536.0,1,-nbitq), 
to_sfixed(1226.0/65536.0,1,-nbitq), 
to_sfixed(39.0/65536.0,1,-nbitq), 
to_sfixed(2622.0/65536.0,1,-nbitq), 
to_sfixed(2357.0/65536.0,1,-nbitq), 
to_sfixed(-2221.0/65536.0,1,-nbitq), 
to_sfixed(-3461.0/65536.0,1,-nbitq), 
to_sfixed(1131.0/65536.0,1,-nbitq), 
to_sfixed(-1960.0/65536.0,1,-nbitq), 
to_sfixed(1381.0/65536.0,1,-nbitq), 
to_sfixed(-301.0/65536.0,1,-nbitq), 
to_sfixed(-103.0/65536.0,1,-nbitq), 
to_sfixed(1969.0/65536.0,1,-nbitq), 
to_sfixed(-3278.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2359.0/65536.0,1,-nbitq), 
to_sfixed(-384.0/65536.0,1,-nbitq), 
to_sfixed(8792.0/65536.0,1,-nbitq), 
to_sfixed(712.0/65536.0,1,-nbitq), 
to_sfixed(-2730.0/65536.0,1,-nbitq), 
to_sfixed(269.0/65536.0,1,-nbitq), 
to_sfixed(2703.0/65536.0,1,-nbitq), 
to_sfixed(8135.0/65536.0,1,-nbitq), 
to_sfixed(662.0/65536.0,1,-nbitq), 
to_sfixed(3132.0/65536.0,1,-nbitq), 
to_sfixed(734.0/65536.0,1,-nbitq), 
to_sfixed(4065.0/65536.0,1,-nbitq), 
to_sfixed(-3291.0/65536.0,1,-nbitq), 
to_sfixed(6735.0/65536.0,1,-nbitq), 
to_sfixed(2403.0/65536.0,1,-nbitq), 
to_sfixed(785.0/65536.0,1,-nbitq), 
to_sfixed(-1472.0/65536.0,1,-nbitq), 
to_sfixed(-2113.0/65536.0,1,-nbitq), 
to_sfixed(5804.0/65536.0,1,-nbitq), 
to_sfixed(812.0/65536.0,1,-nbitq), 
to_sfixed(-3995.0/65536.0,1,-nbitq), 
to_sfixed(-2366.0/65536.0,1,-nbitq), 
to_sfixed(2856.0/65536.0,1,-nbitq), 
to_sfixed(-4409.0/65536.0,1,-nbitq), 
to_sfixed(-3446.0/65536.0,1,-nbitq), 
to_sfixed(1100.0/65536.0,1,-nbitq), 
to_sfixed(-828.0/65536.0,1,-nbitq), 
to_sfixed(1184.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(1829.0/65536.0,1,-nbitq), 
to_sfixed(-1008.0/65536.0,1,-nbitq), 
to_sfixed(5648.0/65536.0,1,-nbitq), 
to_sfixed(1674.0/65536.0,1,-nbitq), 
to_sfixed(10199.0/65536.0,1,-nbitq), 
to_sfixed(-4077.0/65536.0,1,-nbitq), 
to_sfixed(430.0/65536.0,1,-nbitq), 
to_sfixed(-8458.0/65536.0,1,-nbitq), 
to_sfixed(2872.0/65536.0,1,-nbitq), 
to_sfixed(-2835.0/65536.0,1,-nbitq), 
to_sfixed(-5445.0/65536.0,1,-nbitq), 
to_sfixed(-3823.0/65536.0,1,-nbitq), 
to_sfixed(-658.0/65536.0,1,-nbitq), 
to_sfixed(9321.0/65536.0,1,-nbitq), 
to_sfixed(-350.0/65536.0,1,-nbitq), 
to_sfixed(-71.0/65536.0,1,-nbitq), 
to_sfixed(-519.0/65536.0,1,-nbitq), 
to_sfixed(312.0/65536.0,1,-nbitq), 
to_sfixed(-1330.0/65536.0,1,-nbitq), 
to_sfixed(1541.0/65536.0,1,-nbitq), 
to_sfixed(3896.0/65536.0,1,-nbitq), 
to_sfixed(917.0/65536.0,1,-nbitq), 
to_sfixed(-4211.0/65536.0,1,-nbitq), 
to_sfixed(-648.0/65536.0,1,-nbitq), 
to_sfixed(8642.0/65536.0,1,-nbitq), 
to_sfixed(-5167.0/65536.0,1,-nbitq), 
to_sfixed(3246.0/65536.0,1,-nbitq), 
to_sfixed(1206.0/65536.0,1,-nbitq), 
to_sfixed(651.0/65536.0,1,-nbitq), 
to_sfixed(1571.0/65536.0,1,-nbitq), 
to_sfixed(656.0/65536.0,1,-nbitq), 
to_sfixed(-1439.0/65536.0,1,-nbitq), 
to_sfixed(1894.0/65536.0,1,-nbitq), 
to_sfixed(2527.0/65536.0,1,-nbitq), 
to_sfixed(1992.0/65536.0,1,-nbitq), 
to_sfixed(1625.0/65536.0,1,-nbitq), 
to_sfixed(-315.0/65536.0,1,-nbitq), 
to_sfixed(-3887.0/65536.0,1,-nbitq), 
to_sfixed(-3699.0/65536.0,1,-nbitq), 
to_sfixed(-4884.0/65536.0,1,-nbitq), 
to_sfixed(986.0/65536.0,1,-nbitq), 
to_sfixed(-2632.0/65536.0,1,-nbitq), 
to_sfixed(5580.0/65536.0,1,-nbitq), 
to_sfixed(-1333.0/65536.0,1,-nbitq), 
to_sfixed(1654.0/65536.0,1,-nbitq), 
to_sfixed(2151.0/65536.0,1,-nbitq), 
to_sfixed(3808.0/65536.0,1,-nbitq), 
to_sfixed(5510.0/65536.0,1,-nbitq), 
to_sfixed(-973.0/65536.0,1,-nbitq), 
to_sfixed(-2288.0/65536.0,1,-nbitq), 
to_sfixed(1220.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1330.0/65536.0,1,-nbitq), 
to_sfixed(-2649.0/65536.0,1,-nbitq), 
to_sfixed(8296.0/65536.0,1,-nbitq), 
to_sfixed(882.0/65536.0,1,-nbitq), 
to_sfixed(-2281.0/65536.0,1,-nbitq), 
to_sfixed(-542.0/65536.0,1,-nbitq), 
to_sfixed(4321.0/65536.0,1,-nbitq), 
to_sfixed(1953.0/65536.0,1,-nbitq), 
to_sfixed(821.0/65536.0,1,-nbitq), 
to_sfixed(375.0/65536.0,1,-nbitq), 
to_sfixed(5088.0/65536.0,1,-nbitq), 
to_sfixed(7179.0/65536.0,1,-nbitq), 
to_sfixed(1679.0/65536.0,1,-nbitq), 
to_sfixed(4704.0/65536.0,1,-nbitq), 
to_sfixed(-227.0/65536.0,1,-nbitq), 
to_sfixed(706.0/65536.0,1,-nbitq), 
to_sfixed(-1472.0/65536.0,1,-nbitq), 
to_sfixed(-3858.0/65536.0,1,-nbitq), 
to_sfixed(3285.0/65536.0,1,-nbitq), 
to_sfixed(219.0/65536.0,1,-nbitq), 
to_sfixed(-3256.0/65536.0,1,-nbitq), 
to_sfixed(381.0/65536.0,1,-nbitq), 
to_sfixed(2363.0/65536.0,1,-nbitq), 
to_sfixed(-6904.0/65536.0,1,-nbitq), 
to_sfixed(-793.0/65536.0,1,-nbitq), 
to_sfixed(2094.0/65536.0,1,-nbitq), 
to_sfixed(-11315.0/65536.0,1,-nbitq), 
to_sfixed(2112.0/65536.0,1,-nbitq), 
to_sfixed(337.0/65536.0,1,-nbitq), 
to_sfixed(496.0/65536.0,1,-nbitq), 
to_sfixed(1242.0/65536.0,1,-nbitq), 
to_sfixed(6626.0/65536.0,1,-nbitq), 
to_sfixed(-1979.0/65536.0,1,-nbitq), 
to_sfixed(6515.0/65536.0,1,-nbitq), 
to_sfixed(-2213.0/65536.0,1,-nbitq), 
to_sfixed(-1131.0/65536.0,1,-nbitq), 
to_sfixed(-3739.0/65536.0,1,-nbitq), 
to_sfixed(2262.0/65536.0,1,-nbitq), 
to_sfixed(2376.0/65536.0,1,-nbitq), 
to_sfixed(-2386.0/65536.0,1,-nbitq), 
to_sfixed(-5092.0/65536.0,1,-nbitq), 
to_sfixed(2415.0/65536.0,1,-nbitq), 
to_sfixed(9409.0/65536.0,1,-nbitq), 
to_sfixed(1793.0/65536.0,1,-nbitq), 
to_sfixed(755.0/65536.0,1,-nbitq), 
to_sfixed(-9174.0/65536.0,1,-nbitq), 
to_sfixed(-2734.0/65536.0,1,-nbitq), 
to_sfixed(-4498.0/65536.0,1,-nbitq), 
to_sfixed(1904.0/65536.0,1,-nbitq), 
to_sfixed(-149.0/65536.0,1,-nbitq), 
to_sfixed(2794.0/65536.0,1,-nbitq), 
to_sfixed(-6841.0/65536.0,1,-nbitq), 
to_sfixed(1185.0/65536.0,1,-nbitq), 
to_sfixed(2592.0/65536.0,1,-nbitq), 
to_sfixed(-3873.0/65536.0,1,-nbitq), 
to_sfixed(5007.0/65536.0,1,-nbitq), 
to_sfixed(-1651.0/65536.0,1,-nbitq), 
to_sfixed(1017.0/65536.0,1,-nbitq), 
to_sfixed(-1653.0/65536.0,1,-nbitq), 
to_sfixed(-4030.0/65536.0,1,-nbitq), 
to_sfixed(1148.0/65536.0,1,-nbitq), 
to_sfixed(2076.0/65536.0,1,-nbitq), 
to_sfixed(2465.0/65536.0,1,-nbitq), 
to_sfixed(-2721.0/65536.0,1,-nbitq), 
to_sfixed(4735.0/65536.0,1,-nbitq), 
to_sfixed(4205.0/65536.0,1,-nbitq), 
to_sfixed(-3878.0/65536.0,1,-nbitq), 
to_sfixed(-4867.0/65536.0,1,-nbitq), 
to_sfixed(2806.0/65536.0,1,-nbitq), 
to_sfixed(1736.0/65536.0,1,-nbitq), 
to_sfixed(709.0/65536.0,1,-nbitq), 
to_sfixed(4918.0/65536.0,1,-nbitq), 
to_sfixed(-690.0/65536.0,1,-nbitq), 
to_sfixed(-2751.0/65536.0,1,-nbitq), 
to_sfixed(-2481.0/65536.0,1,-nbitq), 
to_sfixed(2371.0/65536.0,1,-nbitq), 
to_sfixed(6932.0/65536.0,1,-nbitq), 
to_sfixed(-991.0/65536.0,1,-nbitq), 
to_sfixed(326.0/65536.0,1,-nbitq), 
to_sfixed(-1183.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3502.0/65536.0,1,-nbitq), 
to_sfixed(-2056.0/65536.0,1,-nbitq), 
to_sfixed(2089.0/65536.0,1,-nbitq), 
to_sfixed(-2386.0/65536.0,1,-nbitq), 
to_sfixed(-1631.0/65536.0,1,-nbitq), 
to_sfixed(-5838.0/65536.0,1,-nbitq), 
to_sfixed(772.0/65536.0,1,-nbitq), 
to_sfixed(1488.0/65536.0,1,-nbitq), 
to_sfixed(-1598.0/65536.0,1,-nbitq), 
to_sfixed(2845.0/65536.0,1,-nbitq), 
to_sfixed(4335.0/65536.0,1,-nbitq), 
to_sfixed(4375.0/65536.0,1,-nbitq), 
to_sfixed(1565.0/65536.0,1,-nbitq), 
to_sfixed(4542.0/65536.0,1,-nbitq), 
to_sfixed(2551.0/65536.0,1,-nbitq), 
to_sfixed(-1459.0/65536.0,1,-nbitq), 
to_sfixed(-2309.0/65536.0,1,-nbitq), 
to_sfixed(-1106.0/65536.0,1,-nbitq), 
to_sfixed(4045.0/65536.0,1,-nbitq), 
to_sfixed(-118.0/65536.0,1,-nbitq), 
to_sfixed(331.0/65536.0,1,-nbitq), 
to_sfixed(3489.0/65536.0,1,-nbitq), 
to_sfixed(1243.0/65536.0,1,-nbitq), 
to_sfixed(-5546.0/65536.0,1,-nbitq), 
to_sfixed(4202.0/65536.0,1,-nbitq), 
to_sfixed(-2167.0/65536.0,1,-nbitq), 
to_sfixed(-9452.0/65536.0,1,-nbitq), 
to_sfixed(-451.0/65536.0,1,-nbitq), 
to_sfixed(-3162.0/65536.0,1,-nbitq), 
to_sfixed(-6911.0/65536.0,1,-nbitq), 
to_sfixed(3651.0/65536.0,1,-nbitq), 
to_sfixed(4456.0/65536.0,1,-nbitq), 
to_sfixed(-4978.0/65536.0,1,-nbitq), 
to_sfixed(9558.0/65536.0,1,-nbitq), 
to_sfixed(1273.0/65536.0,1,-nbitq), 
to_sfixed(-1920.0/65536.0,1,-nbitq), 
to_sfixed(6412.0/65536.0,1,-nbitq), 
to_sfixed(4626.0/65536.0,1,-nbitq), 
to_sfixed(-2297.0/65536.0,1,-nbitq), 
to_sfixed(43.0/65536.0,1,-nbitq), 
to_sfixed(-4727.0/65536.0,1,-nbitq), 
to_sfixed(-2764.0/65536.0,1,-nbitq), 
to_sfixed(10039.0/65536.0,1,-nbitq), 
to_sfixed(-3902.0/65536.0,1,-nbitq), 
to_sfixed(2519.0/65536.0,1,-nbitq), 
to_sfixed(-18605.0/65536.0,1,-nbitq), 
to_sfixed(1493.0/65536.0,1,-nbitq), 
to_sfixed(-719.0/65536.0,1,-nbitq), 
to_sfixed(-626.0/65536.0,1,-nbitq), 
to_sfixed(2823.0/65536.0,1,-nbitq), 
to_sfixed(2389.0/65536.0,1,-nbitq), 
to_sfixed(-6862.0/65536.0,1,-nbitq), 
to_sfixed(1282.0/65536.0,1,-nbitq), 
to_sfixed(-19.0/65536.0,1,-nbitq), 
to_sfixed(-8826.0/65536.0,1,-nbitq), 
to_sfixed(491.0/65536.0,1,-nbitq), 
to_sfixed(-1400.0/65536.0,1,-nbitq), 
to_sfixed(3962.0/65536.0,1,-nbitq), 
to_sfixed(-69.0/65536.0,1,-nbitq), 
to_sfixed(-6885.0/65536.0,1,-nbitq), 
to_sfixed(1050.0/65536.0,1,-nbitq), 
to_sfixed(154.0/65536.0,1,-nbitq), 
to_sfixed(2368.0/65536.0,1,-nbitq), 
to_sfixed(-2590.0/65536.0,1,-nbitq), 
to_sfixed(7612.0/65536.0,1,-nbitq), 
to_sfixed(3315.0/65536.0,1,-nbitq), 
to_sfixed(-6580.0/65536.0,1,-nbitq), 
to_sfixed(2926.0/65536.0,1,-nbitq), 
to_sfixed(3295.0/65536.0,1,-nbitq), 
to_sfixed(4052.0/65536.0,1,-nbitq), 
to_sfixed(-89.0/65536.0,1,-nbitq), 
to_sfixed(5913.0/65536.0,1,-nbitq), 
to_sfixed(-2605.0/65536.0,1,-nbitq), 
to_sfixed(-1602.0/65536.0,1,-nbitq), 
to_sfixed(2747.0/65536.0,1,-nbitq), 
to_sfixed(-1017.0/65536.0,1,-nbitq), 
to_sfixed(1475.0/65536.0,1,-nbitq), 
to_sfixed(-1204.0/65536.0,1,-nbitq), 
to_sfixed(2414.0/65536.0,1,-nbitq), 
to_sfixed(-2453.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2989.0/65536.0,1,-nbitq), 
to_sfixed(3683.0/65536.0,1,-nbitq), 
to_sfixed(-6502.0/65536.0,1,-nbitq), 
to_sfixed(1222.0/65536.0,1,-nbitq), 
to_sfixed(-3989.0/65536.0,1,-nbitq), 
to_sfixed(-6873.0/65536.0,1,-nbitq), 
to_sfixed(41.0/65536.0,1,-nbitq), 
to_sfixed(-3452.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(2483.0/65536.0,1,-nbitq), 
to_sfixed(6592.0/65536.0,1,-nbitq), 
to_sfixed(1628.0/65536.0,1,-nbitq), 
to_sfixed(142.0/65536.0,1,-nbitq), 
to_sfixed(-1200.0/65536.0,1,-nbitq), 
to_sfixed(5383.0/65536.0,1,-nbitq), 
to_sfixed(1533.0/65536.0,1,-nbitq), 
to_sfixed(-1737.0/65536.0,1,-nbitq), 
to_sfixed(5796.0/65536.0,1,-nbitq), 
to_sfixed(3465.0/65536.0,1,-nbitq), 
to_sfixed(689.0/65536.0,1,-nbitq), 
to_sfixed(-3621.0/65536.0,1,-nbitq), 
to_sfixed(6593.0/65536.0,1,-nbitq), 
to_sfixed(-1955.0/65536.0,1,-nbitq), 
to_sfixed(-5628.0/65536.0,1,-nbitq), 
to_sfixed(-631.0/65536.0,1,-nbitq), 
to_sfixed(-2722.0/65536.0,1,-nbitq), 
to_sfixed(-9524.0/65536.0,1,-nbitq), 
to_sfixed(1210.0/65536.0,1,-nbitq), 
to_sfixed(-8629.0/65536.0,1,-nbitq), 
to_sfixed(-3408.0/65536.0,1,-nbitq), 
to_sfixed(613.0/65536.0,1,-nbitq), 
to_sfixed(3721.0/65536.0,1,-nbitq), 
to_sfixed(-2468.0/65536.0,1,-nbitq), 
to_sfixed(5440.0/65536.0,1,-nbitq), 
to_sfixed(3446.0/65536.0,1,-nbitq), 
to_sfixed(2933.0/65536.0,1,-nbitq), 
to_sfixed(8942.0/65536.0,1,-nbitq), 
to_sfixed(-1286.0/65536.0,1,-nbitq), 
to_sfixed(404.0/65536.0,1,-nbitq), 
to_sfixed(95.0/65536.0,1,-nbitq), 
to_sfixed(-3335.0/65536.0,1,-nbitq), 
to_sfixed(2472.0/65536.0,1,-nbitq), 
to_sfixed(9818.0/65536.0,1,-nbitq), 
to_sfixed(-2971.0/65536.0,1,-nbitq), 
to_sfixed(-661.0/65536.0,1,-nbitq), 
to_sfixed(-11795.0/65536.0,1,-nbitq), 
to_sfixed(-960.0/65536.0,1,-nbitq), 
to_sfixed(-2631.0/65536.0,1,-nbitq), 
to_sfixed(-1078.0/65536.0,1,-nbitq), 
to_sfixed(-2267.0/65536.0,1,-nbitq), 
to_sfixed(2744.0/65536.0,1,-nbitq), 
to_sfixed(-4060.0/65536.0,1,-nbitq), 
to_sfixed(5971.0/65536.0,1,-nbitq), 
to_sfixed(-459.0/65536.0,1,-nbitq), 
to_sfixed(-4577.0/65536.0,1,-nbitq), 
to_sfixed(-2679.0/65536.0,1,-nbitq), 
to_sfixed(-506.0/65536.0,1,-nbitq), 
to_sfixed(-1375.0/65536.0,1,-nbitq), 
to_sfixed(-1533.0/65536.0,1,-nbitq), 
to_sfixed(-7730.0/65536.0,1,-nbitq), 
to_sfixed(4981.0/65536.0,1,-nbitq), 
to_sfixed(-1477.0/65536.0,1,-nbitq), 
to_sfixed(-2280.0/65536.0,1,-nbitq), 
to_sfixed(-1150.0/65536.0,1,-nbitq), 
to_sfixed(-587.0/65536.0,1,-nbitq), 
to_sfixed(4502.0/65536.0,1,-nbitq), 
to_sfixed(-7010.0/65536.0,1,-nbitq), 
to_sfixed(5728.0/65536.0,1,-nbitq), 
to_sfixed(-3491.0/65536.0,1,-nbitq), 
to_sfixed(5573.0/65536.0,1,-nbitq), 
to_sfixed(-2594.0/65536.0,1,-nbitq), 
to_sfixed(8828.0/65536.0,1,-nbitq), 
to_sfixed(-3160.0/65536.0,1,-nbitq), 
to_sfixed(-2787.0/65536.0,1,-nbitq), 
to_sfixed(1617.0/65536.0,1,-nbitq), 
to_sfixed(3068.0/65536.0,1,-nbitq), 
to_sfixed(-3297.0/65536.0,1,-nbitq), 
to_sfixed(-6107.0/65536.0,1,-nbitq), 
to_sfixed(-88.0/65536.0,1,-nbitq), 
to_sfixed(-4117.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-875.0/65536.0,1,-nbitq), 
to_sfixed(-595.0/65536.0,1,-nbitq), 
to_sfixed(-9025.0/65536.0,1,-nbitq), 
to_sfixed(-1492.0/65536.0,1,-nbitq), 
to_sfixed(1749.0/65536.0,1,-nbitq), 
to_sfixed(-5370.0/65536.0,1,-nbitq), 
to_sfixed(3125.0/65536.0,1,-nbitq), 
to_sfixed(-3025.0/65536.0,1,-nbitq), 
to_sfixed(-2165.0/65536.0,1,-nbitq), 
to_sfixed(-2357.0/65536.0,1,-nbitq), 
to_sfixed(5056.0/65536.0,1,-nbitq), 
to_sfixed(6497.0/65536.0,1,-nbitq), 
to_sfixed(1892.0/65536.0,1,-nbitq), 
to_sfixed(4635.0/65536.0,1,-nbitq), 
to_sfixed(6632.0/65536.0,1,-nbitq), 
to_sfixed(-2761.0/65536.0,1,-nbitq), 
to_sfixed(700.0/65536.0,1,-nbitq), 
to_sfixed(7156.0/65536.0,1,-nbitq), 
to_sfixed(8719.0/65536.0,1,-nbitq), 
to_sfixed(-800.0/65536.0,1,-nbitq), 
to_sfixed(-7478.0/65536.0,1,-nbitq), 
to_sfixed(3541.0/65536.0,1,-nbitq), 
to_sfixed(8921.0/65536.0,1,-nbitq), 
to_sfixed(-5387.0/65536.0,1,-nbitq), 
to_sfixed(1503.0/65536.0,1,-nbitq), 
to_sfixed(-7926.0/65536.0,1,-nbitq), 
to_sfixed(-10936.0/65536.0,1,-nbitq), 
to_sfixed(-1157.0/65536.0,1,-nbitq), 
to_sfixed(-11374.0/65536.0,1,-nbitq), 
to_sfixed(544.0/65536.0,1,-nbitq), 
to_sfixed(2551.0/65536.0,1,-nbitq), 
to_sfixed(-1370.0/65536.0,1,-nbitq), 
to_sfixed(-1114.0/65536.0,1,-nbitq), 
to_sfixed(-3187.0/65536.0,1,-nbitq), 
to_sfixed(-2484.0/65536.0,1,-nbitq), 
to_sfixed(-376.0/65536.0,1,-nbitq), 
to_sfixed(12136.0/65536.0,1,-nbitq), 
to_sfixed(-4717.0/65536.0,1,-nbitq), 
to_sfixed(5079.0/65536.0,1,-nbitq), 
to_sfixed(1393.0/65536.0,1,-nbitq), 
to_sfixed(-4937.0/65536.0,1,-nbitq), 
to_sfixed(265.0/65536.0,1,-nbitq), 
to_sfixed(510.0/65536.0,1,-nbitq), 
to_sfixed(-4506.0/65536.0,1,-nbitq), 
to_sfixed(1896.0/65536.0,1,-nbitq), 
to_sfixed(-3987.0/65536.0,1,-nbitq), 
to_sfixed(-2044.0/65536.0,1,-nbitq), 
to_sfixed(-1061.0/65536.0,1,-nbitq), 
to_sfixed(-335.0/65536.0,1,-nbitq), 
to_sfixed(1043.0/65536.0,1,-nbitq), 
to_sfixed(-460.0/65536.0,1,-nbitq), 
to_sfixed(-4285.0/65536.0,1,-nbitq), 
to_sfixed(2552.0/65536.0,1,-nbitq), 
to_sfixed(-988.0/65536.0,1,-nbitq), 
to_sfixed(-3899.0/65536.0,1,-nbitq), 
to_sfixed(-3226.0/65536.0,1,-nbitq), 
to_sfixed(-2350.0/65536.0,1,-nbitq), 
to_sfixed(-656.0/65536.0,1,-nbitq), 
to_sfixed(2637.0/65536.0,1,-nbitq), 
to_sfixed(-8076.0/65536.0,1,-nbitq), 
to_sfixed(4171.0/65536.0,1,-nbitq), 
to_sfixed(-2037.0/65536.0,1,-nbitq), 
to_sfixed(-1028.0/65536.0,1,-nbitq), 
to_sfixed(2287.0/65536.0,1,-nbitq), 
to_sfixed(-3392.0/65536.0,1,-nbitq), 
to_sfixed(2910.0/65536.0,1,-nbitq), 
to_sfixed(-3672.0/65536.0,1,-nbitq), 
to_sfixed(4919.0/65536.0,1,-nbitq), 
to_sfixed(-989.0/65536.0,1,-nbitq), 
to_sfixed(7945.0/65536.0,1,-nbitq), 
to_sfixed(-3221.0/65536.0,1,-nbitq), 
to_sfixed(5235.0/65536.0,1,-nbitq), 
to_sfixed(-5309.0/65536.0,1,-nbitq), 
to_sfixed(-1872.0/65536.0,1,-nbitq), 
to_sfixed(-2759.0/65536.0,1,-nbitq), 
to_sfixed(1813.0/65536.0,1,-nbitq), 
to_sfixed(1152.0/65536.0,1,-nbitq), 
to_sfixed(-10047.0/65536.0,1,-nbitq), 
to_sfixed(-837.0/65536.0,1,-nbitq), 
to_sfixed(-10181.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1254.0/65536.0,1,-nbitq), 
to_sfixed(819.0/65536.0,1,-nbitq), 
to_sfixed(-14515.0/65536.0,1,-nbitq), 
to_sfixed(1747.0/65536.0,1,-nbitq), 
to_sfixed(7691.0/65536.0,1,-nbitq), 
to_sfixed(-4626.0/65536.0,1,-nbitq), 
to_sfixed(2070.0/65536.0,1,-nbitq), 
to_sfixed(-1708.0/65536.0,1,-nbitq), 
to_sfixed(-101.0/65536.0,1,-nbitq), 
to_sfixed(1176.0/65536.0,1,-nbitq), 
to_sfixed(5727.0/65536.0,1,-nbitq), 
to_sfixed(57.0/65536.0,1,-nbitq), 
to_sfixed(-226.0/65536.0,1,-nbitq), 
to_sfixed(-296.0/65536.0,1,-nbitq), 
to_sfixed(4971.0/65536.0,1,-nbitq), 
to_sfixed(2686.0/65536.0,1,-nbitq), 
to_sfixed(-952.0/65536.0,1,-nbitq), 
to_sfixed(9899.0/65536.0,1,-nbitq), 
to_sfixed(8866.0/65536.0,1,-nbitq), 
to_sfixed(-2280.0/65536.0,1,-nbitq), 
to_sfixed(-4679.0/65536.0,1,-nbitq), 
to_sfixed(-1507.0/65536.0,1,-nbitq), 
to_sfixed(15891.0/65536.0,1,-nbitq), 
to_sfixed(-1779.0/65536.0,1,-nbitq), 
to_sfixed(-4331.0/65536.0,1,-nbitq), 
to_sfixed(-4826.0/65536.0,1,-nbitq), 
to_sfixed(-4605.0/65536.0,1,-nbitq), 
to_sfixed(87.0/65536.0,1,-nbitq), 
to_sfixed(-2709.0/65536.0,1,-nbitq), 
to_sfixed(-3063.0/65536.0,1,-nbitq), 
to_sfixed(3320.0/65536.0,1,-nbitq), 
to_sfixed(1653.0/65536.0,1,-nbitq), 
to_sfixed(-526.0/65536.0,1,-nbitq), 
to_sfixed(-2945.0/65536.0,1,-nbitq), 
to_sfixed(-1845.0/65536.0,1,-nbitq), 
to_sfixed(-1416.0/65536.0,1,-nbitq), 
to_sfixed(8536.0/65536.0,1,-nbitq), 
to_sfixed(-8127.0/65536.0,1,-nbitq), 
to_sfixed(619.0/65536.0,1,-nbitq), 
to_sfixed(-3256.0/65536.0,1,-nbitq), 
to_sfixed(-4407.0/65536.0,1,-nbitq), 
to_sfixed(905.0/65536.0,1,-nbitq), 
to_sfixed(-4102.0/65536.0,1,-nbitq), 
to_sfixed(-2528.0/65536.0,1,-nbitq), 
to_sfixed(-44.0/65536.0,1,-nbitq), 
to_sfixed(-1581.0/65536.0,1,-nbitq), 
to_sfixed(-1207.0/65536.0,1,-nbitq), 
to_sfixed(963.0/65536.0,1,-nbitq), 
to_sfixed(848.0/65536.0,1,-nbitq), 
to_sfixed(-315.0/65536.0,1,-nbitq), 
to_sfixed(1574.0/65536.0,1,-nbitq), 
to_sfixed(-606.0/65536.0,1,-nbitq), 
to_sfixed(802.0/65536.0,1,-nbitq), 
to_sfixed(-1920.0/65536.0,1,-nbitq), 
to_sfixed(-5534.0/65536.0,1,-nbitq), 
to_sfixed(-2224.0/65536.0,1,-nbitq), 
to_sfixed(488.0/65536.0,1,-nbitq), 
to_sfixed(-1516.0/65536.0,1,-nbitq), 
to_sfixed(1258.0/65536.0,1,-nbitq), 
to_sfixed(-6782.0/65536.0,1,-nbitq), 
to_sfixed(7831.0/65536.0,1,-nbitq), 
to_sfixed(411.0/65536.0,1,-nbitq), 
to_sfixed(-778.0/65536.0,1,-nbitq), 
to_sfixed(-292.0/65536.0,1,-nbitq), 
to_sfixed(-4034.0/65536.0,1,-nbitq), 
to_sfixed(-4341.0/65536.0,1,-nbitq), 
to_sfixed(-1343.0/65536.0,1,-nbitq), 
to_sfixed(10705.0/65536.0,1,-nbitq), 
to_sfixed(-2538.0/65536.0,1,-nbitq), 
to_sfixed(10967.0/65536.0,1,-nbitq), 
to_sfixed(-2257.0/65536.0,1,-nbitq), 
to_sfixed(2234.0/65536.0,1,-nbitq), 
to_sfixed(824.0/65536.0,1,-nbitq), 
to_sfixed(-2971.0/65536.0,1,-nbitq), 
to_sfixed(2599.0/65536.0,1,-nbitq), 
to_sfixed(-5639.0/65536.0,1,-nbitq), 
to_sfixed(631.0/65536.0,1,-nbitq), 
to_sfixed(-6528.0/65536.0,1,-nbitq), 
to_sfixed(-2664.0/65536.0,1,-nbitq), 
to_sfixed(-8811.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2256.0/65536.0,1,-nbitq), 
to_sfixed(371.0/65536.0,1,-nbitq), 
to_sfixed(-18577.0/65536.0,1,-nbitq), 
to_sfixed(2186.0/65536.0,1,-nbitq), 
to_sfixed(4456.0/65536.0,1,-nbitq), 
to_sfixed(-2638.0/65536.0,1,-nbitq), 
to_sfixed(2294.0/65536.0,1,-nbitq), 
to_sfixed(-5929.0/65536.0,1,-nbitq), 
to_sfixed(-5667.0/65536.0,1,-nbitq), 
to_sfixed(36.0/65536.0,1,-nbitq), 
to_sfixed(3173.0/65536.0,1,-nbitq), 
to_sfixed(-3096.0/65536.0,1,-nbitq), 
to_sfixed(2707.0/65536.0,1,-nbitq), 
to_sfixed(-2888.0/65536.0,1,-nbitq), 
to_sfixed(1857.0/65536.0,1,-nbitq), 
to_sfixed(-2125.0/65536.0,1,-nbitq), 
to_sfixed(772.0/65536.0,1,-nbitq), 
to_sfixed(4217.0/65536.0,1,-nbitq), 
to_sfixed(11939.0/65536.0,1,-nbitq), 
to_sfixed(-143.0/65536.0,1,-nbitq), 
to_sfixed(-5494.0/65536.0,1,-nbitq), 
to_sfixed(-525.0/65536.0,1,-nbitq), 
to_sfixed(10818.0/65536.0,1,-nbitq), 
to_sfixed(-1901.0/65536.0,1,-nbitq), 
to_sfixed(-863.0/65536.0,1,-nbitq), 
to_sfixed(235.0/65536.0,1,-nbitq), 
to_sfixed(-2849.0/65536.0,1,-nbitq), 
to_sfixed(901.0/65536.0,1,-nbitq), 
to_sfixed(6116.0/65536.0,1,-nbitq), 
to_sfixed(-2231.0/65536.0,1,-nbitq), 
to_sfixed(1019.0/65536.0,1,-nbitq), 
to_sfixed(549.0/65536.0,1,-nbitq), 
to_sfixed(-3125.0/65536.0,1,-nbitq), 
to_sfixed(-9476.0/65536.0,1,-nbitq), 
to_sfixed(-1659.0/65536.0,1,-nbitq), 
to_sfixed(-1853.0/65536.0,1,-nbitq), 
to_sfixed(10792.0/65536.0,1,-nbitq), 
to_sfixed(-6589.0/65536.0,1,-nbitq), 
to_sfixed(-1817.0/65536.0,1,-nbitq), 
to_sfixed(-880.0/65536.0,1,-nbitq), 
to_sfixed(-7844.0/65536.0,1,-nbitq), 
to_sfixed(2732.0/65536.0,1,-nbitq), 
to_sfixed(-4250.0/65536.0,1,-nbitq), 
to_sfixed(3436.0/65536.0,1,-nbitq), 
to_sfixed(-1776.0/65536.0,1,-nbitq), 
to_sfixed(-4489.0/65536.0,1,-nbitq), 
to_sfixed(-1488.0/65536.0,1,-nbitq), 
to_sfixed(10733.0/65536.0,1,-nbitq), 
to_sfixed(-2105.0/65536.0,1,-nbitq), 
to_sfixed(426.0/65536.0,1,-nbitq), 
to_sfixed(1471.0/65536.0,1,-nbitq), 
to_sfixed(-4567.0/65536.0,1,-nbitq), 
to_sfixed(-1588.0/65536.0,1,-nbitq), 
to_sfixed(-5231.0/65536.0,1,-nbitq), 
to_sfixed(-3533.0/65536.0,1,-nbitq), 
to_sfixed(-6270.0/65536.0,1,-nbitq), 
to_sfixed(1023.0/65536.0,1,-nbitq), 
to_sfixed(-851.0/65536.0,1,-nbitq), 
to_sfixed(381.0/65536.0,1,-nbitq), 
to_sfixed(-5697.0/65536.0,1,-nbitq), 
to_sfixed(6552.0/65536.0,1,-nbitq), 
to_sfixed(-867.0/65536.0,1,-nbitq), 
to_sfixed(275.0/65536.0,1,-nbitq), 
to_sfixed(-1162.0/65536.0,1,-nbitq), 
to_sfixed(-7997.0/65536.0,1,-nbitq), 
to_sfixed(-10112.0/65536.0,1,-nbitq), 
to_sfixed(-2106.0/65536.0,1,-nbitq), 
to_sfixed(7700.0/65536.0,1,-nbitq), 
to_sfixed(153.0/65536.0,1,-nbitq), 
to_sfixed(10566.0/65536.0,1,-nbitq), 
to_sfixed(-2025.0/65536.0,1,-nbitq), 
to_sfixed(2418.0/65536.0,1,-nbitq), 
to_sfixed(-4585.0/65536.0,1,-nbitq), 
to_sfixed(-494.0/65536.0,1,-nbitq), 
to_sfixed(68.0/65536.0,1,-nbitq), 
to_sfixed(-6057.0/65536.0,1,-nbitq), 
to_sfixed(5091.0/65536.0,1,-nbitq), 
to_sfixed(3364.0/65536.0,1,-nbitq), 
to_sfixed(773.0/65536.0,1,-nbitq), 
to_sfixed(-1473.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-173.0/65536.0,1,-nbitq), 
to_sfixed(2456.0/65536.0,1,-nbitq), 
to_sfixed(-14212.0/65536.0,1,-nbitq), 
to_sfixed(-10991.0/65536.0,1,-nbitq), 
to_sfixed(4202.0/65536.0,1,-nbitq), 
to_sfixed(-857.0/65536.0,1,-nbitq), 
to_sfixed(642.0/65536.0,1,-nbitq), 
to_sfixed(225.0/65536.0,1,-nbitq), 
to_sfixed(7843.0/65536.0,1,-nbitq), 
to_sfixed(1709.0/65536.0,1,-nbitq), 
to_sfixed(-1444.0/65536.0,1,-nbitq), 
to_sfixed(-8776.0/65536.0,1,-nbitq), 
to_sfixed(3404.0/65536.0,1,-nbitq), 
to_sfixed(1286.0/65536.0,1,-nbitq), 
to_sfixed(140.0/65536.0,1,-nbitq), 
to_sfixed(2431.0/65536.0,1,-nbitq), 
to_sfixed(-577.0/65536.0,1,-nbitq), 
to_sfixed(-342.0/65536.0,1,-nbitq), 
to_sfixed(4585.0/65536.0,1,-nbitq), 
to_sfixed(-2640.0/65536.0,1,-nbitq), 
to_sfixed(-8597.0/65536.0,1,-nbitq), 
to_sfixed(2854.0/65536.0,1,-nbitq), 
to_sfixed(13019.0/65536.0,1,-nbitq), 
to_sfixed(-703.0/65536.0,1,-nbitq), 
to_sfixed(-992.0/65536.0,1,-nbitq), 
to_sfixed(2210.0/65536.0,1,-nbitq), 
to_sfixed(-10714.0/65536.0,1,-nbitq), 
to_sfixed(1246.0/65536.0,1,-nbitq), 
to_sfixed(7067.0/65536.0,1,-nbitq), 
to_sfixed(2849.0/65536.0,1,-nbitq), 
to_sfixed(-48.0/65536.0,1,-nbitq), 
to_sfixed(-2104.0/65536.0,1,-nbitq), 
to_sfixed(-3201.0/65536.0,1,-nbitq), 
to_sfixed(-4237.0/65536.0,1,-nbitq), 
to_sfixed(4129.0/65536.0,1,-nbitq), 
to_sfixed(794.0/65536.0,1,-nbitq), 
to_sfixed(6387.0/65536.0,1,-nbitq), 
to_sfixed(-5024.0/65536.0,1,-nbitq), 
to_sfixed(3935.0/65536.0,1,-nbitq), 
to_sfixed(-4724.0/65536.0,1,-nbitq), 
to_sfixed(-6983.0/65536.0,1,-nbitq), 
to_sfixed(1235.0/65536.0,1,-nbitq), 
to_sfixed(-6064.0/65536.0,1,-nbitq), 
to_sfixed(1838.0/65536.0,1,-nbitq), 
to_sfixed(344.0/65536.0,1,-nbitq), 
to_sfixed(1183.0/65536.0,1,-nbitq), 
to_sfixed(263.0/65536.0,1,-nbitq), 
to_sfixed(8953.0/65536.0,1,-nbitq), 
to_sfixed(2383.0/65536.0,1,-nbitq), 
to_sfixed(-112.0/65536.0,1,-nbitq), 
to_sfixed(-2579.0/65536.0,1,-nbitq), 
to_sfixed(-7898.0/65536.0,1,-nbitq), 
to_sfixed(-3526.0/65536.0,1,-nbitq), 
to_sfixed(1140.0/65536.0,1,-nbitq), 
to_sfixed(-4912.0/65536.0,1,-nbitq), 
to_sfixed(-5159.0/65536.0,1,-nbitq), 
to_sfixed(-375.0/65536.0,1,-nbitq), 
to_sfixed(-854.0/65536.0,1,-nbitq), 
to_sfixed(-2911.0/65536.0,1,-nbitq), 
to_sfixed(-3557.0/65536.0,1,-nbitq), 
to_sfixed(3439.0/65536.0,1,-nbitq), 
to_sfixed(1300.0/65536.0,1,-nbitq), 
to_sfixed(92.0/65536.0,1,-nbitq), 
to_sfixed(2291.0/65536.0,1,-nbitq), 
to_sfixed(-3010.0/65536.0,1,-nbitq), 
to_sfixed(-9221.0/65536.0,1,-nbitq), 
to_sfixed(-6797.0/65536.0,1,-nbitq), 
to_sfixed(13445.0/65536.0,1,-nbitq), 
to_sfixed(4734.0/65536.0,1,-nbitq), 
to_sfixed(4309.0/65536.0,1,-nbitq), 
to_sfixed(641.0/65536.0,1,-nbitq), 
to_sfixed(6486.0/65536.0,1,-nbitq), 
to_sfixed(-5621.0/65536.0,1,-nbitq), 
to_sfixed(-1476.0/65536.0,1,-nbitq), 
to_sfixed(463.0/65536.0,1,-nbitq), 
to_sfixed(-838.0/65536.0,1,-nbitq), 
to_sfixed(8839.0/65536.0,1,-nbitq), 
to_sfixed(5033.0/65536.0,1,-nbitq), 
to_sfixed(-2938.0/65536.0,1,-nbitq), 
to_sfixed(2831.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-878.0/65536.0,1,-nbitq), 
to_sfixed(1577.0/65536.0,1,-nbitq), 
to_sfixed(-843.0/65536.0,1,-nbitq), 
to_sfixed(-3201.0/65536.0,1,-nbitq), 
to_sfixed(-2452.0/65536.0,1,-nbitq), 
to_sfixed(3218.0/65536.0,1,-nbitq), 
to_sfixed(-2881.0/65536.0,1,-nbitq), 
to_sfixed(-1571.0/65536.0,1,-nbitq), 
to_sfixed(7209.0/65536.0,1,-nbitq), 
to_sfixed(1219.0/65536.0,1,-nbitq), 
to_sfixed(52.0/65536.0,1,-nbitq), 
to_sfixed(-8328.0/65536.0,1,-nbitq), 
to_sfixed(372.0/65536.0,1,-nbitq), 
to_sfixed(3383.0/65536.0,1,-nbitq), 
to_sfixed(-1855.0/65536.0,1,-nbitq), 
to_sfixed(-209.0/65536.0,1,-nbitq), 
to_sfixed(-2157.0/65536.0,1,-nbitq), 
to_sfixed(-5256.0/65536.0,1,-nbitq), 
to_sfixed(1900.0/65536.0,1,-nbitq), 
to_sfixed(-1781.0/65536.0,1,-nbitq), 
to_sfixed(-7746.0/65536.0,1,-nbitq), 
to_sfixed(323.0/65536.0,1,-nbitq), 
to_sfixed(-4447.0/65536.0,1,-nbitq), 
to_sfixed(3542.0/65536.0,1,-nbitq), 
to_sfixed(61.0/65536.0,1,-nbitq), 
to_sfixed(3215.0/65536.0,1,-nbitq), 
to_sfixed(-5974.0/65536.0,1,-nbitq), 
to_sfixed(-654.0/65536.0,1,-nbitq), 
to_sfixed(6226.0/65536.0,1,-nbitq), 
to_sfixed(3394.0/65536.0,1,-nbitq), 
to_sfixed(-3788.0/65536.0,1,-nbitq), 
to_sfixed(-3355.0/65536.0,1,-nbitq), 
to_sfixed(-1656.0/65536.0,1,-nbitq), 
to_sfixed(1124.0/65536.0,1,-nbitq), 
to_sfixed(1817.0/65536.0,1,-nbitq), 
to_sfixed(1922.0/65536.0,1,-nbitq), 
to_sfixed(464.0/65536.0,1,-nbitq), 
to_sfixed(-1693.0/65536.0,1,-nbitq), 
to_sfixed(6085.0/65536.0,1,-nbitq), 
to_sfixed(-1940.0/65536.0,1,-nbitq), 
to_sfixed(-4559.0/65536.0,1,-nbitq), 
to_sfixed(-2670.0/65536.0,1,-nbitq), 
to_sfixed(-28.0/65536.0,1,-nbitq), 
to_sfixed(2533.0/65536.0,1,-nbitq), 
to_sfixed(-313.0/65536.0,1,-nbitq), 
to_sfixed(6374.0/65536.0,1,-nbitq), 
to_sfixed(744.0/65536.0,1,-nbitq), 
to_sfixed(8532.0/65536.0,1,-nbitq), 
to_sfixed(2644.0/65536.0,1,-nbitq), 
to_sfixed(1267.0/65536.0,1,-nbitq), 
to_sfixed(59.0/65536.0,1,-nbitq), 
to_sfixed(-11961.0/65536.0,1,-nbitq), 
to_sfixed(-6762.0/65536.0,1,-nbitq), 
to_sfixed(-6151.0/65536.0,1,-nbitq), 
to_sfixed(-1769.0/65536.0,1,-nbitq), 
to_sfixed(1128.0/65536.0,1,-nbitq), 
to_sfixed(1009.0/65536.0,1,-nbitq), 
to_sfixed(521.0/65536.0,1,-nbitq), 
to_sfixed(1333.0/65536.0,1,-nbitq), 
to_sfixed(-3786.0/65536.0,1,-nbitq), 
to_sfixed(-2001.0/65536.0,1,-nbitq), 
to_sfixed(1592.0/65536.0,1,-nbitq), 
to_sfixed(-747.0/65536.0,1,-nbitq), 
to_sfixed(759.0/65536.0,1,-nbitq), 
to_sfixed(629.0/65536.0,1,-nbitq), 
to_sfixed(-12232.0/65536.0,1,-nbitq), 
to_sfixed(-7994.0/65536.0,1,-nbitq), 
to_sfixed(6957.0/65536.0,1,-nbitq), 
to_sfixed(4272.0/65536.0,1,-nbitq), 
to_sfixed(-5883.0/65536.0,1,-nbitq), 
to_sfixed(-2911.0/65536.0,1,-nbitq), 
to_sfixed(8538.0/65536.0,1,-nbitq), 
to_sfixed(-11215.0/65536.0,1,-nbitq), 
to_sfixed(377.0/65536.0,1,-nbitq), 
to_sfixed(446.0/65536.0,1,-nbitq), 
to_sfixed(408.0/65536.0,1,-nbitq), 
to_sfixed(9863.0/65536.0,1,-nbitq), 
to_sfixed(2838.0/65536.0,1,-nbitq), 
to_sfixed(3163.0/65536.0,1,-nbitq), 
to_sfixed(4289.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2446.0/65536.0,1,-nbitq), 
to_sfixed(3603.0/65536.0,1,-nbitq), 
to_sfixed(2499.0/65536.0,1,-nbitq), 
to_sfixed(-3031.0/65536.0,1,-nbitq), 
to_sfixed(-4072.0/65536.0,1,-nbitq), 
to_sfixed(7230.0/65536.0,1,-nbitq), 
to_sfixed(2279.0/65536.0,1,-nbitq), 
to_sfixed(1908.0/65536.0,1,-nbitq), 
to_sfixed(7612.0/65536.0,1,-nbitq), 
to_sfixed(2434.0/65536.0,1,-nbitq), 
to_sfixed(-2595.0/65536.0,1,-nbitq), 
to_sfixed(-7424.0/65536.0,1,-nbitq), 
to_sfixed(1045.0/65536.0,1,-nbitq), 
to_sfixed(918.0/65536.0,1,-nbitq), 
to_sfixed(-222.0/65536.0,1,-nbitq), 
to_sfixed(-553.0/65536.0,1,-nbitq), 
to_sfixed(1464.0/65536.0,1,-nbitq), 
to_sfixed(-2860.0/65536.0,1,-nbitq), 
to_sfixed(1209.0/65536.0,1,-nbitq), 
to_sfixed(2061.0/65536.0,1,-nbitq), 
to_sfixed(-2903.0/65536.0,1,-nbitq), 
to_sfixed(-157.0/65536.0,1,-nbitq), 
to_sfixed(-7347.0/65536.0,1,-nbitq), 
to_sfixed(5345.0/65536.0,1,-nbitq), 
to_sfixed(-1603.0/65536.0,1,-nbitq), 
to_sfixed(2761.0/65536.0,1,-nbitq), 
to_sfixed(-2348.0/65536.0,1,-nbitq), 
to_sfixed(2115.0/65536.0,1,-nbitq), 
to_sfixed(7527.0/65536.0,1,-nbitq), 
to_sfixed(1889.0/65536.0,1,-nbitq), 
to_sfixed(-847.0/65536.0,1,-nbitq), 
to_sfixed(-7361.0/65536.0,1,-nbitq), 
to_sfixed(-3668.0/65536.0,1,-nbitq), 
to_sfixed(6050.0/65536.0,1,-nbitq), 
to_sfixed(139.0/65536.0,1,-nbitq), 
to_sfixed(4009.0/65536.0,1,-nbitq), 
to_sfixed(1300.0/65536.0,1,-nbitq), 
to_sfixed(600.0/65536.0,1,-nbitq), 
to_sfixed(5501.0/65536.0,1,-nbitq), 
to_sfixed(-508.0/65536.0,1,-nbitq), 
to_sfixed(-3854.0/65536.0,1,-nbitq), 
to_sfixed(-2786.0/65536.0,1,-nbitq), 
to_sfixed(-10446.0/65536.0,1,-nbitq), 
to_sfixed(-984.0/65536.0,1,-nbitq), 
to_sfixed(-2377.0/65536.0,1,-nbitq), 
to_sfixed(3529.0/65536.0,1,-nbitq), 
to_sfixed(-1504.0/65536.0,1,-nbitq), 
to_sfixed(1157.0/65536.0,1,-nbitq), 
to_sfixed(557.0/65536.0,1,-nbitq), 
to_sfixed(1169.0/65536.0,1,-nbitq), 
to_sfixed(-1947.0/65536.0,1,-nbitq), 
to_sfixed(-4077.0/65536.0,1,-nbitq), 
to_sfixed(-4731.0/65536.0,1,-nbitq), 
to_sfixed(-5899.0/65536.0,1,-nbitq), 
to_sfixed(-4091.0/65536.0,1,-nbitq), 
to_sfixed(-4139.0/65536.0,1,-nbitq), 
to_sfixed(-3042.0/65536.0,1,-nbitq), 
to_sfixed(-2952.0/65536.0,1,-nbitq), 
to_sfixed(533.0/65536.0,1,-nbitq), 
to_sfixed(-2956.0/65536.0,1,-nbitq), 
to_sfixed(-2896.0/65536.0,1,-nbitq), 
to_sfixed(2259.0/65536.0,1,-nbitq), 
to_sfixed(1508.0/65536.0,1,-nbitq), 
to_sfixed(-1154.0/65536.0,1,-nbitq), 
to_sfixed(-1051.0/65536.0,1,-nbitq), 
to_sfixed(-6188.0/65536.0,1,-nbitq), 
to_sfixed(-5615.0/65536.0,1,-nbitq), 
to_sfixed(2818.0/65536.0,1,-nbitq), 
to_sfixed(4912.0/65536.0,1,-nbitq), 
to_sfixed(-6117.0/65536.0,1,-nbitq), 
to_sfixed(-4335.0/65536.0,1,-nbitq), 
to_sfixed(2493.0/65536.0,1,-nbitq), 
to_sfixed(-1483.0/65536.0,1,-nbitq), 
to_sfixed(-1470.0/65536.0,1,-nbitq), 
to_sfixed(-834.0/65536.0,1,-nbitq), 
to_sfixed(505.0/65536.0,1,-nbitq), 
to_sfixed(7016.0/65536.0,1,-nbitq), 
to_sfixed(347.0/65536.0,1,-nbitq), 
to_sfixed(2521.0/65536.0,1,-nbitq), 
to_sfixed(6197.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-5704.0/65536.0,1,-nbitq), 
to_sfixed(-1037.0/65536.0,1,-nbitq), 
to_sfixed(4364.0/65536.0,1,-nbitq), 
to_sfixed(-4390.0/65536.0,1,-nbitq), 
to_sfixed(2507.0/65536.0,1,-nbitq), 
to_sfixed(13864.0/65536.0,1,-nbitq), 
to_sfixed(-984.0/65536.0,1,-nbitq), 
to_sfixed(-1784.0/65536.0,1,-nbitq), 
to_sfixed(5832.0/65536.0,1,-nbitq), 
to_sfixed(3176.0/65536.0,1,-nbitq), 
to_sfixed(922.0/65536.0,1,-nbitq), 
to_sfixed(-7919.0/65536.0,1,-nbitq), 
to_sfixed(-842.0/65536.0,1,-nbitq), 
to_sfixed(-2006.0/65536.0,1,-nbitq), 
to_sfixed(303.0/65536.0,1,-nbitq), 
to_sfixed(3027.0/65536.0,1,-nbitq), 
to_sfixed(1009.0/65536.0,1,-nbitq), 
to_sfixed(-2018.0/65536.0,1,-nbitq), 
to_sfixed(1229.0/65536.0,1,-nbitq), 
to_sfixed(1440.0/65536.0,1,-nbitq), 
to_sfixed(-3170.0/65536.0,1,-nbitq), 
to_sfixed(4309.0/65536.0,1,-nbitq), 
to_sfixed(155.0/65536.0,1,-nbitq), 
to_sfixed(1201.0/65536.0,1,-nbitq), 
to_sfixed(-24.0/65536.0,1,-nbitq), 
to_sfixed(20.0/65536.0,1,-nbitq), 
to_sfixed(969.0/65536.0,1,-nbitq), 
to_sfixed(1600.0/65536.0,1,-nbitq), 
to_sfixed(3231.0/65536.0,1,-nbitq), 
to_sfixed(-1189.0/65536.0,1,-nbitq), 
to_sfixed(742.0/65536.0,1,-nbitq), 
to_sfixed(-9749.0/65536.0,1,-nbitq), 
to_sfixed(-6103.0/65536.0,1,-nbitq), 
to_sfixed(4198.0/65536.0,1,-nbitq), 
to_sfixed(-1693.0/65536.0,1,-nbitq), 
to_sfixed(-887.0/65536.0,1,-nbitq), 
to_sfixed(4828.0/65536.0,1,-nbitq), 
to_sfixed(-48.0/65536.0,1,-nbitq), 
to_sfixed(3902.0/65536.0,1,-nbitq), 
to_sfixed(-1976.0/65536.0,1,-nbitq), 
to_sfixed(-1118.0/65536.0,1,-nbitq), 
to_sfixed(-722.0/65536.0,1,-nbitq), 
to_sfixed(-13550.0/65536.0,1,-nbitq), 
to_sfixed(-5900.0/65536.0,1,-nbitq), 
to_sfixed(2613.0/65536.0,1,-nbitq), 
to_sfixed(-4081.0/65536.0,1,-nbitq), 
to_sfixed(1584.0/65536.0,1,-nbitq), 
to_sfixed(1138.0/65536.0,1,-nbitq), 
to_sfixed(-742.0/65536.0,1,-nbitq), 
to_sfixed(-992.0/65536.0,1,-nbitq), 
to_sfixed(55.0/65536.0,1,-nbitq), 
to_sfixed(-2412.0/65536.0,1,-nbitq), 
to_sfixed(-1166.0/65536.0,1,-nbitq), 
to_sfixed(1708.0/65536.0,1,-nbitq), 
to_sfixed(-3147.0/65536.0,1,-nbitq), 
to_sfixed(-9195.0/65536.0,1,-nbitq), 
to_sfixed(-280.0/65536.0,1,-nbitq), 
to_sfixed(-2547.0/65536.0,1,-nbitq), 
to_sfixed(-1218.0/65536.0,1,-nbitq), 
to_sfixed(3684.0/65536.0,1,-nbitq), 
to_sfixed(-1867.0/65536.0,1,-nbitq), 
to_sfixed(1290.0/65536.0,1,-nbitq), 
to_sfixed(2256.0/65536.0,1,-nbitq), 
to_sfixed(-425.0/65536.0,1,-nbitq), 
to_sfixed(1967.0/65536.0,1,-nbitq), 
to_sfixed(-6114.0/65536.0,1,-nbitq), 
to_sfixed(-11145.0/65536.0,1,-nbitq), 
to_sfixed(5198.0/65536.0,1,-nbitq), 
to_sfixed(1938.0/65536.0,1,-nbitq), 
to_sfixed(-4375.0/65536.0,1,-nbitq), 
to_sfixed(-4283.0/65536.0,1,-nbitq), 
to_sfixed(-162.0/65536.0,1,-nbitq), 
to_sfixed(2119.0/65536.0,1,-nbitq), 
to_sfixed(-1288.0/65536.0,1,-nbitq), 
to_sfixed(277.0/65536.0,1,-nbitq), 
to_sfixed(-3353.0/65536.0,1,-nbitq), 
to_sfixed(4889.0/65536.0,1,-nbitq), 
to_sfixed(-1506.0/65536.0,1,-nbitq), 
to_sfixed(2888.0/65536.0,1,-nbitq), 
to_sfixed(2869.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3292.0/65536.0,1,-nbitq), 
to_sfixed(-4118.0/65536.0,1,-nbitq), 
to_sfixed(4212.0/65536.0,1,-nbitq), 
to_sfixed(-5291.0/65536.0,1,-nbitq), 
to_sfixed(8601.0/65536.0,1,-nbitq), 
to_sfixed(13792.0/65536.0,1,-nbitq), 
to_sfixed(1199.0/65536.0,1,-nbitq), 
to_sfixed(1867.0/65536.0,1,-nbitq), 
to_sfixed(6411.0/65536.0,1,-nbitq), 
to_sfixed(2204.0/65536.0,1,-nbitq), 
to_sfixed(-1685.0/65536.0,1,-nbitq), 
to_sfixed(167.0/65536.0,1,-nbitq), 
to_sfixed(-3023.0/65536.0,1,-nbitq), 
to_sfixed(-694.0/65536.0,1,-nbitq), 
to_sfixed(155.0/65536.0,1,-nbitq), 
to_sfixed(897.0/65536.0,1,-nbitq), 
to_sfixed(2561.0/65536.0,1,-nbitq), 
to_sfixed(-2554.0/65536.0,1,-nbitq), 
to_sfixed(134.0/65536.0,1,-nbitq), 
to_sfixed(1156.0/65536.0,1,-nbitq), 
to_sfixed(4692.0/65536.0,1,-nbitq), 
to_sfixed(2306.0/65536.0,1,-nbitq), 
to_sfixed(3829.0/65536.0,1,-nbitq), 
to_sfixed(-3490.0/65536.0,1,-nbitq), 
to_sfixed(509.0/65536.0,1,-nbitq), 
to_sfixed(8289.0/65536.0,1,-nbitq), 
to_sfixed(4241.0/65536.0,1,-nbitq), 
to_sfixed(1033.0/65536.0,1,-nbitq), 
to_sfixed(5501.0/65536.0,1,-nbitq), 
to_sfixed(550.0/65536.0,1,-nbitq), 
to_sfixed(1984.0/65536.0,1,-nbitq), 
to_sfixed(-8185.0/65536.0,1,-nbitq), 
to_sfixed(-1308.0/65536.0,1,-nbitq), 
to_sfixed(6107.0/65536.0,1,-nbitq), 
to_sfixed(750.0/65536.0,1,-nbitq), 
to_sfixed(1714.0/65536.0,1,-nbitq), 
to_sfixed(5984.0/65536.0,1,-nbitq), 
to_sfixed(-4915.0/65536.0,1,-nbitq), 
to_sfixed(-1603.0/65536.0,1,-nbitq), 
to_sfixed(315.0/65536.0,1,-nbitq), 
to_sfixed(-563.0/65536.0,1,-nbitq), 
to_sfixed(883.0/65536.0,1,-nbitq), 
to_sfixed(-9967.0/65536.0,1,-nbitq), 
to_sfixed(-1771.0/65536.0,1,-nbitq), 
to_sfixed(-647.0/65536.0,1,-nbitq), 
to_sfixed(-8395.0/65536.0,1,-nbitq), 
to_sfixed(1040.0/65536.0,1,-nbitq), 
to_sfixed(-3405.0/65536.0,1,-nbitq), 
to_sfixed(1559.0/65536.0,1,-nbitq), 
to_sfixed(3460.0/65536.0,1,-nbitq), 
to_sfixed(2247.0/65536.0,1,-nbitq), 
to_sfixed(-1062.0/65536.0,1,-nbitq), 
to_sfixed(-1450.0/65536.0,1,-nbitq), 
to_sfixed(3262.0/65536.0,1,-nbitq), 
to_sfixed(-1321.0/65536.0,1,-nbitq), 
to_sfixed(-1676.0/65536.0,1,-nbitq), 
to_sfixed(-137.0/65536.0,1,-nbitq), 
to_sfixed(-2151.0/65536.0,1,-nbitq), 
to_sfixed(922.0/65536.0,1,-nbitq), 
to_sfixed(5548.0/65536.0,1,-nbitq), 
to_sfixed(-5144.0/65536.0,1,-nbitq), 
to_sfixed(-1428.0/65536.0,1,-nbitq), 
to_sfixed(893.0/65536.0,1,-nbitq), 
to_sfixed(-2496.0/65536.0,1,-nbitq), 
to_sfixed(-1002.0/65536.0,1,-nbitq), 
to_sfixed(-23.0/65536.0,1,-nbitq), 
to_sfixed(-5494.0/65536.0,1,-nbitq), 
to_sfixed(1862.0/65536.0,1,-nbitq), 
to_sfixed(-2368.0/65536.0,1,-nbitq), 
to_sfixed(-4371.0/65536.0,1,-nbitq), 
to_sfixed(1756.0/65536.0,1,-nbitq), 
to_sfixed(980.0/65536.0,1,-nbitq), 
to_sfixed(8548.0/65536.0,1,-nbitq), 
to_sfixed(-484.0/65536.0,1,-nbitq), 
to_sfixed(2811.0/65536.0,1,-nbitq), 
to_sfixed(657.0/65536.0,1,-nbitq), 
to_sfixed(6203.0/65536.0,1,-nbitq), 
to_sfixed(-4863.0/65536.0,1,-nbitq), 
to_sfixed(2902.0/65536.0,1,-nbitq), 
to_sfixed(2291.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3564.0/65536.0,1,-nbitq), 
to_sfixed(-3259.0/65536.0,1,-nbitq), 
to_sfixed(1140.0/65536.0,1,-nbitq), 
to_sfixed(-1926.0/65536.0,1,-nbitq), 
to_sfixed(8736.0/65536.0,1,-nbitq), 
to_sfixed(10195.0/65536.0,1,-nbitq), 
to_sfixed(2997.0/65536.0,1,-nbitq), 
to_sfixed(-1177.0/65536.0,1,-nbitq), 
to_sfixed(-1475.0/65536.0,1,-nbitq), 
to_sfixed(1177.0/65536.0,1,-nbitq), 
to_sfixed(-4021.0/65536.0,1,-nbitq), 
to_sfixed(-2593.0/65536.0,1,-nbitq), 
to_sfixed(1859.0/65536.0,1,-nbitq), 
to_sfixed(5034.0/65536.0,1,-nbitq), 
to_sfixed(-421.0/65536.0,1,-nbitq), 
to_sfixed(1919.0/65536.0,1,-nbitq), 
to_sfixed(-415.0/65536.0,1,-nbitq), 
to_sfixed(-6317.0/65536.0,1,-nbitq), 
to_sfixed(2896.0/65536.0,1,-nbitq), 
to_sfixed(-1567.0/65536.0,1,-nbitq), 
to_sfixed(3184.0/65536.0,1,-nbitq), 
to_sfixed(-1515.0/65536.0,1,-nbitq), 
to_sfixed(1254.0/65536.0,1,-nbitq), 
to_sfixed(1333.0/65536.0,1,-nbitq), 
to_sfixed(4090.0/65536.0,1,-nbitq), 
to_sfixed(7232.0/65536.0,1,-nbitq), 
to_sfixed(5090.0/65536.0,1,-nbitq), 
to_sfixed(-1618.0/65536.0,1,-nbitq), 
to_sfixed(4837.0/65536.0,1,-nbitq), 
to_sfixed(3314.0/65536.0,1,-nbitq), 
to_sfixed(3061.0/65536.0,1,-nbitq), 
to_sfixed(-5049.0/65536.0,1,-nbitq), 
to_sfixed(2447.0/65536.0,1,-nbitq), 
to_sfixed(8127.0/65536.0,1,-nbitq), 
to_sfixed(-2330.0/65536.0,1,-nbitq), 
to_sfixed(31.0/65536.0,1,-nbitq), 
to_sfixed(7799.0/65536.0,1,-nbitq), 
to_sfixed(-2815.0/65536.0,1,-nbitq), 
to_sfixed(511.0/65536.0,1,-nbitq), 
to_sfixed(-730.0/65536.0,1,-nbitq), 
to_sfixed(4475.0/65536.0,1,-nbitq), 
to_sfixed(-371.0/65536.0,1,-nbitq), 
to_sfixed(-188.0/65536.0,1,-nbitq), 
to_sfixed(-3203.0/65536.0,1,-nbitq), 
to_sfixed(-1158.0/65536.0,1,-nbitq), 
to_sfixed(-4944.0/65536.0,1,-nbitq), 
to_sfixed(882.0/65536.0,1,-nbitq), 
to_sfixed(-8155.0/65536.0,1,-nbitq), 
to_sfixed(-2132.0/65536.0,1,-nbitq), 
to_sfixed(430.0/65536.0,1,-nbitq), 
to_sfixed(-508.0/65536.0,1,-nbitq), 
to_sfixed(-1012.0/65536.0,1,-nbitq), 
to_sfixed(-3162.0/65536.0,1,-nbitq), 
to_sfixed(-2528.0/65536.0,1,-nbitq), 
to_sfixed(2785.0/65536.0,1,-nbitq), 
to_sfixed(1901.0/65536.0,1,-nbitq), 
to_sfixed(-1402.0/65536.0,1,-nbitq), 
to_sfixed(-551.0/65536.0,1,-nbitq), 
to_sfixed(-2438.0/65536.0,1,-nbitq), 
to_sfixed(-2299.0/65536.0,1,-nbitq), 
to_sfixed(-1924.0/65536.0,1,-nbitq), 
to_sfixed(1612.0/65536.0,1,-nbitq), 
to_sfixed(1187.0/65536.0,1,-nbitq), 
to_sfixed(-2712.0/65536.0,1,-nbitq), 
to_sfixed(-962.0/65536.0,1,-nbitq), 
to_sfixed(163.0/65536.0,1,-nbitq), 
to_sfixed(-6154.0/65536.0,1,-nbitq), 
to_sfixed(2080.0/65536.0,1,-nbitq), 
to_sfixed(1553.0/65536.0,1,-nbitq), 
to_sfixed(-8100.0/65536.0,1,-nbitq), 
to_sfixed(-487.0/65536.0,1,-nbitq), 
to_sfixed(5448.0/65536.0,1,-nbitq), 
to_sfixed(3553.0/65536.0,1,-nbitq), 
to_sfixed(-1717.0/65536.0,1,-nbitq), 
to_sfixed(1574.0/65536.0,1,-nbitq), 
to_sfixed(7638.0/65536.0,1,-nbitq), 
to_sfixed(9723.0/65536.0,1,-nbitq), 
to_sfixed(-8055.0/65536.0,1,-nbitq), 
to_sfixed(-1639.0/65536.0,1,-nbitq), 
to_sfixed(-1111.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2953.0/65536.0,1,-nbitq), 
to_sfixed(409.0/65536.0,1,-nbitq), 
to_sfixed(1178.0/65536.0,1,-nbitq), 
to_sfixed(-2537.0/65536.0,1,-nbitq), 
to_sfixed(4997.0/65536.0,1,-nbitq), 
to_sfixed(8938.0/65536.0,1,-nbitq), 
to_sfixed(-170.0/65536.0,1,-nbitq), 
to_sfixed(2107.0/65536.0,1,-nbitq), 
to_sfixed(2431.0/65536.0,1,-nbitq), 
to_sfixed(2072.0/65536.0,1,-nbitq), 
to_sfixed(-2527.0/65536.0,1,-nbitq), 
to_sfixed(-1499.0/65536.0,1,-nbitq), 
to_sfixed(111.0/65536.0,1,-nbitq), 
to_sfixed(10407.0/65536.0,1,-nbitq), 
to_sfixed(-4622.0/65536.0,1,-nbitq), 
to_sfixed(-1517.0/65536.0,1,-nbitq), 
to_sfixed(-500.0/65536.0,1,-nbitq), 
to_sfixed(-484.0/65536.0,1,-nbitq), 
to_sfixed(259.0/65536.0,1,-nbitq), 
to_sfixed(-1028.0/65536.0,1,-nbitq), 
to_sfixed(1474.0/65536.0,1,-nbitq), 
to_sfixed(104.0/65536.0,1,-nbitq), 
to_sfixed(-1924.0/65536.0,1,-nbitq), 
to_sfixed(9834.0/65536.0,1,-nbitq), 
to_sfixed(299.0/65536.0,1,-nbitq), 
to_sfixed(3260.0/65536.0,1,-nbitq), 
to_sfixed(2734.0/65536.0,1,-nbitq), 
to_sfixed(-2176.0/65536.0,1,-nbitq), 
to_sfixed(1401.0/65536.0,1,-nbitq), 
to_sfixed(-5174.0/65536.0,1,-nbitq), 
to_sfixed(1378.0/65536.0,1,-nbitq), 
to_sfixed(-811.0/65536.0,1,-nbitq), 
to_sfixed(1377.0/65536.0,1,-nbitq), 
to_sfixed(4917.0/65536.0,1,-nbitq), 
to_sfixed(-4217.0/65536.0,1,-nbitq), 
to_sfixed(-276.0/65536.0,1,-nbitq), 
to_sfixed(7254.0/65536.0,1,-nbitq), 
to_sfixed(-1898.0/65536.0,1,-nbitq), 
to_sfixed(3558.0/65536.0,1,-nbitq), 
to_sfixed(3121.0/65536.0,1,-nbitq), 
to_sfixed(6994.0/65536.0,1,-nbitq), 
to_sfixed(-1258.0/65536.0,1,-nbitq), 
to_sfixed(3589.0/65536.0,1,-nbitq), 
to_sfixed(-1701.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(-1148.0/65536.0,1,-nbitq), 
to_sfixed(131.0/65536.0,1,-nbitq), 
to_sfixed(-4036.0/65536.0,1,-nbitq), 
to_sfixed(-2274.0/65536.0,1,-nbitq), 
to_sfixed(2129.0/65536.0,1,-nbitq), 
to_sfixed(-2174.0/65536.0,1,-nbitq), 
to_sfixed(-8590.0/65536.0,1,-nbitq), 
to_sfixed(-12046.0/65536.0,1,-nbitq), 
to_sfixed(-2299.0/65536.0,1,-nbitq), 
to_sfixed(8628.0/65536.0,1,-nbitq), 
to_sfixed(6989.0/65536.0,1,-nbitq), 
to_sfixed(1866.0/65536.0,1,-nbitq), 
to_sfixed(375.0/65536.0,1,-nbitq), 
to_sfixed(1801.0/65536.0,1,-nbitq), 
to_sfixed(-3129.0/65536.0,1,-nbitq), 
to_sfixed(-1630.0/65536.0,1,-nbitq), 
to_sfixed(974.0/65536.0,1,-nbitq), 
to_sfixed(-2208.0/65536.0,1,-nbitq), 
to_sfixed(-2378.0/65536.0,1,-nbitq), 
to_sfixed(1216.0/65536.0,1,-nbitq), 
to_sfixed(-4985.0/65536.0,1,-nbitq), 
to_sfixed(-2069.0/65536.0,1,-nbitq), 
to_sfixed(-4035.0/65536.0,1,-nbitq), 
to_sfixed(4319.0/65536.0,1,-nbitq), 
to_sfixed(-6411.0/65536.0,1,-nbitq), 
to_sfixed(2277.0/65536.0,1,-nbitq), 
to_sfixed(8159.0/65536.0,1,-nbitq), 
to_sfixed(4672.0/65536.0,1,-nbitq), 
to_sfixed(-852.0/65536.0,1,-nbitq), 
to_sfixed(1524.0/65536.0,1,-nbitq), 
to_sfixed(1003.0/65536.0,1,-nbitq), 
to_sfixed(9225.0/65536.0,1,-nbitq), 
to_sfixed(-11314.0/65536.0,1,-nbitq), 
to_sfixed(-1860.0/65536.0,1,-nbitq), 
to_sfixed(-5551.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1854.0/65536.0,1,-nbitq), 
to_sfixed(-4422.0/65536.0,1,-nbitq), 
to_sfixed(-926.0/65536.0,1,-nbitq), 
to_sfixed(3829.0/65536.0,1,-nbitq), 
to_sfixed(2176.0/65536.0,1,-nbitq), 
to_sfixed(5457.0/65536.0,1,-nbitq), 
to_sfixed(1296.0/65536.0,1,-nbitq), 
to_sfixed(-616.0/65536.0,1,-nbitq), 
to_sfixed(-561.0/65536.0,1,-nbitq), 
to_sfixed(286.0/65536.0,1,-nbitq), 
to_sfixed(-3981.0/65536.0,1,-nbitq), 
to_sfixed(3659.0/65536.0,1,-nbitq), 
to_sfixed(-3629.0/65536.0,1,-nbitq), 
to_sfixed(6929.0/65536.0,1,-nbitq), 
to_sfixed(-70.0/65536.0,1,-nbitq), 
to_sfixed(-863.0/65536.0,1,-nbitq), 
to_sfixed(-1817.0/65536.0,1,-nbitq), 
to_sfixed(-331.0/65536.0,1,-nbitq), 
to_sfixed(-2139.0/65536.0,1,-nbitq), 
to_sfixed(-992.0/65536.0,1,-nbitq), 
to_sfixed(-793.0/65536.0,1,-nbitq), 
to_sfixed(4387.0/65536.0,1,-nbitq), 
to_sfixed(-3269.0/65536.0,1,-nbitq), 
to_sfixed(12333.0/65536.0,1,-nbitq), 
to_sfixed(-1229.0/65536.0,1,-nbitq), 
to_sfixed(2070.0/65536.0,1,-nbitq), 
to_sfixed(6821.0/65536.0,1,-nbitq), 
to_sfixed(-2432.0/65536.0,1,-nbitq), 
to_sfixed(134.0/65536.0,1,-nbitq), 
to_sfixed(-3218.0/65536.0,1,-nbitq), 
to_sfixed(-2570.0/65536.0,1,-nbitq), 
to_sfixed(3766.0/65536.0,1,-nbitq), 
to_sfixed(2745.0/65536.0,1,-nbitq), 
to_sfixed(-4241.0/65536.0,1,-nbitq), 
to_sfixed(-1084.0/65536.0,1,-nbitq), 
to_sfixed(-4693.0/65536.0,1,-nbitq), 
to_sfixed(4439.0/65536.0,1,-nbitq), 
to_sfixed(-1779.0/65536.0,1,-nbitq), 
to_sfixed(5386.0/65536.0,1,-nbitq), 
to_sfixed(2532.0/65536.0,1,-nbitq), 
to_sfixed(6071.0/65536.0,1,-nbitq), 
to_sfixed(1292.0/65536.0,1,-nbitq), 
to_sfixed(3232.0/65536.0,1,-nbitq), 
to_sfixed(-3405.0/65536.0,1,-nbitq), 
to_sfixed(-841.0/65536.0,1,-nbitq), 
to_sfixed(-2987.0/65536.0,1,-nbitq), 
to_sfixed(-842.0/65536.0,1,-nbitq), 
to_sfixed(-275.0/65536.0,1,-nbitq), 
to_sfixed(-859.0/65536.0,1,-nbitq), 
to_sfixed(3314.0/65536.0,1,-nbitq), 
to_sfixed(-638.0/65536.0,1,-nbitq), 
to_sfixed(-3989.0/65536.0,1,-nbitq), 
to_sfixed(-9081.0/65536.0,1,-nbitq), 
to_sfixed(1947.0/65536.0,1,-nbitq), 
to_sfixed(1668.0/65536.0,1,-nbitq), 
to_sfixed(5396.0/65536.0,1,-nbitq), 
to_sfixed(2457.0/65536.0,1,-nbitq), 
to_sfixed(555.0/65536.0,1,-nbitq), 
to_sfixed(1848.0/65536.0,1,-nbitq), 
to_sfixed(2637.0/65536.0,1,-nbitq), 
to_sfixed(-2194.0/65536.0,1,-nbitq), 
to_sfixed(1517.0/65536.0,1,-nbitq), 
to_sfixed(824.0/65536.0,1,-nbitq), 
to_sfixed(863.0/65536.0,1,-nbitq), 
to_sfixed(-7022.0/65536.0,1,-nbitq), 
to_sfixed(-2324.0/65536.0,1,-nbitq), 
to_sfixed(-5046.0/65536.0,1,-nbitq), 
to_sfixed(-555.0/65536.0,1,-nbitq), 
to_sfixed(-6893.0/65536.0,1,-nbitq), 
to_sfixed(-6088.0/65536.0,1,-nbitq), 
to_sfixed(5233.0/65536.0,1,-nbitq), 
to_sfixed(955.0/65536.0,1,-nbitq), 
to_sfixed(3271.0/65536.0,1,-nbitq), 
to_sfixed(-973.0/65536.0,1,-nbitq), 
to_sfixed(142.0/65536.0,1,-nbitq), 
to_sfixed(1604.0/65536.0,1,-nbitq), 
to_sfixed(7271.0/65536.0,1,-nbitq), 
to_sfixed(-5082.0/65536.0,1,-nbitq), 
to_sfixed(570.0/65536.0,1,-nbitq), 
to_sfixed(-1829.0/65536.0,1,-nbitq)  ), 
( to_sfixed(6280.0/65536.0,1,-nbitq), 
to_sfixed(611.0/65536.0,1,-nbitq), 
to_sfixed(3534.0/65536.0,1,-nbitq), 
to_sfixed(1244.0/65536.0,1,-nbitq), 
to_sfixed(-2486.0/65536.0,1,-nbitq), 
to_sfixed(2854.0/65536.0,1,-nbitq), 
to_sfixed(2734.0/65536.0,1,-nbitq), 
to_sfixed(1728.0/65536.0,1,-nbitq), 
to_sfixed(-1749.0/65536.0,1,-nbitq), 
to_sfixed(-1498.0/65536.0,1,-nbitq), 
to_sfixed(-1799.0/65536.0,1,-nbitq), 
to_sfixed(4432.0/65536.0,1,-nbitq), 
to_sfixed(-2407.0/65536.0,1,-nbitq), 
to_sfixed(3633.0/65536.0,1,-nbitq), 
to_sfixed(1107.0/65536.0,1,-nbitq), 
to_sfixed(1758.0/65536.0,1,-nbitq), 
to_sfixed(212.0/65536.0,1,-nbitq), 
to_sfixed(658.0/65536.0,1,-nbitq), 
to_sfixed(-4037.0/65536.0,1,-nbitq), 
to_sfixed(50.0/65536.0,1,-nbitq), 
to_sfixed(414.0/65536.0,1,-nbitq), 
to_sfixed(1408.0/65536.0,1,-nbitq), 
to_sfixed(-2003.0/65536.0,1,-nbitq), 
to_sfixed(6391.0/65536.0,1,-nbitq), 
to_sfixed(-505.0/65536.0,1,-nbitq), 
to_sfixed(2635.0/65536.0,1,-nbitq), 
to_sfixed(2644.0/65536.0,1,-nbitq), 
to_sfixed(-1128.0/65536.0,1,-nbitq), 
to_sfixed(-1620.0/65536.0,1,-nbitq), 
to_sfixed(901.0/65536.0,1,-nbitq), 
to_sfixed(-2870.0/65536.0,1,-nbitq), 
to_sfixed(-1347.0/65536.0,1,-nbitq), 
to_sfixed(2424.0/65536.0,1,-nbitq), 
to_sfixed(-1722.0/65536.0,1,-nbitq), 
to_sfixed(-236.0/65536.0,1,-nbitq), 
to_sfixed(-620.0/65536.0,1,-nbitq), 
to_sfixed(3229.0/65536.0,1,-nbitq), 
to_sfixed(1967.0/65536.0,1,-nbitq), 
to_sfixed(4792.0/65536.0,1,-nbitq), 
to_sfixed(-1849.0/65536.0,1,-nbitq), 
to_sfixed(3604.0/65536.0,1,-nbitq), 
to_sfixed(-2786.0/65536.0,1,-nbitq), 
to_sfixed(5798.0/65536.0,1,-nbitq), 
to_sfixed(-558.0/65536.0,1,-nbitq), 
to_sfixed(-182.0/65536.0,1,-nbitq), 
to_sfixed(475.0/65536.0,1,-nbitq), 
to_sfixed(1588.0/65536.0,1,-nbitq), 
to_sfixed(2016.0/65536.0,1,-nbitq), 
to_sfixed(2230.0/65536.0,1,-nbitq), 
to_sfixed(1254.0/65536.0,1,-nbitq), 
to_sfixed(2915.0/65536.0,1,-nbitq), 
to_sfixed(-3069.0/65536.0,1,-nbitq), 
to_sfixed(-2139.0/65536.0,1,-nbitq), 
to_sfixed(-3017.0/65536.0,1,-nbitq), 
to_sfixed(6776.0/65536.0,1,-nbitq), 
to_sfixed(1004.0/65536.0,1,-nbitq), 
to_sfixed(-675.0/65536.0,1,-nbitq), 
to_sfixed(2231.0/65536.0,1,-nbitq), 
to_sfixed(-240.0/65536.0,1,-nbitq), 
to_sfixed(4819.0/65536.0,1,-nbitq), 
to_sfixed(-1404.0/65536.0,1,-nbitq), 
to_sfixed(-1294.0/65536.0,1,-nbitq), 
to_sfixed(1583.0/65536.0,1,-nbitq), 
to_sfixed(-2145.0/65536.0,1,-nbitq), 
to_sfixed(-6456.0/65536.0,1,-nbitq), 
to_sfixed(-448.0/65536.0,1,-nbitq), 
to_sfixed(-4949.0/65536.0,1,-nbitq), 
to_sfixed(-3010.0/65536.0,1,-nbitq), 
to_sfixed(-7486.0/65536.0,1,-nbitq), 
to_sfixed(-8316.0/65536.0,1,-nbitq), 
to_sfixed(5339.0/65536.0,1,-nbitq), 
to_sfixed(-4966.0/65536.0,1,-nbitq), 
to_sfixed(467.0/65536.0,1,-nbitq), 
to_sfixed(-1675.0/65536.0,1,-nbitq), 
to_sfixed(-1629.0/65536.0,1,-nbitq), 
to_sfixed(4778.0/65536.0,1,-nbitq), 
to_sfixed(-780.0/65536.0,1,-nbitq), 
to_sfixed(-2199.0/65536.0,1,-nbitq), 
to_sfixed(-82.0/65536.0,1,-nbitq), 
to_sfixed(-1913.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4504.0/65536.0,1,-nbitq), 
to_sfixed(3381.0/65536.0,1,-nbitq), 
to_sfixed(2036.0/65536.0,1,-nbitq), 
to_sfixed(-8.0/65536.0,1,-nbitq), 
to_sfixed(-2628.0/65536.0,1,-nbitq), 
to_sfixed(469.0/65536.0,1,-nbitq), 
to_sfixed(-1746.0/65536.0,1,-nbitq), 
to_sfixed(-164.0/65536.0,1,-nbitq), 
to_sfixed(1589.0/65536.0,1,-nbitq), 
to_sfixed(634.0/65536.0,1,-nbitq), 
to_sfixed(3875.0/65536.0,1,-nbitq), 
to_sfixed(3750.0/65536.0,1,-nbitq), 
to_sfixed(846.0/65536.0,1,-nbitq), 
to_sfixed(817.0/65536.0,1,-nbitq), 
to_sfixed(-4078.0/65536.0,1,-nbitq), 
to_sfixed(2528.0/65536.0,1,-nbitq), 
to_sfixed(-3159.0/65536.0,1,-nbitq), 
to_sfixed(108.0/65536.0,1,-nbitq), 
to_sfixed(-2187.0/65536.0,1,-nbitq), 
to_sfixed(-832.0/65536.0,1,-nbitq), 
to_sfixed(2379.0/65536.0,1,-nbitq), 
to_sfixed(3799.0/65536.0,1,-nbitq), 
to_sfixed(-4918.0/65536.0,1,-nbitq), 
to_sfixed(3997.0/65536.0,1,-nbitq), 
to_sfixed(-2229.0/65536.0,1,-nbitq), 
to_sfixed(3094.0/65536.0,1,-nbitq), 
to_sfixed(4295.0/65536.0,1,-nbitq), 
to_sfixed(928.0/65536.0,1,-nbitq), 
to_sfixed(-154.0/65536.0,1,-nbitq), 
to_sfixed(-2301.0/65536.0,1,-nbitq), 
to_sfixed(675.0/65536.0,1,-nbitq), 
to_sfixed(-1793.0/65536.0,1,-nbitq), 
to_sfixed(9484.0/65536.0,1,-nbitq), 
to_sfixed(-1921.0/65536.0,1,-nbitq), 
to_sfixed(1516.0/65536.0,1,-nbitq), 
to_sfixed(1216.0/65536.0,1,-nbitq), 
to_sfixed(2997.0/65536.0,1,-nbitq), 
to_sfixed(2175.0/65536.0,1,-nbitq), 
to_sfixed(1706.0/65536.0,1,-nbitq), 
to_sfixed(-2292.0/65536.0,1,-nbitq), 
to_sfixed(1605.0/65536.0,1,-nbitq), 
to_sfixed(-1969.0/65536.0,1,-nbitq), 
to_sfixed(2968.0/65536.0,1,-nbitq), 
to_sfixed(-2104.0/65536.0,1,-nbitq), 
to_sfixed(598.0/65536.0,1,-nbitq), 
to_sfixed(-377.0/65536.0,1,-nbitq), 
to_sfixed(1822.0/65536.0,1,-nbitq), 
to_sfixed(-949.0/65536.0,1,-nbitq), 
to_sfixed(132.0/65536.0,1,-nbitq), 
to_sfixed(-1453.0/65536.0,1,-nbitq), 
to_sfixed(-2296.0/65536.0,1,-nbitq), 
to_sfixed(-4591.0/65536.0,1,-nbitq), 
to_sfixed(1116.0/65536.0,1,-nbitq), 
to_sfixed(-1568.0/65536.0,1,-nbitq), 
to_sfixed(8739.0/65536.0,1,-nbitq), 
to_sfixed(1842.0/65536.0,1,-nbitq), 
to_sfixed(1683.0/65536.0,1,-nbitq), 
to_sfixed(-954.0/65536.0,1,-nbitq), 
to_sfixed(-2539.0/65536.0,1,-nbitq), 
to_sfixed(-1076.0/65536.0,1,-nbitq), 
to_sfixed(678.0/65536.0,1,-nbitq), 
to_sfixed(494.0/65536.0,1,-nbitq), 
to_sfixed(2484.0/65536.0,1,-nbitq), 
to_sfixed(-1123.0/65536.0,1,-nbitq), 
to_sfixed(-1668.0/65536.0,1,-nbitq), 
to_sfixed(1055.0/65536.0,1,-nbitq), 
to_sfixed(-2584.0/65536.0,1,-nbitq), 
to_sfixed(-2242.0/65536.0,1,-nbitq), 
to_sfixed(-6080.0/65536.0,1,-nbitq), 
to_sfixed(-4758.0/65536.0,1,-nbitq), 
to_sfixed(64.0/65536.0,1,-nbitq), 
to_sfixed(-3951.0/65536.0,1,-nbitq), 
to_sfixed(345.0/65536.0,1,-nbitq), 
to_sfixed(591.0/65536.0,1,-nbitq), 
to_sfixed(2392.0/65536.0,1,-nbitq), 
to_sfixed(3165.0/65536.0,1,-nbitq), 
to_sfixed(-3126.0/65536.0,1,-nbitq), 
to_sfixed(12.0/65536.0,1,-nbitq), 
to_sfixed(-2570.0/65536.0,1,-nbitq), 
to_sfixed(-5228.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1130.0/65536.0,1,-nbitq), 
to_sfixed(-316.0/65536.0,1,-nbitq), 
to_sfixed(817.0/65536.0,1,-nbitq), 
to_sfixed(291.0/65536.0,1,-nbitq), 
to_sfixed(-1884.0/65536.0,1,-nbitq), 
to_sfixed(3263.0/65536.0,1,-nbitq), 
to_sfixed(-3409.0/65536.0,1,-nbitq), 
to_sfixed(3002.0/65536.0,1,-nbitq), 
to_sfixed(1893.0/65536.0,1,-nbitq), 
to_sfixed(-1232.0/65536.0,1,-nbitq), 
to_sfixed(2057.0/65536.0,1,-nbitq), 
to_sfixed(-1197.0/65536.0,1,-nbitq), 
to_sfixed(1704.0/65536.0,1,-nbitq), 
to_sfixed(-574.0/65536.0,1,-nbitq), 
to_sfixed(-1324.0/65536.0,1,-nbitq), 
to_sfixed(-1581.0/65536.0,1,-nbitq), 
to_sfixed(-674.0/65536.0,1,-nbitq), 
to_sfixed(1052.0/65536.0,1,-nbitq), 
to_sfixed(302.0/65536.0,1,-nbitq), 
to_sfixed(3044.0/65536.0,1,-nbitq), 
to_sfixed(-189.0/65536.0,1,-nbitq), 
to_sfixed(734.0/65536.0,1,-nbitq), 
to_sfixed(-1868.0/65536.0,1,-nbitq), 
to_sfixed(1748.0/65536.0,1,-nbitq), 
to_sfixed(76.0/65536.0,1,-nbitq), 
to_sfixed(4614.0/65536.0,1,-nbitq), 
to_sfixed(2215.0/65536.0,1,-nbitq), 
to_sfixed(2558.0/65536.0,1,-nbitq), 
to_sfixed(2287.0/65536.0,1,-nbitq), 
to_sfixed(1819.0/65536.0,1,-nbitq), 
to_sfixed(-78.0/65536.0,1,-nbitq), 
to_sfixed(1484.0/65536.0,1,-nbitq), 
to_sfixed(9184.0/65536.0,1,-nbitq), 
to_sfixed(1851.0/65536.0,1,-nbitq), 
to_sfixed(2606.0/65536.0,1,-nbitq), 
to_sfixed(1925.0/65536.0,1,-nbitq), 
to_sfixed(-806.0/65536.0,1,-nbitq), 
to_sfixed(4165.0/65536.0,1,-nbitq), 
to_sfixed(-1767.0/65536.0,1,-nbitq), 
to_sfixed(144.0/65536.0,1,-nbitq), 
to_sfixed(-1009.0/65536.0,1,-nbitq), 
to_sfixed(117.0/65536.0,1,-nbitq), 
to_sfixed(5424.0/65536.0,1,-nbitq), 
to_sfixed(-80.0/65536.0,1,-nbitq), 
to_sfixed(-687.0/65536.0,1,-nbitq), 
to_sfixed(-1146.0/65536.0,1,-nbitq), 
to_sfixed(-857.0/65536.0,1,-nbitq), 
to_sfixed(1302.0/65536.0,1,-nbitq), 
to_sfixed(2666.0/65536.0,1,-nbitq), 
to_sfixed(3237.0/65536.0,1,-nbitq), 
to_sfixed(-854.0/65536.0,1,-nbitq), 
to_sfixed(-6497.0/65536.0,1,-nbitq), 
to_sfixed(4755.0/65536.0,1,-nbitq), 
to_sfixed(-6412.0/65536.0,1,-nbitq), 
to_sfixed(8407.0/65536.0,1,-nbitq), 
to_sfixed(-1077.0/65536.0,1,-nbitq), 
to_sfixed(1549.0/65536.0,1,-nbitq), 
to_sfixed(-189.0/65536.0,1,-nbitq), 
to_sfixed(-170.0/65536.0,1,-nbitq), 
to_sfixed(-769.0/65536.0,1,-nbitq), 
to_sfixed(-1833.0/65536.0,1,-nbitq), 
to_sfixed(-463.0/65536.0,1,-nbitq), 
to_sfixed(829.0/65536.0,1,-nbitq), 
to_sfixed(-841.0/65536.0,1,-nbitq), 
to_sfixed(50.0/65536.0,1,-nbitq), 
to_sfixed(1232.0/65536.0,1,-nbitq), 
to_sfixed(-2322.0/65536.0,1,-nbitq), 
to_sfixed(-1739.0/65536.0,1,-nbitq), 
to_sfixed(-6546.0/65536.0,1,-nbitq), 
to_sfixed(-6655.0/65536.0,1,-nbitq), 
to_sfixed(4873.0/65536.0,1,-nbitq), 
to_sfixed(-7444.0/65536.0,1,-nbitq), 
to_sfixed(-1567.0/65536.0,1,-nbitq), 
to_sfixed(-1418.0/65536.0,1,-nbitq), 
to_sfixed(2163.0/65536.0,1,-nbitq), 
to_sfixed(2101.0/65536.0,1,-nbitq), 
to_sfixed(-4144.0/65536.0,1,-nbitq), 
to_sfixed(-2724.0/65536.0,1,-nbitq), 
to_sfixed(1493.0/65536.0,1,-nbitq), 
to_sfixed(-2492.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1310.0/65536.0,1,-nbitq), 
to_sfixed(2349.0/65536.0,1,-nbitq), 
to_sfixed(-363.0/65536.0,1,-nbitq), 
to_sfixed(-355.0/65536.0,1,-nbitq), 
to_sfixed(627.0/65536.0,1,-nbitq), 
to_sfixed(-1922.0/65536.0,1,-nbitq), 
to_sfixed(1669.0/65536.0,1,-nbitq), 
to_sfixed(1143.0/65536.0,1,-nbitq), 
to_sfixed(-1384.0/65536.0,1,-nbitq), 
to_sfixed(669.0/65536.0,1,-nbitq), 
to_sfixed(-3156.0/65536.0,1,-nbitq), 
to_sfixed(-1265.0/65536.0,1,-nbitq), 
to_sfixed(-1473.0/65536.0,1,-nbitq), 
to_sfixed(-3049.0/65536.0,1,-nbitq), 
to_sfixed(302.0/65536.0,1,-nbitq), 
to_sfixed(2449.0/65536.0,1,-nbitq), 
to_sfixed(-1435.0/65536.0,1,-nbitq), 
to_sfixed(-2800.0/65536.0,1,-nbitq), 
to_sfixed(-2654.0/65536.0,1,-nbitq), 
to_sfixed(-714.0/65536.0,1,-nbitq), 
to_sfixed(595.0/65536.0,1,-nbitq), 
to_sfixed(1243.0/65536.0,1,-nbitq), 
to_sfixed(1589.0/65536.0,1,-nbitq), 
to_sfixed(227.0/65536.0,1,-nbitq), 
to_sfixed(4328.0/65536.0,1,-nbitq), 
to_sfixed(3837.0/65536.0,1,-nbitq), 
to_sfixed(491.0/65536.0,1,-nbitq), 
to_sfixed(3080.0/65536.0,1,-nbitq), 
to_sfixed(-1873.0/65536.0,1,-nbitq), 
to_sfixed(3124.0/65536.0,1,-nbitq), 
to_sfixed(208.0/65536.0,1,-nbitq), 
to_sfixed(258.0/65536.0,1,-nbitq), 
to_sfixed(2402.0/65536.0,1,-nbitq), 
to_sfixed(4064.0/65536.0,1,-nbitq), 
to_sfixed(850.0/65536.0,1,-nbitq), 
to_sfixed(2643.0/65536.0,1,-nbitq), 
to_sfixed(1760.0/65536.0,1,-nbitq), 
to_sfixed(-411.0/65536.0,1,-nbitq), 
to_sfixed(94.0/65536.0,1,-nbitq), 
to_sfixed(2162.0/65536.0,1,-nbitq), 
to_sfixed(-3331.0/65536.0,1,-nbitq), 
to_sfixed(715.0/65536.0,1,-nbitq), 
to_sfixed(2004.0/65536.0,1,-nbitq), 
to_sfixed(1021.0/65536.0,1,-nbitq), 
to_sfixed(-1437.0/65536.0,1,-nbitq), 
to_sfixed(2875.0/65536.0,1,-nbitq), 
to_sfixed(870.0/65536.0,1,-nbitq), 
to_sfixed(-3259.0/65536.0,1,-nbitq), 
to_sfixed(3388.0/65536.0,1,-nbitq), 
to_sfixed(757.0/65536.0,1,-nbitq), 
to_sfixed(-1351.0/65536.0,1,-nbitq), 
to_sfixed(-5625.0/65536.0,1,-nbitq), 
to_sfixed(6476.0/65536.0,1,-nbitq), 
to_sfixed(-2967.0/65536.0,1,-nbitq), 
to_sfixed(4279.0/65536.0,1,-nbitq), 
to_sfixed(5318.0/65536.0,1,-nbitq), 
to_sfixed(412.0/65536.0,1,-nbitq), 
to_sfixed(-85.0/65536.0,1,-nbitq), 
to_sfixed(1359.0/65536.0,1,-nbitq), 
to_sfixed(-394.0/65536.0,1,-nbitq), 
to_sfixed(-2020.0/65536.0,1,-nbitq), 
to_sfixed(-339.0/65536.0,1,-nbitq), 
to_sfixed(-2126.0/65536.0,1,-nbitq), 
to_sfixed(1041.0/65536.0,1,-nbitq), 
to_sfixed(792.0/65536.0,1,-nbitq), 
to_sfixed(-1262.0/65536.0,1,-nbitq), 
to_sfixed(-3025.0/65536.0,1,-nbitq), 
to_sfixed(-2585.0/65536.0,1,-nbitq), 
to_sfixed(-6780.0/65536.0,1,-nbitq), 
to_sfixed(-3253.0/65536.0,1,-nbitq), 
to_sfixed(2293.0/65536.0,1,-nbitq), 
to_sfixed(-2899.0/65536.0,1,-nbitq), 
to_sfixed(-1986.0/65536.0,1,-nbitq), 
to_sfixed(1911.0/65536.0,1,-nbitq), 
to_sfixed(267.0/65536.0,1,-nbitq), 
to_sfixed(5541.0/65536.0,1,-nbitq), 
to_sfixed(-1338.0/65536.0,1,-nbitq), 
to_sfixed(260.0/65536.0,1,-nbitq), 
to_sfixed(-401.0/65536.0,1,-nbitq), 
to_sfixed(-1809.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-723.0/65536.0,1,-nbitq), 
to_sfixed(2045.0/65536.0,1,-nbitq), 
to_sfixed(-1014.0/65536.0,1,-nbitq), 
to_sfixed(1509.0/65536.0,1,-nbitq), 
to_sfixed(-2708.0/65536.0,1,-nbitq), 
to_sfixed(-2794.0/65536.0,1,-nbitq), 
to_sfixed(867.0/65536.0,1,-nbitq), 
to_sfixed(-2678.0/65536.0,1,-nbitq), 
to_sfixed(421.0/65536.0,1,-nbitq), 
to_sfixed(676.0/65536.0,1,-nbitq), 
to_sfixed(-3601.0/65536.0,1,-nbitq), 
to_sfixed(3374.0/65536.0,1,-nbitq), 
to_sfixed(3650.0/65536.0,1,-nbitq), 
to_sfixed(-1995.0/65536.0,1,-nbitq), 
to_sfixed(-1642.0/65536.0,1,-nbitq), 
to_sfixed(-2296.0/65536.0,1,-nbitq), 
to_sfixed(-2531.0/65536.0,1,-nbitq), 
to_sfixed(-1399.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(2323.0/65536.0,1,-nbitq), 
to_sfixed(635.0/65536.0,1,-nbitq), 
to_sfixed(-634.0/65536.0,1,-nbitq), 
to_sfixed(1399.0/65536.0,1,-nbitq), 
to_sfixed(1438.0/65536.0,1,-nbitq), 
to_sfixed(1654.0/65536.0,1,-nbitq), 
to_sfixed(-1007.0/65536.0,1,-nbitq), 
to_sfixed(3705.0/65536.0,1,-nbitq), 
to_sfixed(-2195.0/65536.0,1,-nbitq), 
to_sfixed(-2437.0/65536.0,1,-nbitq), 
to_sfixed(-2300.0/65536.0,1,-nbitq), 
to_sfixed(3072.0/65536.0,1,-nbitq), 
to_sfixed(2035.0/65536.0,1,-nbitq), 
to_sfixed(26.0/65536.0,1,-nbitq), 
to_sfixed(1486.0/65536.0,1,-nbitq), 
to_sfixed(1155.0/65536.0,1,-nbitq), 
to_sfixed(-2529.0/65536.0,1,-nbitq), 
to_sfixed(-1244.0/65536.0,1,-nbitq), 
to_sfixed(-1612.0/65536.0,1,-nbitq), 
to_sfixed(740.0/65536.0,1,-nbitq), 
to_sfixed(-1929.0/65536.0,1,-nbitq), 
to_sfixed(-2807.0/65536.0,1,-nbitq), 
to_sfixed(968.0/65536.0,1,-nbitq), 
to_sfixed(-1664.0/65536.0,1,-nbitq), 
to_sfixed(2744.0/65536.0,1,-nbitq), 
to_sfixed(2492.0/65536.0,1,-nbitq), 
to_sfixed(3584.0/65536.0,1,-nbitq), 
to_sfixed(-1033.0/65536.0,1,-nbitq), 
to_sfixed(1304.0/65536.0,1,-nbitq), 
to_sfixed(2991.0/65536.0,1,-nbitq), 
to_sfixed(337.0/65536.0,1,-nbitq), 
to_sfixed(2997.0/65536.0,1,-nbitq), 
to_sfixed(-6332.0/65536.0,1,-nbitq), 
to_sfixed(116.0/65536.0,1,-nbitq), 
to_sfixed(-5011.0/65536.0,1,-nbitq), 
to_sfixed(-913.0/65536.0,1,-nbitq), 
to_sfixed(1223.0/65536.0,1,-nbitq), 
to_sfixed(2395.0/65536.0,1,-nbitq), 
to_sfixed(-1699.0/65536.0,1,-nbitq), 
to_sfixed(-1508.0/65536.0,1,-nbitq), 
to_sfixed(3205.0/65536.0,1,-nbitq), 
to_sfixed(-3447.0/65536.0,1,-nbitq), 
to_sfixed(816.0/65536.0,1,-nbitq), 
to_sfixed(2500.0/65536.0,1,-nbitq), 
to_sfixed(2151.0/65536.0,1,-nbitq), 
to_sfixed(2377.0/65536.0,1,-nbitq), 
to_sfixed(3272.0/65536.0,1,-nbitq), 
to_sfixed(2006.0/65536.0,1,-nbitq), 
to_sfixed(-153.0/65536.0,1,-nbitq), 
to_sfixed(-4103.0/65536.0,1,-nbitq), 
to_sfixed(-841.0/65536.0,1,-nbitq), 
to_sfixed(-295.0/65536.0,1,-nbitq), 
to_sfixed(-2403.0/65536.0,1,-nbitq), 
to_sfixed(438.0/65536.0,1,-nbitq), 
to_sfixed(1415.0/65536.0,1,-nbitq), 
to_sfixed(438.0/65536.0,1,-nbitq), 
to_sfixed(-1165.0/65536.0,1,-nbitq), 
to_sfixed(1254.0/65536.0,1,-nbitq), 
to_sfixed(-83.0/65536.0,1,-nbitq), 
to_sfixed(-2066.0/65536.0,1,-nbitq), 
to_sfixed(3249.0/65536.0,1,-nbitq)  ), 
( to_sfixed(823.0/65536.0,1,-nbitq), 
to_sfixed(-1695.0/65536.0,1,-nbitq), 
to_sfixed(-386.0/65536.0,1,-nbitq), 
to_sfixed(-1978.0/65536.0,1,-nbitq), 
to_sfixed(133.0/65536.0,1,-nbitq), 
to_sfixed(984.0/65536.0,1,-nbitq), 
to_sfixed(-1418.0/65536.0,1,-nbitq), 
to_sfixed(-1082.0/65536.0,1,-nbitq), 
to_sfixed(-2234.0/65536.0,1,-nbitq), 
to_sfixed(2553.0/65536.0,1,-nbitq), 
to_sfixed(-1640.0/65536.0,1,-nbitq), 
to_sfixed(442.0/65536.0,1,-nbitq), 
to_sfixed(-927.0/65536.0,1,-nbitq), 
to_sfixed(-288.0/65536.0,1,-nbitq), 
to_sfixed(2333.0/65536.0,1,-nbitq), 
to_sfixed(233.0/65536.0,1,-nbitq), 
to_sfixed(-1629.0/65536.0,1,-nbitq), 
to_sfixed(-1026.0/65536.0,1,-nbitq), 
to_sfixed(-1505.0/65536.0,1,-nbitq), 
to_sfixed(1169.0/65536.0,1,-nbitq), 
to_sfixed(-3913.0/65536.0,1,-nbitq), 
to_sfixed(-681.0/65536.0,1,-nbitq), 
to_sfixed(-1668.0/65536.0,1,-nbitq), 
to_sfixed(1376.0/65536.0,1,-nbitq), 
to_sfixed(-1883.0/65536.0,1,-nbitq), 
to_sfixed(2599.0/65536.0,1,-nbitq), 
to_sfixed(-1628.0/65536.0,1,-nbitq), 
to_sfixed(3266.0/65536.0,1,-nbitq), 
to_sfixed(1638.0/65536.0,1,-nbitq), 
to_sfixed(-447.0/65536.0,1,-nbitq), 
to_sfixed(2917.0/65536.0,1,-nbitq), 
to_sfixed(-994.0/65536.0,1,-nbitq), 
to_sfixed(-1294.0/65536.0,1,-nbitq), 
to_sfixed(1018.0/65536.0,1,-nbitq), 
to_sfixed(2760.0/65536.0,1,-nbitq), 
to_sfixed(722.0/65536.0,1,-nbitq), 
to_sfixed(-3028.0/65536.0,1,-nbitq), 
to_sfixed(905.0/65536.0,1,-nbitq), 
to_sfixed(-1250.0/65536.0,1,-nbitq), 
to_sfixed(1552.0/65536.0,1,-nbitq), 
to_sfixed(1690.0/65536.0,1,-nbitq), 
to_sfixed(-2233.0/65536.0,1,-nbitq), 
to_sfixed(-4107.0/65536.0,1,-nbitq), 
to_sfixed(1002.0/65536.0,1,-nbitq), 
to_sfixed(-1407.0/65536.0,1,-nbitq), 
to_sfixed(3125.0/65536.0,1,-nbitq), 
to_sfixed(1904.0/65536.0,1,-nbitq), 
to_sfixed(833.0/65536.0,1,-nbitq), 
to_sfixed(891.0/65536.0,1,-nbitq), 
to_sfixed(80.0/65536.0,1,-nbitq), 
to_sfixed(-799.0/65536.0,1,-nbitq), 
to_sfixed(-2264.0/65536.0,1,-nbitq), 
to_sfixed(2978.0/65536.0,1,-nbitq), 
to_sfixed(575.0/65536.0,1,-nbitq), 
to_sfixed(2021.0/65536.0,1,-nbitq), 
to_sfixed(-2437.0/65536.0,1,-nbitq), 
to_sfixed(-219.0/65536.0,1,-nbitq), 
to_sfixed(785.0/65536.0,1,-nbitq), 
to_sfixed(-2886.0/65536.0,1,-nbitq), 
to_sfixed(4588.0/65536.0,1,-nbitq), 
to_sfixed(-680.0/65536.0,1,-nbitq), 
to_sfixed(-2567.0/65536.0,1,-nbitq), 
to_sfixed(560.0/65536.0,1,-nbitq), 
to_sfixed(-2508.0/65536.0,1,-nbitq), 
to_sfixed(-288.0/65536.0,1,-nbitq), 
to_sfixed(2413.0/65536.0,1,-nbitq), 
to_sfixed(-911.0/65536.0,1,-nbitq), 
to_sfixed(-1792.0/65536.0,1,-nbitq), 
to_sfixed(-3445.0/65536.0,1,-nbitq), 
to_sfixed(818.0/65536.0,1,-nbitq), 
to_sfixed(-1114.0/65536.0,1,-nbitq), 
to_sfixed(1787.0/65536.0,1,-nbitq), 
to_sfixed(-1738.0/65536.0,1,-nbitq), 
to_sfixed(-212.0/65536.0,1,-nbitq), 
to_sfixed(-3149.0/65536.0,1,-nbitq), 
to_sfixed(2843.0/65536.0,1,-nbitq), 
to_sfixed(-2230.0/65536.0,1,-nbitq), 
to_sfixed(4956.0/65536.0,1,-nbitq), 
to_sfixed(-1001.0/65536.0,1,-nbitq), 
to_sfixed(1293.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1706.0/65536.0,1,-nbitq), 
to_sfixed(-1724.0/65536.0,1,-nbitq), 
to_sfixed(1298.0/65536.0,1,-nbitq), 
to_sfixed(2001.0/65536.0,1,-nbitq), 
to_sfixed(-3167.0/65536.0,1,-nbitq), 
to_sfixed(-1132.0/65536.0,1,-nbitq), 
to_sfixed(1416.0/65536.0,1,-nbitq), 
to_sfixed(987.0/65536.0,1,-nbitq), 
to_sfixed(-67.0/65536.0,1,-nbitq), 
to_sfixed(1165.0/65536.0,1,-nbitq), 
to_sfixed(1910.0/65536.0,1,-nbitq), 
to_sfixed(-2548.0/65536.0,1,-nbitq), 
to_sfixed(3049.0/65536.0,1,-nbitq), 
to_sfixed(-2452.0/65536.0,1,-nbitq), 
to_sfixed(999.0/65536.0,1,-nbitq), 
to_sfixed(-1902.0/65536.0,1,-nbitq), 
to_sfixed(556.0/65536.0,1,-nbitq), 
to_sfixed(2087.0/65536.0,1,-nbitq), 
to_sfixed(-1153.0/65536.0,1,-nbitq), 
to_sfixed(200.0/65536.0,1,-nbitq), 
to_sfixed(398.0/65536.0,1,-nbitq), 
to_sfixed(2155.0/65536.0,1,-nbitq), 
to_sfixed(-2370.0/65536.0,1,-nbitq), 
to_sfixed(1098.0/65536.0,1,-nbitq), 
to_sfixed(3220.0/65536.0,1,-nbitq), 
to_sfixed(701.0/65536.0,1,-nbitq), 
to_sfixed(-3305.0/65536.0,1,-nbitq), 
to_sfixed(1354.0/65536.0,1,-nbitq), 
to_sfixed(1176.0/65536.0,1,-nbitq), 
to_sfixed(-70.0/65536.0,1,-nbitq), 
to_sfixed(-2219.0/65536.0,1,-nbitq), 
to_sfixed(-772.0/65536.0,1,-nbitq), 
to_sfixed(-1213.0/65536.0,1,-nbitq), 
to_sfixed(-1694.0/65536.0,1,-nbitq), 
to_sfixed(-2071.0/65536.0,1,-nbitq), 
to_sfixed(1433.0/65536.0,1,-nbitq), 
to_sfixed(-230.0/65536.0,1,-nbitq), 
to_sfixed(1885.0/65536.0,1,-nbitq), 
to_sfixed(1510.0/65536.0,1,-nbitq), 
to_sfixed(2756.0/65536.0,1,-nbitq), 
to_sfixed(-3305.0/65536.0,1,-nbitq), 
to_sfixed(-743.0/65536.0,1,-nbitq), 
to_sfixed(-3541.0/65536.0,1,-nbitq), 
to_sfixed(3127.0/65536.0,1,-nbitq), 
to_sfixed(581.0/65536.0,1,-nbitq), 
to_sfixed(425.0/65536.0,1,-nbitq), 
to_sfixed(-1846.0/65536.0,1,-nbitq), 
to_sfixed(2757.0/65536.0,1,-nbitq), 
to_sfixed(-809.0/65536.0,1,-nbitq), 
to_sfixed(3788.0/65536.0,1,-nbitq), 
to_sfixed(-1204.0/65536.0,1,-nbitq), 
to_sfixed(1089.0/65536.0,1,-nbitq), 
to_sfixed(-1694.0/65536.0,1,-nbitq), 
to_sfixed(-3321.0/65536.0,1,-nbitq), 
to_sfixed(1636.0/65536.0,1,-nbitq), 
to_sfixed(-682.0/65536.0,1,-nbitq), 
to_sfixed(2765.0/65536.0,1,-nbitq), 
to_sfixed(-2858.0/65536.0,1,-nbitq), 
to_sfixed(2203.0/65536.0,1,-nbitq), 
to_sfixed(2205.0/65536.0,1,-nbitq), 
to_sfixed(1767.0/65536.0,1,-nbitq), 
to_sfixed(-1660.0/65536.0,1,-nbitq), 
to_sfixed(-2645.0/65536.0,1,-nbitq), 
to_sfixed(1839.0/65536.0,1,-nbitq), 
to_sfixed(761.0/65536.0,1,-nbitq), 
to_sfixed(890.0/65536.0,1,-nbitq), 
to_sfixed(-561.0/65536.0,1,-nbitq), 
to_sfixed(1796.0/65536.0,1,-nbitq), 
to_sfixed(-2621.0/65536.0,1,-nbitq), 
to_sfixed(62.0/65536.0,1,-nbitq), 
to_sfixed(1452.0/65536.0,1,-nbitq), 
to_sfixed(-2555.0/65536.0,1,-nbitq), 
to_sfixed(1488.0/65536.0,1,-nbitq), 
to_sfixed(-1137.0/65536.0,1,-nbitq), 
to_sfixed(1096.0/65536.0,1,-nbitq), 
to_sfixed(-1712.0/65536.0,1,-nbitq), 
to_sfixed(472.0/65536.0,1,-nbitq), 
to_sfixed(115.0/65536.0,1,-nbitq), 
to_sfixed(1535.0/65536.0,1,-nbitq), 
to_sfixed(2115.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(157.0/65536.0,1,-nbitq), 
to_sfixed(-2516.0/65536.0,1,-nbitq), 
to_sfixed(2359.0/65536.0,1,-nbitq), 
to_sfixed(-1207.0/65536.0,1,-nbitq), 
to_sfixed(-1705.0/65536.0,1,-nbitq), 
to_sfixed(-4980.0/65536.0,1,-nbitq), 
to_sfixed(1753.0/65536.0,1,-nbitq), 
to_sfixed(2524.0/65536.0,1,-nbitq), 
to_sfixed(1466.0/65536.0,1,-nbitq), 
to_sfixed(1851.0/65536.0,1,-nbitq), 
to_sfixed(-3140.0/65536.0,1,-nbitq), 
to_sfixed(-1363.0/65536.0,1,-nbitq), 
to_sfixed(2426.0/65536.0,1,-nbitq), 
to_sfixed(2404.0/65536.0,1,-nbitq), 
to_sfixed(2700.0/65536.0,1,-nbitq), 
to_sfixed(193.0/65536.0,1,-nbitq), 
to_sfixed(671.0/65536.0,1,-nbitq), 
to_sfixed(-1682.0/65536.0,1,-nbitq), 
to_sfixed(1016.0/65536.0,1,-nbitq), 
to_sfixed(-2491.0/65536.0,1,-nbitq), 
to_sfixed(-1061.0/65536.0,1,-nbitq), 
to_sfixed(-454.0/65536.0,1,-nbitq), 
to_sfixed(1937.0/65536.0,1,-nbitq), 
to_sfixed(3128.0/65536.0,1,-nbitq), 
to_sfixed(-2315.0/65536.0,1,-nbitq), 
to_sfixed(-1138.0/65536.0,1,-nbitq), 
to_sfixed(-933.0/65536.0,1,-nbitq), 
to_sfixed(562.0/65536.0,1,-nbitq), 
to_sfixed(-2146.0/65536.0,1,-nbitq), 
to_sfixed(-2297.0/65536.0,1,-nbitq), 
to_sfixed(633.0/65536.0,1,-nbitq), 
to_sfixed(-580.0/65536.0,1,-nbitq), 
to_sfixed(-2332.0/65536.0,1,-nbitq), 
to_sfixed(-5359.0/65536.0,1,-nbitq), 
to_sfixed(-88.0/65536.0,1,-nbitq), 
to_sfixed(-1119.0/65536.0,1,-nbitq), 
to_sfixed(-2430.0/65536.0,1,-nbitq), 
to_sfixed(-1272.0/65536.0,1,-nbitq), 
to_sfixed(-1668.0/65536.0,1,-nbitq), 
to_sfixed(1601.0/65536.0,1,-nbitq), 
to_sfixed(-24.0/65536.0,1,-nbitq), 
to_sfixed(-2519.0/65536.0,1,-nbitq), 
to_sfixed(-3829.0/65536.0,1,-nbitq), 
to_sfixed(-1134.0/65536.0,1,-nbitq), 
to_sfixed(589.0/65536.0,1,-nbitq), 
to_sfixed(114.0/65536.0,1,-nbitq), 
to_sfixed(-1340.0/65536.0,1,-nbitq), 
to_sfixed(-149.0/65536.0,1,-nbitq), 
to_sfixed(-1104.0/65536.0,1,-nbitq), 
to_sfixed(4000.0/65536.0,1,-nbitq), 
to_sfixed(822.0/65536.0,1,-nbitq), 
to_sfixed(747.0/65536.0,1,-nbitq), 
to_sfixed(378.0/65536.0,1,-nbitq), 
to_sfixed(498.0/65536.0,1,-nbitq), 
to_sfixed(-132.0/65536.0,1,-nbitq), 
to_sfixed(-806.0/65536.0,1,-nbitq), 
to_sfixed(1936.0/65536.0,1,-nbitq), 
to_sfixed(2305.0/65536.0,1,-nbitq), 
to_sfixed(695.0/65536.0,1,-nbitq), 
to_sfixed(2494.0/65536.0,1,-nbitq), 
to_sfixed(-3996.0/65536.0,1,-nbitq), 
to_sfixed(-2529.0/65536.0,1,-nbitq), 
to_sfixed(1721.0/65536.0,1,-nbitq), 
to_sfixed(-755.0/65536.0,1,-nbitq), 
to_sfixed(1977.0/65536.0,1,-nbitq), 
to_sfixed(3759.0/65536.0,1,-nbitq), 
to_sfixed(-1083.0/65536.0,1,-nbitq), 
to_sfixed(-3751.0/65536.0,1,-nbitq), 
to_sfixed(168.0/65536.0,1,-nbitq), 
to_sfixed(-444.0/65536.0,1,-nbitq), 
to_sfixed(-1353.0/65536.0,1,-nbitq), 
to_sfixed(101.0/65536.0,1,-nbitq), 
to_sfixed(604.0/65536.0,1,-nbitq), 
to_sfixed(-1608.0/65536.0,1,-nbitq), 
to_sfixed(19.0/65536.0,1,-nbitq), 
to_sfixed(1089.0/65536.0,1,-nbitq), 
to_sfixed(-1900.0/65536.0,1,-nbitq), 
to_sfixed(2182.0/65536.0,1,-nbitq), 
to_sfixed(-2555.0/65536.0,1,-nbitq), 
to_sfixed(1370.0/65536.0,1,-nbitq)  ), 
( to_sfixed(891.0/65536.0,1,-nbitq), 
to_sfixed(-339.0/65536.0,1,-nbitq), 
to_sfixed(-999.0/65536.0,1,-nbitq), 
to_sfixed(-4601.0/65536.0,1,-nbitq), 
to_sfixed(-324.0/65536.0,1,-nbitq), 
to_sfixed(-3529.0/65536.0,1,-nbitq), 
to_sfixed(115.0/65536.0,1,-nbitq), 
to_sfixed(2503.0/65536.0,1,-nbitq), 
to_sfixed(-458.0/65536.0,1,-nbitq), 
to_sfixed(-2252.0/65536.0,1,-nbitq), 
to_sfixed(-2618.0/65536.0,1,-nbitq), 
to_sfixed(1687.0/65536.0,1,-nbitq), 
to_sfixed(-2767.0/65536.0,1,-nbitq), 
to_sfixed(548.0/65536.0,1,-nbitq), 
to_sfixed(-2435.0/65536.0,1,-nbitq), 
to_sfixed(291.0/65536.0,1,-nbitq), 
to_sfixed(-1474.0/65536.0,1,-nbitq), 
to_sfixed(1530.0/65536.0,1,-nbitq), 
to_sfixed(38.0/65536.0,1,-nbitq), 
to_sfixed(-56.0/65536.0,1,-nbitq), 
to_sfixed(-3512.0/65536.0,1,-nbitq), 
to_sfixed(-417.0/65536.0,1,-nbitq), 
to_sfixed(1100.0/65536.0,1,-nbitq), 
to_sfixed(485.0/65536.0,1,-nbitq), 
to_sfixed(435.0/65536.0,1,-nbitq), 
to_sfixed(2315.0/65536.0,1,-nbitq), 
to_sfixed(-4459.0/65536.0,1,-nbitq), 
to_sfixed(-2490.0/65536.0,1,-nbitq), 
to_sfixed(430.0/65536.0,1,-nbitq), 
to_sfixed(292.0/65536.0,1,-nbitq), 
to_sfixed(1988.0/65536.0,1,-nbitq), 
to_sfixed(143.0/65536.0,1,-nbitq), 
to_sfixed(-1108.0/65536.0,1,-nbitq), 
to_sfixed(-2661.0/65536.0,1,-nbitq), 
to_sfixed(2417.0/65536.0,1,-nbitq), 
to_sfixed(-2345.0/65536.0,1,-nbitq), 
to_sfixed(669.0/65536.0,1,-nbitq), 
to_sfixed(235.0/65536.0,1,-nbitq), 
to_sfixed(443.0/65536.0,1,-nbitq), 
to_sfixed(2665.0/65536.0,1,-nbitq), 
to_sfixed(678.0/65536.0,1,-nbitq), 
to_sfixed(-346.0/65536.0,1,-nbitq), 
to_sfixed(-2988.0/65536.0,1,-nbitq), 
to_sfixed(3103.0/65536.0,1,-nbitq), 
to_sfixed(-2099.0/65536.0,1,-nbitq), 
to_sfixed(1956.0/65536.0,1,-nbitq), 
to_sfixed(3117.0/65536.0,1,-nbitq), 
to_sfixed(519.0/65536.0,1,-nbitq), 
to_sfixed(2302.0/65536.0,1,-nbitq), 
to_sfixed(970.0/65536.0,1,-nbitq), 
to_sfixed(699.0/65536.0,1,-nbitq), 
to_sfixed(2423.0/65536.0,1,-nbitq), 
to_sfixed(2824.0/65536.0,1,-nbitq), 
to_sfixed(-591.0/65536.0,1,-nbitq), 
to_sfixed(-1623.0/65536.0,1,-nbitq), 
to_sfixed(1564.0/65536.0,1,-nbitq), 
to_sfixed(313.0/65536.0,1,-nbitq), 
to_sfixed(-1044.0/65536.0,1,-nbitq), 
to_sfixed(1781.0/65536.0,1,-nbitq), 
to_sfixed(1593.0/65536.0,1,-nbitq), 
to_sfixed(709.0/65536.0,1,-nbitq), 
to_sfixed(2542.0/65536.0,1,-nbitq), 
to_sfixed(2418.0/65536.0,1,-nbitq), 
to_sfixed(-1441.0/65536.0,1,-nbitq), 
to_sfixed(1754.0/65536.0,1,-nbitq), 
to_sfixed(-595.0/65536.0,1,-nbitq), 
to_sfixed(2752.0/65536.0,1,-nbitq), 
to_sfixed(-2325.0/65536.0,1,-nbitq), 
to_sfixed(991.0/65536.0,1,-nbitq), 
to_sfixed(-838.0/65536.0,1,-nbitq), 
to_sfixed(1592.0/65536.0,1,-nbitq), 
to_sfixed(749.0/65536.0,1,-nbitq), 
to_sfixed(1493.0/65536.0,1,-nbitq), 
to_sfixed(604.0/65536.0,1,-nbitq), 
to_sfixed(2748.0/65536.0,1,-nbitq), 
to_sfixed(1939.0/65536.0,1,-nbitq), 
to_sfixed(1030.0/65536.0,1,-nbitq), 
to_sfixed(4611.0/65536.0,1,-nbitq), 
to_sfixed(-1895.0/65536.0,1,-nbitq), 
to_sfixed(1526.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3148.0/65536.0,1,-nbitq), 
to_sfixed(974.0/65536.0,1,-nbitq), 
to_sfixed(-1194.0/65536.0,1,-nbitq), 
to_sfixed(-4423.0/65536.0,1,-nbitq), 
to_sfixed(-2240.0/65536.0,1,-nbitq), 
to_sfixed(-568.0/65536.0,1,-nbitq), 
to_sfixed(-1494.0/65536.0,1,-nbitq), 
to_sfixed(-25.0/65536.0,1,-nbitq), 
to_sfixed(388.0/65536.0,1,-nbitq), 
to_sfixed(749.0/65536.0,1,-nbitq), 
to_sfixed(-3261.0/65536.0,1,-nbitq), 
to_sfixed(-1916.0/65536.0,1,-nbitq), 
to_sfixed(-1037.0/65536.0,1,-nbitq), 
to_sfixed(1623.0/65536.0,1,-nbitq), 
to_sfixed(-4888.0/65536.0,1,-nbitq), 
to_sfixed(-1929.0/65536.0,1,-nbitq), 
to_sfixed(2671.0/65536.0,1,-nbitq), 
to_sfixed(2454.0/65536.0,1,-nbitq), 
to_sfixed(-2664.0/65536.0,1,-nbitq), 
to_sfixed(-562.0/65536.0,1,-nbitq), 
to_sfixed(-1480.0/65536.0,1,-nbitq), 
to_sfixed(2029.0/65536.0,1,-nbitq), 
to_sfixed(3079.0/65536.0,1,-nbitq), 
to_sfixed(1699.0/65536.0,1,-nbitq), 
to_sfixed(1132.0/65536.0,1,-nbitq), 
to_sfixed(-1746.0/65536.0,1,-nbitq), 
to_sfixed(-5363.0/65536.0,1,-nbitq), 
to_sfixed(-1731.0/65536.0,1,-nbitq), 
to_sfixed(-2475.0/65536.0,1,-nbitq), 
to_sfixed(-3246.0/65536.0,1,-nbitq), 
to_sfixed(-2282.0/65536.0,1,-nbitq), 
to_sfixed(-1992.0/65536.0,1,-nbitq), 
to_sfixed(-1409.0/65536.0,1,-nbitq), 
to_sfixed(263.0/65536.0,1,-nbitq), 
to_sfixed(2615.0/65536.0,1,-nbitq), 
to_sfixed(2842.0/65536.0,1,-nbitq), 
to_sfixed(1006.0/65536.0,1,-nbitq), 
to_sfixed(1233.0/65536.0,1,-nbitq), 
to_sfixed(2728.0/65536.0,1,-nbitq), 
to_sfixed(19.0/65536.0,1,-nbitq), 
to_sfixed(-3125.0/65536.0,1,-nbitq), 
to_sfixed(-1240.0/65536.0,1,-nbitq), 
to_sfixed(-3900.0/65536.0,1,-nbitq), 
to_sfixed(21.0/65536.0,1,-nbitq), 
to_sfixed(-641.0/65536.0,1,-nbitq), 
to_sfixed(54.0/65536.0,1,-nbitq), 
to_sfixed(1395.0/65536.0,1,-nbitq), 
to_sfixed(-79.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(-989.0/65536.0,1,-nbitq), 
to_sfixed(-736.0/65536.0,1,-nbitq), 
to_sfixed(-1563.0/65536.0,1,-nbitq), 
to_sfixed(126.0/65536.0,1,-nbitq), 
to_sfixed(-2802.0/65536.0,1,-nbitq), 
to_sfixed(10.0/65536.0,1,-nbitq), 
to_sfixed(1444.0/65536.0,1,-nbitq), 
to_sfixed(-846.0/65536.0,1,-nbitq), 
to_sfixed(4564.0/65536.0,1,-nbitq), 
to_sfixed(2867.0/65536.0,1,-nbitq), 
to_sfixed(4050.0/65536.0,1,-nbitq), 
to_sfixed(-722.0/65536.0,1,-nbitq), 
to_sfixed(-2677.0/65536.0,1,-nbitq), 
to_sfixed(-1687.0/65536.0,1,-nbitq), 
to_sfixed(-421.0/65536.0,1,-nbitq), 
to_sfixed(-2104.0/65536.0,1,-nbitq), 
to_sfixed(1569.0/65536.0,1,-nbitq), 
to_sfixed(2158.0/65536.0,1,-nbitq), 
to_sfixed(-758.0/65536.0,1,-nbitq), 
to_sfixed(542.0/65536.0,1,-nbitq), 
to_sfixed(2093.0/65536.0,1,-nbitq), 
to_sfixed(971.0/65536.0,1,-nbitq), 
to_sfixed(-1437.0/65536.0,1,-nbitq), 
to_sfixed(131.0/65536.0,1,-nbitq), 
to_sfixed(-1556.0/65536.0,1,-nbitq), 
to_sfixed(2191.0/65536.0,1,-nbitq), 
to_sfixed(1799.0/65536.0,1,-nbitq), 
to_sfixed(723.0/65536.0,1,-nbitq), 
to_sfixed(1665.0/65536.0,1,-nbitq), 
to_sfixed(2115.0/65536.0,1,-nbitq), 
to_sfixed(1737.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-967.0/65536.0,1,-nbitq), 
to_sfixed(-2275.0/65536.0,1,-nbitq), 
to_sfixed(-6346.0/65536.0,1,-nbitq), 
to_sfixed(-2214.0/65536.0,1,-nbitq), 
to_sfixed(3321.0/65536.0,1,-nbitq), 
to_sfixed(-2330.0/65536.0,1,-nbitq), 
to_sfixed(750.0/65536.0,1,-nbitq), 
to_sfixed(-1940.0/65536.0,1,-nbitq), 
to_sfixed(-2161.0/65536.0,1,-nbitq), 
to_sfixed(1376.0/65536.0,1,-nbitq), 
to_sfixed(-4283.0/65536.0,1,-nbitq), 
to_sfixed(4398.0/65536.0,1,-nbitq), 
to_sfixed(-1245.0/65536.0,1,-nbitq), 
to_sfixed(5468.0/65536.0,1,-nbitq), 
to_sfixed(-2254.0/65536.0,1,-nbitq), 
to_sfixed(221.0/65536.0,1,-nbitq), 
to_sfixed(-2468.0/65536.0,1,-nbitq), 
to_sfixed(-1059.0/65536.0,1,-nbitq), 
to_sfixed(-4319.0/65536.0,1,-nbitq), 
to_sfixed(3409.0/65536.0,1,-nbitq), 
to_sfixed(534.0/65536.0,1,-nbitq), 
to_sfixed(2104.0/65536.0,1,-nbitq), 
to_sfixed(2084.0/65536.0,1,-nbitq), 
to_sfixed(-5180.0/65536.0,1,-nbitq), 
to_sfixed(-2516.0/65536.0,1,-nbitq), 
to_sfixed(-8208.0/65536.0,1,-nbitq), 
to_sfixed(-1015.0/65536.0,1,-nbitq), 
to_sfixed(-1245.0/65536.0,1,-nbitq), 
to_sfixed(-3843.0/65536.0,1,-nbitq), 
to_sfixed(-629.0/65536.0,1,-nbitq), 
to_sfixed(1187.0/65536.0,1,-nbitq), 
to_sfixed(-2592.0/65536.0,1,-nbitq), 
to_sfixed(-2103.0/65536.0,1,-nbitq), 
to_sfixed(5993.0/65536.0,1,-nbitq), 
to_sfixed(2213.0/65536.0,1,-nbitq), 
to_sfixed(2232.0/65536.0,1,-nbitq), 
to_sfixed(-1193.0/65536.0,1,-nbitq), 
to_sfixed(-2340.0/65536.0,1,-nbitq), 
to_sfixed(2284.0/65536.0,1,-nbitq), 
to_sfixed(-116.0/65536.0,1,-nbitq), 
to_sfixed(-815.0/65536.0,1,-nbitq), 
to_sfixed(-2812.0/65536.0,1,-nbitq), 
to_sfixed(349.0/65536.0,1,-nbitq), 
to_sfixed(3085.0/65536.0,1,-nbitq), 
to_sfixed(514.0/65536.0,1,-nbitq), 
to_sfixed(-1704.0/65536.0,1,-nbitq), 
to_sfixed(1872.0/65536.0,1,-nbitq), 
to_sfixed(-3534.0/65536.0,1,-nbitq), 
to_sfixed(3785.0/65536.0,1,-nbitq), 
to_sfixed(4861.0/65536.0,1,-nbitq), 
to_sfixed(3074.0/65536.0,1,-nbitq), 
to_sfixed(-2747.0/65536.0,1,-nbitq), 
to_sfixed(-1374.0/65536.0,1,-nbitq), 
to_sfixed(-4008.0/65536.0,1,-nbitq), 
to_sfixed(385.0/65536.0,1,-nbitq), 
to_sfixed(-2814.0/65536.0,1,-nbitq), 
to_sfixed(-2413.0/65536.0,1,-nbitq), 
to_sfixed(4644.0/65536.0,1,-nbitq), 
to_sfixed(116.0/65536.0,1,-nbitq), 
to_sfixed(2127.0/65536.0,1,-nbitq), 
to_sfixed(-438.0/65536.0,1,-nbitq), 
to_sfixed(-295.0/65536.0,1,-nbitq), 
to_sfixed(2941.0/65536.0,1,-nbitq), 
to_sfixed(-997.0/65536.0,1,-nbitq), 
to_sfixed(2392.0/65536.0,1,-nbitq), 
to_sfixed(-1406.0/65536.0,1,-nbitq), 
to_sfixed(445.0/65536.0,1,-nbitq), 
to_sfixed(-2361.0/65536.0,1,-nbitq), 
to_sfixed(2512.0/65536.0,1,-nbitq), 
to_sfixed(2783.0/65536.0,1,-nbitq), 
to_sfixed(-1600.0/65536.0,1,-nbitq), 
to_sfixed(4243.0/65536.0,1,-nbitq), 
to_sfixed(-98.0/65536.0,1,-nbitq), 
to_sfixed(1375.0/65536.0,1,-nbitq), 
to_sfixed(-1622.0/65536.0,1,-nbitq), 
to_sfixed(2231.0/65536.0,1,-nbitq), 
to_sfixed(2297.0/65536.0,1,-nbitq), 
to_sfixed(-29.0/65536.0,1,-nbitq), 
to_sfixed(2485.0/65536.0,1,-nbitq), 
to_sfixed(-600.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2067.0/65536.0,1,-nbitq), 
to_sfixed(-3636.0/65536.0,1,-nbitq), 
to_sfixed(-2144.0/65536.0,1,-nbitq), 
to_sfixed(-2706.0/65536.0,1,-nbitq), 
to_sfixed(5318.0/65536.0,1,-nbitq), 
to_sfixed(-1322.0/65536.0,1,-nbitq), 
to_sfixed(-797.0/65536.0,1,-nbitq), 
to_sfixed(-2873.0/65536.0,1,-nbitq), 
to_sfixed(-634.0/65536.0,1,-nbitq), 
to_sfixed(-558.0/65536.0,1,-nbitq), 
to_sfixed(-2935.0/65536.0,1,-nbitq), 
to_sfixed(7154.0/65536.0,1,-nbitq), 
to_sfixed(1686.0/65536.0,1,-nbitq), 
to_sfixed(5580.0/65536.0,1,-nbitq), 
to_sfixed(2811.0/65536.0,1,-nbitq), 
to_sfixed(-1244.0/65536.0,1,-nbitq), 
to_sfixed(-2810.0/65536.0,1,-nbitq), 
to_sfixed(-5354.0/65536.0,1,-nbitq), 
to_sfixed(-4890.0/65536.0,1,-nbitq), 
to_sfixed(1633.0/65536.0,1,-nbitq), 
to_sfixed(-5318.0/65536.0,1,-nbitq), 
to_sfixed(-1413.0/65536.0,1,-nbitq), 
to_sfixed(1669.0/65536.0,1,-nbitq), 
to_sfixed(-177.0/65536.0,1,-nbitq), 
to_sfixed(-1852.0/65536.0,1,-nbitq), 
to_sfixed(30.0/65536.0,1,-nbitq), 
to_sfixed(-1838.0/65536.0,1,-nbitq), 
to_sfixed(1323.0/65536.0,1,-nbitq), 
to_sfixed(-2468.0/65536.0,1,-nbitq), 
to_sfixed(1941.0/65536.0,1,-nbitq), 
to_sfixed(-895.0/65536.0,1,-nbitq), 
to_sfixed(1946.0/65536.0,1,-nbitq), 
to_sfixed(2759.0/65536.0,1,-nbitq), 
to_sfixed(3299.0/65536.0,1,-nbitq), 
to_sfixed(550.0/65536.0,1,-nbitq), 
to_sfixed(1426.0/65536.0,1,-nbitq), 
to_sfixed(-277.0/65536.0,1,-nbitq), 
to_sfixed(-4552.0/65536.0,1,-nbitq), 
to_sfixed(4100.0/65536.0,1,-nbitq), 
to_sfixed(-828.0/65536.0,1,-nbitq), 
to_sfixed(-3229.0/65536.0,1,-nbitq), 
to_sfixed(2003.0/65536.0,1,-nbitq), 
to_sfixed(5389.0/65536.0,1,-nbitq), 
to_sfixed(3109.0/65536.0,1,-nbitq), 
to_sfixed(-493.0/65536.0,1,-nbitq), 
to_sfixed(1028.0/65536.0,1,-nbitq), 
to_sfixed(1286.0/65536.0,1,-nbitq), 
to_sfixed(-237.0/65536.0,1,-nbitq), 
to_sfixed(3890.0/65536.0,1,-nbitq), 
to_sfixed(2106.0/65536.0,1,-nbitq), 
to_sfixed(1824.0/65536.0,1,-nbitq), 
to_sfixed(-936.0/65536.0,1,-nbitq), 
to_sfixed(1539.0/65536.0,1,-nbitq), 
to_sfixed(-2212.0/65536.0,1,-nbitq), 
to_sfixed(-2873.0/65536.0,1,-nbitq), 
to_sfixed(1980.0/65536.0,1,-nbitq), 
to_sfixed(-1583.0/65536.0,1,-nbitq), 
to_sfixed(3671.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(-625.0/65536.0,1,-nbitq), 
to_sfixed(-1245.0/65536.0,1,-nbitq), 
to_sfixed(-2642.0/65536.0,1,-nbitq), 
to_sfixed(742.0/65536.0,1,-nbitq), 
to_sfixed(189.0/65536.0,1,-nbitq), 
to_sfixed(2920.0/65536.0,1,-nbitq), 
to_sfixed(-977.0/65536.0,1,-nbitq), 
to_sfixed(1436.0/65536.0,1,-nbitq), 
to_sfixed(-552.0/65536.0,1,-nbitq), 
to_sfixed(-678.0/65536.0,1,-nbitq), 
to_sfixed(2378.0/65536.0,1,-nbitq), 
to_sfixed(1054.0/65536.0,1,-nbitq), 
to_sfixed(562.0/65536.0,1,-nbitq), 
to_sfixed(-1504.0/65536.0,1,-nbitq), 
to_sfixed(87.0/65536.0,1,-nbitq), 
to_sfixed(-754.0/65536.0,1,-nbitq), 
to_sfixed(-882.0/65536.0,1,-nbitq), 
to_sfixed(4578.0/65536.0,1,-nbitq), 
to_sfixed(-540.0/65536.0,1,-nbitq), 
to_sfixed(-729.0/65536.0,1,-nbitq), 
to_sfixed(-2354.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1760.0/65536.0,1,-nbitq), 
to_sfixed(-3127.0/65536.0,1,-nbitq), 
to_sfixed(2066.0/65536.0,1,-nbitq), 
to_sfixed(-849.0/65536.0,1,-nbitq), 
to_sfixed(-103.0/65536.0,1,-nbitq), 
to_sfixed(-2352.0/65536.0,1,-nbitq), 
to_sfixed(735.0/65536.0,1,-nbitq), 
to_sfixed(-891.0/65536.0,1,-nbitq), 
to_sfixed(-2407.0/65536.0,1,-nbitq), 
to_sfixed(-1067.0/65536.0,1,-nbitq), 
to_sfixed(-5322.0/65536.0,1,-nbitq), 
to_sfixed(9188.0/65536.0,1,-nbitq), 
to_sfixed(-2783.0/65536.0,1,-nbitq), 
to_sfixed(3758.0/65536.0,1,-nbitq), 
to_sfixed(2379.0/65536.0,1,-nbitq), 
to_sfixed(-196.0/65536.0,1,-nbitq), 
to_sfixed(-1868.0/65536.0,1,-nbitq), 
to_sfixed(-3590.0/65536.0,1,-nbitq), 
to_sfixed(439.0/65536.0,1,-nbitq), 
to_sfixed(19.0/65536.0,1,-nbitq), 
to_sfixed(-6401.0/65536.0,1,-nbitq), 
to_sfixed(1065.0/65536.0,1,-nbitq), 
to_sfixed(4050.0/65536.0,1,-nbitq), 
to_sfixed(-934.0/65536.0,1,-nbitq), 
to_sfixed(-2745.0/65536.0,1,-nbitq), 
to_sfixed(-3645.0/65536.0,1,-nbitq), 
to_sfixed(27.0/65536.0,1,-nbitq), 
to_sfixed(-1849.0/65536.0,1,-nbitq), 
to_sfixed(-3127.0/65536.0,1,-nbitq), 
to_sfixed(591.0/65536.0,1,-nbitq), 
to_sfixed(-781.0/65536.0,1,-nbitq), 
to_sfixed(1171.0/65536.0,1,-nbitq), 
to_sfixed(-1006.0/65536.0,1,-nbitq), 
to_sfixed(10301.0/65536.0,1,-nbitq), 
to_sfixed(-4537.0/65536.0,1,-nbitq), 
to_sfixed(2028.0/65536.0,1,-nbitq), 
to_sfixed(-5118.0/65536.0,1,-nbitq), 
to_sfixed(3492.0/65536.0,1,-nbitq), 
to_sfixed(2884.0/65536.0,1,-nbitq), 
to_sfixed(-4380.0/65536.0,1,-nbitq), 
to_sfixed(-3224.0/65536.0,1,-nbitq), 
to_sfixed(287.0/65536.0,1,-nbitq), 
to_sfixed(7140.0/65536.0,1,-nbitq), 
to_sfixed(3062.0/65536.0,1,-nbitq), 
to_sfixed(-198.0/65536.0,1,-nbitq), 
to_sfixed(-1767.0/65536.0,1,-nbitq), 
to_sfixed(728.0/65536.0,1,-nbitq), 
to_sfixed(-4794.0/65536.0,1,-nbitq), 
to_sfixed(387.0/65536.0,1,-nbitq), 
to_sfixed(4087.0/65536.0,1,-nbitq), 
to_sfixed(-320.0/65536.0,1,-nbitq), 
to_sfixed(-1290.0/65536.0,1,-nbitq), 
to_sfixed(2517.0/65536.0,1,-nbitq), 
to_sfixed(-911.0/65536.0,1,-nbitq), 
to_sfixed(211.0/65536.0,1,-nbitq), 
to_sfixed(-3714.0/65536.0,1,-nbitq), 
to_sfixed(-836.0/65536.0,1,-nbitq), 
to_sfixed(-1752.0/65536.0,1,-nbitq), 
to_sfixed(2513.0/65536.0,1,-nbitq), 
to_sfixed(2325.0/65536.0,1,-nbitq), 
to_sfixed(-2208.0/65536.0,1,-nbitq), 
to_sfixed(-3167.0/65536.0,1,-nbitq), 
to_sfixed(-813.0/65536.0,1,-nbitq), 
to_sfixed(1290.0/65536.0,1,-nbitq), 
to_sfixed(1070.0/65536.0,1,-nbitq), 
to_sfixed(362.0/65536.0,1,-nbitq), 
to_sfixed(-3624.0/65536.0,1,-nbitq), 
to_sfixed(4047.0/65536.0,1,-nbitq), 
to_sfixed(1371.0/65536.0,1,-nbitq), 
to_sfixed(2844.0/65536.0,1,-nbitq), 
to_sfixed(1279.0/65536.0,1,-nbitq), 
to_sfixed(3282.0/65536.0,1,-nbitq), 
to_sfixed(1796.0/65536.0,1,-nbitq), 
to_sfixed(2137.0/65536.0,1,-nbitq), 
to_sfixed(-2269.0/65536.0,1,-nbitq), 
to_sfixed(3667.0/65536.0,1,-nbitq), 
to_sfixed(3857.0/65536.0,1,-nbitq), 
to_sfixed(-803.0/65536.0,1,-nbitq), 
to_sfixed(2149.0/65536.0,1,-nbitq), 
to_sfixed(-1666.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1120.0/65536.0,1,-nbitq), 
to_sfixed(741.0/65536.0,1,-nbitq), 
to_sfixed(2973.0/65536.0,1,-nbitq), 
to_sfixed(-3154.0/65536.0,1,-nbitq), 
to_sfixed(-5300.0/65536.0,1,-nbitq), 
to_sfixed(2555.0/65536.0,1,-nbitq), 
to_sfixed(1565.0/65536.0,1,-nbitq), 
to_sfixed(4385.0/65536.0,1,-nbitq), 
to_sfixed(1479.0/65536.0,1,-nbitq), 
to_sfixed(-379.0/65536.0,1,-nbitq), 
to_sfixed(-3198.0/65536.0,1,-nbitq), 
to_sfixed(8113.0/65536.0,1,-nbitq), 
to_sfixed(1577.0/65536.0,1,-nbitq), 
to_sfixed(4142.0/65536.0,1,-nbitq), 
to_sfixed(2531.0/65536.0,1,-nbitq), 
to_sfixed(232.0/65536.0,1,-nbitq), 
to_sfixed(2991.0/65536.0,1,-nbitq), 
to_sfixed(1184.0/65536.0,1,-nbitq), 
to_sfixed(-503.0/65536.0,1,-nbitq), 
to_sfixed(-2468.0/65536.0,1,-nbitq), 
to_sfixed(-6199.0/65536.0,1,-nbitq), 
to_sfixed(-4105.0/65536.0,1,-nbitq), 
to_sfixed(570.0/65536.0,1,-nbitq), 
to_sfixed(-4846.0/65536.0,1,-nbitq), 
to_sfixed(-145.0/65536.0,1,-nbitq), 
to_sfixed(-7401.0/65536.0,1,-nbitq), 
to_sfixed(-5663.0/65536.0,1,-nbitq), 
to_sfixed(291.0/65536.0,1,-nbitq), 
to_sfixed(166.0/65536.0,1,-nbitq), 
to_sfixed(-2442.0/65536.0,1,-nbitq), 
to_sfixed(978.0/65536.0,1,-nbitq), 
to_sfixed(-381.0/65536.0,1,-nbitq), 
to_sfixed(2729.0/65536.0,1,-nbitq), 
to_sfixed(9552.0/65536.0,1,-nbitq), 
to_sfixed(-2793.0/65536.0,1,-nbitq), 
to_sfixed(-1182.0/65536.0,1,-nbitq), 
to_sfixed(-382.0/65536.0,1,-nbitq), 
to_sfixed(4648.0/65536.0,1,-nbitq), 
to_sfixed(2543.0/65536.0,1,-nbitq), 
to_sfixed(-937.0/65536.0,1,-nbitq), 
to_sfixed(-4423.0/65536.0,1,-nbitq), 
to_sfixed(1481.0/65536.0,1,-nbitq), 
to_sfixed(9164.0/65536.0,1,-nbitq), 
to_sfixed(5086.0/65536.0,1,-nbitq), 
to_sfixed(-1075.0/65536.0,1,-nbitq), 
to_sfixed(-6106.0/65536.0,1,-nbitq), 
to_sfixed(2080.0/65536.0,1,-nbitq), 
to_sfixed(-2818.0/65536.0,1,-nbitq), 
to_sfixed(2099.0/65536.0,1,-nbitq), 
to_sfixed(5477.0/65536.0,1,-nbitq), 
to_sfixed(-389.0/65536.0,1,-nbitq), 
to_sfixed(-8309.0/65536.0,1,-nbitq), 
to_sfixed(-3240.0/65536.0,1,-nbitq), 
to_sfixed(-1873.0/65536.0,1,-nbitq), 
to_sfixed(-5183.0/65536.0,1,-nbitq), 
to_sfixed(1306.0/65536.0,1,-nbitq), 
to_sfixed(3084.0/65536.0,1,-nbitq), 
to_sfixed(4282.0/65536.0,1,-nbitq), 
to_sfixed(-2491.0/65536.0,1,-nbitq), 
to_sfixed(-5855.0/65536.0,1,-nbitq), 
to_sfixed(76.0/65536.0,1,-nbitq), 
to_sfixed(2407.0/65536.0,1,-nbitq), 
to_sfixed(334.0/65536.0,1,-nbitq), 
to_sfixed(-2204.0/65536.0,1,-nbitq), 
to_sfixed(776.0/65536.0,1,-nbitq), 
to_sfixed(-2330.0/65536.0,1,-nbitq), 
to_sfixed(-2120.0/65536.0,1,-nbitq), 
to_sfixed(4758.0/65536.0,1,-nbitq), 
to_sfixed(-1531.0/65536.0,1,-nbitq), 
to_sfixed(1555.0/65536.0,1,-nbitq), 
to_sfixed(-577.0/65536.0,1,-nbitq), 
to_sfixed(5976.0/65536.0,1,-nbitq), 
to_sfixed(2087.0/65536.0,1,-nbitq), 
to_sfixed(-276.0/65536.0,1,-nbitq), 
to_sfixed(-882.0/65536.0,1,-nbitq), 
to_sfixed(1581.0/65536.0,1,-nbitq), 
to_sfixed(6892.0/65536.0,1,-nbitq), 
to_sfixed(2356.0/65536.0,1,-nbitq), 
to_sfixed(2331.0/65536.0,1,-nbitq), 
to_sfixed(-2389.0/65536.0,1,-nbitq)  ), 
( to_sfixed(573.0/65536.0,1,-nbitq), 
to_sfixed(572.0/65536.0,1,-nbitq), 
to_sfixed(3680.0/65536.0,1,-nbitq), 
to_sfixed(-3382.0/65536.0,1,-nbitq), 
to_sfixed(-2438.0/65536.0,1,-nbitq), 
to_sfixed(-2768.0/65536.0,1,-nbitq), 
to_sfixed(3294.0/65536.0,1,-nbitq), 
to_sfixed(3809.0/65536.0,1,-nbitq), 
to_sfixed(3742.0/65536.0,1,-nbitq), 
to_sfixed(2537.0/65536.0,1,-nbitq), 
to_sfixed(-1921.0/65536.0,1,-nbitq), 
to_sfixed(2505.0/65536.0,1,-nbitq), 
to_sfixed(237.0/65536.0,1,-nbitq), 
to_sfixed(-4687.0/65536.0,1,-nbitq), 
to_sfixed(3292.0/65536.0,1,-nbitq), 
to_sfixed(-289.0/65536.0,1,-nbitq), 
to_sfixed(-1584.0/65536.0,1,-nbitq), 
to_sfixed(6775.0/65536.0,1,-nbitq), 
to_sfixed(414.0/65536.0,1,-nbitq), 
to_sfixed(512.0/65536.0,1,-nbitq), 
to_sfixed(-4134.0/65536.0,1,-nbitq), 
to_sfixed(2317.0/65536.0,1,-nbitq), 
to_sfixed(-3837.0/65536.0,1,-nbitq), 
to_sfixed(-8045.0/65536.0,1,-nbitq), 
to_sfixed(-968.0/65536.0,1,-nbitq), 
to_sfixed(-5657.0/65536.0,1,-nbitq), 
to_sfixed(-5348.0/65536.0,1,-nbitq), 
to_sfixed(-2342.0/65536.0,1,-nbitq), 
to_sfixed(-5096.0/65536.0,1,-nbitq), 
to_sfixed(86.0/65536.0,1,-nbitq), 
to_sfixed(4038.0/65536.0,1,-nbitq), 
to_sfixed(778.0/65536.0,1,-nbitq), 
to_sfixed(2409.0/65536.0,1,-nbitq), 
to_sfixed(2543.0/65536.0,1,-nbitq), 
to_sfixed(-960.0/65536.0,1,-nbitq), 
to_sfixed(1637.0/65536.0,1,-nbitq), 
to_sfixed(4985.0/65536.0,1,-nbitq), 
to_sfixed(3909.0/65536.0,1,-nbitq), 
to_sfixed(-1160.0/65536.0,1,-nbitq), 
to_sfixed(1715.0/65536.0,1,-nbitq), 
to_sfixed(3170.0/65536.0,1,-nbitq), 
to_sfixed(-1682.0/65536.0,1,-nbitq), 
to_sfixed(7306.0/65536.0,1,-nbitq), 
to_sfixed(1096.0/65536.0,1,-nbitq), 
to_sfixed(-115.0/65536.0,1,-nbitq), 
to_sfixed(-7822.0/65536.0,1,-nbitq), 
to_sfixed(2805.0/65536.0,1,-nbitq), 
to_sfixed(-2820.0/65536.0,1,-nbitq), 
to_sfixed(3393.0/65536.0,1,-nbitq), 
to_sfixed(2880.0/65536.0,1,-nbitq), 
to_sfixed(1536.0/65536.0,1,-nbitq), 
to_sfixed(-7459.0/65536.0,1,-nbitq), 
to_sfixed(3466.0/65536.0,1,-nbitq), 
to_sfixed(-1024.0/65536.0,1,-nbitq), 
to_sfixed(-2262.0/65536.0,1,-nbitq), 
to_sfixed(2030.0/65536.0,1,-nbitq), 
to_sfixed(-2469.0/65536.0,1,-nbitq), 
to_sfixed(-2423.0/65536.0,1,-nbitq), 
to_sfixed(1981.0/65536.0,1,-nbitq), 
to_sfixed(-10627.0/65536.0,1,-nbitq), 
to_sfixed(-738.0/65536.0,1,-nbitq), 
to_sfixed(-684.0/65536.0,1,-nbitq), 
to_sfixed(3291.0/65536.0,1,-nbitq), 
to_sfixed(2596.0/65536.0,1,-nbitq), 
to_sfixed(5273.0/65536.0,1,-nbitq), 
to_sfixed(699.0/65536.0,1,-nbitq), 
to_sfixed(-2197.0/65536.0,1,-nbitq), 
to_sfixed(8880.0/65536.0,1,-nbitq), 
to_sfixed(636.0/65536.0,1,-nbitq), 
to_sfixed(3283.0/65536.0,1,-nbitq), 
to_sfixed(-3382.0/65536.0,1,-nbitq), 
to_sfixed(8814.0/65536.0,1,-nbitq), 
to_sfixed(-777.0/65536.0,1,-nbitq), 
to_sfixed(-955.0/65536.0,1,-nbitq), 
to_sfixed(-1658.0/65536.0,1,-nbitq), 
to_sfixed(371.0/65536.0,1,-nbitq), 
to_sfixed(6593.0/65536.0,1,-nbitq), 
to_sfixed(-1768.0/65536.0,1,-nbitq), 
to_sfixed(2871.0/65536.0,1,-nbitq), 
to_sfixed(-1699.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-489.0/65536.0,1,-nbitq), 
to_sfixed(-4096.0/65536.0,1,-nbitq), 
to_sfixed(-364.0/65536.0,1,-nbitq), 
to_sfixed(-3071.0/65536.0,1,-nbitq), 
to_sfixed(-2100.0/65536.0,1,-nbitq), 
to_sfixed(-5273.0/65536.0,1,-nbitq), 
to_sfixed(-536.0/65536.0,1,-nbitq), 
to_sfixed(-2995.0/65536.0,1,-nbitq), 
to_sfixed(1221.0/65536.0,1,-nbitq), 
to_sfixed(-427.0/65536.0,1,-nbitq), 
to_sfixed(4829.0/65536.0,1,-nbitq), 
to_sfixed(-323.0/65536.0,1,-nbitq), 
to_sfixed(1407.0/65536.0,1,-nbitq), 
to_sfixed(351.0/65536.0,1,-nbitq), 
to_sfixed(6374.0/65536.0,1,-nbitq), 
to_sfixed(-1134.0/65536.0,1,-nbitq), 
to_sfixed(-2294.0/65536.0,1,-nbitq), 
to_sfixed(4766.0/65536.0,1,-nbitq), 
to_sfixed(4395.0/65536.0,1,-nbitq), 
to_sfixed(1854.0/65536.0,1,-nbitq), 
to_sfixed(-6065.0/65536.0,1,-nbitq), 
to_sfixed(3245.0/65536.0,1,-nbitq), 
to_sfixed(621.0/65536.0,1,-nbitq), 
to_sfixed(-8271.0/65536.0,1,-nbitq), 
to_sfixed(3292.0/65536.0,1,-nbitq), 
to_sfixed(-7333.0/65536.0,1,-nbitq), 
to_sfixed(-2275.0/65536.0,1,-nbitq), 
to_sfixed(1433.0/65536.0,1,-nbitq), 
to_sfixed(-9875.0/65536.0,1,-nbitq), 
to_sfixed(-528.0/65536.0,1,-nbitq), 
to_sfixed(430.0/65536.0,1,-nbitq), 
to_sfixed(-2904.0/65536.0,1,-nbitq), 
to_sfixed(3166.0/65536.0,1,-nbitq), 
to_sfixed(1284.0/65536.0,1,-nbitq), 
to_sfixed(-828.0/65536.0,1,-nbitq), 
to_sfixed(-2430.0/65536.0,1,-nbitq), 
to_sfixed(7922.0/65536.0,1,-nbitq), 
to_sfixed(6878.0/65536.0,1,-nbitq), 
to_sfixed(2524.0/65536.0,1,-nbitq), 
to_sfixed(2712.0/65536.0,1,-nbitq), 
to_sfixed(784.0/65536.0,1,-nbitq), 
to_sfixed(1304.0/65536.0,1,-nbitq), 
to_sfixed(7358.0/65536.0,1,-nbitq), 
to_sfixed(5291.0/65536.0,1,-nbitq), 
to_sfixed(-1579.0/65536.0,1,-nbitq), 
to_sfixed(-7999.0/65536.0,1,-nbitq), 
to_sfixed(508.0/65536.0,1,-nbitq), 
to_sfixed(-214.0/65536.0,1,-nbitq), 
to_sfixed(1366.0/65536.0,1,-nbitq), 
to_sfixed(2674.0/65536.0,1,-nbitq), 
to_sfixed(-1432.0/65536.0,1,-nbitq), 
to_sfixed(-1320.0/65536.0,1,-nbitq), 
to_sfixed(3752.0/65536.0,1,-nbitq), 
to_sfixed(683.0/65536.0,1,-nbitq), 
to_sfixed(-3177.0/65536.0,1,-nbitq), 
to_sfixed(1797.0/65536.0,1,-nbitq), 
to_sfixed(-1136.0/65536.0,1,-nbitq), 
to_sfixed(1835.0/65536.0,1,-nbitq), 
to_sfixed(-494.0/65536.0,1,-nbitq), 
to_sfixed(-12437.0/65536.0,1,-nbitq), 
to_sfixed(3099.0/65536.0,1,-nbitq), 
to_sfixed(-1647.0/65536.0,1,-nbitq), 
to_sfixed(-1885.0/65536.0,1,-nbitq), 
to_sfixed(222.0/65536.0,1,-nbitq), 
to_sfixed(4009.0/65536.0,1,-nbitq), 
to_sfixed(4389.0/65536.0,1,-nbitq), 
to_sfixed(-1723.0/65536.0,1,-nbitq), 
to_sfixed(8393.0/65536.0,1,-nbitq), 
to_sfixed(-1342.0/65536.0,1,-nbitq), 
to_sfixed(1877.0/65536.0,1,-nbitq), 
to_sfixed(-2902.0/65536.0,1,-nbitq), 
to_sfixed(5371.0/65536.0,1,-nbitq), 
to_sfixed(-5444.0/65536.0,1,-nbitq), 
to_sfixed(1846.0/65536.0,1,-nbitq), 
to_sfixed(-3065.0/65536.0,1,-nbitq), 
to_sfixed(-1752.0/65536.0,1,-nbitq), 
to_sfixed(926.0/65536.0,1,-nbitq), 
to_sfixed(-5440.0/65536.0,1,-nbitq), 
to_sfixed(-2616.0/65536.0,1,-nbitq), 
to_sfixed(-6235.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-790.0/65536.0,1,-nbitq), 
to_sfixed(-335.0/65536.0,1,-nbitq), 
to_sfixed(-7434.0/65536.0,1,-nbitq), 
to_sfixed(-2602.0/65536.0,1,-nbitq), 
to_sfixed(9741.0/65536.0,1,-nbitq), 
to_sfixed(-4679.0/65536.0,1,-nbitq), 
to_sfixed(-1858.0/65536.0,1,-nbitq), 
to_sfixed(-1406.0/65536.0,1,-nbitq), 
to_sfixed(631.0/65536.0,1,-nbitq), 
to_sfixed(-2318.0/65536.0,1,-nbitq), 
to_sfixed(11012.0/65536.0,1,-nbitq), 
to_sfixed(1171.0/65536.0,1,-nbitq), 
to_sfixed(-1461.0/65536.0,1,-nbitq), 
to_sfixed(79.0/65536.0,1,-nbitq), 
to_sfixed(5340.0/65536.0,1,-nbitq), 
to_sfixed(2662.0/65536.0,1,-nbitq), 
to_sfixed(691.0/65536.0,1,-nbitq), 
to_sfixed(6730.0/65536.0,1,-nbitq), 
to_sfixed(4447.0/65536.0,1,-nbitq), 
to_sfixed(871.0/65536.0,1,-nbitq), 
to_sfixed(-7492.0/65536.0,1,-nbitq), 
to_sfixed(858.0/65536.0,1,-nbitq), 
to_sfixed(7556.0/65536.0,1,-nbitq), 
to_sfixed(-3592.0/65536.0,1,-nbitq), 
to_sfixed(-1017.0/65536.0,1,-nbitq), 
to_sfixed(-4198.0/65536.0,1,-nbitq), 
to_sfixed(-1537.0/65536.0,1,-nbitq), 
to_sfixed(865.0/65536.0,1,-nbitq), 
to_sfixed(-6964.0/65536.0,1,-nbitq), 
to_sfixed(-2876.0/65536.0,1,-nbitq), 
to_sfixed(2995.0/65536.0,1,-nbitq), 
to_sfixed(464.0/65536.0,1,-nbitq), 
to_sfixed(-1148.0/65536.0,1,-nbitq), 
to_sfixed(-4808.0/65536.0,1,-nbitq), 
to_sfixed(-1563.0/65536.0,1,-nbitq), 
to_sfixed(421.0/65536.0,1,-nbitq), 
to_sfixed(8324.0/65536.0,1,-nbitq), 
to_sfixed(-2492.0/65536.0,1,-nbitq), 
to_sfixed(3560.0/65536.0,1,-nbitq), 
to_sfixed(4103.0/65536.0,1,-nbitq), 
to_sfixed(18.0/65536.0,1,-nbitq), 
to_sfixed(2205.0/65536.0,1,-nbitq), 
to_sfixed(268.0/65536.0,1,-nbitq), 
to_sfixed(1697.0/65536.0,1,-nbitq), 
to_sfixed(2757.0/65536.0,1,-nbitq), 
to_sfixed(-6944.0/65536.0,1,-nbitq), 
to_sfixed(1944.0/65536.0,1,-nbitq), 
to_sfixed(-1574.0/65536.0,1,-nbitq), 
to_sfixed(34.0/65536.0,1,-nbitq), 
to_sfixed(-1406.0/65536.0,1,-nbitq), 
to_sfixed(-1224.0/65536.0,1,-nbitq), 
to_sfixed(1534.0/65536.0,1,-nbitq), 
to_sfixed(397.0/65536.0,1,-nbitq), 
to_sfixed(-3738.0/65536.0,1,-nbitq), 
to_sfixed(-4672.0/65536.0,1,-nbitq), 
to_sfixed(-475.0/65536.0,1,-nbitq), 
to_sfixed(-1058.0/65536.0,1,-nbitq), 
to_sfixed(-62.0/65536.0,1,-nbitq), 
to_sfixed(-965.0/65536.0,1,-nbitq), 
to_sfixed(-12747.0/65536.0,1,-nbitq), 
to_sfixed(5909.0/65536.0,1,-nbitq), 
to_sfixed(1618.0/65536.0,1,-nbitq), 
to_sfixed(2588.0/65536.0,1,-nbitq), 
to_sfixed(1990.0/65536.0,1,-nbitq), 
to_sfixed(1999.0/65536.0,1,-nbitq), 
to_sfixed(-166.0/65536.0,1,-nbitq), 
to_sfixed(-3314.0/65536.0,1,-nbitq), 
to_sfixed(6362.0/65536.0,1,-nbitq), 
to_sfixed(-3.0/65536.0,1,-nbitq), 
to_sfixed(12208.0/65536.0,1,-nbitq), 
to_sfixed(847.0/65536.0,1,-nbitq), 
to_sfixed(-2498.0/65536.0,1,-nbitq), 
to_sfixed(-2053.0/65536.0,1,-nbitq), 
to_sfixed(-2028.0/65536.0,1,-nbitq), 
to_sfixed(855.0/65536.0,1,-nbitq), 
to_sfixed(4993.0/65536.0,1,-nbitq), 
to_sfixed(-1323.0/65536.0,1,-nbitq), 
to_sfixed(-2894.0/65536.0,1,-nbitq), 
to_sfixed(-2686.0/65536.0,1,-nbitq), 
to_sfixed(-6059.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-848.0/65536.0,1,-nbitq), 
to_sfixed(-2658.0/65536.0,1,-nbitq), 
to_sfixed(-15193.0/65536.0,1,-nbitq), 
to_sfixed(-5095.0/65536.0,1,-nbitq), 
to_sfixed(5497.0/65536.0,1,-nbitq), 
to_sfixed(-7779.0/65536.0,1,-nbitq), 
to_sfixed(-603.0/65536.0,1,-nbitq), 
to_sfixed(-5895.0/65536.0,1,-nbitq), 
to_sfixed(-1186.0/65536.0,1,-nbitq), 
to_sfixed(-2746.0/65536.0,1,-nbitq), 
to_sfixed(6544.0/65536.0,1,-nbitq), 
to_sfixed(-4920.0/65536.0,1,-nbitq), 
to_sfixed(1643.0/65536.0,1,-nbitq), 
to_sfixed(-8353.0/65536.0,1,-nbitq), 
to_sfixed(1211.0/65536.0,1,-nbitq), 
to_sfixed(-1811.0/65536.0,1,-nbitq), 
to_sfixed(-1247.0/65536.0,1,-nbitq), 
to_sfixed(3755.0/65536.0,1,-nbitq), 
to_sfixed(4890.0/65536.0,1,-nbitq), 
to_sfixed(-950.0/65536.0,1,-nbitq), 
to_sfixed(-6872.0/65536.0,1,-nbitq), 
to_sfixed(7834.0/65536.0,1,-nbitq), 
to_sfixed(14194.0/65536.0,1,-nbitq), 
to_sfixed(-6039.0/65536.0,1,-nbitq), 
to_sfixed(-2898.0/65536.0,1,-nbitq), 
to_sfixed(-4722.0/65536.0,1,-nbitq), 
to_sfixed(221.0/65536.0,1,-nbitq), 
to_sfixed(2453.0/65536.0,1,-nbitq), 
to_sfixed(4095.0/65536.0,1,-nbitq), 
to_sfixed(-3138.0/65536.0,1,-nbitq), 
to_sfixed(2801.0/65536.0,1,-nbitq), 
to_sfixed(-2183.0/65536.0,1,-nbitq), 
to_sfixed(-800.0/65536.0,1,-nbitq), 
to_sfixed(-9421.0/65536.0,1,-nbitq), 
to_sfixed(-2262.0/65536.0,1,-nbitq), 
to_sfixed(-2280.0/65536.0,1,-nbitq), 
to_sfixed(12206.0/65536.0,1,-nbitq), 
to_sfixed(-5030.0/65536.0,1,-nbitq), 
to_sfixed(8006.0/65536.0,1,-nbitq), 
to_sfixed(2294.0/65536.0,1,-nbitq), 
to_sfixed(-3142.0/65536.0,1,-nbitq), 
to_sfixed(1357.0/65536.0,1,-nbitq), 
to_sfixed(-4176.0/65536.0,1,-nbitq), 
to_sfixed(7166.0/65536.0,1,-nbitq), 
to_sfixed(2437.0/65536.0,1,-nbitq), 
to_sfixed(-5496.0/65536.0,1,-nbitq), 
to_sfixed(-1365.0/65536.0,1,-nbitq), 
to_sfixed(4329.0/65536.0,1,-nbitq), 
to_sfixed(3372.0/65536.0,1,-nbitq), 
to_sfixed(-462.0/65536.0,1,-nbitq), 
to_sfixed(-883.0/65536.0,1,-nbitq), 
to_sfixed(-2013.0/65536.0,1,-nbitq), 
to_sfixed(-3349.0/65536.0,1,-nbitq), 
to_sfixed(-9954.0/65536.0,1,-nbitq), 
to_sfixed(-839.0/65536.0,1,-nbitq), 
to_sfixed(1050.0/65536.0,1,-nbitq), 
to_sfixed(1587.0/65536.0,1,-nbitq), 
to_sfixed(364.0/65536.0,1,-nbitq), 
to_sfixed(750.0/65536.0,1,-nbitq), 
to_sfixed(-10834.0/65536.0,1,-nbitq), 
to_sfixed(168.0/65536.0,1,-nbitq), 
to_sfixed(2068.0/65536.0,1,-nbitq), 
to_sfixed(-1065.0/65536.0,1,-nbitq), 
to_sfixed(2752.0/65536.0,1,-nbitq), 
to_sfixed(-867.0/65536.0,1,-nbitq), 
to_sfixed(-5574.0/65536.0,1,-nbitq), 
to_sfixed(-715.0/65536.0,1,-nbitq), 
to_sfixed(4939.0/65536.0,1,-nbitq), 
to_sfixed(315.0/65536.0,1,-nbitq), 
to_sfixed(13121.0/65536.0,1,-nbitq), 
to_sfixed(-3584.0/65536.0,1,-nbitq), 
to_sfixed(-623.0/65536.0,1,-nbitq), 
to_sfixed(-4745.0/65536.0,1,-nbitq), 
to_sfixed(163.0/65536.0,1,-nbitq), 
to_sfixed(-3187.0/65536.0,1,-nbitq), 
to_sfixed(-4213.0/65536.0,1,-nbitq), 
to_sfixed(4234.0/65536.0,1,-nbitq), 
to_sfixed(488.0/65536.0,1,-nbitq), 
to_sfixed(-126.0/65536.0,1,-nbitq), 
to_sfixed(-4407.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2759.0/65536.0,1,-nbitq), 
to_sfixed(3076.0/65536.0,1,-nbitq), 
to_sfixed(-14466.0/65536.0,1,-nbitq), 
to_sfixed(-7624.0/65536.0,1,-nbitq), 
to_sfixed(-2328.0/65536.0,1,-nbitq), 
to_sfixed(1830.0/65536.0,1,-nbitq), 
to_sfixed(1432.0/65536.0,1,-nbitq), 
to_sfixed(-2802.0/65536.0,1,-nbitq), 
to_sfixed(-906.0/65536.0,1,-nbitq), 
to_sfixed(599.0/65536.0,1,-nbitq), 
to_sfixed(5646.0/65536.0,1,-nbitq), 
to_sfixed(-10384.0/65536.0,1,-nbitq), 
to_sfixed(-2879.0/65536.0,1,-nbitq), 
to_sfixed(-5542.0/65536.0,1,-nbitq), 
to_sfixed(2506.0/65536.0,1,-nbitq), 
to_sfixed(1336.0/65536.0,1,-nbitq), 
to_sfixed(-2066.0/65536.0,1,-nbitq), 
to_sfixed(-410.0/65536.0,1,-nbitq), 
to_sfixed(5359.0/65536.0,1,-nbitq), 
to_sfixed(2230.0/65536.0,1,-nbitq), 
to_sfixed(-11042.0/65536.0,1,-nbitq), 
to_sfixed(8384.0/65536.0,1,-nbitq), 
to_sfixed(18684.0/65536.0,1,-nbitq), 
to_sfixed(5963.0/65536.0,1,-nbitq), 
to_sfixed(-3596.0/65536.0,1,-nbitq), 
to_sfixed(4037.0/65536.0,1,-nbitq), 
to_sfixed(-1866.0/65536.0,1,-nbitq), 
to_sfixed(-2058.0/65536.0,1,-nbitq), 
to_sfixed(-666.0/65536.0,1,-nbitq), 
to_sfixed(-123.0/65536.0,1,-nbitq), 
to_sfixed(8187.0/65536.0,1,-nbitq), 
to_sfixed(-6932.0/65536.0,1,-nbitq), 
to_sfixed(-3505.0/65536.0,1,-nbitq), 
to_sfixed(-7122.0/65536.0,1,-nbitq), 
to_sfixed(-1597.0/65536.0,1,-nbitq), 
to_sfixed(-1573.0/65536.0,1,-nbitq), 
to_sfixed(12746.0/65536.0,1,-nbitq), 
to_sfixed(-3495.0/65536.0,1,-nbitq), 
to_sfixed(6695.0/65536.0,1,-nbitq), 
to_sfixed(-1209.0/65536.0,1,-nbitq), 
to_sfixed(-4351.0/65536.0,1,-nbitq), 
to_sfixed(1129.0/65536.0,1,-nbitq), 
to_sfixed(-4448.0/65536.0,1,-nbitq), 
to_sfixed(1520.0/65536.0,1,-nbitq), 
to_sfixed(1291.0/65536.0,1,-nbitq), 
to_sfixed(-3778.0/65536.0,1,-nbitq), 
to_sfixed(1862.0/65536.0,1,-nbitq), 
to_sfixed(7756.0/65536.0,1,-nbitq), 
to_sfixed(-1160.0/65536.0,1,-nbitq), 
to_sfixed(-716.0/65536.0,1,-nbitq), 
to_sfixed(-2352.0/65536.0,1,-nbitq), 
to_sfixed(-8003.0/65536.0,1,-nbitq), 
to_sfixed(-3550.0/65536.0,1,-nbitq), 
to_sfixed(-3632.0/65536.0,1,-nbitq), 
to_sfixed(-2320.0/65536.0,1,-nbitq), 
to_sfixed(-2681.0/65536.0,1,-nbitq), 
to_sfixed(-2231.0/65536.0,1,-nbitq), 
to_sfixed(-1654.0/65536.0,1,-nbitq), 
to_sfixed(-3742.0/65536.0,1,-nbitq), 
to_sfixed(-14283.0/65536.0,1,-nbitq), 
to_sfixed(979.0/65536.0,1,-nbitq), 
to_sfixed(2155.0/65536.0,1,-nbitq), 
to_sfixed(1573.0/65536.0,1,-nbitq), 
to_sfixed(-2372.0/65536.0,1,-nbitq), 
to_sfixed(296.0/65536.0,1,-nbitq), 
to_sfixed(-3611.0/65536.0,1,-nbitq), 
to_sfixed(-3091.0/65536.0,1,-nbitq), 
to_sfixed(4372.0/65536.0,1,-nbitq), 
to_sfixed(3180.0/65536.0,1,-nbitq), 
to_sfixed(9177.0/65536.0,1,-nbitq), 
to_sfixed(-1033.0/65536.0,1,-nbitq), 
to_sfixed(4882.0/65536.0,1,-nbitq), 
to_sfixed(-8281.0/65536.0,1,-nbitq), 
to_sfixed(847.0/65536.0,1,-nbitq), 
to_sfixed(2295.0/65536.0,1,-nbitq), 
to_sfixed(-4038.0/65536.0,1,-nbitq), 
to_sfixed(1942.0/65536.0,1,-nbitq), 
to_sfixed(6657.0/65536.0,1,-nbitq), 
to_sfixed(-3286.0/65536.0,1,-nbitq), 
to_sfixed(1062.0/65536.0,1,-nbitq)  ), 
( to_sfixed(556.0/65536.0,1,-nbitq), 
to_sfixed(4323.0/65536.0,1,-nbitq), 
to_sfixed(-12336.0/65536.0,1,-nbitq), 
to_sfixed(-5555.0/65536.0,1,-nbitq), 
to_sfixed(803.0/65536.0,1,-nbitq), 
to_sfixed(4067.0/65536.0,1,-nbitq), 
to_sfixed(-1175.0/65536.0,1,-nbitq), 
to_sfixed(-4273.0/65536.0,1,-nbitq), 
to_sfixed(5693.0/65536.0,1,-nbitq), 
to_sfixed(-150.0/65536.0,1,-nbitq), 
to_sfixed(5601.0/65536.0,1,-nbitq), 
to_sfixed(-4487.0/65536.0,1,-nbitq), 
to_sfixed(-136.0/65536.0,1,-nbitq), 
to_sfixed(-713.0/65536.0,1,-nbitq), 
to_sfixed(-63.0/65536.0,1,-nbitq), 
to_sfixed(1883.0/65536.0,1,-nbitq), 
to_sfixed(3049.0/65536.0,1,-nbitq), 
to_sfixed(868.0/65536.0,1,-nbitq), 
to_sfixed(3381.0/65536.0,1,-nbitq), 
to_sfixed(-1128.0/65536.0,1,-nbitq), 
to_sfixed(-7819.0/65536.0,1,-nbitq), 
to_sfixed(10587.0/65536.0,1,-nbitq), 
to_sfixed(9427.0/65536.0,1,-nbitq), 
to_sfixed(8367.0/65536.0,1,-nbitq), 
to_sfixed(-6577.0/65536.0,1,-nbitq), 
to_sfixed(-2530.0/65536.0,1,-nbitq), 
to_sfixed(1009.0/65536.0,1,-nbitq), 
to_sfixed(2645.0/65536.0,1,-nbitq), 
to_sfixed(5412.0/65536.0,1,-nbitq), 
to_sfixed(-2429.0/65536.0,1,-nbitq), 
to_sfixed(6278.0/65536.0,1,-nbitq), 
to_sfixed(-8049.0/65536.0,1,-nbitq), 
to_sfixed(2746.0/65536.0,1,-nbitq), 
to_sfixed(49.0/65536.0,1,-nbitq), 
to_sfixed(2573.0/65536.0,1,-nbitq), 
to_sfixed(401.0/65536.0,1,-nbitq), 
to_sfixed(8685.0/65536.0,1,-nbitq), 
to_sfixed(506.0/65536.0,1,-nbitq), 
to_sfixed(6125.0/65536.0,1,-nbitq), 
to_sfixed(-1926.0/65536.0,1,-nbitq), 
to_sfixed(-6027.0/65536.0,1,-nbitq), 
to_sfixed(-2399.0/65536.0,1,-nbitq), 
to_sfixed(-1007.0/65536.0,1,-nbitq), 
to_sfixed(2066.0/65536.0,1,-nbitq), 
to_sfixed(-2513.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(-1743.0/65536.0,1,-nbitq), 
to_sfixed(5155.0/65536.0,1,-nbitq), 
to_sfixed(1789.0/65536.0,1,-nbitq), 
to_sfixed(719.0/65536.0,1,-nbitq), 
to_sfixed(-1404.0/65536.0,1,-nbitq), 
to_sfixed(-6127.0/65536.0,1,-nbitq), 
to_sfixed(-3741.0/65536.0,1,-nbitq), 
to_sfixed(-1159.0/65536.0,1,-nbitq), 
to_sfixed(-2291.0/65536.0,1,-nbitq), 
to_sfixed(-6882.0/65536.0,1,-nbitq), 
to_sfixed(-1702.0/65536.0,1,-nbitq), 
to_sfixed(-1307.0/65536.0,1,-nbitq), 
to_sfixed(-429.0/65536.0,1,-nbitq), 
to_sfixed(-3549.0/65536.0,1,-nbitq), 
to_sfixed(8138.0/65536.0,1,-nbitq), 
to_sfixed(1334.0/65536.0,1,-nbitq), 
to_sfixed(910.0/65536.0,1,-nbitq), 
to_sfixed(2249.0/65536.0,1,-nbitq), 
to_sfixed(1407.0/65536.0,1,-nbitq), 
to_sfixed(-7925.0/65536.0,1,-nbitq), 
to_sfixed(-7499.0/65536.0,1,-nbitq), 
to_sfixed(8201.0/65536.0,1,-nbitq), 
to_sfixed(2985.0/65536.0,1,-nbitq), 
to_sfixed(3369.0/65536.0,1,-nbitq), 
to_sfixed(-31.0/65536.0,1,-nbitq), 
to_sfixed(3611.0/65536.0,1,-nbitq), 
to_sfixed(-6472.0/65536.0,1,-nbitq), 
to_sfixed(-2364.0/65536.0,1,-nbitq), 
to_sfixed(643.0/65536.0,1,-nbitq), 
to_sfixed(-3112.0/65536.0,1,-nbitq), 
to_sfixed(5232.0/65536.0,1,-nbitq), 
to_sfixed(2200.0/65536.0,1,-nbitq), 
to_sfixed(-2711.0/65536.0,1,-nbitq), 
to_sfixed(384.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-104.0/65536.0,1,-nbitq), 
to_sfixed(3831.0/65536.0,1,-nbitq), 
to_sfixed(-4522.0/65536.0,1,-nbitq), 
to_sfixed(-2324.0/65536.0,1,-nbitq), 
to_sfixed(-1184.0/65536.0,1,-nbitq), 
to_sfixed(5044.0/65536.0,1,-nbitq), 
to_sfixed(1378.0/65536.0,1,-nbitq), 
to_sfixed(-2866.0/65536.0,1,-nbitq), 
to_sfixed(4809.0/65536.0,1,-nbitq), 
to_sfixed(330.0/65536.0,1,-nbitq), 
to_sfixed(6005.0/65536.0,1,-nbitq), 
to_sfixed(-7764.0/65536.0,1,-nbitq), 
to_sfixed(-31.0/65536.0,1,-nbitq), 
to_sfixed(3168.0/65536.0,1,-nbitq), 
to_sfixed(436.0/65536.0,1,-nbitq), 
to_sfixed(-638.0/65536.0,1,-nbitq), 
to_sfixed(-3180.0/65536.0,1,-nbitq), 
to_sfixed(-1549.0/65536.0,1,-nbitq), 
to_sfixed(1950.0/65536.0,1,-nbitq), 
to_sfixed(1096.0/65536.0,1,-nbitq), 
to_sfixed(-6941.0/65536.0,1,-nbitq), 
to_sfixed(696.0/65536.0,1,-nbitq), 
to_sfixed(-4579.0/65536.0,1,-nbitq), 
to_sfixed(9595.0/65536.0,1,-nbitq), 
to_sfixed(-2367.0/65536.0,1,-nbitq), 
to_sfixed(4848.0/65536.0,1,-nbitq), 
to_sfixed(-936.0/65536.0,1,-nbitq), 
to_sfixed(1385.0/65536.0,1,-nbitq), 
to_sfixed(4305.0/65536.0,1,-nbitq), 
to_sfixed(-1421.0/65536.0,1,-nbitq), 
to_sfixed(3022.0/65536.0,1,-nbitq), 
to_sfixed(-7458.0/65536.0,1,-nbitq), 
to_sfixed(-2031.0/65536.0,1,-nbitq), 
to_sfixed(-2366.0/65536.0,1,-nbitq), 
to_sfixed(-16.0/65536.0,1,-nbitq), 
to_sfixed(-974.0/65536.0,1,-nbitq), 
to_sfixed(4070.0/65536.0,1,-nbitq), 
to_sfixed(1448.0/65536.0,1,-nbitq), 
to_sfixed(-3265.0/65536.0,1,-nbitq), 
to_sfixed(695.0/65536.0,1,-nbitq), 
to_sfixed(-5985.0/65536.0,1,-nbitq), 
to_sfixed(-228.0/65536.0,1,-nbitq), 
to_sfixed(1902.0/65536.0,1,-nbitq), 
to_sfixed(1220.0/65536.0,1,-nbitq), 
to_sfixed(2860.0/65536.0,1,-nbitq), 
to_sfixed(2966.0/65536.0,1,-nbitq), 
to_sfixed(1022.0/65536.0,1,-nbitq), 
to_sfixed(6809.0/65536.0,1,-nbitq), 
to_sfixed(1688.0/65536.0,1,-nbitq), 
to_sfixed(2517.0/65536.0,1,-nbitq), 
to_sfixed(989.0/65536.0,1,-nbitq), 
to_sfixed(-4082.0/65536.0,1,-nbitq), 
to_sfixed(-5682.0/65536.0,1,-nbitq), 
to_sfixed(-7467.0/65536.0,1,-nbitq), 
to_sfixed(-6095.0/65536.0,1,-nbitq), 
to_sfixed(-3371.0/65536.0,1,-nbitq), 
to_sfixed(284.0/65536.0,1,-nbitq), 
to_sfixed(-1662.0/65536.0,1,-nbitq), 
to_sfixed(-132.0/65536.0,1,-nbitq), 
to_sfixed(1517.0/65536.0,1,-nbitq), 
to_sfixed(1932.0/65536.0,1,-nbitq), 
to_sfixed(824.0/65536.0,1,-nbitq), 
to_sfixed(3226.0/65536.0,1,-nbitq), 
to_sfixed(2437.0/65536.0,1,-nbitq), 
to_sfixed(192.0/65536.0,1,-nbitq), 
to_sfixed(-8441.0/65536.0,1,-nbitq), 
to_sfixed(-4974.0/65536.0,1,-nbitq), 
to_sfixed(5019.0/65536.0,1,-nbitq), 
to_sfixed(7162.0/65536.0,1,-nbitq), 
to_sfixed(-377.0/65536.0,1,-nbitq), 
to_sfixed(-3313.0/65536.0,1,-nbitq), 
to_sfixed(243.0/65536.0,1,-nbitq), 
to_sfixed(-1084.0/65536.0,1,-nbitq), 
to_sfixed(1474.0/65536.0,1,-nbitq), 
to_sfixed(2671.0/65536.0,1,-nbitq), 
to_sfixed(-3027.0/65536.0,1,-nbitq), 
to_sfixed(4150.0/65536.0,1,-nbitq), 
to_sfixed(-1531.0/65536.0,1,-nbitq), 
to_sfixed(187.0/65536.0,1,-nbitq), 
to_sfixed(3455.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2061.0/65536.0,1,-nbitq), 
to_sfixed(1713.0/65536.0,1,-nbitq), 
to_sfixed(768.0/65536.0,1,-nbitq), 
to_sfixed(-2784.0/65536.0,1,-nbitq), 
to_sfixed(1090.0/65536.0,1,-nbitq), 
to_sfixed(8305.0/65536.0,1,-nbitq), 
to_sfixed(-1899.0/65536.0,1,-nbitq), 
to_sfixed(-5416.0/65536.0,1,-nbitq), 
to_sfixed(6959.0/65536.0,1,-nbitq), 
to_sfixed(1945.0/65536.0,1,-nbitq), 
to_sfixed(2257.0/65536.0,1,-nbitq), 
to_sfixed(-15622.0/65536.0,1,-nbitq), 
to_sfixed(-1826.0/65536.0,1,-nbitq), 
to_sfixed(5384.0/65536.0,1,-nbitq), 
to_sfixed(-2965.0/65536.0,1,-nbitq), 
to_sfixed(-609.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(85.0/65536.0,1,-nbitq), 
to_sfixed(5265.0/65536.0,1,-nbitq), 
to_sfixed(-635.0/65536.0,1,-nbitq), 
to_sfixed(-11969.0/65536.0,1,-nbitq), 
to_sfixed(-947.0/65536.0,1,-nbitq), 
to_sfixed(-5079.0/65536.0,1,-nbitq), 
to_sfixed(6707.0/65536.0,1,-nbitq), 
to_sfixed(-191.0/65536.0,1,-nbitq), 
to_sfixed(4310.0/65536.0,1,-nbitq), 
to_sfixed(988.0/65536.0,1,-nbitq), 
to_sfixed(3012.0/65536.0,1,-nbitq), 
to_sfixed(3534.0/65536.0,1,-nbitq), 
to_sfixed(-3191.0/65536.0,1,-nbitq), 
to_sfixed(3275.0/65536.0,1,-nbitq), 
to_sfixed(-10389.0/65536.0,1,-nbitq), 
to_sfixed(-9053.0/65536.0,1,-nbitq), 
to_sfixed(-3977.0/65536.0,1,-nbitq), 
to_sfixed(401.0/65536.0,1,-nbitq), 
to_sfixed(3496.0/65536.0,1,-nbitq), 
to_sfixed(1035.0/65536.0,1,-nbitq), 
to_sfixed(-657.0/65536.0,1,-nbitq), 
to_sfixed(219.0/65536.0,1,-nbitq), 
to_sfixed(2311.0/65536.0,1,-nbitq), 
to_sfixed(83.0/65536.0,1,-nbitq), 
to_sfixed(-1996.0/65536.0,1,-nbitq), 
to_sfixed(-12042.0/65536.0,1,-nbitq), 
to_sfixed(-265.0/65536.0,1,-nbitq), 
to_sfixed(3111.0/65536.0,1,-nbitq), 
to_sfixed(-3336.0/65536.0,1,-nbitq), 
to_sfixed(-3032.0/65536.0,1,-nbitq), 
to_sfixed(11.0/65536.0,1,-nbitq), 
to_sfixed(1819.0/65536.0,1,-nbitq), 
to_sfixed(-1530.0/65536.0,1,-nbitq), 
to_sfixed(-2693.0/65536.0,1,-nbitq), 
to_sfixed(-2696.0/65536.0,1,-nbitq), 
to_sfixed(-2669.0/65536.0,1,-nbitq), 
to_sfixed(-6473.0/65536.0,1,-nbitq), 
to_sfixed(-5680.0/65536.0,1,-nbitq), 
to_sfixed(-2036.0/65536.0,1,-nbitq), 
to_sfixed(555.0/65536.0,1,-nbitq), 
to_sfixed(-298.0/65536.0,1,-nbitq), 
to_sfixed(527.0/65536.0,1,-nbitq), 
to_sfixed(-1873.0/65536.0,1,-nbitq), 
to_sfixed(-4145.0/65536.0,1,-nbitq), 
to_sfixed(-795.0/65536.0,1,-nbitq), 
to_sfixed(245.0/65536.0,1,-nbitq), 
to_sfixed(1503.0/65536.0,1,-nbitq), 
to_sfixed(-2680.0/65536.0,1,-nbitq), 
to_sfixed(-7004.0/65536.0,1,-nbitq), 
to_sfixed(-2357.0/65536.0,1,-nbitq), 
to_sfixed(8017.0/65536.0,1,-nbitq), 
to_sfixed(6053.0/65536.0,1,-nbitq), 
to_sfixed(-4777.0/65536.0,1,-nbitq), 
to_sfixed(-1601.0/65536.0,1,-nbitq), 
to_sfixed(800.0/65536.0,1,-nbitq), 
to_sfixed(-1084.0/65536.0,1,-nbitq), 
to_sfixed(2508.0/65536.0,1,-nbitq), 
to_sfixed(-519.0/65536.0,1,-nbitq), 
to_sfixed(-8572.0/65536.0,1,-nbitq), 
to_sfixed(567.0/65536.0,1,-nbitq), 
to_sfixed(-2440.0/65536.0,1,-nbitq), 
to_sfixed(-1206.0/65536.0,1,-nbitq), 
to_sfixed(4142.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1236.0/65536.0,1,-nbitq), 
to_sfixed(2216.0/65536.0,1,-nbitq), 
to_sfixed(5618.0/65536.0,1,-nbitq), 
to_sfixed(1379.0/65536.0,1,-nbitq), 
to_sfixed(4628.0/65536.0,1,-nbitq), 
to_sfixed(9533.0/65536.0,1,-nbitq), 
to_sfixed(-411.0/65536.0,1,-nbitq), 
to_sfixed(-4219.0/65536.0,1,-nbitq), 
to_sfixed(2606.0/65536.0,1,-nbitq), 
to_sfixed(1581.0/65536.0,1,-nbitq), 
to_sfixed(2798.0/65536.0,1,-nbitq), 
to_sfixed(-11909.0/65536.0,1,-nbitq), 
to_sfixed(-1752.0/65536.0,1,-nbitq), 
to_sfixed(-2104.0/65536.0,1,-nbitq), 
to_sfixed(172.0/65536.0,1,-nbitq), 
to_sfixed(-1295.0/65536.0,1,-nbitq), 
to_sfixed(189.0/65536.0,1,-nbitq), 
to_sfixed(1042.0/65536.0,1,-nbitq), 
to_sfixed(1934.0/65536.0,1,-nbitq), 
to_sfixed(1596.0/65536.0,1,-nbitq), 
to_sfixed(-490.0/65536.0,1,-nbitq), 
to_sfixed(-1264.0/65536.0,1,-nbitq), 
to_sfixed(1960.0/65536.0,1,-nbitq), 
to_sfixed(1108.0/65536.0,1,-nbitq), 
to_sfixed(-428.0/65536.0,1,-nbitq), 
to_sfixed(6088.0/65536.0,1,-nbitq), 
to_sfixed(5638.0/65536.0,1,-nbitq), 
to_sfixed(2283.0/65536.0,1,-nbitq), 
to_sfixed(6932.0/65536.0,1,-nbitq), 
to_sfixed(-4708.0/65536.0,1,-nbitq), 
to_sfixed(1770.0/65536.0,1,-nbitq), 
to_sfixed(-4418.0/65536.0,1,-nbitq), 
to_sfixed(-6757.0/65536.0,1,-nbitq), 
to_sfixed(1716.0/65536.0,1,-nbitq), 
to_sfixed(1821.0/65536.0,1,-nbitq), 
to_sfixed(-126.0/65536.0,1,-nbitq), 
to_sfixed(6818.0/65536.0,1,-nbitq), 
to_sfixed(2018.0/65536.0,1,-nbitq), 
to_sfixed(5714.0/65536.0,1,-nbitq), 
to_sfixed(-1605.0/65536.0,1,-nbitq), 
to_sfixed(-6531.0/65536.0,1,-nbitq), 
to_sfixed(-2568.0/65536.0,1,-nbitq), 
to_sfixed(-10715.0/65536.0,1,-nbitq), 
to_sfixed(-4970.0/65536.0,1,-nbitq), 
to_sfixed(2595.0/65536.0,1,-nbitq), 
to_sfixed(-5311.0/65536.0,1,-nbitq), 
to_sfixed(-2409.0/65536.0,1,-nbitq), 
to_sfixed(-418.0/65536.0,1,-nbitq), 
to_sfixed(-1366.0/65536.0,1,-nbitq), 
to_sfixed(3111.0/65536.0,1,-nbitq), 
to_sfixed(2654.0/65536.0,1,-nbitq), 
to_sfixed(-7059.0/65536.0,1,-nbitq), 
to_sfixed(-1781.0/65536.0,1,-nbitq), 
to_sfixed(3146.0/65536.0,1,-nbitq), 
to_sfixed(-5465.0/65536.0,1,-nbitq), 
to_sfixed(-3383.0/65536.0,1,-nbitq), 
to_sfixed(773.0/65536.0,1,-nbitq), 
to_sfixed(-1937.0/65536.0,1,-nbitq), 
to_sfixed(664.0/65536.0,1,-nbitq), 
to_sfixed(3691.0/65536.0,1,-nbitq), 
to_sfixed(-2858.0/65536.0,1,-nbitq), 
to_sfixed(-2653.0/65536.0,1,-nbitq), 
to_sfixed(540.0/65536.0,1,-nbitq), 
to_sfixed(2314.0/65536.0,1,-nbitq), 
to_sfixed(-2880.0/65536.0,1,-nbitq), 
to_sfixed(1118.0/65536.0,1,-nbitq), 
to_sfixed(-4436.0/65536.0,1,-nbitq), 
to_sfixed(9604.0/65536.0,1,-nbitq), 
to_sfixed(5829.0/65536.0,1,-nbitq), 
to_sfixed(-5569.0/65536.0,1,-nbitq), 
to_sfixed(-4952.0/65536.0,1,-nbitq), 
to_sfixed(-1409.0/65536.0,1,-nbitq), 
to_sfixed(2833.0/65536.0,1,-nbitq), 
to_sfixed(2245.0/65536.0,1,-nbitq), 
to_sfixed(-1604.0/65536.0,1,-nbitq), 
to_sfixed(-2311.0/65536.0,1,-nbitq), 
to_sfixed(2731.0/65536.0,1,-nbitq), 
to_sfixed(-3190.0/65536.0,1,-nbitq), 
to_sfixed(-1179.0/65536.0,1,-nbitq), 
to_sfixed(-254.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1534.0/65536.0,1,-nbitq), 
to_sfixed(-531.0/65536.0,1,-nbitq), 
to_sfixed(4380.0/65536.0,1,-nbitq), 
to_sfixed(2179.0/65536.0,1,-nbitq), 
to_sfixed(8902.0/65536.0,1,-nbitq), 
to_sfixed(7177.0/65536.0,1,-nbitq), 
to_sfixed(207.0/65536.0,1,-nbitq), 
to_sfixed(-2925.0/65536.0,1,-nbitq), 
to_sfixed(1608.0/65536.0,1,-nbitq), 
to_sfixed(-1574.0/65536.0,1,-nbitq), 
to_sfixed(-361.0/65536.0,1,-nbitq), 
to_sfixed(3636.0/65536.0,1,-nbitq), 
to_sfixed(2795.0/65536.0,1,-nbitq), 
to_sfixed(284.0/65536.0,1,-nbitq), 
to_sfixed(-2041.0/65536.0,1,-nbitq), 
to_sfixed(-1747.0/65536.0,1,-nbitq), 
to_sfixed(-1597.0/65536.0,1,-nbitq), 
to_sfixed(1911.0/65536.0,1,-nbitq), 
to_sfixed(4555.0/65536.0,1,-nbitq), 
to_sfixed(-2535.0/65536.0,1,-nbitq), 
to_sfixed(1006.0/65536.0,1,-nbitq), 
to_sfixed(-742.0/65536.0,1,-nbitq), 
to_sfixed(-466.0/65536.0,1,-nbitq), 
to_sfixed(-1325.0/65536.0,1,-nbitq), 
to_sfixed(-646.0/65536.0,1,-nbitq), 
to_sfixed(5549.0/65536.0,1,-nbitq), 
to_sfixed(200.0/65536.0,1,-nbitq), 
to_sfixed(-2697.0/65536.0,1,-nbitq), 
to_sfixed(6596.0/65536.0,1,-nbitq), 
to_sfixed(1409.0/65536.0,1,-nbitq), 
to_sfixed(3617.0/65536.0,1,-nbitq), 
to_sfixed(-3187.0/65536.0,1,-nbitq), 
to_sfixed(1006.0/65536.0,1,-nbitq), 
to_sfixed(5524.0/65536.0,1,-nbitq), 
to_sfixed(1155.0/65536.0,1,-nbitq), 
to_sfixed(-1425.0/65536.0,1,-nbitq), 
to_sfixed(7562.0/65536.0,1,-nbitq), 
to_sfixed(-2416.0/65536.0,1,-nbitq), 
to_sfixed(-5465.0/65536.0,1,-nbitq), 
to_sfixed(1154.0/65536.0,1,-nbitq), 
to_sfixed(-5717.0/65536.0,1,-nbitq), 
to_sfixed(-701.0/65536.0,1,-nbitq), 
to_sfixed(-6620.0/65536.0,1,-nbitq), 
to_sfixed(1053.0/65536.0,1,-nbitq), 
to_sfixed(-28.0/65536.0,1,-nbitq), 
to_sfixed(-7917.0/65536.0,1,-nbitq), 
to_sfixed(-35.0/65536.0,1,-nbitq), 
to_sfixed(-5892.0/65536.0,1,-nbitq), 
to_sfixed(-2436.0/65536.0,1,-nbitq), 
to_sfixed(-430.0/65536.0,1,-nbitq), 
to_sfixed(1645.0/65536.0,1,-nbitq), 
to_sfixed(-7255.0/65536.0,1,-nbitq), 
to_sfixed(-6099.0/65536.0,1,-nbitq), 
to_sfixed(5873.0/65536.0,1,-nbitq), 
to_sfixed(-3120.0/65536.0,1,-nbitq), 
to_sfixed(-3610.0/65536.0,1,-nbitq), 
to_sfixed(1193.0/65536.0,1,-nbitq), 
to_sfixed(578.0/65536.0,1,-nbitq), 
to_sfixed(1238.0/65536.0,1,-nbitq), 
to_sfixed(7953.0/65536.0,1,-nbitq), 
to_sfixed(-1607.0/65536.0,1,-nbitq), 
to_sfixed(1005.0/65536.0,1,-nbitq), 
to_sfixed(1979.0/65536.0,1,-nbitq), 
to_sfixed(-3423.0/65536.0,1,-nbitq), 
to_sfixed(-633.0/65536.0,1,-nbitq), 
to_sfixed(634.0/65536.0,1,-nbitq), 
to_sfixed(-1331.0/65536.0,1,-nbitq), 
to_sfixed(4705.0/65536.0,1,-nbitq), 
to_sfixed(2814.0/65536.0,1,-nbitq), 
to_sfixed(-685.0/65536.0,1,-nbitq), 
to_sfixed(-5495.0/65536.0,1,-nbitq), 
to_sfixed(-2903.0/65536.0,1,-nbitq), 
to_sfixed(7987.0/65536.0,1,-nbitq), 
to_sfixed(1073.0/65536.0,1,-nbitq), 
to_sfixed(1846.0/65536.0,1,-nbitq), 
to_sfixed(2521.0/65536.0,1,-nbitq), 
to_sfixed(5745.0/65536.0,1,-nbitq), 
to_sfixed(-5624.0/65536.0,1,-nbitq), 
to_sfixed(-291.0/65536.0,1,-nbitq), 
to_sfixed(51.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1726.0/65536.0,1,-nbitq), 
to_sfixed(1569.0/65536.0,1,-nbitq), 
to_sfixed(3440.0/65536.0,1,-nbitq), 
to_sfixed(-2389.0/65536.0,1,-nbitq), 
to_sfixed(4543.0/65536.0,1,-nbitq), 
to_sfixed(10268.0/65536.0,1,-nbitq), 
to_sfixed(3861.0/65536.0,1,-nbitq), 
to_sfixed(-3453.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(2489.0/65536.0,1,-nbitq), 
to_sfixed(4338.0/65536.0,1,-nbitq), 
to_sfixed(452.0/65536.0,1,-nbitq), 
to_sfixed(-302.0/65536.0,1,-nbitq), 
to_sfixed(1473.0/65536.0,1,-nbitq), 
to_sfixed(-1576.0/65536.0,1,-nbitq), 
to_sfixed(-1030.0/65536.0,1,-nbitq), 
to_sfixed(-2433.0/65536.0,1,-nbitq), 
to_sfixed(-3457.0/65536.0,1,-nbitq), 
to_sfixed(2236.0/65536.0,1,-nbitq), 
to_sfixed(823.0/65536.0,1,-nbitq), 
to_sfixed(-301.0/65536.0,1,-nbitq), 
to_sfixed(-383.0/65536.0,1,-nbitq), 
to_sfixed(2987.0/65536.0,1,-nbitq), 
to_sfixed(3091.0/65536.0,1,-nbitq), 
to_sfixed(-1203.0/65536.0,1,-nbitq), 
to_sfixed(3848.0/65536.0,1,-nbitq), 
to_sfixed(-5217.0/65536.0,1,-nbitq), 
to_sfixed(1562.0/65536.0,1,-nbitq), 
to_sfixed(5086.0/65536.0,1,-nbitq), 
to_sfixed(1790.0/65536.0,1,-nbitq), 
to_sfixed(6167.0/65536.0,1,-nbitq), 
to_sfixed(1937.0/65536.0,1,-nbitq), 
to_sfixed(1110.0/65536.0,1,-nbitq), 
to_sfixed(7207.0/65536.0,1,-nbitq), 
to_sfixed(792.0/65536.0,1,-nbitq), 
to_sfixed(-2270.0/65536.0,1,-nbitq), 
to_sfixed(7080.0/65536.0,1,-nbitq), 
to_sfixed(2218.0/65536.0,1,-nbitq), 
to_sfixed(-2372.0/65536.0,1,-nbitq), 
to_sfixed(-742.0/65536.0,1,-nbitq), 
to_sfixed(2192.0/65536.0,1,-nbitq), 
to_sfixed(1510.0/65536.0,1,-nbitq), 
to_sfixed(3031.0/65536.0,1,-nbitq), 
to_sfixed(-610.0/65536.0,1,-nbitq), 
to_sfixed(454.0/65536.0,1,-nbitq), 
to_sfixed(-6016.0/65536.0,1,-nbitq), 
to_sfixed(-2446.0/65536.0,1,-nbitq), 
to_sfixed(-8954.0/65536.0,1,-nbitq), 
to_sfixed(-299.0/65536.0,1,-nbitq), 
to_sfixed(-142.0/65536.0,1,-nbitq), 
to_sfixed(2270.0/65536.0,1,-nbitq), 
to_sfixed(-10706.0/65536.0,1,-nbitq), 
to_sfixed(-5790.0/65536.0,1,-nbitq), 
to_sfixed(-4462.0/65536.0,1,-nbitq), 
to_sfixed(5848.0/65536.0,1,-nbitq), 
to_sfixed(5425.0/65536.0,1,-nbitq), 
to_sfixed(1930.0/65536.0,1,-nbitq), 
to_sfixed(-1334.0/65536.0,1,-nbitq), 
to_sfixed(-451.0/65536.0,1,-nbitq), 
to_sfixed(153.0/65536.0,1,-nbitq), 
to_sfixed(-863.0/65536.0,1,-nbitq), 
to_sfixed(2250.0/65536.0,1,-nbitq), 
to_sfixed(1332.0/65536.0,1,-nbitq), 
to_sfixed(1134.0/65536.0,1,-nbitq), 
to_sfixed(3263.0/65536.0,1,-nbitq), 
to_sfixed(-2134.0/65536.0,1,-nbitq), 
to_sfixed(-4010.0/65536.0,1,-nbitq), 
to_sfixed(2356.0/65536.0,1,-nbitq), 
to_sfixed(1631.0/65536.0,1,-nbitq), 
to_sfixed(-5086.0/65536.0,1,-nbitq), 
to_sfixed(34.0/65536.0,1,-nbitq), 
to_sfixed(-3862.0/65536.0,1,-nbitq), 
to_sfixed(-169.0/65536.0,1,-nbitq), 
to_sfixed(1576.0/65536.0,1,-nbitq), 
to_sfixed(1900.0/65536.0,1,-nbitq), 
to_sfixed(1887.0/65536.0,1,-nbitq), 
to_sfixed(9239.0/65536.0,1,-nbitq), 
to_sfixed(-10441.0/65536.0,1,-nbitq), 
to_sfixed(-1692.0/65536.0,1,-nbitq), 
to_sfixed(-2606.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3226.0/65536.0,1,-nbitq), 
to_sfixed(1828.0/65536.0,1,-nbitq), 
to_sfixed(3619.0/65536.0,1,-nbitq), 
to_sfixed(-3279.0/65536.0,1,-nbitq), 
to_sfixed(1457.0/65536.0,1,-nbitq), 
to_sfixed(7846.0/65536.0,1,-nbitq), 
to_sfixed(1527.0/65536.0,1,-nbitq), 
to_sfixed(1557.0/65536.0,1,-nbitq), 
to_sfixed(3293.0/65536.0,1,-nbitq), 
to_sfixed(-2174.0/65536.0,1,-nbitq), 
to_sfixed(5390.0/65536.0,1,-nbitq), 
to_sfixed(-8521.0/65536.0,1,-nbitq), 
to_sfixed(1817.0/65536.0,1,-nbitq), 
to_sfixed(5428.0/65536.0,1,-nbitq), 
to_sfixed(-3786.0/65536.0,1,-nbitq), 
to_sfixed(-2827.0/65536.0,1,-nbitq), 
to_sfixed(-1721.0/65536.0,1,-nbitq), 
to_sfixed(-3278.0/65536.0,1,-nbitq), 
to_sfixed(1764.0/65536.0,1,-nbitq), 
to_sfixed(-1285.0/65536.0,1,-nbitq), 
to_sfixed(18.0/65536.0,1,-nbitq), 
to_sfixed(151.0/65536.0,1,-nbitq), 
to_sfixed(5723.0/65536.0,1,-nbitq), 
to_sfixed(8162.0/65536.0,1,-nbitq), 
to_sfixed(643.0/65536.0,1,-nbitq), 
to_sfixed(1473.0/65536.0,1,-nbitq), 
to_sfixed(-1597.0/65536.0,1,-nbitq), 
to_sfixed(-2493.0/65536.0,1,-nbitq), 
to_sfixed(-314.0/65536.0,1,-nbitq), 
to_sfixed(-374.0/65536.0,1,-nbitq), 
to_sfixed(3907.0/65536.0,1,-nbitq), 
to_sfixed(3647.0/65536.0,1,-nbitq), 
to_sfixed(3518.0/65536.0,1,-nbitq), 
to_sfixed(3838.0/65536.0,1,-nbitq), 
to_sfixed(-958.0/65536.0,1,-nbitq), 
to_sfixed(-185.0/65536.0,1,-nbitq), 
to_sfixed(3715.0/65536.0,1,-nbitq), 
to_sfixed(3135.0/65536.0,1,-nbitq), 
to_sfixed(179.0/65536.0,1,-nbitq), 
to_sfixed(943.0/65536.0,1,-nbitq), 
to_sfixed(9098.0/65536.0,1,-nbitq), 
to_sfixed(625.0/65536.0,1,-nbitq), 
to_sfixed(-10.0/65536.0,1,-nbitq), 
to_sfixed(-4098.0/65536.0,1,-nbitq), 
to_sfixed(-1666.0/65536.0,1,-nbitq), 
to_sfixed(-260.0/65536.0,1,-nbitq), 
to_sfixed(-1183.0/65536.0,1,-nbitq), 
to_sfixed(-6552.0/65536.0,1,-nbitq), 
to_sfixed(1590.0/65536.0,1,-nbitq), 
to_sfixed(-1321.0/65536.0,1,-nbitq), 
to_sfixed(2123.0/65536.0,1,-nbitq), 
to_sfixed(-10635.0/65536.0,1,-nbitq), 
to_sfixed(-11158.0/65536.0,1,-nbitq), 
to_sfixed(-6113.0/65536.0,1,-nbitq), 
to_sfixed(2480.0/65536.0,1,-nbitq), 
to_sfixed(7520.0/65536.0,1,-nbitq), 
to_sfixed(2553.0/65536.0,1,-nbitq), 
to_sfixed(-3886.0/65536.0,1,-nbitq), 
to_sfixed(474.0/65536.0,1,-nbitq), 
to_sfixed(-4514.0/65536.0,1,-nbitq), 
to_sfixed(-1127.0/65536.0,1,-nbitq), 
to_sfixed(-306.0/65536.0,1,-nbitq), 
to_sfixed(277.0/65536.0,1,-nbitq), 
to_sfixed(2200.0/65536.0,1,-nbitq), 
to_sfixed(-343.0/65536.0,1,-nbitq), 
to_sfixed(-4025.0/65536.0,1,-nbitq), 
to_sfixed(-3833.0/65536.0,1,-nbitq), 
to_sfixed(-2336.0/65536.0,1,-nbitq), 
to_sfixed(5397.0/65536.0,1,-nbitq), 
to_sfixed(-4623.0/65536.0,1,-nbitq), 
to_sfixed(-1352.0/65536.0,1,-nbitq), 
to_sfixed(-1286.0/65536.0,1,-nbitq), 
to_sfixed(2789.0/65536.0,1,-nbitq), 
to_sfixed(980.0/65536.0,1,-nbitq), 
to_sfixed(-2432.0/65536.0,1,-nbitq), 
to_sfixed(2275.0/65536.0,1,-nbitq), 
to_sfixed(11161.0/65536.0,1,-nbitq), 
to_sfixed(-6307.0/65536.0,1,-nbitq), 
to_sfixed(-1118.0/65536.0,1,-nbitq), 
to_sfixed(1125.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1426.0/65536.0,1,-nbitq), 
to_sfixed(335.0/65536.0,1,-nbitq), 
to_sfixed(-419.0/65536.0,1,-nbitq), 
to_sfixed(700.0/65536.0,1,-nbitq), 
to_sfixed(5386.0/65536.0,1,-nbitq), 
to_sfixed(4382.0/65536.0,1,-nbitq), 
to_sfixed(193.0/65536.0,1,-nbitq), 
to_sfixed(-1817.0/65536.0,1,-nbitq), 
to_sfixed(-853.0/65536.0,1,-nbitq), 
to_sfixed(-2510.0/65536.0,1,-nbitq), 
to_sfixed(4555.0/65536.0,1,-nbitq), 
to_sfixed(-2236.0/65536.0,1,-nbitq), 
to_sfixed(1684.0/65536.0,1,-nbitq), 
to_sfixed(8265.0/65536.0,1,-nbitq), 
to_sfixed(621.0/65536.0,1,-nbitq), 
to_sfixed(533.0/65536.0,1,-nbitq), 
to_sfixed(156.0/65536.0,1,-nbitq), 
to_sfixed(-2808.0/65536.0,1,-nbitq), 
to_sfixed(-1303.0/65536.0,1,-nbitq), 
to_sfixed(179.0/65536.0,1,-nbitq), 
to_sfixed(-490.0/65536.0,1,-nbitq), 
to_sfixed(1035.0/65536.0,1,-nbitq), 
to_sfixed(4535.0/65536.0,1,-nbitq), 
to_sfixed(8565.0/65536.0,1,-nbitq), 
to_sfixed(-506.0/65536.0,1,-nbitq), 
to_sfixed(5265.0/65536.0,1,-nbitq), 
to_sfixed(-291.0/65536.0,1,-nbitq), 
to_sfixed(-738.0/65536.0,1,-nbitq), 
to_sfixed(-703.0/65536.0,1,-nbitq), 
to_sfixed(2006.0/65536.0,1,-nbitq), 
to_sfixed(-2132.0/65536.0,1,-nbitq), 
to_sfixed(654.0/65536.0,1,-nbitq), 
to_sfixed(1143.0/65536.0,1,-nbitq), 
to_sfixed(-5433.0/65536.0,1,-nbitq), 
to_sfixed(-3269.0/65536.0,1,-nbitq), 
to_sfixed(-3796.0/65536.0,1,-nbitq), 
to_sfixed(1262.0/65536.0,1,-nbitq), 
to_sfixed(595.0/65536.0,1,-nbitq), 
to_sfixed(4977.0/65536.0,1,-nbitq), 
to_sfixed(2436.0/65536.0,1,-nbitq), 
to_sfixed(8310.0/65536.0,1,-nbitq), 
to_sfixed(-975.0/65536.0,1,-nbitq), 
to_sfixed(1843.0/65536.0,1,-nbitq), 
to_sfixed(-408.0/65536.0,1,-nbitq), 
to_sfixed(-2376.0/65536.0,1,-nbitq), 
to_sfixed(413.0/65536.0,1,-nbitq), 
to_sfixed(-2477.0/65536.0,1,-nbitq), 
to_sfixed(3163.0/65536.0,1,-nbitq), 
to_sfixed(2020.0/65536.0,1,-nbitq), 
to_sfixed(197.0/65536.0,1,-nbitq), 
to_sfixed(3062.0/65536.0,1,-nbitq), 
to_sfixed(-4925.0/65536.0,1,-nbitq), 
to_sfixed(-7225.0/65536.0,1,-nbitq), 
to_sfixed(199.0/65536.0,1,-nbitq), 
to_sfixed(1414.0/65536.0,1,-nbitq), 
to_sfixed(5994.0/65536.0,1,-nbitq), 
to_sfixed(-2010.0/65536.0,1,-nbitq), 
to_sfixed(1120.0/65536.0,1,-nbitq), 
to_sfixed(362.0/65536.0,1,-nbitq), 
to_sfixed(-1951.0/65536.0,1,-nbitq), 
to_sfixed(-4213.0/65536.0,1,-nbitq), 
to_sfixed(839.0/65536.0,1,-nbitq), 
to_sfixed(-157.0/65536.0,1,-nbitq), 
to_sfixed(-1550.0/65536.0,1,-nbitq), 
to_sfixed(-4079.0/65536.0,1,-nbitq), 
to_sfixed(-3692.0/65536.0,1,-nbitq), 
to_sfixed(-5970.0/65536.0,1,-nbitq), 
to_sfixed(-3104.0/65536.0,1,-nbitq), 
to_sfixed(-4533.0/65536.0,1,-nbitq), 
to_sfixed(-3710.0/65536.0,1,-nbitq), 
to_sfixed(-1571.0/65536.0,1,-nbitq), 
to_sfixed(-1783.0/65536.0,1,-nbitq), 
to_sfixed(1101.0/65536.0,1,-nbitq), 
to_sfixed(-643.0/65536.0,1,-nbitq), 
to_sfixed(-1105.0/65536.0,1,-nbitq), 
to_sfixed(1133.0/65536.0,1,-nbitq), 
to_sfixed(9043.0/65536.0,1,-nbitq), 
to_sfixed(-6152.0/65536.0,1,-nbitq), 
to_sfixed(1929.0/65536.0,1,-nbitq), 
to_sfixed(-2171.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4885.0/65536.0,1,-nbitq), 
to_sfixed(2138.0/65536.0,1,-nbitq), 
to_sfixed(3818.0/65536.0,1,-nbitq), 
to_sfixed(2317.0/65536.0,1,-nbitq), 
to_sfixed(3067.0/65536.0,1,-nbitq), 
to_sfixed(2236.0/65536.0,1,-nbitq), 
to_sfixed(-509.0/65536.0,1,-nbitq), 
to_sfixed(-1443.0/65536.0,1,-nbitq), 
to_sfixed(1279.0/65536.0,1,-nbitq), 
to_sfixed(2023.0/65536.0,1,-nbitq), 
to_sfixed(2380.0/65536.0,1,-nbitq), 
to_sfixed(3004.0/65536.0,1,-nbitq), 
to_sfixed(1146.0/65536.0,1,-nbitq), 
to_sfixed(4907.0/65536.0,1,-nbitq), 
to_sfixed(-470.0/65536.0,1,-nbitq), 
to_sfixed(1281.0/65536.0,1,-nbitq), 
to_sfixed(2713.0/65536.0,1,-nbitq), 
to_sfixed(-197.0/65536.0,1,-nbitq), 
to_sfixed(-1505.0/65536.0,1,-nbitq), 
to_sfixed(2695.0/65536.0,1,-nbitq), 
to_sfixed(-3068.0/65536.0,1,-nbitq), 
to_sfixed(1775.0/65536.0,1,-nbitq), 
to_sfixed(-1265.0/65536.0,1,-nbitq), 
to_sfixed(1520.0/65536.0,1,-nbitq), 
to_sfixed(90.0/65536.0,1,-nbitq), 
to_sfixed(4625.0/65536.0,1,-nbitq), 
to_sfixed(3041.0/65536.0,1,-nbitq), 
to_sfixed(2115.0/65536.0,1,-nbitq), 
to_sfixed(-3054.0/65536.0,1,-nbitq), 
to_sfixed(-1825.0/65536.0,1,-nbitq), 
to_sfixed(773.0/65536.0,1,-nbitq), 
to_sfixed(-3004.0/65536.0,1,-nbitq), 
to_sfixed(4789.0/65536.0,1,-nbitq), 
to_sfixed(-2445.0/65536.0,1,-nbitq), 
to_sfixed(-3344.0/65536.0,1,-nbitq), 
to_sfixed(633.0/65536.0,1,-nbitq), 
to_sfixed(795.0/65536.0,1,-nbitq), 
to_sfixed(-2872.0/65536.0,1,-nbitq), 
to_sfixed(7281.0/65536.0,1,-nbitq), 
to_sfixed(-242.0/65536.0,1,-nbitq), 
to_sfixed(8375.0/65536.0,1,-nbitq), 
to_sfixed(-1994.0/65536.0,1,-nbitq), 
to_sfixed(-462.0/65536.0,1,-nbitq), 
to_sfixed(195.0/65536.0,1,-nbitq), 
to_sfixed(2726.0/65536.0,1,-nbitq), 
to_sfixed(1996.0/65536.0,1,-nbitq), 
to_sfixed(-86.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(800.0/65536.0,1,-nbitq), 
to_sfixed(1145.0/65536.0,1,-nbitq), 
to_sfixed(-1124.0/65536.0,1,-nbitq), 
to_sfixed(-5198.0/65536.0,1,-nbitq), 
to_sfixed(-5201.0/65536.0,1,-nbitq), 
to_sfixed(-815.0/65536.0,1,-nbitq), 
to_sfixed(2113.0/65536.0,1,-nbitq), 
to_sfixed(1644.0/65536.0,1,-nbitq), 
to_sfixed(-951.0/65536.0,1,-nbitq), 
to_sfixed(1711.0/65536.0,1,-nbitq), 
to_sfixed(2057.0/65536.0,1,-nbitq), 
to_sfixed(4739.0/65536.0,1,-nbitq), 
to_sfixed(2776.0/65536.0,1,-nbitq), 
to_sfixed(2014.0/65536.0,1,-nbitq), 
to_sfixed(-295.0/65536.0,1,-nbitq), 
to_sfixed(-1777.0/65536.0,1,-nbitq), 
to_sfixed(-3205.0/65536.0,1,-nbitq), 
to_sfixed(-1379.0/65536.0,1,-nbitq), 
to_sfixed(-5323.0/65536.0,1,-nbitq), 
to_sfixed(-9224.0/65536.0,1,-nbitq), 
to_sfixed(-5759.0/65536.0,1,-nbitq), 
to_sfixed(-7379.0/65536.0,1,-nbitq), 
to_sfixed(-55.0/65536.0,1,-nbitq), 
to_sfixed(-5211.0/65536.0,1,-nbitq), 
to_sfixed(4846.0/65536.0,1,-nbitq), 
to_sfixed(-2776.0/65536.0,1,-nbitq), 
to_sfixed(2021.0/65536.0,1,-nbitq), 
to_sfixed(-2433.0/65536.0,1,-nbitq), 
to_sfixed(1986.0/65536.0,1,-nbitq), 
to_sfixed(-4554.0/65536.0,1,-nbitq), 
to_sfixed(606.0/65536.0,1,-nbitq), 
to_sfixed(-692.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2266.0/65536.0,1,-nbitq), 
to_sfixed(-1627.0/65536.0,1,-nbitq), 
to_sfixed(1733.0/65536.0,1,-nbitq), 
to_sfixed(3284.0/65536.0,1,-nbitq), 
to_sfixed(3320.0/65536.0,1,-nbitq), 
to_sfixed(2064.0/65536.0,1,-nbitq), 
to_sfixed(-2296.0/65536.0,1,-nbitq), 
to_sfixed(-1467.0/65536.0,1,-nbitq), 
to_sfixed(-2333.0/65536.0,1,-nbitq), 
to_sfixed(1773.0/65536.0,1,-nbitq), 
to_sfixed(-91.0/65536.0,1,-nbitq), 
to_sfixed(3625.0/65536.0,1,-nbitq), 
to_sfixed(-1771.0/65536.0,1,-nbitq), 
to_sfixed(5423.0/65536.0,1,-nbitq), 
to_sfixed(1233.0/65536.0,1,-nbitq), 
to_sfixed(2498.0/65536.0,1,-nbitq), 
to_sfixed(1671.0/65536.0,1,-nbitq), 
to_sfixed(589.0/65536.0,1,-nbitq), 
to_sfixed(-662.0/65536.0,1,-nbitq), 
to_sfixed(-2194.0/65536.0,1,-nbitq), 
to_sfixed(-3688.0/65536.0,1,-nbitq), 
to_sfixed(2795.0/65536.0,1,-nbitq), 
to_sfixed(1317.0/65536.0,1,-nbitq), 
to_sfixed(2181.0/65536.0,1,-nbitq), 
to_sfixed(-1499.0/65536.0,1,-nbitq), 
to_sfixed(-248.0/65536.0,1,-nbitq), 
to_sfixed(23.0/65536.0,1,-nbitq), 
to_sfixed(2320.0/65536.0,1,-nbitq), 
to_sfixed(-1514.0/65536.0,1,-nbitq), 
to_sfixed(518.0/65536.0,1,-nbitq), 
to_sfixed(-248.0/65536.0,1,-nbitq), 
to_sfixed(363.0/65536.0,1,-nbitq), 
to_sfixed(5551.0/65536.0,1,-nbitq), 
to_sfixed(465.0/65536.0,1,-nbitq), 
to_sfixed(-1762.0/65536.0,1,-nbitq), 
to_sfixed(2170.0/65536.0,1,-nbitq), 
to_sfixed(-327.0/65536.0,1,-nbitq), 
to_sfixed(1463.0/65536.0,1,-nbitq), 
to_sfixed(-938.0/65536.0,1,-nbitq), 
to_sfixed(1151.0/65536.0,1,-nbitq), 
to_sfixed(2433.0/65536.0,1,-nbitq), 
to_sfixed(799.0/65536.0,1,-nbitq), 
to_sfixed(1047.0/65536.0,1,-nbitq), 
to_sfixed(373.0/65536.0,1,-nbitq), 
to_sfixed(3355.0/65536.0,1,-nbitq), 
to_sfixed(2634.0/65536.0,1,-nbitq), 
to_sfixed(220.0/65536.0,1,-nbitq), 
to_sfixed(-843.0/65536.0,1,-nbitq), 
to_sfixed(-1766.0/65536.0,1,-nbitq), 
to_sfixed(215.0/65536.0,1,-nbitq), 
to_sfixed(1240.0/65536.0,1,-nbitq), 
to_sfixed(-6394.0/65536.0,1,-nbitq), 
to_sfixed(1682.0/65536.0,1,-nbitq), 
to_sfixed(-3322.0/65536.0,1,-nbitq), 
to_sfixed(1874.0/65536.0,1,-nbitq), 
to_sfixed(-1377.0/65536.0,1,-nbitq), 
to_sfixed(389.0/65536.0,1,-nbitq), 
to_sfixed(2731.0/65536.0,1,-nbitq), 
to_sfixed(2661.0/65536.0,1,-nbitq), 
to_sfixed(384.0/65536.0,1,-nbitq), 
to_sfixed(-1346.0/65536.0,1,-nbitq), 
to_sfixed(-1714.0/65536.0,1,-nbitq), 
to_sfixed(2088.0/65536.0,1,-nbitq), 
to_sfixed(-256.0/65536.0,1,-nbitq), 
to_sfixed(371.0/65536.0,1,-nbitq), 
to_sfixed(-2007.0/65536.0,1,-nbitq), 
to_sfixed(-6602.0/65536.0,1,-nbitq), 
to_sfixed(-2227.0/65536.0,1,-nbitq), 
to_sfixed(-5426.0/65536.0,1,-nbitq), 
to_sfixed(-5182.0/65536.0,1,-nbitq), 
to_sfixed(-511.0/65536.0,1,-nbitq), 
to_sfixed(-3210.0/65536.0,1,-nbitq), 
to_sfixed(378.0/65536.0,1,-nbitq), 
to_sfixed(792.0/65536.0,1,-nbitq), 
to_sfixed(-941.0/65536.0,1,-nbitq), 
to_sfixed(3671.0/65536.0,1,-nbitq), 
to_sfixed(-4009.0/65536.0,1,-nbitq), 
to_sfixed(-3809.0/65536.0,1,-nbitq), 
to_sfixed(1405.0/65536.0,1,-nbitq), 
to_sfixed(-4000.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1856.0/65536.0,1,-nbitq), 
to_sfixed(-3237.0/65536.0,1,-nbitq), 
to_sfixed(663.0/65536.0,1,-nbitq), 
to_sfixed(-1304.0/65536.0,1,-nbitq), 
to_sfixed(-390.0/65536.0,1,-nbitq), 
to_sfixed(-762.0/65536.0,1,-nbitq), 
to_sfixed(1095.0/65536.0,1,-nbitq), 
to_sfixed(-241.0/65536.0,1,-nbitq), 
to_sfixed(-281.0/65536.0,1,-nbitq), 
to_sfixed(2997.0/65536.0,1,-nbitq), 
to_sfixed(-1024.0/65536.0,1,-nbitq), 
to_sfixed(3027.0/65536.0,1,-nbitq), 
to_sfixed(2075.0/65536.0,1,-nbitq), 
to_sfixed(-281.0/65536.0,1,-nbitq), 
to_sfixed(138.0/65536.0,1,-nbitq), 
to_sfixed(1998.0/65536.0,1,-nbitq), 
to_sfixed(1972.0/65536.0,1,-nbitq), 
to_sfixed(-2362.0/65536.0,1,-nbitq), 
to_sfixed(-3217.0/65536.0,1,-nbitq), 
to_sfixed(655.0/65536.0,1,-nbitq), 
to_sfixed(871.0/65536.0,1,-nbitq), 
to_sfixed(-677.0/65536.0,1,-nbitq), 
to_sfixed(2161.0/65536.0,1,-nbitq), 
to_sfixed(4294.0/65536.0,1,-nbitq), 
to_sfixed(909.0/65536.0,1,-nbitq), 
to_sfixed(1994.0/65536.0,1,-nbitq), 
to_sfixed(-189.0/65536.0,1,-nbitq), 
to_sfixed(3212.0/65536.0,1,-nbitq), 
to_sfixed(-3333.0/65536.0,1,-nbitq), 
to_sfixed(3611.0/65536.0,1,-nbitq), 
to_sfixed(-1131.0/65536.0,1,-nbitq), 
to_sfixed(2514.0/65536.0,1,-nbitq), 
to_sfixed(4717.0/65536.0,1,-nbitq), 
to_sfixed(5511.0/65536.0,1,-nbitq), 
to_sfixed(-538.0/65536.0,1,-nbitq), 
to_sfixed(-1640.0/65536.0,1,-nbitq), 
to_sfixed(1378.0/65536.0,1,-nbitq), 
to_sfixed(1262.0/65536.0,1,-nbitq), 
to_sfixed(605.0/65536.0,1,-nbitq), 
to_sfixed(-1304.0/65536.0,1,-nbitq), 
to_sfixed(-5855.0/65536.0,1,-nbitq), 
to_sfixed(-531.0/65536.0,1,-nbitq), 
to_sfixed(2254.0/65536.0,1,-nbitq), 
to_sfixed(-33.0/65536.0,1,-nbitq), 
to_sfixed(309.0/65536.0,1,-nbitq), 
to_sfixed(2365.0/65536.0,1,-nbitq), 
to_sfixed(-1383.0/65536.0,1,-nbitq), 
to_sfixed(-2922.0/65536.0,1,-nbitq), 
to_sfixed(1327.0/65536.0,1,-nbitq), 
to_sfixed(1767.0/65536.0,1,-nbitq), 
to_sfixed(3084.0/65536.0,1,-nbitq), 
to_sfixed(-6051.0/65536.0,1,-nbitq), 
to_sfixed(4219.0/65536.0,1,-nbitq), 
to_sfixed(-3240.0/65536.0,1,-nbitq), 
to_sfixed(2081.0/65536.0,1,-nbitq), 
to_sfixed(2859.0/65536.0,1,-nbitq), 
to_sfixed(-349.0/65536.0,1,-nbitq), 
to_sfixed(1746.0/65536.0,1,-nbitq), 
to_sfixed(-1733.0/65536.0,1,-nbitq), 
to_sfixed(3167.0/65536.0,1,-nbitq), 
to_sfixed(-1370.0/65536.0,1,-nbitq), 
to_sfixed(-2606.0/65536.0,1,-nbitq), 
to_sfixed(-121.0/65536.0,1,-nbitq), 
to_sfixed(726.0/65536.0,1,-nbitq), 
to_sfixed(-1420.0/65536.0,1,-nbitq), 
to_sfixed(-376.0/65536.0,1,-nbitq), 
to_sfixed(-1178.0/65536.0,1,-nbitq), 
to_sfixed(-98.0/65536.0,1,-nbitq), 
to_sfixed(-5927.0/65536.0,1,-nbitq), 
to_sfixed(-1390.0/65536.0,1,-nbitq), 
to_sfixed(-352.0/65536.0,1,-nbitq), 
to_sfixed(-4659.0/65536.0,1,-nbitq), 
to_sfixed(2037.0/65536.0,1,-nbitq), 
to_sfixed(-3243.0/65536.0,1,-nbitq), 
to_sfixed(386.0/65536.0,1,-nbitq), 
to_sfixed(5553.0/65536.0,1,-nbitq), 
to_sfixed(-2227.0/65536.0,1,-nbitq), 
to_sfixed(1815.0/65536.0,1,-nbitq), 
to_sfixed(-2392.0/65536.0,1,-nbitq), 
to_sfixed(-671.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3916.0/65536.0,1,-nbitq), 
to_sfixed(-2618.0/65536.0,1,-nbitq), 
to_sfixed(-978.0/65536.0,1,-nbitq), 
to_sfixed(1187.0/65536.0,1,-nbitq), 
to_sfixed(1235.0/65536.0,1,-nbitq), 
to_sfixed(-1859.0/65536.0,1,-nbitq), 
to_sfixed(-3354.0/65536.0,1,-nbitq), 
to_sfixed(1588.0/65536.0,1,-nbitq), 
to_sfixed(1771.0/65536.0,1,-nbitq), 
to_sfixed(-1363.0/65536.0,1,-nbitq), 
to_sfixed(-398.0/65536.0,1,-nbitq), 
to_sfixed(3038.0/65536.0,1,-nbitq), 
to_sfixed(105.0/65536.0,1,-nbitq), 
to_sfixed(-1967.0/65536.0,1,-nbitq), 
to_sfixed(1650.0/65536.0,1,-nbitq), 
to_sfixed(1286.0/65536.0,1,-nbitq), 
to_sfixed(-2741.0/65536.0,1,-nbitq), 
to_sfixed(-2996.0/65536.0,1,-nbitq), 
to_sfixed(1616.0/65536.0,1,-nbitq), 
to_sfixed(-2488.0/65536.0,1,-nbitq), 
to_sfixed(323.0/65536.0,1,-nbitq), 
to_sfixed(1327.0/65536.0,1,-nbitq), 
to_sfixed(1926.0/65536.0,1,-nbitq), 
to_sfixed(32.0/65536.0,1,-nbitq), 
to_sfixed(3047.0/65536.0,1,-nbitq), 
to_sfixed(125.0/65536.0,1,-nbitq), 
to_sfixed(3366.0/65536.0,1,-nbitq), 
to_sfixed(-1209.0/65536.0,1,-nbitq), 
to_sfixed(-281.0/65536.0,1,-nbitq), 
to_sfixed(-1153.0/65536.0,1,-nbitq), 
to_sfixed(437.0/65536.0,1,-nbitq), 
to_sfixed(2336.0/65536.0,1,-nbitq), 
to_sfixed(-440.0/65536.0,1,-nbitq), 
to_sfixed(2373.0/65536.0,1,-nbitq), 
to_sfixed(704.0/65536.0,1,-nbitq), 
to_sfixed(-2134.0/65536.0,1,-nbitq), 
to_sfixed(2601.0/65536.0,1,-nbitq), 
to_sfixed(815.0/65536.0,1,-nbitq), 
to_sfixed(246.0/65536.0,1,-nbitq), 
to_sfixed(1800.0/65536.0,1,-nbitq), 
to_sfixed(-3892.0/65536.0,1,-nbitq), 
to_sfixed(-2926.0/65536.0,1,-nbitq), 
to_sfixed(-1378.0/65536.0,1,-nbitq), 
to_sfixed(-2671.0/65536.0,1,-nbitq), 
to_sfixed(722.0/65536.0,1,-nbitq), 
to_sfixed(1087.0/65536.0,1,-nbitq), 
to_sfixed(-296.0/65536.0,1,-nbitq), 
to_sfixed(-295.0/65536.0,1,-nbitq), 
to_sfixed(3095.0/65536.0,1,-nbitq), 
to_sfixed(-476.0/65536.0,1,-nbitq), 
to_sfixed(1605.0/65536.0,1,-nbitq), 
to_sfixed(-6623.0/65536.0,1,-nbitq), 
to_sfixed(965.0/65536.0,1,-nbitq), 
to_sfixed(-1841.0/65536.0,1,-nbitq), 
to_sfixed(954.0/65536.0,1,-nbitq), 
to_sfixed(1642.0/65536.0,1,-nbitq), 
to_sfixed(-1477.0/65536.0,1,-nbitq), 
to_sfixed(-336.0/65536.0,1,-nbitq), 
to_sfixed(2912.0/65536.0,1,-nbitq), 
to_sfixed(1588.0/65536.0,1,-nbitq), 
to_sfixed(2733.0/65536.0,1,-nbitq), 
to_sfixed(1009.0/65536.0,1,-nbitq), 
to_sfixed(1789.0/65536.0,1,-nbitq), 
to_sfixed(-1366.0/65536.0,1,-nbitq), 
to_sfixed(-1004.0/65536.0,1,-nbitq), 
to_sfixed(3108.0/65536.0,1,-nbitq), 
to_sfixed(-4229.0/65536.0,1,-nbitq), 
to_sfixed(-868.0/65536.0,1,-nbitq), 
to_sfixed(-1086.0/65536.0,1,-nbitq), 
to_sfixed(-244.0/65536.0,1,-nbitq), 
to_sfixed(-471.0/65536.0,1,-nbitq), 
to_sfixed(-4796.0/65536.0,1,-nbitq), 
to_sfixed(-1975.0/65536.0,1,-nbitq), 
to_sfixed(-1236.0/65536.0,1,-nbitq), 
to_sfixed(-721.0/65536.0,1,-nbitq), 
to_sfixed(1372.0/65536.0,1,-nbitq), 
to_sfixed(88.0/65536.0,1,-nbitq), 
to_sfixed(3568.0/65536.0,1,-nbitq), 
to_sfixed(-3251.0/65536.0,1,-nbitq), 
to_sfixed(-785.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-904.0/65536.0,1,-nbitq), 
to_sfixed(-639.0/65536.0,1,-nbitq), 
to_sfixed(-2810.0/65536.0,1,-nbitq), 
to_sfixed(2301.0/65536.0,1,-nbitq), 
to_sfixed(1831.0/65536.0,1,-nbitq), 
to_sfixed(398.0/65536.0,1,-nbitq), 
to_sfixed(-992.0/65536.0,1,-nbitq), 
to_sfixed(-3059.0/65536.0,1,-nbitq), 
to_sfixed(1464.0/65536.0,1,-nbitq), 
to_sfixed(1884.0/65536.0,1,-nbitq), 
to_sfixed(-372.0/65536.0,1,-nbitq), 
to_sfixed(-1303.0/65536.0,1,-nbitq), 
to_sfixed(3299.0/65536.0,1,-nbitq), 
to_sfixed(-3773.0/65536.0,1,-nbitq), 
to_sfixed(1328.0/65536.0,1,-nbitq), 
to_sfixed(-702.0/65536.0,1,-nbitq), 
to_sfixed(-3073.0/65536.0,1,-nbitq), 
to_sfixed(-485.0/65536.0,1,-nbitq), 
to_sfixed(-1491.0/65536.0,1,-nbitq), 
to_sfixed(3072.0/65536.0,1,-nbitq), 
to_sfixed(103.0/65536.0,1,-nbitq), 
to_sfixed(-2875.0/65536.0,1,-nbitq), 
to_sfixed(-1884.0/65536.0,1,-nbitq), 
to_sfixed(1727.0/65536.0,1,-nbitq), 
to_sfixed(1319.0/65536.0,1,-nbitq), 
to_sfixed(2431.0/65536.0,1,-nbitq), 
to_sfixed(-2377.0/65536.0,1,-nbitq), 
to_sfixed(821.0/65536.0,1,-nbitq), 
to_sfixed(-447.0/65536.0,1,-nbitq), 
to_sfixed(-1077.0/65536.0,1,-nbitq), 
to_sfixed(2546.0/65536.0,1,-nbitq), 
to_sfixed(-1196.0/65536.0,1,-nbitq), 
to_sfixed(-102.0/65536.0,1,-nbitq), 
to_sfixed(-2231.0/65536.0,1,-nbitq), 
to_sfixed(1406.0/65536.0,1,-nbitq), 
to_sfixed(-1721.0/65536.0,1,-nbitq), 
to_sfixed(479.0/65536.0,1,-nbitq), 
to_sfixed(-3359.0/65536.0,1,-nbitq), 
to_sfixed(-3941.0/65536.0,1,-nbitq), 
to_sfixed(-1777.0/65536.0,1,-nbitq), 
to_sfixed(-1653.0/65536.0,1,-nbitq), 
to_sfixed(-25.0/65536.0,1,-nbitq), 
to_sfixed(-1673.0/65536.0,1,-nbitq), 
to_sfixed(-1435.0/65536.0,1,-nbitq), 
to_sfixed(-708.0/65536.0,1,-nbitq), 
to_sfixed(-444.0/65536.0,1,-nbitq), 
to_sfixed(-2510.0/65536.0,1,-nbitq), 
to_sfixed(-3564.0/65536.0,1,-nbitq), 
to_sfixed(1096.0/65536.0,1,-nbitq), 
to_sfixed(1926.0/65536.0,1,-nbitq), 
to_sfixed(902.0/65536.0,1,-nbitq), 
to_sfixed(-3242.0/65536.0,1,-nbitq), 
to_sfixed(3148.0/65536.0,1,-nbitq), 
to_sfixed(-856.0/65536.0,1,-nbitq), 
to_sfixed(1980.0/65536.0,1,-nbitq), 
to_sfixed(2972.0/65536.0,1,-nbitq), 
to_sfixed(-1534.0/65536.0,1,-nbitq), 
to_sfixed(-632.0/65536.0,1,-nbitq), 
to_sfixed(-2465.0/65536.0,1,-nbitq), 
to_sfixed(4530.0/65536.0,1,-nbitq), 
to_sfixed(1240.0/65536.0,1,-nbitq), 
to_sfixed(-2271.0/65536.0,1,-nbitq), 
to_sfixed(-165.0/65536.0,1,-nbitq), 
to_sfixed(2577.0/65536.0,1,-nbitq), 
to_sfixed(229.0/65536.0,1,-nbitq), 
to_sfixed(1119.0/65536.0,1,-nbitq), 
to_sfixed(1430.0/65536.0,1,-nbitq), 
to_sfixed(1982.0/65536.0,1,-nbitq), 
to_sfixed(-3497.0/65536.0,1,-nbitq), 
to_sfixed(1124.0/65536.0,1,-nbitq), 
to_sfixed(320.0/65536.0,1,-nbitq), 
to_sfixed(-3179.0/65536.0,1,-nbitq), 
to_sfixed(-2463.0/65536.0,1,-nbitq), 
to_sfixed(-3240.0/65536.0,1,-nbitq), 
to_sfixed(-76.0/65536.0,1,-nbitq), 
to_sfixed(231.0/65536.0,1,-nbitq), 
to_sfixed(-1232.0/65536.0,1,-nbitq), 
to_sfixed(4266.0/65536.0,1,-nbitq), 
to_sfixed(-1960.0/65536.0,1,-nbitq), 
to_sfixed(2860.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2933.0/65536.0,1,-nbitq), 
to_sfixed(1062.0/65536.0,1,-nbitq), 
to_sfixed(3326.0/65536.0,1,-nbitq), 
to_sfixed(-1049.0/65536.0,1,-nbitq), 
to_sfixed(2424.0/65536.0,1,-nbitq), 
to_sfixed(-1032.0/65536.0,1,-nbitq), 
to_sfixed(-1104.0/65536.0,1,-nbitq), 
to_sfixed(899.0/65536.0,1,-nbitq), 
to_sfixed(-2381.0/65536.0,1,-nbitq), 
to_sfixed(-1766.0/65536.0,1,-nbitq), 
to_sfixed(922.0/65536.0,1,-nbitq), 
to_sfixed(777.0/65536.0,1,-nbitq), 
to_sfixed(-2338.0/65536.0,1,-nbitq), 
to_sfixed(-46.0/65536.0,1,-nbitq), 
to_sfixed(531.0/65536.0,1,-nbitq), 
to_sfixed(-1922.0/65536.0,1,-nbitq), 
to_sfixed(-2904.0/65536.0,1,-nbitq), 
to_sfixed(187.0/65536.0,1,-nbitq), 
to_sfixed(-1744.0/65536.0,1,-nbitq), 
to_sfixed(956.0/65536.0,1,-nbitq), 
to_sfixed(-3766.0/65536.0,1,-nbitq), 
to_sfixed(1022.0/65536.0,1,-nbitq), 
to_sfixed(-2610.0/65536.0,1,-nbitq), 
to_sfixed(-1005.0/65536.0,1,-nbitq), 
to_sfixed(2831.0/65536.0,1,-nbitq), 
to_sfixed(823.0/65536.0,1,-nbitq), 
to_sfixed(-3830.0/65536.0,1,-nbitq), 
to_sfixed(1100.0/65536.0,1,-nbitq), 
to_sfixed(-2292.0/65536.0,1,-nbitq), 
to_sfixed(-1419.0/65536.0,1,-nbitq), 
to_sfixed(-1236.0/65536.0,1,-nbitq), 
to_sfixed(-2153.0/65536.0,1,-nbitq), 
to_sfixed(-4341.0/65536.0,1,-nbitq), 
to_sfixed(-4725.0/65536.0,1,-nbitq), 
to_sfixed(1777.0/65536.0,1,-nbitq), 
to_sfixed(-571.0/65536.0,1,-nbitq), 
to_sfixed(100.0/65536.0,1,-nbitq), 
to_sfixed(-2119.0/65536.0,1,-nbitq), 
to_sfixed(-3184.0/65536.0,1,-nbitq), 
to_sfixed(471.0/65536.0,1,-nbitq), 
to_sfixed(1084.0/65536.0,1,-nbitq), 
to_sfixed(-525.0/65536.0,1,-nbitq), 
to_sfixed(19.0/65536.0,1,-nbitq), 
to_sfixed(1714.0/65536.0,1,-nbitq), 
to_sfixed(1595.0/65536.0,1,-nbitq), 
to_sfixed(433.0/65536.0,1,-nbitq), 
to_sfixed(-1196.0/65536.0,1,-nbitq), 
to_sfixed(1366.0/65536.0,1,-nbitq), 
to_sfixed(2101.0/65536.0,1,-nbitq), 
to_sfixed(1972.0/65536.0,1,-nbitq), 
to_sfixed(1714.0/65536.0,1,-nbitq), 
to_sfixed(-245.0/65536.0,1,-nbitq), 
to_sfixed(-2107.0/65536.0,1,-nbitq), 
to_sfixed(-3594.0/65536.0,1,-nbitq), 
to_sfixed(2272.0/65536.0,1,-nbitq), 
to_sfixed(2511.0/65536.0,1,-nbitq), 
to_sfixed(110.0/65536.0,1,-nbitq), 
to_sfixed(-231.0/65536.0,1,-nbitq), 
to_sfixed(1619.0/65536.0,1,-nbitq), 
to_sfixed(2332.0/65536.0,1,-nbitq), 
to_sfixed(-1339.0/65536.0,1,-nbitq), 
to_sfixed(-2159.0/65536.0,1,-nbitq), 
to_sfixed(510.0/65536.0,1,-nbitq), 
to_sfixed(-3131.0/65536.0,1,-nbitq), 
to_sfixed(1475.0/65536.0,1,-nbitq), 
to_sfixed(3712.0/65536.0,1,-nbitq), 
to_sfixed(1218.0/65536.0,1,-nbitq), 
to_sfixed(-3327.0/65536.0,1,-nbitq), 
to_sfixed(-1765.0/65536.0,1,-nbitq), 
to_sfixed(-817.0/65536.0,1,-nbitq), 
to_sfixed(3037.0/65536.0,1,-nbitq), 
to_sfixed(1650.0/65536.0,1,-nbitq), 
to_sfixed(1705.0/65536.0,1,-nbitq), 
to_sfixed(74.0/65536.0,1,-nbitq), 
to_sfixed(138.0/65536.0,1,-nbitq), 
to_sfixed(3950.0/65536.0,1,-nbitq), 
to_sfixed(759.0/65536.0,1,-nbitq), 
to_sfixed(1474.0/65536.0,1,-nbitq), 
to_sfixed(-3080.0/65536.0,1,-nbitq), 
to_sfixed(5055.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-635.0/65536.0,1,-nbitq), 
to_sfixed(332.0/65536.0,1,-nbitq), 
to_sfixed(2985.0/65536.0,1,-nbitq), 
to_sfixed(-3864.0/65536.0,1,-nbitq), 
to_sfixed(1304.0/65536.0,1,-nbitq), 
to_sfixed(-1198.0/65536.0,1,-nbitq), 
to_sfixed(2465.0/65536.0,1,-nbitq), 
to_sfixed(-2620.0/65536.0,1,-nbitq), 
to_sfixed(-1326.0/65536.0,1,-nbitq), 
to_sfixed(2945.0/65536.0,1,-nbitq), 
to_sfixed(681.0/65536.0,1,-nbitq), 
to_sfixed(455.0/65536.0,1,-nbitq), 
to_sfixed(1246.0/65536.0,1,-nbitq), 
to_sfixed(-2877.0/65536.0,1,-nbitq), 
to_sfixed(2757.0/65536.0,1,-nbitq), 
to_sfixed(2440.0/65536.0,1,-nbitq), 
to_sfixed(-2845.0/65536.0,1,-nbitq), 
to_sfixed(2824.0/65536.0,1,-nbitq), 
to_sfixed(-1078.0/65536.0,1,-nbitq), 
to_sfixed(2118.0/65536.0,1,-nbitq), 
to_sfixed(412.0/65536.0,1,-nbitq), 
to_sfixed(-2918.0/65536.0,1,-nbitq), 
to_sfixed(-557.0/65536.0,1,-nbitq), 
to_sfixed(-229.0/65536.0,1,-nbitq), 
to_sfixed(423.0/65536.0,1,-nbitq), 
to_sfixed(1936.0/65536.0,1,-nbitq), 
to_sfixed(-1126.0/65536.0,1,-nbitq), 
to_sfixed(-1241.0/65536.0,1,-nbitq), 
to_sfixed(-2517.0/65536.0,1,-nbitq), 
to_sfixed(-2223.0/65536.0,1,-nbitq), 
to_sfixed(-501.0/65536.0,1,-nbitq), 
to_sfixed(-1367.0/65536.0,1,-nbitq), 
to_sfixed(-5489.0/65536.0,1,-nbitq), 
to_sfixed(-4245.0/65536.0,1,-nbitq), 
to_sfixed(-1953.0/65536.0,1,-nbitq), 
to_sfixed(-2703.0/65536.0,1,-nbitq), 
to_sfixed(609.0/65536.0,1,-nbitq), 
to_sfixed(-2810.0/65536.0,1,-nbitq), 
to_sfixed(1302.0/65536.0,1,-nbitq), 
to_sfixed(-1746.0/65536.0,1,-nbitq), 
to_sfixed(-1575.0/65536.0,1,-nbitq), 
to_sfixed(-835.0/65536.0,1,-nbitq), 
to_sfixed(-1592.0/65536.0,1,-nbitq), 
to_sfixed(702.0/65536.0,1,-nbitq), 
to_sfixed(2785.0/65536.0,1,-nbitq), 
to_sfixed(-137.0/65536.0,1,-nbitq), 
to_sfixed(1180.0/65536.0,1,-nbitq), 
to_sfixed(3051.0/65536.0,1,-nbitq), 
to_sfixed(1450.0/65536.0,1,-nbitq), 
to_sfixed(2139.0/65536.0,1,-nbitq), 
to_sfixed(456.0/65536.0,1,-nbitq), 
to_sfixed(-529.0/65536.0,1,-nbitq), 
to_sfixed(2447.0/65536.0,1,-nbitq), 
to_sfixed(182.0/65536.0,1,-nbitq), 
to_sfixed(2353.0/65536.0,1,-nbitq), 
to_sfixed(2948.0/65536.0,1,-nbitq), 
to_sfixed(-1464.0/65536.0,1,-nbitq), 
to_sfixed(1881.0/65536.0,1,-nbitq), 
to_sfixed(-1990.0/65536.0,1,-nbitq), 
to_sfixed(2453.0/65536.0,1,-nbitq), 
to_sfixed(-2067.0/65536.0,1,-nbitq), 
to_sfixed(689.0/65536.0,1,-nbitq), 
to_sfixed(3086.0/65536.0,1,-nbitq), 
to_sfixed(632.0/65536.0,1,-nbitq), 
to_sfixed(-1526.0/65536.0,1,-nbitq), 
to_sfixed(784.0/65536.0,1,-nbitq), 
to_sfixed(-2380.0/65536.0,1,-nbitq), 
to_sfixed(-2078.0/65536.0,1,-nbitq), 
to_sfixed(-250.0/65536.0,1,-nbitq), 
to_sfixed(2781.0/65536.0,1,-nbitq), 
to_sfixed(-824.0/65536.0,1,-nbitq), 
to_sfixed(1175.0/65536.0,1,-nbitq), 
to_sfixed(2753.0/65536.0,1,-nbitq), 
to_sfixed(-2029.0/65536.0,1,-nbitq), 
to_sfixed(-872.0/65536.0,1,-nbitq), 
to_sfixed(-1462.0/65536.0,1,-nbitq), 
to_sfixed(-2345.0/65536.0,1,-nbitq), 
to_sfixed(3563.0/65536.0,1,-nbitq), 
to_sfixed(1089.0/65536.0,1,-nbitq), 
to_sfixed(1687.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3452.0/65536.0,1,-nbitq), 
to_sfixed(-1134.0/65536.0,1,-nbitq), 
to_sfixed(2150.0/65536.0,1,-nbitq), 
to_sfixed(-1257.0/65536.0,1,-nbitq), 
to_sfixed(-2175.0/65536.0,1,-nbitq), 
to_sfixed(667.0/65536.0,1,-nbitq), 
to_sfixed(-1977.0/65536.0,1,-nbitq), 
to_sfixed(-295.0/65536.0,1,-nbitq), 
to_sfixed(769.0/65536.0,1,-nbitq), 
to_sfixed(3000.0/65536.0,1,-nbitq), 
to_sfixed(1032.0/65536.0,1,-nbitq), 
to_sfixed(-610.0/65536.0,1,-nbitq), 
to_sfixed(-1922.0/65536.0,1,-nbitq), 
to_sfixed(-3234.0/65536.0,1,-nbitq), 
to_sfixed(580.0/65536.0,1,-nbitq), 
to_sfixed(-1431.0/65536.0,1,-nbitq), 
to_sfixed(-555.0/65536.0,1,-nbitq), 
to_sfixed(-1321.0/65536.0,1,-nbitq), 
to_sfixed(3319.0/65536.0,1,-nbitq), 
to_sfixed(296.0/65536.0,1,-nbitq), 
to_sfixed(-1477.0/65536.0,1,-nbitq), 
to_sfixed(-1700.0/65536.0,1,-nbitq), 
to_sfixed(2166.0/65536.0,1,-nbitq), 
to_sfixed(1503.0/65536.0,1,-nbitq), 
to_sfixed(500.0/65536.0,1,-nbitq), 
to_sfixed(1318.0/65536.0,1,-nbitq), 
to_sfixed(-1136.0/65536.0,1,-nbitq), 
to_sfixed(895.0/65536.0,1,-nbitq), 
to_sfixed(-3358.0/65536.0,1,-nbitq), 
to_sfixed(1041.0/65536.0,1,-nbitq), 
to_sfixed(-2201.0/65536.0,1,-nbitq), 
to_sfixed(364.0/65536.0,1,-nbitq), 
to_sfixed(-4053.0/65536.0,1,-nbitq), 
to_sfixed(-869.0/65536.0,1,-nbitq), 
to_sfixed(685.0/65536.0,1,-nbitq), 
to_sfixed(-1077.0/65536.0,1,-nbitq), 
to_sfixed(-2301.0/65536.0,1,-nbitq), 
to_sfixed(-2610.0/65536.0,1,-nbitq), 
to_sfixed(-1339.0/65536.0,1,-nbitq), 
to_sfixed(-757.0/65536.0,1,-nbitq), 
to_sfixed(-3737.0/65536.0,1,-nbitq), 
to_sfixed(-140.0/65536.0,1,-nbitq), 
to_sfixed(361.0/65536.0,1,-nbitq), 
to_sfixed(801.0/65536.0,1,-nbitq), 
to_sfixed(186.0/65536.0,1,-nbitq), 
to_sfixed(2126.0/65536.0,1,-nbitq), 
to_sfixed(3032.0/65536.0,1,-nbitq), 
to_sfixed(-2322.0/65536.0,1,-nbitq), 
to_sfixed(2375.0/65536.0,1,-nbitq), 
to_sfixed(989.0/65536.0,1,-nbitq), 
to_sfixed(1033.0/65536.0,1,-nbitq), 
to_sfixed(406.0/65536.0,1,-nbitq), 
to_sfixed(452.0/65536.0,1,-nbitq), 
to_sfixed(-1658.0/65536.0,1,-nbitq), 
to_sfixed(3498.0/65536.0,1,-nbitq), 
to_sfixed(-1584.0/65536.0,1,-nbitq), 
to_sfixed(-1614.0/65536.0,1,-nbitq), 
to_sfixed(2201.0/65536.0,1,-nbitq), 
to_sfixed(-2231.0/65536.0,1,-nbitq), 
to_sfixed(4449.0/65536.0,1,-nbitq), 
to_sfixed(-3910.0/65536.0,1,-nbitq), 
to_sfixed(-758.0/65536.0,1,-nbitq), 
to_sfixed(-1926.0/65536.0,1,-nbitq), 
to_sfixed(-353.0/65536.0,1,-nbitq), 
to_sfixed(-1434.0/65536.0,1,-nbitq), 
to_sfixed(330.0/65536.0,1,-nbitq), 
to_sfixed(2922.0/65536.0,1,-nbitq), 
to_sfixed(-2515.0/65536.0,1,-nbitq), 
to_sfixed(-994.0/65536.0,1,-nbitq), 
to_sfixed(2803.0/65536.0,1,-nbitq), 
to_sfixed(2810.0/65536.0,1,-nbitq), 
to_sfixed(-1554.0/65536.0,1,-nbitq), 
to_sfixed(-1505.0/65536.0,1,-nbitq), 
to_sfixed(-993.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(769.0/65536.0,1,-nbitq), 
to_sfixed(16.0/65536.0,1,-nbitq), 
to_sfixed(3415.0/65536.0,1,-nbitq), 
to_sfixed(-2247.0/65536.0,1,-nbitq), 
to_sfixed(3577.0/65536.0,1,-nbitq)  ), 
( to_sfixed(25.0/65536.0,1,-nbitq), 
to_sfixed(1888.0/65536.0,1,-nbitq), 
to_sfixed(2538.0/65536.0,1,-nbitq), 
to_sfixed(-6107.0/65536.0,1,-nbitq), 
to_sfixed(-533.0/65536.0,1,-nbitq), 
to_sfixed(-4010.0/65536.0,1,-nbitq), 
to_sfixed(-2855.0/65536.0,1,-nbitq), 
to_sfixed(1323.0/65536.0,1,-nbitq), 
to_sfixed(1660.0/65536.0,1,-nbitq), 
to_sfixed(-76.0/65536.0,1,-nbitq), 
to_sfixed(-2992.0/65536.0,1,-nbitq), 
to_sfixed(-804.0/65536.0,1,-nbitq), 
to_sfixed(64.0/65536.0,1,-nbitq), 
to_sfixed(-1747.0/65536.0,1,-nbitq), 
to_sfixed(-2864.0/65536.0,1,-nbitq), 
to_sfixed(1730.0/65536.0,1,-nbitq), 
to_sfixed(-1615.0/65536.0,1,-nbitq), 
to_sfixed(-1932.0/65536.0,1,-nbitq), 
to_sfixed(-82.0/65536.0,1,-nbitq), 
to_sfixed(-1182.0/65536.0,1,-nbitq), 
to_sfixed(-1063.0/65536.0,1,-nbitq), 
to_sfixed(3267.0/65536.0,1,-nbitq), 
to_sfixed(-587.0/65536.0,1,-nbitq), 
to_sfixed(3377.0/65536.0,1,-nbitq), 
to_sfixed(482.0/65536.0,1,-nbitq), 
to_sfixed(-1991.0/65536.0,1,-nbitq), 
to_sfixed(-1766.0/65536.0,1,-nbitq), 
to_sfixed(-944.0/65536.0,1,-nbitq), 
to_sfixed(-472.0/65536.0,1,-nbitq), 
to_sfixed(-1086.0/65536.0,1,-nbitq), 
to_sfixed(-2928.0/65536.0,1,-nbitq), 
to_sfixed(1396.0/65536.0,1,-nbitq), 
to_sfixed(-4650.0/65536.0,1,-nbitq), 
to_sfixed(-998.0/65536.0,1,-nbitq), 
to_sfixed(-870.0/65536.0,1,-nbitq), 
to_sfixed(-159.0/65536.0,1,-nbitq), 
to_sfixed(-2992.0/65536.0,1,-nbitq), 
to_sfixed(-2876.0/65536.0,1,-nbitq), 
to_sfixed(1110.0/65536.0,1,-nbitq), 
to_sfixed(3019.0/65536.0,1,-nbitq), 
to_sfixed(-997.0/65536.0,1,-nbitq), 
to_sfixed(-3203.0/65536.0,1,-nbitq), 
to_sfixed(-665.0/65536.0,1,-nbitq), 
to_sfixed(-1651.0/65536.0,1,-nbitq), 
to_sfixed(-1287.0/65536.0,1,-nbitq), 
to_sfixed(2106.0/65536.0,1,-nbitq), 
to_sfixed(806.0/65536.0,1,-nbitq), 
to_sfixed(-455.0/65536.0,1,-nbitq), 
to_sfixed(1017.0/65536.0,1,-nbitq), 
to_sfixed(4283.0/65536.0,1,-nbitq), 
to_sfixed(-2127.0/65536.0,1,-nbitq), 
to_sfixed(-2270.0/65536.0,1,-nbitq), 
to_sfixed(1839.0/65536.0,1,-nbitq), 
to_sfixed(52.0/65536.0,1,-nbitq), 
to_sfixed(-1083.0/65536.0,1,-nbitq), 
to_sfixed(671.0/65536.0,1,-nbitq), 
to_sfixed(-2220.0/65536.0,1,-nbitq), 
to_sfixed(3033.0/65536.0,1,-nbitq), 
to_sfixed(1682.0/65536.0,1,-nbitq), 
to_sfixed(1081.0/65536.0,1,-nbitq), 
to_sfixed(-751.0/65536.0,1,-nbitq), 
to_sfixed(2183.0/65536.0,1,-nbitq), 
to_sfixed(-788.0/65536.0,1,-nbitq), 
to_sfixed(21.0/65536.0,1,-nbitq), 
to_sfixed(1892.0/65536.0,1,-nbitq), 
to_sfixed(2504.0/65536.0,1,-nbitq), 
to_sfixed(2674.0/65536.0,1,-nbitq), 
to_sfixed(803.0/65536.0,1,-nbitq), 
to_sfixed(3327.0/65536.0,1,-nbitq), 
to_sfixed(3482.0/65536.0,1,-nbitq), 
to_sfixed(2932.0/65536.0,1,-nbitq), 
to_sfixed(-669.0/65536.0,1,-nbitq), 
to_sfixed(3699.0/65536.0,1,-nbitq), 
to_sfixed(-2446.0/65536.0,1,-nbitq), 
to_sfixed(1527.0/65536.0,1,-nbitq), 
to_sfixed(-2898.0/65536.0,1,-nbitq), 
to_sfixed(-2660.0/65536.0,1,-nbitq), 
to_sfixed(1138.0/65536.0,1,-nbitq), 
to_sfixed(-1768.0/65536.0,1,-nbitq), 
to_sfixed(1548.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1444.0/65536.0,1,-nbitq), 
to_sfixed(-3086.0/65536.0,1,-nbitq), 
to_sfixed(-1582.0/65536.0,1,-nbitq), 
to_sfixed(-987.0/65536.0,1,-nbitq), 
to_sfixed(-806.0/65536.0,1,-nbitq), 
to_sfixed(-432.0/65536.0,1,-nbitq), 
to_sfixed(2794.0/65536.0,1,-nbitq), 
to_sfixed(1154.0/65536.0,1,-nbitq), 
to_sfixed(-1841.0/65536.0,1,-nbitq), 
to_sfixed(2555.0/65536.0,1,-nbitq), 
to_sfixed(273.0/65536.0,1,-nbitq), 
to_sfixed(1291.0/65536.0,1,-nbitq), 
to_sfixed(-446.0/65536.0,1,-nbitq), 
to_sfixed(-2313.0/65536.0,1,-nbitq), 
to_sfixed(-4018.0/65536.0,1,-nbitq), 
to_sfixed(-1580.0/65536.0,1,-nbitq), 
to_sfixed(-290.0/65536.0,1,-nbitq), 
to_sfixed(-1065.0/65536.0,1,-nbitq), 
to_sfixed(-1.0/65536.0,1,-nbitq), 
to_sfixed(2336.0/65536.0,1,-nbitq), 
to_sfixed(-3742.0/65536.0,1,-nbitq), 
to_sfixed(-126.0/65536.0,1,-nbitq), 
to_sfixed(3980.0/65536.0,1,-nbitq), 
to_sfixed(749.0/65536.0,1,-nbitq), 
to_sfixed(-1545.0/65536.0,1,-nbitq), 
to_sfixed(412.0/65536.0,1,-nbitq), 
to_sfixed(-63.0/65536.0,1,-nbitq), 
to_sfixed(-2445.0/65536.0,1,-nbitq), 
to_sfixed(-1488.0/65536.0,1,-nbitq), 
to_sfixed(-1877.0/65536.0,1,-nbitq), 
to_sfixed(-612.0/65536.0,1,-nbitq), 
to_sfixed(-1514.0/65536.0,1,-nbitq), 
to_sfixed(-2450.0/65536.0,1,-nbitq), 
to_sfixed(767.0/65536.0,1,-nbitq), 
to_sfixed(-3030.0/65536.0,1,-nbitq), 
to_sfixed(-797.0/65536.0,1,-nbitq), 
to_sfixed(-1019.0/65536.0,1,-nbitq), 
to_sfixed(461.0/65536.0,1,-nbitq), 
to_sfixed(-882.0/65536.0,1,-nbitq), 
to_sfixed(-1510.0/65536.0,1,-nbitq), 
to_sfixed(-2477.0/65536.0,1,-nbitq), 
to_sfixed(-3075.0/65536.0,1,-nbitq), 
to_sfixed(-4081.0/65536.0,1,-nbitq), 
to_sfixed(-1086.0/65536.0,1,-nbitq), 
to_sfixed(1112.0/65536.0,1,-nbitq), 
to_sfixed(1182.0/65536.0,1,-nbitq), 
to_sfixed(-1658.0/65536.0,1,-nbitq), 
to_sfixed(1490.0/65536.0,1,-nbitq), 
to_sfixed(-2010.0/65536.0,1,-nbitq), 
to_sfixed(316.0/65536.0,1,-nbitq), 
to_sfixed(2157.0/65536.0,1,-nbitq), 
to_sfixed(2501.0/65536.0,1,-nbitq), 
to_sfixed(2043.0/65536.0,1,-nbitq), 
to_sfixed(275.0/65536.0,1,-nbitq), 
to_sfixed(3242.0/65536.0,1,-nbitq), 
to_sfixed(-1659.0/65536.0,1,-nbitq), 
to_sfixed(-1329.0/65536.0,1,-nbitq), 
to_sfixed(965.0/65536.0,1,-nbitq), 
to_sfixed(1127.0/65536.0,1,-nbitq), 
to_sfixed(1069.0/65536.0,1,-nbitq), 
to_sfixed(-3249.0/65536.0,1,-nbitq), 
to_sfixed(-107.0/65536.0,1,-nbitq), 
to_sfixed(2690.0/65536.0,1,-nbitq), 
to_sfixed(-2757.0/65536.0,1,-nbitq), 
to_sfixed(-1060.0/65536.0,1,-nbitq), 
to_sfixed(1269.0/65536.0,1,-nbitq), 
to_sfixed(-2590.0/65536.0,1,-nbitq), 
to_sfixed(99.0/65536.0,1,-nbitq), 
to_sfixed(-952.0/65536.0,1,-nbitq), 
to_sfixed(304.0/65536.0,1,-nbitq), 
to_sfixed(2287.0/65536.0,1,-nbitq), 
to_sfixed(3598.0/65536.0,1,-nbitq), 
to_sfixed(226.0/65536.0,1,-nbitq), 
to_sfixed(417.0/65536.0,1,-nbitq), 
to_sfixed(-1412.0/65536.0,1,-nbitq), 
to_sfixed(77.0/65536.0,1,-nbitq), 
to_sfixed(706.0/65536.0,1,-nbitq), 
to_sfixed(-1093.0/65536.0,1,-nbitq), 
to_sfixed(-234.0/65536.0,1,-nbitq), 
to_sfixed(2661.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1956.0/65536.0,1,-nbitq), 
to_sfixed(-2020.0/65536.0,1,-nbitq), 
to_sfixed(-5427.0/65536.0,1,-nbitq), 
to_sfixed(-4393.0/65536.0,1,-nbitq), 
to_sfixed(2581.0/65536.0,1,-nbitq), 
to_sfixed(-3479.0/65536.0,1,-nbitq), 
to_sfixed(3149.0/65536.0,1,-nbitq), 
to_sfixed(-3348.0/65536.0,1,-nbitq), 
to_sfixed(-1984.0/65536.0,1,-nbitq), 
to_sfixed(-2036.0/65536.0,1,-nbitq), 
to_sfixed(129.0/65536.0,1,-nbitq), 
to_sfixed(5448.0/65536.0,1,-nbitq), 
to_sfixed(1002.0/65536.0,1,-nbitq), 
to_sfixed(5072.0/65536.0,1,-nbitq), 
to_sfixed(-1511.0/65536.0,1,-nbitq), 
to_sfixed(-1502.0/65536.0,1,-nbitq), 
to_sfixed(-2150.0/65536.0,1,-nbitq), 
to_sfixed(-3388.0/65536.0,1,-nbitq), 
to_sfixed(-4893.0/65536.0,1,-nbitq), 
to_sfixed(1133.0/65536.0,1,-nbitq), 
to_sfixed(-1729.0/65536.0,1,-nbitq), 
to_sfixed(-1507.0/65536.0,1,-nbitq), 
to_sfixed(2481.0/65536.0,1,-nbitq), 
to_sfixed(-1316.0/65536.0,1,-nbitq), 
to_sfixed(-2845.0/65536.0,1,-nbitq), 
to_sfixed(-4303.0/65536.0,1,-nbitq), 
to_sfixed(-4539.0/65536.0,1,-nbitq), 
to_sfixed(-2401.0/65536.0,1,-nbitq), 
to_sfixed(-2300.0/65536.0,1,-nbitq), 
to_sfixed(1548.0/65536.0,1,-nbitq), 
to_sfixed(2506.0/65536.0,1,-nbitq), 
to_sfixed(-3979.0/65536.0,1,-nbitq), 
to_sfixed(-49.0/65536.0,1,-nbitq), 
to_sfixed(1851.0/65536.0,1,-nbitq), 
to_sfixed(-1173.0/65536.0,1,-nbitq), 
to_sfixed(339.0/65536.0,1,-nbitq), 
to_sfixed(-1443.0/65536.0,1,-nbitq), 
to_sfixed(-2927.0/65536.0,1,-nbitq), 
to_sfixed(5063.0/65536.0,1,-nbitq), 
to_sfixed(-220.0/65536.0,1,-nbitq), 
to_sfixed(-636.0/65536.0,1,-nbitq), 
to_sfixed(1649.0/65536.0,1,-nbitq), 
to_sfixed(-1203.0/65536.0,1,-nbitq), 
to_sfixed(2119.0/65536.0,1,-nbitq), 
to_sfixed(356.0/65536.0,1,-nbitq), 
to_sfixed(-1017.0/65536.0,1,-nbitq), 
to_sfixed(-3546.0/65536.0,1,-nbitq), 
to_sfixed(-617.0/65536.0,1,-nbitq), 
to_sfixed(401.0/65536.0,1,-nbitq), 
to_sfixed(3651.0/65536.0,1,-nbitq), 
to_sfixed(2947.0/65536.0,1,-nbitq), 
to_sfixed(-976.0/65536.0,1,-nbitq), 
to_sfixed(607.0/65536.0,1,-nbitq), 
to_sfixed(-1582.0/65536.0,1,-nbitq), 
to_sfixed(2802.0/65536.0,1,-nbitq), 
to_sfixed(854.0/65536.0,1,-nbitq), 
to_sfixed(-2190.0/65536.0,1,-nbitq), 
to_sfixed(-306.0/65536.0,1,-nbitq), 
to_sfixed(-2389.0/65536.0,1,-nbitq), 
to_sfixed(-564.0/65536.0,1,-nbitq), 
to_sfixed(-316.0/65536.0,1,-nbitq), 
to_sfixed(868.0/65536.0,1,-nbitq), 
to_sfixed(631.0/65536.0,1,-nbitq), 
to_sfixed(2059.0/65536.0,1,-nbitq), 
to_sfixed(2237.0/65536.0,1,-nbitq), 
to_sfixed(-3498.0/65536.0,1,-nbitq), 
to_sfixed(1721.0/65536.0,1,-nbitq), 
to_sfixed(-2934.0/65536.0,1,-nbitq), 
to_sfixed(-173.0/65536.0,1,-nbitq), 
to_sfixed(1132.0/65536.0,1,-nbitq), 
to_sfixed(-1888.0/65536.0,1,-nbitq), 
to_sfixed(627.0/65536.0,1,-nbitq), 
to_sfixed(-1376.0/65536.0,1,-nbitq), 
to_sfixed(-1571.0/65536.0,1,-nbitq), 
to_sfixed(-701.0/65536.0,1,-nbitq), 
to_sfixed(52.0/65536.0,1,-nbitq), 
to_sfixed(1213.0/65536.0,1,-nbitq), 
to_sfixed(-815.0/65536.0,1,-nbitq), 
to_sfixed(2443.0/65536.0,1,-nbitq), 
to_sfixed(2793.0/65536.0,1,-nbitq)  ), 
( to_sfixed(747.0/65536.0,1,-nbitq), 
to_sfixed(-2793.0/65536.0,1,-nbitq), 
to_sfixed(220.0/65536.0,1,-nbitq), 
to_sfixed(-1344.0/65536.0,1,-nbitq), 
to_sfixed(3804.0/65536.0,1,-nbitq), 
to_sfixed(-782.0/65536.0,1,-nbitq), 
to_sfixed(-503.0/65536.0,1,-nbitq), 
to_sfixed(-2026.0/65536.0,1,-nbitq), 
to_sfixed(-299.0/65536.0,1,-nbitq), 
to_sfixed(-2236.0/65536.0,1,-nbitq), 
to_sfixed(1536.0/65536.0,1,-nbitq), 
to_sfixed(7382.0/65536.0,1,-nbitq), 
to_sfixed(-725.0/65536.0,1,-nbitq), 
to_sfixed(6293.0/65536.0,1,-nbitq), 
to_sfixed(3234.0/65536.0,1,-nbitq), 
to_sfixed(1443.0/65536.0,1,-nbitq), 
to_sfixed(149.0/65536.0,1,-nbitq), 
to_sfixed(-2365.0/65536.0,1,-nbitq), 
to_sfixed(1731.0/65536.0,1,-nbitq), 
to_sfixed(-37.0/65536.0,1,-nbitq), 
to_sfixed(-4265.0/65536.0,1,-nbitq), 
to_sfixed(-2901.0/65536.0,1,-nbitq), 
to_sfixed(830.0/65536.0,1,-nbitq), 
to_sfixed(-3427.0/65536.0,1,-nbitq), 
to_sfixed(309.0/65536.0,1,-nbitq), 
to_sfixed(-1326.0/65536.0,1,-nbitq), 
to_sfixed(-46.0/65536.0,1,-nbitq), 
to_sfixed(-1766.0/65536.0,1,-nbitq), 
to_sfixed(-1812.0/65536.0,1,-nbitq), 
to_sfixed(-1362.0/65536.0,1,-nbitq), 
to_sfixed(-1580.0/65536.0,1,-nbitq), 
to_sfixed(-5088.0/65536.0,1,-nbitq), 
to_sfixed(-1715.0/65536.0,1,-nbitq), 
to_sfixed(5622.0/65536.0,1,-nbitq), 
to_sfixed(447.0/65536.0,1,-nbitq), 
to_sfixed(851.0/65536.0,1,-nbitq), 
to_sfixed(1526.0/65536.0,1,-nbitq), 
to_sfixed(1580.0/65536.0,1,-nbitq), 
to_sfixed(6363.0/65536.0,1,-nbitq), 
to_sfixed(-905.0/65536.0,1,-nbitq), 
to_sfixed(-206.0/65536.0,1,-nbitq), 
to_sfixed(-2647.0/65536.0,1,-nbitq), 
to_sfixed(2182.0/65536.0,1,-nbitq), 
to_sfixed(4200.0/65536.0,1,-nbitq), 
to_sfixed(1841.0/65536.0,1,-nbitq), 
to_sfixed(-772.0/65536.0,1,-nbitq), 
to_sfixed(-872.0/65536.0,1,-nbitq), 
to_sfixed(-1303.0/65536.0,1,-nbitq), 
to_sfixed(1128.0/65536.0,1,-nbitq), 
to_sfixed(4599.0/65536.0,1,-nbitq), 
to_sfixed(1735.0/65536.0,1,-nbitq), 
to_sfixed(-2944.0/65536.0,1,-nbitq), 
to_sfixed(-2662.0/65536.0,1,-nbitq), 
to_sfixed(-7047.0/65536.0,1,-nbitq), 
to_sfixed(1424.0/65536.0,1,-nbitq), 
to_sfixed(-262.0/65536.0,1,-nbitq), 
to_sfixed(3715.0/65536.0,1,-nbitq), 
to_sfixed(1666.0/65536.0,1,-nbitq), 
to_sfixed(-2386.0/65536.0,1,-nbitq), 
to_sfixed(-1372.0/65536.0,1,-nbitq), 
to_sfixed(1819.0/65536.0,1,-nbitq), 
to_sfixed(-1989.0/65536.0,1,-nbitq), 
to_sfixed(506.0/65536.0,1,-nbitq), 
to_sfixed(-2455.0/65536.0,1,-nbitq), 
to_sfixed(3794.0/65536.0,1,-nbitq), 
to_sfixed(-1940.0/65536.0,1,-nbitq), 
to_sfixed(-3567.0/65536.0,1,-nbitq), 
to_sfixed(3019.0/65536.0,1,-nbitq), 
to_sfixed(2397.0/65536.0,1,-nbitq), 
to_sfixed(1413.0/65536.0,1,-nbitq), 
to_sfixed(-1734.0/65536.0,1,-nbitq), 
to_sfixed(3334.0/65536.0,1,-nbitq), 
to_sfixed(256.0/65536.0,1,-nbitq), 
to_sfixed(-1483.0/65536.0,1,-nbitq), 
to_sfixed(633.0/65536.0,1,-nbitq), 
to_sfixed(-908.0/65536.0,1,-nbitq), 
to_sfixed(1925.0/65536.0,1,-nbitq), 
to_sfixed(134.0/65536.0,1,-nbitq), 
to_sfixed(-1053.0/65536.0,1,-nbitq), 
to_sfixed(-158.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-102.0/65536.0,1,-nbitq), 
to_sfixed(-2617.0/65536.0,1,-nbitq), 
to_sfixed(3390.0/65536.0,1,-nbitq), 
to_sfixed(-3535.0/65536.0,1,-nbitq), 
to_sfixed(-7079.0/65536.0,1,-nbitq), 
to_sfixed(-2566.0/65536.0,1,-nbitq), 
to_sfixed(4108.0/65536.0,1,-nbitq), 
to_sfixed(1274.0/65536.0,1,-nbitq), 
to_sfixed(4312.0/65536.0,1,-nbitq), 
to_sfixed(1461.0/65536.0,1,-nbitq), 
to_sfixed(1642.0/65536.0,1,-nbitq), 
to_sfixed(8033.0/65536.0,1,-nbitq), 
to_sfixed(1167.0/65536.0,1,-nbitq), 
to_sfixed(897.0/65536.0,1,-nbitq), 
to_sfixed(4354.0/65536.0,1,-nbitq), 
to_sfixed(-2902.0/65536.0,1,-nbitq), 
to_sfixed(-2490.0/65536.0,1,-nbitq), 
to_sfixed(194.0/65536.0,1,-nbitq), 
to_sfixed(-3608.0/65536.0,1,-nbitq), 
to_sfixed(1030.0/65536.0,1,-nbitq), 
to_sfixed(-1222.0/65536.0,1,-nbitq), 
to_sfixed(1395.0/65536.0,1,-nbitq), 
to_sfixed(-6.0/65536.0,1,-nbitq), 
to_sfixed(-1302.0/65536.0,1,-nbitq), 
to_sfixed(1541.0/65536.0,1,-nbitq), 
to_sfixed(-7280.0/65536.0,1,-nbitq), 
to_sfixed(1279.0/65536.0,1,-nbitq), 
to_sfixed(1362.0/65536.0,1,-nbitq), 
to_sfixed(415.0/65536.0,1,-nbitq), 
to_sfixed(-541.0/65536.0,1,-nbitq), 
to_sfixed(2299.0/65536.0,1,-nbitq), 
to_sfixed(-4898.0/65536.0,1,-nbitq), 
to_sfixed(747.0/65536.0,1,-nbitq), 
to_sfixed(4851.0/65536.0,1,-nbitq), 
to_sfixed(-2803.0/65536.0,1,-nbitq), 
to_sfixed(-932.0/65536.0,1,-nbitq), 
to_sfixed(1151.0/65536.0,1,-nbitq), 
to_sfixed(9306.0/65536.0,1,-nbitq), 
to_sfixed(6357.0/65536.0,1,-nbitq), 
to_sfixed(1566.0/65536.0,1,-nbitq), 
to_sfixed(-2194.0/65536.0,1,-nbitq), 
to_sfixed(-855.0/65536.0,1,-nbitq), 
to_sfixed(8090.0/65536.0,1,-nbitq), 
to_sfixed(4864.0/65536.0,1,-nbitq), 
to_sfixed(2905.0/65536.0,1,-nbitq), 
to_sfixed(-10153.0/65536.0,1,-nbitq), 
to_sfixed(-2441.0/65536.0,1,-nbitq), 
to_sfixed(3574.0/65536.0,1,-nbitq), 
to_sfixed(531.0/65536.0,1,-nbitq), 
to_sfixed(5176.0/65536.0,1,-nbitq), 
to_sfixed(2287.0/65536.0,1,-nbitq), 
to_sfixed(-8379.0/65536.0,1,-nbitq), 
to_sfixed(-1664.0/65536.0,1,-nbitq), 
to_sfixed(-7834.0/65536.0,1,-nbitq), 
to_sfixed(-1804.0/65536.0,1,-nbitq), 
to_sfixed(-951.0/65536.0,1,-nbitq), 
to_sfixed(-328.0/65536.0,1,-nbitq), 
to_sfixed(-1709.0/65536.0,1,-nbitq), 
to_sfixed(1443.0/65536.0,1,-nbitq), 
to_sfixed(-4760.0/65536.0,1,-nbitq), 
to_sfixed(-1526.0/65536.0,1,-nbitq), 
to_sfixed(-449.0/65536.0,1,-nbitq), 
to_sfixed(2396.0/65536.0,1,-nbitq), 
to_sfixed(-683.0/65536.0,1,-nbitq), 
to_sfixed(4913.0/65536.0,1,-nbitq), 
to_sfixed(-6528.0/65536.0,1,-nbitq), 
to_sfixed(1534.0/65536.0,1,-nbitq), 
to_sfixed(9164.0/65536.0,1,-nbitq), 
to_sfixed(5070.0/65536.0,1,-nbitq), 
to_sfixed(3374.0/65536.0,1,-nbitq), 
to_sfixed(996.0/65536.0,1,-nbitq), 
to_sfixed(6670.0/65536.0,1,-nbitq), 
to_sfixed(690.0/65536.0,1,-nbitq), 
to_sfixed(1552.0/65536.0,1,-nbitq), 
to_sfixed(1721.0/65536.0,1,-nbitq), 
to_sfixed(-2214.0/65536.0,1,-nbitq), 
to_sfixed(4699.0/65536.0,1,-nbitq), 
to_sfixed(1001.0/65536.0,1,-nbitq), 
to_sfixed(-2447.0/65536.0,1,-nbitq), 
to_sfixed(-3432.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1323.0/65536.0,1,-nbitq), 
to_sfixed(-3364.0/65536.0,1,-nbitq), 
to_sfixed(1378.0/65536.0,1,-nbitq), 
to_sfixed(-4756.0/65536.0,1,-nbitq), 
to_sfixed(-9122.0/65536.0,1,-nbitq), 
to_sfixed(-3087.0/65536.0,1,-nbitq), 
to_sfixed(4089.0/65536.0,1,-nbitq), 
to_sfixed(5000.0/65536.0,1,-nbitq), 
to_sfixed(-1622.0/65536.0,1,-nbitq), 
to_sfixed(-612.0/65536.0,1,-nbitq), 
to_sfixed(-4146.0/65536.0,1,-nbitq), 
to_sfixed(3030.0/65536.0,1,-nbitq), 
to_sfixed(227.0/65536.0,1,-nbitq), 
to_sfixed(2317.0/65536.0,1,-nbitq), 
to_sfixed(-428.0/65536.0,1,-nbitq), 
to_sfixed(2644.0/65536.0,1,-nbitq), 
to_sfixed(832.0/65536.0,1,-nbitq), 
to_sfixed(2905.0/65536.0,1,-nbitq), 
to_sfixed(1667.0/65536.0,1,-nbitq), 
to_sfixed(-207.0/65536.0,1,-nbitq), 
to_sfixed(-4721.0/65536.0,1,-nbitq), 
to_sfixed(1317.0/65536.0,1,-nbitq), 
to_sfixed(-1763.0/65536.0,1,-nbitq), 
to_sfixed(-4232.0/65536.0,1,-nbitq), 
to_sfixed(511.0/65536.0,1,-nbitq), 
to_sfixed(-9436.0/65536.0,1,-nbitq), 
to_sfixed(872.0/65536.0,1,-nbitq), 
to_sfixed(-2340.0/65536.0,1,-nbitq), 
to_sfixed(-3879.0/65536.0,1,-nbitq), 
to_sfixed(208.0/65536.0,1,-nbitq), 
to_sfixed(1281.0/65536.0,1,-nbitq), 
to_sfixed(-8670.0/65536.0,1,-nbitq), 
to_sfixed(1415.0/65536.0,1,-nbitq), 
to_sfixed(4081.0/65536.0,1,-nbitq), 
to_sfixed(-2931.0/65536.0,1,-nbitq), 
to_sfixed(2286.0/65536.0,1,-nbitq), 
to_sfixed(2908.0/65536.0,1,-nbitq), 
to_sfixed(6725.0/65536.0,1,-nbitq), 
to_sfixed(9507.0/65536.0,1,-nbitq), 
to_sfixed(-691.0/65536.0,1,-nbitq), 
to_sfixed(2164.0/65536.0,1,-nbitq), 
to_sfixed(543.0/65536.0,1,-nbitq), 
to_sfixed(3998.0/65536.0,1,-nbitq), 
to_sfixed(4824.0/65536.0,1,-nbitq), 
to_sfixed(390.0/65536.0,1,-nbitq), 
to_sfixed(-7178.0/65536.0,1,-nbitq), 
to_sfixed(1097.0/65536.0,1,-nbitq), 
to_sfixed(2716.0/65536.0,1,-nbitq), 
to_sfixed(1119.0/65536.0,1,-nbitq), 
to_sfixed(1290.0/65536.0,1,-nbitq), 
to_sfixed(-2034.0/65536.0,1,-nbitq), 
to_sfixed(-8588.0/65536.0,1,-nbitq), 
to_sfixed(491.0/65536.0,1,-nbitq), 
to_sfixed(-5450.0/65536.0,1,-nbitq), 
to_sfixed(-2418.0/65536.0,1,-nbitq), 
to_sfixed(-4322.0/65536.0,1,-nbitq), 
to_sfixed(3230.0/65536.0,1,-nbitq), 
to_sfixed(-4224.0/65536.0,1,-nbitq), 
to_sfixed(1619.0/65536.0,1,-nbitq), 
to_sfixed(-6445.0/65536.0,1,-nbitq), 
to_sfixed(-131.0/65536.0,1,-nbitq), 
to_sfixed(1338.0/65536.0,1,-nbitq), 
to_sfixed(559.0/65536.0,1,-nbitq), 
to_sfixed(-1922.0/65536.0,1,-nbitq), 
to_sfixed(3941.0/65536.0,1,-nbitq), 
to_sfixed(-5540.0/65536.0,1,-nbitq), 
to_sfixed(3476.0/65536.0,1,-nbitq), 
to_sfixed(10948.0/65536.0,1,-nbitq), 
to_sfixed(2562.0/65536.0,1,-nbitq), 
to_sfixed(5301.0/65536.0,1,-nbitq), 
to_sfixed(-610.0/65536.0,1,-nbitq), 
to_sfixed(8821.0/65536.0,1,-nbitq), 
to_sfixed(-4556.0/65536.0,1,-nbitq), 
to_sfixed(-166.0/65536.0,1,-nbitq), 
to_sfixed(-1809.0/65536.0,1,-nbitq), 
to_sfixed(-2286.0/65536.0,1,-nbitq), 
to_sfixed(10067.0/65536.0,1,-nbitq), 
to_sfixed(-2432.0/65536.0,1,-nbitq), 
to_sfixed(-1852.0/65536.0,1,-nbitq), 
to_sfixed(-1595.0/65536.0,1,-nbitq)  ), 
( to_sfixed(151.0/65536.0,1,-nbitq), 
to_sfixed(-1122.0/65536.0,1,-nbitq), 
to_sfixed(-4360.0/65536.0,1,-nbitq), 
to_sfixed(-593.0/65536.0,1,-nbitq), 
to_sfixed(-9186.0/65536.0,1,-nbitq), 
to_sfixed(-270.0/65536.0,1,-nbitq), 
to_sfixed(-716.0/65536.0,1,-nbitq), 
to_sfixed(2392.0/65536.0,1,-nbitq), 
to_sfixed(-1064.0/65536.0,1,-nbitq), 
to_sfixed(-1964.0/65536.0,1,-nbitq), 
to_sfixed(71.0/65536.0,1,-nbitq), 
to_sfixed(-5347.0/65536.0,1,-nbitq), 
to_sfixed(-1673.0/65536.0,1,-nbitq), 
to_sfixed(1531.0/65536.0,1,-nbitq), 
to_sfixed(1869.0/65536.0,1,-nbitq), 
to_sfixed(-1976.0/65536.0,1,-nbitq), 
to_sfixed(1675.0/65536.0,1,-nbitq), 
to_sfixed(1020.0/65536.0,1,-nbitq), 
to_sfixed(1343.0/65536.0,1,-nbitq), 
to_sfixed(41.0/65536.0,1,-nbitq), 
to_sfixed(-10361.0/65536.0,1,-nbitq), 
to_sfixed(-1711.0/65536.0,1,-nbitq), 
to_sfixed(4603.0/65536.0,1,-nbitq), 
to_sfixed(-7935.0/65536.0,1,-nbitq), 
to_sfixed(-2303.0/65536.0,1,-nbitq), 
to_sfixed(-9716.0/65536.0,1,-nbitq), 
to_sfixed(2781.0/65536.0,1,-nbitq), 
to_sfixed(1767.0/65536.0,1,-nbitq), 
to_sfixed(-5901.0/65536.0,1,-nbitq), 
to_sfixed(-2258.0/65536.0,1,-nbitq), 
to_sfixed(4678.0/65536.0,1,-nbitq), 
to_sfixed(-6871.0/65536.0,1,-nbitq), 
to_sfixed(373.0/65536.0,1,-nbitq), 
to_sfixed(-839.0/65536.0,1,-nbitq), 
to_sfixed(2596.0/65536.0,1,-nbitq), 
to_sfixed(2694.0/65536.0,1,-nbitq), 
to_sfixed(5927.0/65536.0,1,-nbitq), 
to_sfixed(12367.0/65536.0,1,-nbitq), 
to_sfixed(13279.0/65536.0,1,-nbitq), 
to_sfixed(1973.0/65536.0,1,-nbitq), 
to_sfixed(4459.0/65536.0,1,-nbitq), 
to_sfixed(1010.0/65536.0,1,-nbitq), 
to_sfixed(2010.0/65536.0,1,-nbitq), 
to_sfixed(1786.0/65536.0,1,-nbitq), 
to_sfixed(144.0/65536.0,1,-nbitq), 
to_sfixed(-6632.0/65536.0,1,-nbitq), 
to_sfixed(-1250.0/65536.0,1,-nbitq), 
to_sfixed(-5297.0/65536.0,1,-nbitq), 
to_sfixed(494.0/65536.0,1,-nbitq), 
to_sfixed(3646.0/65536.0,1,-nbitq), 
to_sfixed(2904.0/65536.0,1,-nbitq), 
to_sfixed(-4273.0/65536.0,1,-nbitq), 
to_sfixed(3525.0/65536.0,1,-nbitq), 
to_sfixed(-4935.0/65536.0,1,-nbitq), 
to_sfixed(457.0/65536.0,1,-nbitq), 
to_sfixed(-4029.0/65536.0,1,-nbitq), 
to_sfixed(1091.0/65536.0,1,-nbitq), 
to_sfixed(-3872.0/65536.0,1,-nbitq), 
to_sfixed(3504.0/65536.0,1,-nbitq), 
to_sfixed(-10285.0/65536.0,1,-nbitq), 
to_sfixed(1338.0/65536.0,1,-nbitq), 
to_sfixed(608.0/65536.0,1,-nbitq), 
to_sfixed(1413.0/65536.0,1,-nbitq), 
to_sfixed(-412.0/65536.0,1,-nbitq), 
to_sfixed(7748.0/65536.0,1,-nbitq), 
to_sfixed(-4696.0/65536.0,1,-nbitq), 
to_sfixed(5183.0/65536.0,1,-nbitq), 
to_sfixed(11546.0/65536.0,1,-nbitq), 
to_sfixed(3301.0/65536.0,1,-nbitq), 
to_sfixed(9426.0/65536.0,1,-nbitq), 
to_sfixed(-4251.0/65536.0,1,-nbitq), 
to_sfixed(3461.0/65536.0,1,-nbitq), 
to_sfixed(-3067.0/65536.0,1,-nbitq), 
to_sfixed(-1786.0/65536.0,1,-nbitq), 
to_sfixed(1251.0/65536.0,1,-nbitq), 
to_sfixed(-2869.0/65536.0,1,-nbitq), 
to_sfixed(3227.0/65536.0,1,-nbitq), 
to_sfixed(-4935.0/65536.0,1,-nbitq), 
to_sfixed(-2813.0/65536.0,1,-nbitq), 
to_sfixed(-3342.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1510.0/65536.0,1,-nbitq), 
to_sfixed(2081.0/65536.0,1,-nbitq), 
to_sfixed(-11443.0/65536.0,1,-nbitq), 
to_sfixed(-5758.0/65536.0,1,-nbitq), 
to_sfixed(-426.0/65536.0,1,-nbitq), 
to_sfixed(-2303.0/65536.0,1,-nbitq), 
to_sfixed(2016.0/65536.0,1,-nbitq), 
to_sfixed(-1294.0/65536.0,1,-nbitq), 
to_sfixed(2069.0/65536.0,1,-nbitq), 
to_sfixed(1551.0/65536.0,1,-nbitq), 
to_sfixed(896.0/65536.0,1,-nbitq), 
to_sfixed(-4862.0/65536.0,1,-nbitq), 
to_sfixed(2261.0/65536.0,1,-nbitq), 
to_sfixed(-3343.0/65536.0,1,-nbitq), 
to_sfixed(793.0/65536.0,1,-nbitq), 
to_sfixed(-756.0/65536.0,1,-nbitq), 
to_sfixed(1339.0/65536.0,1,-nbitq), 
to_sfixed(4116.0/65536.0,1,-nbitq), 
to_sfixed(1663.0/65536.0,1,-nbitq), 
to_sfixed(-895.0/65536.0,1,-nbitq), 
to_sfixed(-3899.0/65536.0,1,-nbitq), 
to_sfixed(2877.0/65536.0,1,-nbitq), 
to_sfixed(5564.0/65536.0,1,-nbitq), 
to_sfixed(-403.0/65536.0,1,-nbitq), 
to_sfixed(-266.0/65536.0,1,-nbitq), 
to_sfixed(-5676.0/65536.0,1,-nbitq), 
to_sfixed(1373.0/65536.0,1,-nbitq), 
to_sfixed(1687.0/65536.0,1,-nbitq), 
to_sfixed(-8781.0/65536.0,1,-nbitq), 
to_sfixed(-2086.0/65536.0,1,-nbitq), 
to_sfixed(4228.0/65536.0,1,-nbitq), 
to_sfixed(-4481.0/65536.0,1,-nbitq), 
to_sfixed(4071.0/65536.0,1,-nbitq), 
to_sfixed(-493.0/65536.0,1,-nbitq), 
to_sfixed(2272.0/65536.0,1,-nbitq), 
to_sfixed(-1596.0/65536.0,1,-nbitq), 
to_sfixed(5171.0/65536.0,1,-nbitq), 
to_sfixed(4172.0/65536.0,1,-nbitq), 
to_sfixed(9239.0/65536.0,1,-nbitq), 
to_sfixed(2001.0/65536.0,1,-nbitq), 
to_sfixed(1149.0/65536.0,1,-nbitq), 
to_sfixed(538.0/65536.0,1,-nbitq), 
to_sfixed(3359.0/65536.0,1,-nbitq), 
to_sfixed(-584.0/65536.0,1,-nbitq), 
to_sfixed(-1963.0/65536.0,1,-nbitq), 
to_sfixed(-3894.0/65536.0,1,-nbitq), 
to_sfixed(1738.0/65536.0,1,-nbitq), 
to_sfixed(-2296.0/65536.0,1,-nbitq), 
to_sfixed(1153.0/65536.0,1,-nbitq), 
to_sfixed(4160.0/65536.0,1,-nbitq), 
to_sfixed(-1687.0/65536.0,1,-nbitq), 
to_sfixed(-2254.0/65536.0,1,-nbitq), 
to_sfixed(-3480.0/65536.0,1,-nbitq), 
to_sfixed(-7801.0/65536.0,1,-nbitq), 
to_sfixed(-1503.0/65536.0,1,-nbitq), 
to_sfixed(-3021.0/65536.0,1,-nbitq), 
to_sfixed(910.0/65536.0,1,-nbitq), 
to_sfixed(-2286.0/65536.0,1,-nbitq), 
to_sfixed(-1976.0/65536.0,1,-nbitq), 
to_sfixed(-14444.0/65536.0,1,-nbitq), 
to_sfixed(287.0/65536.0,1,-nbitq), 
to_sfixed(883.0/65536.0,1,-nbitq), 
to_sfixed(-2104.0/65536.0,1,-nbitq), 
to_sfixed(325.0/65536.0,1,-nbitq), 
to_sfixed(7012.0/65536.0,1,-nbitq), 
to_sfixed(-7974.0/65536.0,1,-nbitq), 
to_sfixed(-496.0/65536.0,1,-nbitq), 
to_sfixed(11327.0/65536.0,1,-nbitq), 
to_sfixed(-1269.0/65536.0,1,-nbitq), 
to_sfixed(11130.0/65536.0,1,-nbitq), 
to_sfixed(-3100.0/65536.0,1,-nbitq), 
to_sfixed(1022.0/65536.0,1,-nbitq), 
to_sfixed(-5887.0/65536.0,1,-nbitq), 
to_sfixed(523.0/65536.0,1,-nbitq), 
to_sfixed(-343.0/65536.0,1,-nbitq), 
to_sfixed(4283.0/65536.0,1,-nbitq), 
to_sfixed(5485.0/65536.0,1,-nbitq), 
to_sfixed(-4724.0/65536.0,1,-nbitq), 
to_sfixed(518.0/65536.0,1,-nbitq), 
to_sfixed(-2955.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-360.0/65536.0,1,-nbitq), 
to_sfixed(1497.0/65536.0,1,-nbitq), 
to_sfixed(-13723.0/65536.0,1,-nbitq), 
to_sfixed(-6693.0/65536.0,1,-nbitq), 
to_sfixed(-2929.0/65536.0,1,-nbitq), 
to_sfixed(-2603.0/65536.0,1,-nbitq), 
to_sfixed(2600.0/65536.0,1,-nbitq), 
to_sfixed(-4109.0/65536.0,1,-nbitq), 
to_sfixed(5951.0/65536.0,1,-nbitq), 
to_sfixed(3027.0/65536.0,1,-nbitq), 
to_sfixed(4273.0/65536.0,1,-nbitq), 
to_sfixed(-9071.0/65536.0,1,-nbitq), 
to_sfixed(1225.0/65536.0,1,-nbitq), 
to_sfixed(-1209.0/65536.0,1,-nbitq), 
to_sfixed(2369.0/65536.0,1,-nbitq), 
to_sfixed(-2307.0/65536.0,1,-nbitq), 
to_sfixed(346.0/65536.0,1,-nbitq), 
to_sfixed(1628.0/65536.0,1,-nbitq), 
to_sfixed(7280.0/65536.0,1,-nbitq), 
to_sfixed(-2062.0/65536.0,1,-nbitq), 
to_sfixed(-8751.0/65536.0,1,-nbitq), 
to_sfixed(6103.0/65536.0,1,-nbitq), 
to_sfixed(12123.0/65536.0,1,-nbitq), 
to_sfixed(2713.0/65536.0,1,-nbitq), 
to_sfixed(-1469.0/65536.0,1,-nbitq), 
to_sfixed(-6938.0/65536.0,1,-nbitq), 
to_sfixed(3546.0/65536.0,1,-nbitq), 
to_sfixed(156.0/65536.0,1,-nbitq), 
to_sfixed(-1558.0/65536.0,1,-nbitq), 
to_sfixed(-2219.0/65536.0,1,-nbitq), 
to_sfixed(2607.0/65536.0,1,-nbitq), 
to_sfixed(-4532.0/65536.0,1,-nbitq), 
to_sfixed(3473.0/65536.0,1,-nbitq), 
to_sfixed(-1881.0/65536.0,1,-nbitq), 
to_sfixed(-94.0/65536.0,1,-nbitq), 
to_sfixed(-1458.0/65536.0,1,-nbitq), 
to_sfixed(11530.0/65536.0,1,-nbitq), 
to_sfixed(1801.0/65536.0,1,-nbitq), 
to_sfixed(7923.0/65536.0,1,-nbitq), 
to_sfixed(1212.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(-2500.0/65536.0,1,-nbitq), 
to_sfixed(1292.0/65536.0,1,-nbitq), 
to_sfixed(1761.0/65536.0,1,-nbitq), 
to_sfixed(2608.0/65536.0,1,-nbitq), 
to_sfixed(-1555.0/65536.0,1,-nbitq), 
to_sfixed(263.0/65536.0,1,-nbitq), 
to_sfixed(4984.0/65536.0,1,-nbitq), 
to_sfixed(2167.0/65536.0,1,-nbitq), 
to_sfixed(-204.0/65536.0,1,-nbitq), 
to_sfixed(-2432.0/65536.0,1,-nbitq), 
to_sfixed(-4483.0/65536.0,1,-nbitq), 
to_sfixed(-6747.0/65536.0,1,-nbitq), 
to_sfixed(-8587.0/65536.0,1,-nbitq), 
to_sfixed(-1301.0/65536.0,1,-nbitq), 
to_sfixed(-5054.0/65536.0,1,-nbitq), 
to_sfixed(2954.0/65536.0,1,-nbitq), 
to_sfixed(95.0/65536.0,1,-nbitq), 
to_sfixed(-567.0/65536.0,1,-nbitq), 
to_sfixed(-14814.0/65536.0,1,-nbitq), 
to_sfixed(4486.0/65536.0,1,-nbitq), 
to_sfixed(-252.0/65536.0,1,-nbitq), 
to_sfixed(2166.0/65536.0,1,-nbitq), 
to_sfixed(-3048.0/65536.0,1,-nbitq), 
to_sfixed(5092.0/65536.0,1,-nbitq), 
to_sfixed(-4317.0/65536.0,1,-nbitq), 
to_sfixed(1832.0/65536.0,1,-nbitq), 
to_sfixed(14992.0/65536.0,1,-nbitq), 
to_sfixed(-73.0/65536.0,1,-nbitq), 
to_sfixed(9153.0/65536.0,1,-nbitq), 
to_sfixed(-414.0/65536.0,1,-nbitq), 
to_sfixed(-3140.0/65536.0,1,-nbitq), 
to_sfixed(-5388.0/65536.0,1,-nbitq), 
to_sfixed(1558.0/65536.0,1,-nbitq), 
to_sfixed(-1556.0/65536.0,1,-nbitq), 
to_sfixed(4857.0/65536.0,1,-nbitq), 
to_sfixed(8378.0/65536.0,1,-nbitq), 
to_sfixed(3788.0/65536.0,1,-nbitq), 
to_sfixed(-2109.0/65536.0,1,-nbitq), 
to_sfixed(-2110.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1541.0/65536.0,1,-nbitq), 
to_sfixed(6549.0/65536.0,1,-nbitq), 
to_sfixed(-17018.0/65536.0,1,-nbitq), 
to_sfixed(-11747.0/65536.0,1,-nbitq), 
to_sfixed(-4018.0/65536.0,1,-nbitq), 
to_sfixed(-193.0/65536.0,1,-nbitq), 
to_sfixed(-1951.0/65536.0,1,-nbitq), 
to_sfixed(-2763.0/65536.0,1,-nbitq), 
to_sfixed(5971.0/65536.0,1,-nbitq), 
to_sfixed(2989.0/65536.0,1,-nbitq), 
to_sfixed(5771.0/65536.0,1,-nbitq), 
to_sfixed(-11018.0/65536.0,1,-nbitq), 
to_sfixed(-944.0/65536.0,1,-nbitq), 
to_sfixed(-6125.0/65536.0,1,-nbitq), 
to_sfixed(4048.0/65536.0,1,-nbitq), 
to_sfixed(1273.0/65536.0,1,-nbitq), 
to_sfixed(-1314.0/65536.0,1,-nbitq), 
to_sfixed(-96.0/65536.0,1,-nbitq), 
to_sfixed(5123.0/65536.0,1,-nbitq), 
to_sfixed(-303.0/65536.0,1,-nbitq), 
to_sfixed(-4910.0/65536.0,1,-nbitq), 
to_sfixed(6590.0/65536.0,1,-nbitq), 
to_sfixed(11506.0/65536.0,1,-nbitq), 
to_sfixed(10303.0/65536.0,1,-nbitq), 
to_sfixed(-5541.0/65536.0,1,-nbitq), 
to_sfixed(-5020.0/65536.0,1,-nbitq), 
to_sfixed(1307.0/65536.0,1,-nbitq), 
to_sfixed(1436.0/65536.0,1,-nbitq), 
to_sfixed(3185.0/65536.0,1,-nbitq), 
to_sfixed(-2284.0/65536.0,1,-nbitq), 
to_sfixed(4372.0/65536.0,1,-nbitq), 
to_sfixed(-13290.0/65536.0,1,-nbitq), 
to_sfixed(2237.0/65536.0,1,-nbitq), 
to_sfixed(-790.0/65536.0,1,-nbitq), 
to_sfixed(-1434.0/65536.0,1,-nbitq), 
to_sfixed(-2390.0/65536.0,1,-nbitq), 
to_sfixed(10978.0/65536.0,1,-nbitq), 
to_sfixed(-3454.0/65536.0,1,-nbitq), 
to_sfixed(6955.0/65536.0,1,-nbitq), 
to_sfixed(-2145.0/65536.0,1,-nbitq), 
to_sfixed(-3451.0/65536.0,1,-nbitq), 
to_sfixed(-2822.0/65536.0,1,-nbitq), 
to_sfixed(-409.0/65536.0,1,-nbitq), 
to_sfixed(2506.0/65536.0,1,-nbitq), 
to_sfixed(1055.0/65536.0,1,-nbitq), 
to_sfixed(-5474.0/65536.0,1,-nbitq), 
to_sfixed(2285.0/65536.0,1,-nbitq), 
to_sfixed(2630.0/65536.0,1,-nbitq), 
to_sfixed(2946.0/65536.0,1,-nbitq), 
to_sfixed(1690.0/65536.0,1,-nbitq), 
to_sfixed(-2719.0/65536.0,1,-nbitq), 
to_sfixed(-4548.0/65536.0,1,-nbitq), 
to_sfixed(-9263.0/65536.0,1,-nbitq), 
to_sfixed(-10056.0/65536.0,1,-nbitq), 
to_sfixed(-3524.0/65536.0,1,-nbitq), 
to_sfixed(-4746.0/65536.0,1,-nbitq), 
to_sfixed(1136.0/65536.0,1,-nbitq), 
to_sfixed(-1384.0/65536.0,1,-nbitq), 
to_sfixed(2369.0/65536.0,1,-nbitq), 
to_sfixed(-12773.0/65536.0,1,-nbitq), 
to_sfixed(820.0/65536.0,1,-nbitq), 
to_sfixed(-1469.0/65536.0,1,-nbitq), 
to_sfixed(-1772.0/65536.0,1,-nbitq), 
to_sfixed(-1095.0/65536.0,1,-nbitq), 
to_sfixed(1648.0/65536.0,1,-nbitq), 
to_sfixed(-1159.0/65536.0,1,-nbitq), 
to_sfixed(4094.0/65536.0,1,-nbitq), 
to_sfixed(12175.0/65536.0,1,-nbitq), 
to_sfixed(686.0/65536.0,1,-nbitq), 
to_sfixed(9937.0/65536.0,1,-nbitq), 
to_sfixed(-396.0/65536.0,1,-nbitq), 
to_sfixed(-3342.0/65536.0,1,-nbitq), 
to_sfixed(-7265.0/65536.0,1,-nbitq), 
to_sfixed(-921.0/65536.0,1,-nbitq), 
to_sfixed(435.0/65536.0,1,-nbitq), 
to_sfixed(-607.0/65536.0,1,-nbitq), 
to_sfixed(3258.0/65536.0,1,-nbitq), 
to_sfixed(4427.0/65536.0,1,-nbitq), 
to_sfixed(-3150.0/65536.0,1,-nbitq), 
to_sfixed(-2654.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3452.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(-9757.0/65536.0,1,-nbitq), 
to_sfixed(-7752.0/65536.0,1,-nbitq), 
to_sfixed(-1681.0/65536.0,1,-nbitq), 
to_sfixed(4692.0/65536.0,1,-nbitq), 
to_sfixed(-499.0/65536.0,1,-nbitq), 
to_sfixed(-3875.0/65536.0,1,-nbitq), 
to_sfixed(4261.0/65536.0,1,-nbitq), 
to_sfixed(2879.0/65536.0,1,-nbitq), 
to_sfixed(5557.0/65536.0,1,-nbitq), 
to_sfixed(-12138.0/65536.0,1,-nbitq), 
to_sfixed(-4614.0/65536.0,1,-nbitq), 
to_sfixed(1116.0/65536.0,1,-nbitq), 
to_sfixed(1126.0/65536.0,1,-nbitq), 
to_sfixed(1730.0/65536.0,1,-nbitq), 
to_sfixed(-1850.0/65536.0,1,-nbitq), 
to_sfixed(-1946.0/65536.0,1,-nbitq), 
to_sfixed(4640.0/65536.0,1,-nbitq), 
to_sfixed(-2205.0/65536.0,1,-nbitq), 
to_sfixed(-10383.0/65536.0,1,-nbitq), 
to_sfixed(8067.0/65536.0,1,-nbitq), 
to_sfixed(7463.0/65536.0,1,-nbitq), 
to_sfixed(11342.0/65536.0,1,-nbitq), 
to_sfixed(-2312.0/65536.0,1,-nbitq), 
to_sfixed(-1548.0/65536.0,1,-nbitq), 
to_sfixed(480.0/65536.0,1,-nbitq), 
to_sfixed(-616.0/65536.0,1,-nbitq), 
to_sfixed(1055.0/65536.0,1,-nbitq), 
to_sfixed(1450.0/65536.0,1,-nbitq), 
to_sfixed(6698.0/65536.0,1,-nbitq), 
to_sfixed(-10798.0/65536.0,1,-nbitq), 
to_sfixed(61.0/65536.0,1,-nbitq), 
to_sfixed(-396.0/65536.0,1,-nbitq), 
to_sfixed(-2865.0/65536.0,1,-nbitq), 
to_sfixed(2491.0/65536.0,1,-nbitq), 
to_sfixed(4211.0/65536.0,1,-nbitq), 
to_sfixed(3453.0/65536.0,1,-nbitq), 
to_sfixed(4481.0/65536.0,1,-nbitq), 
to_sfixed(-2967.0/65536.0,1,-nbitq), 
to_sfixed(-4114.0/65536.0,1,-nbitq), 
to_sfixed(-2793.0/65536.0,1,-nbitq), 
to_sfixed(-2660.0/65536.0,1,-nbitq), 
to_sfixed(1679.0/65536.0,1,-nbitq), 
to_sfixed(-2464.0/65536.0,1,-nbitq), 
to_sfixed(-2630.0/65536.0,1,-nbitq), 
to_sfixed(-599.0/65536.0,1,-nbitq), 
to_sfixed(2694.0/65536.0,1,-nbitq), 
to_sfixed(2570.0/65536.0,1,-nbitq), 
to_sfixed(145.0/65536.0,1,-nbitq), 
to_sfixed(-460.0/65536.0,1,-nbitq), 
to_sfixed(-6161.0/65536.0,1,-nbitq), 
to_sfixed(-7149.0/65536.0,1,-nbitq), 
to_sfixed(-2175.0/65536.0,1,-nbitq), 
to_sfixed(-2471.0/65536.0,1,-nbitq), 
to_sfixed(-8174.0/65536.0,1,-nbitq), 
to_sfixed(1921.0/65536.0,1,-nbitq), 
to_sfixed(-4383.0/65536.0,1,-nbitq), 
to_sfixed(-1624.0/65536.0,1,-nbitq), 
to_sfixed(-7523.0/65536.0,1,-nbitq), 
to_sfixed(5286.0/65536.0,1,-nbitq), 
to_sfixed(-249.0/65536.0,1,-nbitq), 
to_sfixed(-623.0/65536.0,1,-nbitq), 
to_sfixed(2265.0/65536.0,1,-nbitq), 
to_sfixed(3592.0/65536.0,1,-nbitq), 
to_sfixed(-3306.0/65536.0,1,-nbitq), 
to_sfixed(-108.0/65536.0,1,-nbitq), 
to_sfixed(8323.0/65536.0,1,-nbitq), 
to_sfixed(-1728.0/65536.0,1,-nbitq), 
to_sfixed(3925.0/65536.0,1,-nbitq), 
to_sfixed(-1643.0/65536.0,1,-nbitq), 
to_sfixed(1647.0/65536.0,1,-nbitq), 
to_sfixed(-4560.0/65536.0,1,-nbitq), 
to_sfixed(425.0/65536.0,1,-nbitq), 
to_sfixed(1060.0/65536.0,1,-nbitq), 
to_sfixed(1680.0/65536.0,1,-nbitq), 
to_sfixed(6208.0/65536.0,1,-nbitq), 
to_sfixed(966.0/65536.0,1,-nbitq), 
to_sfixed(-1810.0/65536.0,1,-nbitq), 
to_sfixed(-1219.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4825.0/65536.0,1,-nbitq), 
to_sfixed(3087.0/65536.0,1,-nbitq), 
to_sfixed(-6101.0/65536.0,1,-nbitq), 
to_sfixed(-5307.0/65536.0,1,-nbitq), 
to_sfixed(-1573.0/65536.0,1,-nbitq), 
to_sfixed(-727.0/65536.0,1,-nbitq), 
to_sfixed(1242.0/65536.0,1,-nbitq), 
to_sfixed(-3149.0/65536.0,1,-nbitq), 
to_sfixed(3731.0/65536.0,1,-nbitq), 
to_sfixed(-1723.0/65536.0,1,-nbitq), 
to_sfixed(2686.0/65536.0,1,-nbitq), 
to_sfixed(-10858.0/65536.0,1,-nbitq), 
to_sfixed(941.0/65536.0,1,-nbitq), 
to_sfixed(5781.0/65536.0,1,-nbitq), 
to_sfixed(-1812.0/65536.0,1,-nbitq), 
to_sfixed(-2219.0/65536.0,1,-nbitq), 
to_sfixed(-2158.0/65536.0,1,-nbitq), 
to_sfixed(-3379.0/65536.0,1,-nbitq), 
to_sfixed(1701.0/65536.0,1,-nbitq), 
to_sfixed(-191.0/65536.0,1,-nbitq), 
to_sfixed(-9234.0/65536.0,1,-nbitq), 
to_sfixed(9287.0/65536.0,1,-nbitq), 
to_sfixed(-664.0/65536.0,1,-nbitq), 
to_sfixed(6703.0/65536.0,1,-nbitq), 
to_sfixed(-2133.0/65536.0,1,-nbitq), 
to_sfixed(2171.0/65536.0,1,-nbitq), 
to_sfixed(-780.0/65536.0,1,-nbitq), 
to_sfixed(-1073.0/65536.0,1,-nbitq), 
to_sfixed(1230.0/65536.0,1,-nbitq), 
to_sfixed(1208.0/65536.0,1,-nbitq), 
to_sfixed(6281.0/65536.0,1,-nbitq), 
to_sfixed(-8409.0/65536.0,1,-nbitq), 
to_sfixed(2311.0/65536.0,1,-nbitq), 
to_sfixed(796.0/65536.0,1,-nbitq), 
to_sfixed(2343.0/65536.0,1,-nbitq), 
to_sfixed(43.0/65536.0,1,-nbitq), 
to_sfixed(8809.0/65536.0,1,-nbitq), 
to_sfixed(1179.0/65536.0,1,-nbitq), 
to_sfixed(4822.0/65536.0,1,-nbitq), 
to_sfixed(2341.0/65536.0,1,-nbitq), 
to_sfixed(-10967.0/65536.0,1,-nbitq), 
to_sfixed(2111.0/65536.0,1,-nbitq), 
to_sfixed(-4574.0/65536.0,1,-nbitq), 
to_sfixed(-3284.0/65536.0,1,-nbitq), 
to_sfixed(-168.0/65536.0,1,-nbitq), 
to_sfixed(-492.0/65536.0,1,-nbitq), 
to_sfixed(299.0/65536.0,1,-nbitq), 
to_sfixed(1958.0/65536.0,1,-nbitq), 
to_sfixed(1147.0/65536.0,1,-nbitq), 
to_sfixed(468.0/65536.0,1,-nbitq), 
to_sfixed(-2066.0/65536.0,1,-nbitq), 
to_sfixed(-5482.0/65536.0,1,-nbitq), 
to_sfixed(-2942.0/65536.0,1,-nbitq), 
to_sfixed(-2000.0/65536.0,1,-nbitq), 
to_sfixed(-937.0/65536.0,1,-nbitq), 
to_sfixed(-8505.0/65536.0,1,-nbitq), 
to_sfixed(-1250.0/65536.0,1,-nbitq), 
to_sfixed(470.0/65536.0,1,-nbitq), 
to_sfixed(1100.0/65536.0,1,-nbitq), 
to_sfixed(-6487.0/65536.0,1,-nbitq), 
to_sfixed(3438.0/65536.0,1,-nbitq), 
to_sfixed(-294.0/65536.0,1,-nbitq), 
to_sfixed(-1460.0/65536.0,1,-nbitq), 
to_sfixed(2192.0/65536.0,1,-nbitq), 
to_sfixed(995.0/65536.0,1,-nbitq), 
to_sfixed(-4827.0/65536.0,1,-nbitq), 
to_sfixed(2010.0/65536.0,1,-nbitq), 
to_sfixed(151.0/65536.0,1,-nbitq), 
to_sfixed(3234.0/65536.0,1,-nbitq), 
to_sfixed(-1334.0/65536.0,1,-nbitq), 
to_sfixed(-4874.0/65536.0,1,-nbitq), 
to_sfixed(-2455.0/65536.0,1,-nbitq), 
to_sfixed(-687.0/65536.0,1,-nbitq), 
to_sfixed(-2625.0/65536.0,1,-nbitq), 
to_sfixed(162.0/65536.0,1,-nbitq), 
to_sfixed(-2741.0/65536.0,1,-nbitq), 
to_sfixed(1851.0/65536.0,1,-nbitq), 
to_sfixed(-2302.0/65536.0,1,-nbitq), 
to_sfixed(-873.0/65536.0,1,-nbitq), 
to_sfixed(473.0/65536.0,1,-nbitq)  ), 
( to_sfixed(903.0/65536.0,1,-nbitq), 
to_sfixed(2496.0/65536.0,1,-nbitq), 
to_sfixed(3350.0/65536.0,1,-nbitq), 
to_sfixed(-2303.0/65536.0,1,-nbitq), 
to_sfixed(3565.0/65536.0,1,-nbitq), 
to_sfixed(1232.0/65536.0,1,-nbitq), 
to_sfixed(3263.0/65536.0,1,-nbitq), 
to_sfixed(-2359.0/65536.0,1,-nbitq), 
to_sfixed(-1118.0/65536.0,1,-nbitq), 
to_sfixed(1386.0/65536.0,1,-nbitq), 
to_sfixed(7208.0/65536.0,1,-nbitq), 
to_sfixed(-10531.0/65536.0,1,-nbitq), 
to_sfixed(607.0/65536.0,1,-nbitq), 
to_sfixed(3660.0/65536.0,1,-nbitq), 
to_sfixed(158.0/65536.0,1,-nbitq), 
to_sfixed(-2809.0/65536.0,1,-nbitq), 
to_sfixed(471.0/65536.0,1,-nbitq), 
to_sfixed(-4298.0/65536.0,1,-nbitq), 
to_sfixed(721.0/65536.0,1,-nbitq), 
to_sfixed(483.0/65536.0,1,-nbitq), 
to_sfixed(-8181.0/65536.0,1,-nbitq), 
to_sfixed(-2963.0/65536.0,1,-nbitq), 
to_sfixed(-420.0/65536.0,1,-nbitq), 
to_sfixed(1858.0/65536.0,1,-nbitq), 
to_sfixed(-556.0/65536.0,1,-nbitq), 
to_sfixed(3378.0/65536.0,1,-nbitq), 
to_sfixed(-387.0/65536.0,1,-nbitq), 
to_sfixed(-2778.0/65536.0,1,-nbitq), 
to_sfixed(1970.0/65536.0,1,-nbitq), 
to_sfixed(-5181.0/65536.0,1,-nbitq), 
to_sfixed(6132.0/65536.0,1,-nbitq), 
to_sfixed(-2671.0/65536.0,1,-nbitq), 
to_sfixed(-6328.0/65536.0,1,-nbitq), 
to_sfixed(-1201.0/65536.0,1,-nbitq), 
to_sfixed(-1894.0/65536.0,1,-nbitq), 
to_sfixed(-665.0/65536.0,1,-nbitq), 
to_sfixed(6699.0/65536.0,1,-nbitq), 
to_sfixed(3898.0/65536.0,1,-nbitq), 
to_sfixed(7609.0/65536.0,1,-nbitq), 
to_sfixed(-2551.0/65536.0,1,-nbitq), 
to_sfixed(-7673.0/65536.0,1,-nbitq), 
to_sfixed(314.0/65536.0,1,-nbitq), 
to_sfixed(-11385.0/65536.0,1,-nbitq), 
to_sfixed(-8076.0/65536.0,1,-nbitq), 
to_sfixed(-2431.0/65536.0,1,-nbitq), 
to_sfixed(-8702.0/65536.0,1,-nbitq), 
to_sfixed(575.0/65536.0,1,-nbitq), 
to_sfixed(-7575.0/65536.0,1,-nbitq), 
to_sfixed(3245.0/65536.0,1,-nbitq), 
to_sfixed(-220.0/65536.0,1,-nbitq), 
to_sfixed(1327.0/65536.0,1,-nbitq), 
to_sfixed(-7049.0/65536.0,1,-nbitq), 
to_sfixed(3013.0/65536.0,1,-nbitq), 
to_sfixed(1248.0/65536.0,1,-nbitq), 
to_sfixed(-2617.0/65536.0,1,-nbitq), 
to_sfixed(-8114.0/65536.0,1,-nbitq), 
to_sfixed(-1606.0/65536.0,1,-nbitq), 
to_sfixed(-837.0/65536.0,1,-nbitq), 
to_sfixed(2194.0/65536.0,1,-nbitq), 
to_sfixed(-4197.0/65536.0,1,-nbitq), 
to_sfixed(-335.0/65536.0,1,-nbitq), 
to_sfixed(2342.0/65536.0,1,-nbitq), 
to_sfixed(3102.0/65536.0,1,-nbitq), 
to_sfixed(-1127.0/65536.0,1,-nbitq), 
to_sfixed(-982.0/65536.0,1,-nbitq), 
to_sfixed(-3859.0/65536.0,1,-nbitq), 
to_sfixed(1027.0/65536.0,1,-nbitq), 
to_sfixed(4773.0/65536.0,1,-nbitq), 
to_sfixed(2864.0/65536.0,1,-nbitq), 
to_sfixed(-4718.0/65536.0,1,-nbitq), 
to_sfixed(-1116.0/65536.0,1,-nbitq), 
to_sfixed(-2142.0/65536.0,1,-nbitq), 
to_sfixed(-1694.0/65536.0,1,-nbitq), 
to_sfixed(545.0/65536.0,1,-nbitq), 
to_sfixed(2188.0/65536.0,1,-nbitq), 
to_sfixed(-8097.0/65536.0,1,-nbitq), 
to_sfixed(-3091.0/65536.0,1,-nbitq), 
to_sfixed(-10822.0/65536.0,1,-nbitq), 
to_sfixed(-311.0/65536.0,1,-nbitq), 
to_sfixed(2303.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3260.0/65536.0,1,-nbitq), 
to_sfixed(244.0/65536.0,1,-nbitq), 
to_sfixed(2655.0/65536.0,1,-nbitq), 
to_sfixed(4872.0/65536.0,1,-nbitq), 
to_sfixed(7207.0/65536.0,1,-nbitq), 
to_sfixed(5664.0/65536.0,1,-nbitq), 
to_sfixed(1823.0/65536.0,1,-nbitq), 
to_sfixed(-5230.0/65536.0,1,-nbitq), 
to_sfixed(4118.0/65536.0,1,-nbitq), 
to_sfixed(404.0/65536.0,1,-nbitq), 
to_sfixed(6370.0/65536.0,1,-nbitq), 
to_sfixed(-8788.0/65536.0,1,-nbitq), 
to_sfixed(542.0/65536.0,1,-nbitq), 
to_sfixed(1314.0/65536.0,1,-nbitq), 
to_sfixed(-1707.0/65536.0,1,-nbitq), 
to_sfixed(-29.0/65536.0,1,-nbitq), 
to_sfixed(552.0/65536.0,1,-nbitq), 
to_sfixed(679.0/65536.0,1,-nbitq), 
to_sfixed(-1386.0/65536.0,1,-nbitq), 
to_sfixed(571.0/65536.0,1,-nbitq), 
to_sfixed(-1622.0/65536.0,1,-nbitq), 
to_sfixed(1922.0/65536.0,1,-nbitq), 
to_sfixed(454.0/65536.0,1,-nbitq), 
to_sfixed(-1493.0/65536.0,1,-nbitq), 
to_sfixed(1945.0/65536.0,1,-nbitq), 
to_sfixed(3241.0/65536.0,1,-nbitq), 
to_sfixed(-1477.0/65536.0,1,-nbitq), 
to_sfixed(1835.0/65536.0,1,-nbitq), 
to_sfixed(5640.0/65536.0,1,-nbitq), 
to_sfixed(-5625.0/65536.0,1,-nbitq), 
to_sfixed(6437.0/65536.0,1,-nbitq), 
to_sfixed(-5103.0/65536.0,1,-nbitq), 
to_sfixed(10.0/65536.0,1,-nbitq), 
to_sfixed(1239.0/65536.0,1,-nbitq), 
to_sfixed(65.0/65536.0,1,-nbitq), 
to_sfixed(549.0/65536.0,1,-nbitq), 
to_sfixed(7343.0/65536.0,1,-nbitq), 
to_sfixed(-783.0/65536.0,1,-nbitq), 
to_sfixed(3175.0/65536.0,1,-nbitq), 
to_sfixed(-1339.0/65536.0,1,-nbitq), 
to_sfixed(-9351.0/65536.0,1,-nbitq), 
to_sfixed(-3210.0/65536.0,1,-nbitq), 
to_sfixed(-12326.0/65536.0,1,-nbitq), 
to_sfixed(-4733.0/65536.0,1,-nbitq), 
to_sfixed(3148.0/65536.0,1,-nbitq), 
to_sfixed(-6243.0/65536.0,1,-nbitq), 
to_sfixed(-939.0/65536.0,1,-nbitq), 
to_sfixed(-3925.0/65536.0,1,-nbitq), 
to_sfixed(-556.0/65536.0,1,-nbitq), 
to_sfixed(-1239.0/65536.0,1,-nbitq), 
to_sfixed(1758.0/65536.0,1,-nbitq), 
to_sfixed(-3576.0/65536.0,1,-nbitq), 
to_sfixed(-2555.0/65536.0,1,-nbitq), 
to_sfixed(4311.0/65536.0,1,-nbitq), 
to_sfixed(-5429.0/65536.0,1,-nbitq), 
to_sfixed(-749.0/65536.0,1,-nbitq), 
to_sfixed(-2246.0/65536.0,1,-nbitq), 
to_sfixed(642.0/65536.0,1,-nbitq), 
to_sfixed(-2008.0/65536.0,1,-nbitq), 
to_sfixed(3121.0/65536.0,1,-nbitq), 
to_sfixed(-1355.0/65536.0,1,-nbitq), 
to_sfixed(-1490.0/65536.0,1,-nbitq), 
to_sfixed(-2129.0/65536.0,1,-nbitq), 
to_sfixed(734.0/65536.0,1,-nbitq), 
to_sfixed(-1761.0/65536.0,1,-nbitq), 
to_sfixed(-4205.0/65536.0,1,-nbitq), 
to_sfixed(-865.0/65536.0,1,-nbitq), 
to_sfixed(10638.0/65536.0,1,-nbitq), 
to_sfixed(1634.0/65536.0,1,-nbitq), 
to_sfixed(-1294.0/65536.0,1,-nbitq), 
to_sfixed(-6642.0/65536.0,1,-nbitq), 
to_sfixed(-5372.0/65536.0,1,-nbitq), 
to_sfixed(-2677.0/65536.0,1,-nbitq), 
to_sfixed(2570.0/65536.0,1,-nbitq), 
to_sfixed(-961.0/65536.0,1,-nbitq), 
to_sfixed(-5949.0/65536.0,1,-nbitq), 
to_sfixed(2286.0/65536.0,1,-nbitq), 
to_sfixed(-6192.0/65536.0,1,-nbitq), 
to_sfixed(-1820.0/65536.0,1,-nbitq), 
to_sfixed(2664.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1175.0/65536.0,1,-nbitq), 
to_sfixed(2223.0/65536.0,1,-nbitq), 
to_sfixed(6436.0/65536.0,1,-nbitq), 
to_sfixed(2973.0/65536.0,1,-nbitq), 
to_sfixed(10898.0/65536.0,1,-nbitq), 
to_sfixed(6100.0/65536.0,1,-nbitq), 
to_sfixed(3843.0/65536.0,1,-nbitq), 
to_sfixed(-6050.0/65536.0,1,-nbitq), 
to_sfixed(-843.0/65536.0,1,-nbitq), 
to_sfixed(1722.0/65536.0,1,-nbitq), 
to_sfixed(5653.0/65536.0,1,-nbitq), 
to_sfixed(3463.0/65536.0,1,-nbitq), 
to_sfixed(1805.0/65536.0,1,-nbitq), 
to_sfixed(-458.0/65536.0,1,-nbitq), 
to_sfixed(-1822.0/65536.0,1,-nbitq), 
to_sfixed(1080.0/65536.0,1,-nbitq), 
to_sfixed(679.0/65536.0,1,-nbitq), 
to_sfixed(3783.0/65536.0,1,-nbitq), 
to_sfixed(2166.0/65536.0,1,-nbitq), 
to_sfixed(1986.0/65536.0,1,-nbitq), 
to_sfixed(-1919.0/65536.0,1,-nbitq), 
to_sfixed(-3283.0/65536.0,1,-nbitq), 
to_sfixed(-1930.0/65536.0,1,-nbitq), 
to_sfixed(4067.0/65536.0,1,-nbitq), 
to_sfixed(-1600.0/65536.0,1,-nbitq), 
to_sfixed(8745.0/65536.0,1,-nbitq), 
to_sfixed(-500.0/65536.0,1,-nbitq), 
to_sfixed(2716.0/65536.0,1,-nbitq), 
to_sfixed(3014.0/65536.0,1,-nbitq), 
to_sfixed(211.0/65536.0,1,-nbitq), 
to_sfixed(4343.0/65536.0,1,-nbitq), 
to_sfixed(-344.0/65536.0,1,-nbitq), 
to_sfixed(3468.0/65536.0,1,-nbitq), 
to_sfixed(4246.0/65536.0,1,-nbitq), 
to_sfixed(-3378.0/65536.0,1,-nbitq), 
to_sfixed(-584.0/65536.0,1,-nbitq), 
to_sfixed(5298.0/65536.0,1,-nbitq), 
to_sfixed(-1296.0/65536.0,1,-nbitq), 
to_sfixed(-8354.0/65536.0,1,-nbitq), 
to_sfixed(1766.0/65536.0,1,-nbitq), 
to_sfixed(-4123.0/65536.0,1,-nbitq), 
to_sfixed(1827.0/65536.0,1,-nbitq), 
to_sfixed(-5528.0/65536.0,1,-nbitq), 
to_sfixed(-1182.0/65536.0,1,-nbitq), 
to_sfixed(958.0/65536.0,1,-nbitq), 
to_sfixed(-1481.0/65536.0,1,-nbitq), 
to_sfixed(916.0/65536.0,1,-nbitq), 
to_sfixed(-5394.0/65536.0,1,-nbitq), 
to_sfixed(1568.0/65536.0,1,-nbitq), 
to_sfixed(2137.0/65536.0,1,-nbitq), 
to_sfixed(840.0/65536.0,1,-nbitq), 
to_sfixed(-3819.0/65536.0,1,-nbitq), 
to_sfixed(-5076.0/65536.0,1,-nbitq), 
to_sfixed(-1667.0/65536.0,1,-nbitq), 
to_sfixed(955.0/65536.0,1,-nbitq), 
to_sfixed(3651.0/65536.0,1,-nbitq), 
to_sfixed(387.0/65536.0,1,-nbitq), 
to_sfixed(-2551.0/65536.0,1,-nbitq), 
to_sfixed(-2878.0/65536.0,1,-nbitq), 
to_sfixed(2742.0/65536.0,1,-nbitq), 
to_sfixed(-1754.0/65536.0,1,-nbitq), 
to_sfixed(1818.0/65536.0,1,-nbitq), 
to_sfixed(-1542.0/65536.0,1,-nbitq), 
to_sfixed(995.0/65536.0,1,-nbitq), 
to_sfixed(-938.0/65536.0,1,-nbitq), 
to_sfixed(-962.0/65536.0,1,-nbitq), 
to_sfixed(-5402.0/65536.0,1,-nbitq), 
to_sfixed(3233.0/65536.0,1,-nbitq), 
to_sfixed(1255.0/65536.0,1,-nbitq), 
to_sfixed(-3571.0/65536.0,1,-nbitq), 
to_sfixed(-3323.0/65536.0,1,-nbitq), 
to_sfixed(-4757.0/65536.0,1,-nbitq), 
to_sfixed(5222.0/65536.0,1,-nbitq), 
to_sfixed(1309.0/65536.0,1,-nbitq), 
to_sfixed(-1237.0/65536.0,1,-nbitq), 
to_sfixed(2561.0/65536.0,1,-nbitq), 
to_sfixed(7537.0/65536.0,1,-nbitq), 
to_sfixed(-9873.0/65536.0,1,-nbitq), 
to_sfixed(662.0/65536.0,1,-nbitq), 
to_sfixed(-751.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-969.0/65536.0,1,-nbitq), 
to_sfixed(966.0/65536.0,1,-nbitq), 
to_sfixed(10559.0/65536.0,1,-nbitq), 
to_sfixed(-303.0/65536.0,1,-nbitq), 
to_sfixed(7964.0/65536.0,1,-nbitq), 
to_sfixed(8245.0/65536.0,1,-nbitq), 
to_sfixed(2999.0/65536.0,1,-nbitq), 
to_sfixed(-3994.0/65536.0,1,-nbitq), 
to_sfixed(3110.0/65536.0,1,-nbitq), 
to_sfixed(-1632.0/65536.0,1,-nbitq), 
to_sfixed(7172.0/65536.0,1,-nbitq), 
to_sfixed(-1268.0/65536.0,1,-nbitq), 
to_sfixed(-444.0/65536.0,1,-nbitq), 
to_sfixed(3569.0/65536.0,1,-nbitq), 
to_sfixed(-1131.0/65536.0,1,-nbitq), 
to_sfixed(-730.0/65536.0,1,-nbitq), 
to_sfixed(2432.0/65536.0,1,-nbitq), 
to_sfixed(-1248.0/65536.0,1,-nbitq), 
to_sfixed(858.0/65536.0,1,-nbitq), 
to_sfixed(1436.0/65536.0,1,-nbitq), 
to_sfixed(-594.0/65536.0,1,-nbitq), 
to_sfixed(2006.0/65536.0,1,-nbitq), 
to_sfixed(1276.0/65536.0,1,-nbitq), 
to_sfixed(5795.0/65536.0,1,-nbitq), 
to_sfixed(1465.0/65536.0,1,-nbitq), 
to_sfixed(7982.0/65536.0,1,-nbitq), 
to_sfixed(156.0/65536.0,1,-nbitq), 
to_sfixed(-1723.0/65536.0,1,-nbitq), 
to_sfixed(1860.0/65536.0,1,-nbitq), 
to_sfixed(-179.0/65536.0,1,-nbitq), 
to_sfixed(3408.0/65536.0,1,-nbitq), 
to_sfixed(3812.0/65536.0,1,-nbitq), 
to_sfixed(1232.0/65536.0,1,-nbitq), 
to_sfixed(3249.0/65536.0,1,-nbitq), 
to_sfixed(-3789.0/65536.0,1,-nbitq), 
to_sfixed(-977.0/65536.0,1,-nbitq), 
to_sfixed(5752.0/65536.0,1,-nbitq), 
to_sfixed(566.0/65536.0,1,-nbitq), 
to_sfixed(-8368.0/65536.0,1,-nbitq), 
to_sfixed(2145.0/65536.0,1,-nbitq), 
to_sfixed(274.0/65536.0,1,-nbitq), 
to_sfixed(-2359.0/65536.0,1,-nbitq), 
to_sfixed(-4334.0/65536.0,1,-nbitq), 
to_sfixed(-2461.0/65536.0,1,-nbitq), 
to_sfixed(-1030.0/65536.0,1,-nbitq), 
to_sfixed(-646.0/65536.0,1,-nbitq), 
to_sfixed(-3508.0/65536.0,1,-nbitq), 
to_sfixed(-6899.0/65536.0,1,-nbitq), 
to_sfixed(-3001.0/65536.0,1,-nbitq), 
to_sfixed(3196.0/65536.0,1,-nbitq), 
to_sfixed(-2374.0/65536.0,1,-nbitq), 
to_sfixed(-8767.0/65536.0,1,-nbitq), 
to_sfixed(-9351.0/65536.0,1,-nbitq), 
to_sfixed(-7026.0/65536.0,1,-nbitq), 
to_sfixed(933.0/65536.0,1,-nbitq), 
to_sfixed(4781.0/65536.0,1,-nbitq), 
to_sfixed(-2074.0/65536.0,1,-nbitq), 
to_sfixed(581.0/65536.0,1,-nbitq), 
to_sfixed(-754.0/65536.0,1,-nbitq), 
to_sfixed(-4502.0/65536.0,1,-nbitq), 
to_sfixed(-1275.0/65536.0,1,-nbitq), 
to_sfixed(425.0/65536.0,1,-nbitq), 
to_sfixed(-1248.0/65536.0,1,-nbitq), 
to_sfixed(-3153.0/65536.0,1,-nbitq), 
to_sfixed(-29.0/65536.0,1,-nbitq), 
to_sfixed(-2353.0/65536.0,1,-nbitq), 
to_sfixed(-5057.0/65536.0,1,-nbitq), 
to_sfixed(5252.0/65536.0,1,-nbitq), 
to_sfixed(8410.0/65536.0,1,-nbitq), 
to_sfixed(-5558.0/65536.0,1,-nbitq), 
to_sfixed(-2606.0/65536.0,1,-nbitq), 
to_sfixed(-3115.0/65536.0,1,-nbitq), 
to_sfixed(6924.0/65536.0,1,-nbitq), 
to_sfixed(1711.0/65536.0,1,-nbitq), 
to_sfixed(1792.0/65536.0,1,-nbitq), 
to_sfixed(4988.0/65536.0,1,-nbitq), 
to_sfixed(9442.0/65536.0,1,-nbitq), 
to_sfixed(-4609.0/65536.0,1,-nbitq), 
to_sfixed(-2646.0/65536.0,1,-nbitq), 
to_sfixed(-1159.0/65536.0,1,-nbitq)  ), 
( to_sfixed(495.0/65536.0,1,-nbitq), 
to_sfixed(-1996.0/65536.0,1,-nbitq), 
to_sfixed(11010.0/65536.0,1,-nbitq), 
to_sfixed(1038.0/65536.0,1,-nbitq), 
to_sfixed(9047.0/65536.0,1,-nbitq), 
to_sfixed(3485.0/65536.0,1,-nbitq), 
to_sfixed(272.0/65536.0,1,-nbitq), 
to_sfixed(-246.0/65536.0,1,-nbitq), 
to_sfixed(-94.0/65536.0,1,-nbitq), 
to_sfixed(-2506.0/65536.0,1,-nbitq), 
to_sfixed(5937.0/65536.0,1,-nbitq), 
to_sfixed(-7999.0/65536.0,1,-nbitq), 
to_sfixed(826.0/65536.0,1,-nbitq), 
to_sfixed(4962.0/65536.0,1,-nbitq), 
to_sfixed(-3390.0/65536.0,1,-nbitq), 
to_sfixed(-692.0/65536.0,1,-nbitq), 
to_sfixed(-3367.0/65536.0,1,-nbitq), 
to_sfixed(2714.0/65536.0,1,-nbitq), 
to_sfixed(852.0/65536.0,1,-nbitq), 
to_sfixed(-1423.0/65536.0,1,-nbitq), 
to_sfixed(313.0/65536.0,1,-nbitq), 
to_sfixed(4584.0/65536.0,1,-nbitq), 
to_sfixed(8527.0/65536.0,1,-nbitq), 
to_sfixed(11251.0/65536.0,1,-nbitq), 
to_sfixed(714.0/65536.0,1,-nbitq), 
to_sfixed(5808.0/65536.0,1,-nbitq), 
to_sfixed(1436.0/65536.0,1,-nbitq), 
to_sfixed(-2901.0/65536.0,1,-nbitq), 
to_sfixed(808.0/65536.0,1,-nbitq), 
to_sfixed(-370.0/65536.0,1,-nbitq), 
to_sfixed(1456.0/65536.0,1,-nbitq), 
to_sfixed(458.0/65536.0,1,-nbitq), 
to_sfixed(3104.0/65536.0,1,-nbitq), 
to_sfixed(733.0/65536.0,1,-nbitq), 
to_sfixed(-38.0/65536.0,1,-nbitq), 
to_sfixed(1430.0/65536.0,1,-nbitq), 
to_sfixed(1826.0/65536.0,1,-nbitq), 
to_sfixed(1595.0/65536.0,1,-nbitq), 
to_sfixed(-118.0/65536.0,1,-nbitq), 
to_sfixed(-1123.0/65536.0,1,-nbitq), 
to_sfixed(5342.0/65536.0,1,-nbitq), 
to_sfixed(-2985.0/65536.0,1,-nbitq), 
to_sfixed(-2198.0/65536.0,1,-nbitq), 
to_sfixed(-7426.0/65536.0,1,-nbitq), 
to_sfixed(-506.0/65536.0,1,-nbitq), 
to_sfixed(2687.0/65536.0,1,-nbitq), 
to_sfixed(-1247.0/65536.0,1,-nbitq), 
to_sfixed(693.0/65536.0,1,-nbitq), 
to_sfixed(-2560.0/65536.0,1,-nbitq), 
to_sfixed(2892.0/65536.0,1,-nbitq), 
to_sfixed(2391.0/65536.0,1,-nbitq), 
to_sfixed(-9619.0/65536.0,1,-nbitq), 
to_sfixed(-9122.0/65536.0,1,-nbitq), 
to_sfixed(272.0/65536.0,1,-nbitq), 
to_sfixed(7147.0/65536.0,1,-nbitq), 
to_sfixed(4121.0/65536.0,1,-nbitq), 
to_sfixed(1996.0/65536.0,1,-nbitq), 
to_sfixed(2010.0/65536.0,1,-nbitq), 
to_sfixed(774.0/65536.0,1,-nbitq), 
to_sfixed(-3823.0/65536.0,1,-nbitq), 
to_sfixed(-3976.0/65536.0,1,-nbitq), 
to_sfixed(-476.0/65536.0,1,-nbitq), 
to_sfixed(1918.0/65536.0,1,-nbitq), 
to_sfixed(-1503.0/65536.0,1,-nbitq), 
to_sfixed(-1439.0/65536.0,1,-nbitq), 
to_sfixed(538.0/65536.0,1,-nbitq), 
to_sfixed(-6025.0/65536.0,1,-nbitq), 
to_sfixed(-500.0/65536.0,1,-nbitq), 
to_sfixed(6239.0/65536.0,1,-nbitq), 
to_sfixed(-8775.0/65536.0,1,-nbitq), 
to_sfixed(-3168.0/65536.0,1,-nbitq), 
to_sfixed(2939.0/65536.0,1,-nbitq), 
to_sfixed(4744.0/65536.0,1,-nbitq), 
to_sfixed(2464.0/65536.0,1,-nbitq), 
to_sfixed(-1306.0/65536.0,1,-nbitq), 
to_sfixed(845.0/65536.0,1,-nbitq), 
to_sfixed(10229.0/65536.0,1,-nbitq), 
to_sfixed(-3422.0/65536.0,1,-nbitq), 
to_sfixed(-1760.0/65536.0,1,-nbitq), 
to_sfixed(-1208.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3294.0/65536.0,1,-nbitq), 
to_sfixed(-3859.0/65536.0,1,-nbitq), 
to_sfixed(781.0/65536.0,1,-nbitq), 
to_sfixed(-168.0/65536.0,1,-nbitq), 
to_sfixed(10035.0/65536.0,1,-nbitq), 
to_sfixed(2908.0/65536.0,1,-nbitq), 
to_sfixed(1597.0/65536.0,1,-nbitq), 
to_sfixed(-3224.0/65536.0,1,-nbitq), 
to_sfixed(2890.0/65536.0,1,-nbitq), 
to_sfixed(337.0/65536.0,1,-nbitq), 
to_sfixed(1832.0/65536.0,1,-nbitq), 
to_sfixed(-1829.0/65536.0,1,-nbitq), 
to_sfixed(-814.0/65536.0,1,-nbitq), 
to_sfixed(5355.0/65536.0,1,-nbitq), 
to_sfixed(-1405.0/65536.0,1,-nbitq), 
to_sfixed(1211.0/65536.0,1,-nbitq), 
to_sfixed(-656.0/65536.0,1,-nbitq), 
to_sfixed(747.0/65536.0,1,-nbitq), 
to_sfixed(-3381.0/65536.0,1,-nbitq), 
to_sfixed(-476.0/65536.0,1,-nbitq), 
to_sfixed(-628.0/65536.0,1,-nbitq), 
to_sfixed(3132.0/65536.0,1,-nbitq), 
to_sfixed(1542.0/65536.0,1,-nbitq), 
to_sfixed(7305.0/65536.0,1,-nbitq), 
to_sfixed(-2928.0/65536.0,1,-nbitq), 
to_sfixed(3438.0/65536.0,1,-nbitq), 
to_sfixed(2477.0/65536.0,1,-nbitq), 
to_sfixed(1162.0/65536.0,1,-nbitq), 
to_sfixed(-1623.0/65536.0,1,-nbitq), 
to_sfixed(2394.0/65536.0,1,-nbitq), 
to_sfixed(-740.0/65536.0,1,-nbitq), 
to_sfixed(2841.0/65536.0,1,-nbitq), 
to_sfixed(718.0/65536.0,1,-nbitq), 
to_sfixed(-1415.0/65536.0,1,-nbitq), 
to_sfixed(-1388.0/65536.0,1,-nbitq), 
to_sfixed(-1569.0/65536.0,1,-nbitq), 
to_sfixed(6265.0/65536.0,1,-nbitq), 
to_sfixed(-486.0/65536.0,1,-nbitq), 
to_sfixed(1039.0/65536.0,1,-nbitq), 
to_sfixed(366.0/65536.0,1,-nbitq), 
to_sfixed(6381.0/65536.0,1,-nbitq), 
to_sfixed(2619.0/65536.0,1,-nbitq), 
to_sfixed(-2705.0/65536.0,1,-nbitq), 
to_sfixed(-2818.0/65536.0,1,-nbitq), 
to_sfixed(1329.0/65536.0,1,-nbitq), 
to_sfixed(5377.0/65536.0,1,-nbitq), 
to_sfixed(671.0/65536.0,1,-nbitq), 
to_sfixed(1230.0/65536.0,1,-nbitq), 
to_sfixed(1151.0/65536.0,1,-nbitq), 
to_sfixed(-906.0/65536.0,1,-nbitq), 
to_sfixed(451.0/65536.0,1,-nbitq), 
to_sfixed(-5547.0/65536.0,1,-nbitq), 
to_sfixed(-6040.0/65536.0,1,-nbitq), 
to_sfixed(29.0/65536.0,1,-nbitq), 
to_sfixed(7835.0/65536.0,1,-nbitq), 
to_sfixed(1822.0/65536.0,1,-nbitq), 
to_sfixed(-527.0/65536.0,1,-nbitq), 
to_sfixed(-1857.0/65536.0,1,-nbitq), 
to_sfixed(-353.0/65536.0,1,-nbitq), 
to_sfixed(3785.0/65536.0,1,-nbitq), 
to_sfixed(596.0/65536.0,1,-nbitq), 
to_sfixed(-1502.0/65536.0,1,-nbitq), 
to_sfixed(-952.0/65536.0,1,-nbitq), 
to_sfixed(-1959.0/65536.0,1,-nbitq), 
to_sfixed(-3443.0/65536.0,1,-nbitq), 
to_sfixed(2628.0/65536.0,1,-nbitq), 
to_sfixed(-4918.0/65536.0,1,-nbitq), 
to_sfixed(-3436.0/65536.0,1,-nbitq), 
to_sfixed(1364.0/65536.0,1,-nbitq), 
to_sfixed(-9356.0/65536.0,1,-nbitq), 
to_sfixed(-1341.0/65536.0,1,-nbitq), 
to_sfixed(-653.0/65536.0,1,-nbitq), 
to_sfixed(777.0/65536.0,1,-nbitq), 
to_sfixed(-1453.0/65536.0,1,-nbitq), 
to_sfixed(-3011.0/65536.0,1,-nbitq), 
to_sfixed(-656.0/65536.0,1,-nbitq), 
to_sfixed(10130.0/65536.0,1,-nbitq), 
to_sfixed(-2615.0/65536.0,1,-nbitq), 
to_sfixed(2075.0/65536.0,1,-nbitq), 
to_sfixed(307.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2640.0/65536.0,1,-nbitq), 
to_sfixed(-3047.0/65536.0,1,-nbitq), 
to_sfixed(3680.0/65536.0,1,-nbitq), 
to_sfixed(-2235.0/65536.0,1,-nbitq), 
to_sfixed(3444.0/65536.0,1,-nbitq), 
to_sfixed(-1809.0/65536.0,1,-nbitq), 
to_sfixed(-323.0/65536.0,1,-nbitq), 
to_sfixed(-905.0/65536.0,1,-nbitq), 
to_sfixed(-716.0/65536.0,1,-nbitq), 
to_sfixed(-1478.0/65536.0,1,-nbitq), 
to_sfixed(-3502.0/65536.0,1,-nbitq), 
to_sfixed(-587.0/65536.0,1,-nbitq), 
to_sfixed(1772.0/65536.0,1,-nbitq), 
to_sfixed(3132.0/65536.0,1,-nbitq), 
to_sfixed(2682.0/65536.0,1,-nbitq), 
to_sfixed(1214.0/65536.0,1,-nbitq), 
to_sfixed(2649.0/65536.0,1,-nbitq), 
to_sfixed(1268.0/65536.0,1,-nbitq), 
to_sfixed(-2051.0/65536.0,1,-nbitq), 
to_sfixed(-1766.0/65536.0,1,-nbitq), 
to_sfixed(-1262.0/65536.0,1,-nbitq), 
to_sfixed(5615.0/65536.0,1,-nbitq), 
to_sfixed(-1907.0/65536.0,1,-nbitq), 
to_sfixed(8640.0/65536.0,1,-nbitq), 
to_sfixed(1902.0/65536.0,1,-nbitq), 
to_sfixed(2288.0/65536.0,1,-nbitq), 
to_sfixed(-722.0/65536.0,1,-nbitq), 
to_sfixed(739.0/65536.0,1,-nbitq), 
to_sfixed(-4109.0/65536.0,1,-nbitq), 
to_sfixed(1064.0/65536.0,1,-nbitq), 
to_sfixed(263.0/65536.0,1,-nbitq), 
to_sfixed(-1706.0/65536.0,1,-nbitq), 
to_sfixed(2133.0/65536.0,1,-nbitq), 
to_sfixed(2016.0/65536.0,1,-nbitq), 
to_sfixed(-1390.0/65536.0,1,-nbitq), 
to_sfixed(1285.0/65536.0,1,-nbitq), 
to_sfixed(2709.0/65536.0,1,-nbitq), 
to_sfixed(-638.0/65536.0,1,-nbitq), 
to_sfixed(3865.0/65536.0,1,-nbitq), 
to_sfixed(638.0/65536.0,1,-nbitq), 
to_sfixed(2788.0/65536.0,1,-nbitq), 
to_sfixed(-750.0/65536.0,1,-nbitq), 
to_sfixed(1067.0/65536.0,1,-nbitq), 
to_sfixed(-5947.0/65536.0,1,-nbitq), 
to_sfixed(-1644.0/65536.0,1,-nbitq), 
to_sfixed(4356.0/65536.0,1,-nbitq), 
to_sfixed(-3083.0/65536.0,1,-nbitq), 
to_sfixed(4043.0/65536.0,1,-nbitq), 
to_sfixed(978.0/65536.0,1,-nbitq), 
to_sfixed(-257.0/65536.0,1,-nbitq), 
to_sfixed(-1064.0/65536.0,1,-nbitq), 
to_sfixed(-8366.0/65536.0,1,-nbitq), 
to_sfixed(-4170.0/65536.0,1,-nbitq), 
to_sfixed(-4395.0/65536.0,1,-nbitq), 
to_sfixed(1701.0/65536.0,1,-nbitq), 
to_sfixed(-167.0/65536.0,1,-nbitq), 
to_sfixed(-2274.0/65536.0,1,-nbitq), 
to_sfixed(-2470.0/65536.0,1,-nbitq), 
to_sfixed(256.0/65536.0,1,-nbitq), 
to_sfixed(4390.0/65536.0,1,-nbitq), 
to_sfixed(-906.0/65536.0,1,-nbitq), 
to_sfixed(-109.0/65536.0,1,-nbitq), 
to_sfixed(446.0/65536.0,1,-nbitq), 
to_sfixed(1921.0/65536.0,1,-nbitq), 
to_sfixed(-321.0/65536.0,1,-nbitq), 
to_sfixed(-1252.0/65536.0,1,-nbitq), 
to_sfixed(-5769.0/65536.0,1,-nbitq), 
to_sfixed(-5716.0/65536.0,1,-nbitq), 
to_sfixed(-5973.0/65536.0,1,-nbitq), 
to_sfixed(-8015.0/65536.0,1,-nbitq), 
to_sfixed(2307.0/65536.0,1,-nbitq), 
to_sfixed(-3439.0/65536.0,1,-nbitq), 
to_sfixed(823.0/65536.0,1,-nbitq), 
to_sfixed(-3013.0/65536.0,1,-nbitq), 
to_sfixed(220.0/65536.0,1,-nbitq), 
to_sfixed(990.0/65536.0,1,-nbitq), 
to_sfixed(3217.0/65536.0,1,-nbitq), 
to_sfixed(2081.0/65536.0,1,-nbitq), 
to_sfixed(-686.0/65536.0,1,-nbitq), 
to_sfixed(-3142.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2701.0/65536.0,1,-nbitq), 
to_sfixed(1742.0/65536.0,1,-nbitq), 
to_sfixed(2283.0/65536.0,1,-nbitq), 
to_sfixed(-2216.0/65536.0,1,-nbitq), 
to_sfixed(4322.0/65536.0,1,-nbitq), 
to_sfixed(-14.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(-38.0/65536.0,1,-nbitq), 
to_sfixed(1314.0/65536.0,1,-nbitq), 
to_sfixed(2942.0/65536.0,1,-nbitq), 
to_sfixed(2517.0/65536.0,1,-nbitq), 
to_sfixed(3587.0/65536.0,1,-nbitq), 
to_sfixed(-1528.0/65536.0,1,-nbitq), 
to_sfixed(2540.0/65536.0,1,-nbitq), 
to_sfixed(-958.0/65536.0,1,-nbitq), 
to_sfixed(2336.0/65536.0,1,-nbitq), 
to_sfixed(-3100.0/65536.0,1,-nbitq), 
to_sfixed(-4126.0/65536.0,1,-nbitq), 
to_sfixed(-2549.0/65536.0,1,-nbitq), 
to_sfixed(385.0/65536.0,1,-nbitq), 
to_sfixed(-4456.0/65536.0,1,-nbitq), 
to_sfixed(-781.0/65536.0,1,-nbitq), 
to_sfixed(-2247.0/65536.0,1,-nbitq), 
to_sfixed(3273.0/65536.0,1,-nbitq), 
to_sfixed(1916.0/65536.0,1,-nbitq), 
to_sfixed(4570.0/65536.0,1,-nbitq), 
to_sfixed(-377.0/65536.0,1,-nbitq), 
to_sfixed(2859.0/65536.0,1,-nbitq), 
to_sfixed(-226.0/65536.0,1,-nbitq), 
to_sfixed(-832.0/65536.0,1,-nbitq), 
to_sfixed(-2719.0/65536.0,1,-nbitq), 
to_sfixed(-1169.0/65536.0,1,-nbitq), 
to_sfixed(2876.0/65536.0,1,-nbitq), 
to_sfixed(2157.0/65536.0,1,-nbitq), 
to_sfixed(-2473.0/65536.0,1,-nbitq), 
to_sfixed(2814.0/65536.0,1,-nbitq), 
to_sfixed(200.0/65536.0,1,-nbitq), 
to_sfixed(-3174.0/65536.0,1,-nbitq), 
to_sfixed(-4188.0/65536.0,1,-nbitq), 
to_sfixed(-1442.0/65536.0,1,-nbitq), 
to_sfixed(-1016.0/65536.0,1,-nbitq), 
to_sfixed(998.0/65536.0,1,-nbitq), 
to_sfixed(-928.0/65536.0,1,-nbitq), 
to_sfixed(-2420.0/65536.0,1,-nbitq), 
to_sfixed(800.0/65536.0,1,-nbitq), 
to_sfixed(2133.0/65536.0,1,-nbitq), 
to_sfixed(-1026.0/65536.0,1,-nbitq), 
to_sfixed(3094.0/65536.0,1,-nbitq), 
to_sfixed(3073.0/65536.0,1,-nbitq), 
to_sfixed(1794.0/65536.0,1,-nbitq), 
to_sfixed(1822.0/65536.0,1,-nbitq), 
to_sfixed(-6320.0/65536.0,1,-nbitq), 
to_sfixed(4325.0/65536.0,1,-nbitq), 
to_sfixed(-1880.0/65536.0,1,-nbitq), 
to_sfixed(2606.0/65536.0,1,-nbitq), 
to_sfixed(2765.0/65536.0,1,-nbitq), 
to_sfixed(-1483.0/65536.0,1,-nbitq), 
to_sfixed(-1452.0/65536.0,1,-nbitq), 
to_sfixed(543.0/65536.0,1,-nbitq), 
to_sfixed(4850.0/65536.0,1,-nbitq), 
to_sfixed(3326.0/65536.0,1,-nbitq), 
to_sfixed(-1218.0/65536.0,1,-nbitq), 
to_sfixed(1723.0/65536.0,1,-nbitq), 
to_sfixed(-2732.0/65536.0,1,-nbitq), 
to_sfixed(725.0/65536.0,1,-nbitq), 
to_sfixed(-978.0/65536.0,1,-nbitq), 
to_sfixed(-6663.0/65536.0,1,-nbitq), 
to_sfixed(-3447.0/65536.0,1,-nbitq), 
to_sfixed(-1743.0/65536.0,1,-nbitq), 
to_sfixed(-7260.0/65536.0,1,-nbitq), 
to_sfixed(3566.0/65536.0,1,-nbitq), 
to_sfixed(-4632.0/65536.0,1,-nbitq), 
to_sfixed(3602.0/65536.0,1,-nbitq), 
to_sfixed(-364.0/65536.0,1,-nbitq), 
to_sfixed(2348.0/65536.0,1,-nbitq), 
to_sfixed(-536.0/65536.0,1,-nbitq), 
to_sfixed(-2642.0/65536.0,1,-nbitq), 
to_sfixed(1738.0/65536.0,1,-nbitq), 
to_sfixed(-353.0/65536.0,1,-nbitq), 
to_sfixed(990.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3139.0/65536.0,1,-nbitq), 
to_sfixed(-3082.0/65536.0,1,-nbitq), 
to_sfixed(-1.0/65536.0,1,-nbitq), 
to_sfixed(-1506.0/65536.0,1,-nbitq), 
to_sfixed(-1753.0/65536.0,1,-nbitq), 
to_sfixed(-2320.0/65536.0,1,-nbitq), 
to_sfixed(2181.0/65536.0,1,-nbitq), 
to_sfixed(-2551.0/65536.0,1,-nbitq), 
to_sfixed(-913.0/65536.0,1,-nbitq), 
to_sfixed(-108.0/65536.0,1,-nbitq), 
to_sfixed(-1386.0/65536.0,1,-nbitq), 
to_sfixed(132.0/65536.0,1,-nbitq), 
to_sfixed(-2044.0/65536.0,1,-nbitq), 
to_sfixed(-513.0/65536.0,1,-nbitq), 
to_sfixed(296.0/65536.0,1,-nbitq), 
to_sfixed(642.0/65536.0,1,-nbitq), 
to_sfixed(1172.0/65536.0,1,-nbitq), 
to_sfixed(1254.0/65536.0,1,-nbitq), 
to_sfixed(-2718.0/65536.0,1,-nbitq), 
to_sfixed(199.0/65536.0,1,-nbitq), 
to_sfixed(-4479.0/65536.0,1,-nbitq), 
to_sfixed(486.0/65536.0,1,-nbitq), 
to_sfixed(2788.0/65536.0,1,-nbitq), 
to_sfixed(-594.0/65536.0,1,-nbitq), 
to_sfixed(1206.0/65536.0,1,-nbitq), 
to_sfixed(4181.0/65536.0,1,-nbitq), 
to_sfixed(2214.0/65536.0,1,-nbitq), 
to_sfixed(326.0/65536.0,1,-nbitq), 
to_sfixed(2041.0/65536.0,1,-nbitq), 
to_sfixed(3396.0/65536.0,1,-nbitq), 
to_sfixed(-507.0/65536.0,1,-nbitq), 
to_sfixed(2805.0/65536.0,1,-nbitq), 
to_sfixed(3043.0/65536.0,1,-nbitq), 
to_sfixed(-696.0/65536.0,1,-nbitq), 
to_sfixed(-439.0/65536.0,1,-nbitq), 
to_sfixed(1887.0/65536.0,1,-nbitq), 
to_sfixed(-349.0/65536.0,1,-nbitq), 
to_sfixed(-1115.0/65536.0,1,-nbitq), 
to_sfixed(1046.0/65536.0,1,-nbitq), 
to_sfixed(-2135.0/65536.0,1,-nbitq), 
to_sfixed(-6600.0/65536.0,1,-nbitq), 
to_sfixed(576.0/65536.0,1,-nbitq), 
to_sfixed(156.0/65536.0,1,-nbitq), 
to_sfixed(235.0/65536.0,1,-nbitq), 
to_sfixed(-1284.0/65536.0,1,-nbitq), 
to_sfixed(5070.0/65536.0,1,-nbitq), 
to_sfixed(845.0/65536.0,1,-nbitq), 
to_sfixed(-2280.0/65536.0,1,-nbitq), 
to_sfixed(1741.0/65536.0,1,-nbitq), 
to_sfixed(-353.0/65536.0,1,-nbitq), 
to_sfixed(-2020.0/65536.0,1,-nbitq), 
to_sfixed(-4751.0/65536.0,1,-nbitq), 
to_sfixed(-1061.0/65536.0,1,-nbitq), 
to_sfixed(-1843.0/65536.0,1,-nbitq), 
to_sfixed(438.0/65536.0,1,-nbitq), 
to_sfixed(3019.0/65536.0,1,-nbitq), 
to_sfixed(-1461.0/65536.0,1,-nbitq), 
to_sfixed(-235.0/65536.0,1,-nbitq), 
to_sfixed(-1053.0/65536.0,1,-nbitq), 
to_sfixed(2967.0/65536.0,1,-nbitq), 
to_sfixed(-849.0/65536.0,1,-nbitq), 
to_sfixed(-2335.0/65536.0,1,-nbitq), 
to_sfixed(-1070.0/65536.0,1,-nbitq), 
to_sfixed(-3007.0/65536.0,1,-nbitq), 
to_sfixed(-679.0/65536.0,1,-nbitq), 
to_sfixed(1181.0/65536.0,1,-nbitq), 
to_sfixed(-6109.0/65536.0,1,-nbitq), 
to_sfixed(949.0/65536.0,1,-nbitq), 
to_sfixed(-2941.0/65536.0,1,-nbitq), 
to_sfixed(-2581.0/65536.0,1,-nbitq), 
to_sfixed(846.0/65536.0,1,-nbitq), 
to_sfixed(-5441.0/65536.0,1,-nbitq), 
to_sfixed(117.0/65536.0,1,-nbitq), 
to_sfixed(2614.0/65536.0,1,-nbitq), 
to_sfixed(-2634.0/65536.0,1,-nbitq), 
to_sfixed(2455.0/65536.0,1,-nbitq), 
to_sfixed(2217.0/65536.0,1,-nbitq), 
to_sfixed(2536.0/65536.0,1,-nbitq), 
to_sfixed(-1712.0/65536.0,1,-nbitq), 
to_sfixed(411.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3418.0/65536.0,1,-nbitq), 
to_sfixed(1687.0/65536.0,1,-nbitq), 
to_sfixed(687.0/65536.0,1,-nbitq), 
to_sfixed(-585.0/65536.0,1,-nbitq), 
to_sfixed(-2356.0/65536.0,1,-nbitq), 
to_sfixed(-2094.0/65536.0,1,-nbitq), 
to_sfixed(-337.0/65536.0,1,-nbitq), 
to_sfixed(177.0/65536.0,1,-nbitq), 
to_sfixed(-479.0/65536.0,1,-nbitq), 
to_sfixed(-1072.0/65536.0,1,-nbitq), 
to_sfixed(47.0/65536.0,1,-nbitq), 
to_sfixed(2459.0/65536.0,1,-nbitq), 
to_sfixed(341.0/65536.0,1,-nbitq), 
to_sfixed(855.0/65536.0,1,-nbitq), 
to_sfixed(-2544.0/65536.0,1,-nbitq), 
to_sfixed(-1739.0/65536.0,1,-nbitq), 
to_sfixed(1594.0/65536.0,1,-nbitq), 
to_sfixed(-3672.0/65536.0,1,-nbitq), 
to_sfixed(1532.0/65536.0,1,-nbitq), 
to_sfixed(2664.0/65536.0,1,-nbitq), 
to_sfixed(-2243.0/65536.0,1,-nbitq), 
to_sfixed(-3294.0/65536.0,1,-nbitq), 
to_sfixed(1059.0/65536.0,1,-nbitq), 
to_sfixed(1534.0/65536.0,1,-nbitq), 
to_sfixed(294.0/65536.0,1,-nbitq), 
to_sfixed(2485.0/65536.0,1,-nbitq), 
to_sfixed(-3393.0/65536.0,1,-nbitq), 
to_sfixed(3155.0/65536.0,1,-nbitq), 
to_sfixed(1862.0/65536.0,1,-nbitq), 
to_sfixed(3759.0/65536.0,1,-nbitq), 
to_sfixed(750.0/65536.0,1,-nbitq), 
to_sfixed(-1321.0/65536.0,1,-nbitq), 
to_sfixed(1808.0/65536.0,1,-nbitq), 
to_sfixed(1184.0/65536.0,1,-nbitq), 
to_sfixed(-2636.0/65536.0,1,-nbitq), 
to_sfixed(-732.0/65536.0,1,-nbitq), 
to_sfixed(809.0/65536.0,1,-nbitq), 
to_sfixed(-902.0/65536.0,1,-nbitq), 
to_sfixed(-798.0/65536.0,1,-nbitq), 
to_sfixed(-1431.0/65536.0,1,-nbitq), 
to_sfixed(-5065.0/65536.0,1,-nbitq), 
to_sfixed(-3266.0/65536.0,1,-nbitq), 
to_sfixed(-4157.0/65536.0,1,-nbitq), 
to_sfixed(-486.0/65536.0,1,-nbitq), 
to_sfixed(-168.0/65536.0,1,-nbitq), 
to_sfixed(4474.0/65536.0,1,-nbitq), 
to_sfixed(1158.0/65536.0,1,-nbitq), 
to_sfixed(1119.0/65536.0,1,-nbitq), 
to_sfixed(2056.0/65536.0,1,-nbitq), 
to_sfixed(3313.0/65536.0,1,-nbitq), 
to_sfixed(-828.0/65536.0,1,-nbitq), 
to_sfixed(1563.0/65536.0,1,-nbitq), 
to_sfixed(4144.0/65536.0,1,-nbitq), 
to_sfixed(324.0/65536.0,1,-nbitq), 
to_sfixed(1476.0/65536.0,1,-nbitq), 
to_sfixed(-296.0/65536.0,1,-nbitq), 
to_sfixed(903.0/65536.0,1,-nbitq), 
to_sfixed(1059.0/65536.0,1,-nbitq), 
to_sfixed(-2368.0/65536.0,1,-nbitq), 
to_sfixed(5901.0/65536.0,1,-nbitq), 
to_sfixed(2339.0/65536.0,1,-nbitq), 
to_sfixed(1274.0/65536.0,1,-nbitq), 
to_sfixed(-709.0/65536.0,1,-nbitq), 
to_sfixed(904.0/65536.0,1,-nbitq), 
to_sfixed(1492.0/65536.0,1,-nbitq), 
to_sfixed(2954.0/65536.0,1,-nbitq), 
to_sfixed(-802.0/65536.0,1,-nbitq), 
to_sfixed(-2531.0/65536.0,1,-nbitq), 
to_sfixed(-2259.0/65536.0,1,-nbitq), 
to_sfixed(310.0/65536.0,1,-nbitq), 
to_sfixed(2330.0/65536.0,1,-nbitq), 
to_sfixed(-1323.0/65536.0,1,-nbitq), 
to_sfixed(909.0/65536.0,1,-nbitq), 
to_sfixed(1528.0/65536.0,1,-nbitq), 
to_sfixed(431.0/65536.0,1,-nbitq), 
to_sfixed(4260.0/65536.0,1,-nbitq), 
to_sfixed(-1667.0/65536.0,1,-nbitq), 
to_sfixed(3401.0/65536.0,1,-nbitq), 
to_sfixed(-1171.0/65536.0,1,-nbitq), 
to_sfixed(265.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-917.0/65536.0,1,-nbitq), 
to_sfixed(996.0/65536.0,1,-nbitq), 
to_sfixed(1614.0/65536.0,1,-nbitq), 
to_sfixed(-4000.0/65536.0,1,-nbitq), 
to_sfixed(927.0/65536.0,1,-nbitq), 
to_sfixed(-1613.0/65536.0,1,-nbitq), 
to_sfixed(-1831.0/65536.0,1,-nbitq), 
to_sfixed(2131.0/65536.0,1,-nbitq), 
to_sfixed(-3586.0/65536.0,1,-nbitq), 
to_sfixed(-1923.0/65536.0,1,-nbitq), 
to_sfixed(-329.0/65536.0,1,-nbitq), 
to_sfixed(1605.0/65536.0,1,-nbitq), 
to_sfixed(-2085.0/65536.0,1,-nbitq), 
to_sfixed(-3298.0/65536.0,1,-nbitq), 
to_sfixed(-1394.0/65536.0,1,-nbitq), 
to_sfixed(-1627.0/65536.0,1,-nbitq), 
to_sfixed(-774.0/65536.0,1,-nbitq), 
to_sfixed(-98.0/65536.0,1,-nbitq), 
to_sfixed(-1635.0/65536.0,1,-nbitq), 
to_sfixed(2169.0/65536.0,1,-nbitq), 
to_sfixed(-1335.0/65536.0,1,-nbitq), 
to_sfixed(-1289.0/65536.0,1,-nbitq), 
to_sfixed(1641.0/65536.0,1,-nbitq), 
to_sfixed(950.0/65536.0,1,-nbitq), 
to_sfixed(1166.0/65536.0,1,-nbitq), 
to_sfixed(-1872.0/65536.0,1,-nbitq), 
to_sfixed(-3812.0/65536.0,1,-nbitq), 
to_sfixed(2581.0/65536.0,1,-nbitq), 
to_sfixed(-396.0/65536.0,1,-nbitq), 
to_sfixed(-1263.0/65536.0,1,-nbitq), 
to_sfixed(536.0/65536.0,1,-nbitq), 
to_sfixed(2962.0/65536.0,1,-nbitq), 
to_sfixed(-4027.0/65536.0,1,-nbitq), 
to_sfixed(-4872.0/65536.0,1,-nbitq), 
to_sfixed(-266.0/65536.0,1,-nbitq), 
to_sfixed(-3093.0/65536.0,1,-nbitq), 
to_sfixed(50.0/65536.0,1,-nbitq), 
to_sfixed(-357.0/65536.0,1,-nbitq), 
to_sfixed(-2292.0/65536.0,1,-nbitq), 
to_sfixed(2279.0/65536.0,1,-nbitq), 
to_sfixed(-311.0/65536.0,1,-nbitq), 
to_sfixed(91.0/65536.0,1,-nbitq), 
to_sfixed(-3500.0/65536.0,1,-nbitq), 
to_sfixed(-1004.0/65536.0,1,-nbitq), 
to_sfixed(-2336.0/65536.0,1,-nbitq), 
to_sfixed(1179.0/65536.0,1,-nbitq), 
to_sfixed(-145.0/65536.0,1,-nbitq), 
to_sfixed(298.0/65536.0,1,-nbitq), 
to_sfixed(3497.0/65536.0,1,-nbitq), 
to_sfixed(332.0/65536.0,1,-nbitq), 
to_sfixed(3355.0/65536.0,1,-nbitq), 
to_sfixed(484.0/65536.0,1,-nbitq), 
to_sfixed(892.0/65536.0,1,-nbitq), 
to_sfixed(1235.0/65536.0,1,-nbitq), 
to_sfixed(4066.0/65536.0,1,-nbitq), 
to_sfixed(495.0/65536.0,1,-nbitq), 
to_sfixed(-838.0/65536.0,1,-nbitq), 
to_sfixed(271.0/65536.0,1,-nbitq), 
to_sfixed(304.0/65536.0,1,-nbitq), 
to_sfixed(5794.0/65536.0,1,-nbitq), 
to_sfixed(1707.0/65536.0,1,-nbitq), 
to_sfixed(2607.0/65536.0,1,-nbitq), 
to_sfixed(-203.0/65536.0,1,-nbitq), 
to_sfixed(1608.0/65536.0,1,-nbitq), 
to_sfixed(547.0/65536.0,1,-nbitq), 
to_sfixed(1472.0/65536.0,1,-nbitq), 
to_sfixed(-87.0/65536.0,1,-nbitq), 
to_sfixed(-1091.0/65536.0,1,-nbitq), 
to_sfixed(-2135.0/65536.0,1,-nbitq), 
to_sfixed(-422.0/65536.0,1,-nbitq), 
to_sfixed(556.0/65536.0,1,-nbitq), 
to_sfixed(-2202.0/65536.0,1,-nbitq), 
to_sfixed(94.0/65536.0,1,-nbitq), 
to_sfixed(-1185.0/65536.0,1,-nbitq), 
to_sfixed(2358.0/65536.0,1,-nbitq), 
to_sfixed(2023.0/65536.0,1,-nbitq), 
to_sfixed(-2617.0/65536.0,1,-nbitq), 
to_sfixed(-858.0/65536.0,1,-nbitq), 
to_sfixed(1990.0/65536.0,1,-nbitq), 
to_sfixed(4754.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3015.0/65536.0,1,-nbitq), 
to_sfixed(-482.0/65536.0,1,-nbitq), 
to_sfixed(1208.0/65536.0,1,-nbitq), 
to_sfixed(-109.0/65536.0,1,-nbitq), 
to_sfixed(-2256.0/65536.0,1,-nbitq), 
to_sfixed(398.0/65536.0,1,-nbitq), 
to_sfixed(-41.0/65536.0,1,-nbitq), 
to_sfixed(352.0/65536.0,1,-nbitq), 
to_sfixed(-2663.0/65536.0,1,-nbitq), 
to_sfixed(-301.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(380.0/65536.0,1,-nbitq), 
to_sfixed(2480.0/65536.0,1,-nbitq), 
to_sfixed(-988.0/65536.0,1,-nbitq), 
to_sfixed(648.0/65536.0,1,-nbitq), 
to_sfixed(-1734.0/65536.0,1,-nbitq), 
to_sfixed(2758.0/65536.0,1,-nbitq), 
to_sfixed(1078.0/65536.0,1,-nbitq), 
to_sfixed(4287.0/65536.0,1,-nbitq), 
to_sfixed(-245.0/65536.0,1,-nbitq), 
to_sfixed(-4187.0/65536.0,1,-nbitq), 
to_sfixed(-617.0/65536.0,1,-nbitq), 
to_sfixed(1260.0/65536.0,1,-nbitq), 
to_sfixed(-436.0/65536.0,1,-nbitq), 
to_sfixed(1947.0/65536.0,1,-nbitq), 
to_sfixed(-520.0/65536.0,1,-nbitq), 
to_sfixed(-2380.0/65536.0,1,-nbitq), 
to_sfixed(-2220.0/65536.0,1,-nbitq), 
to_sfixed(-308.0/65536.0,1,-nbitq), 
to_sfixed(-2182.0/65536.0,1,-nbitq), 
to_sfixed(2205.0/65536.0,1,-nbitq), 
to_sfixed(2599.0/65536.0,1,-nbitq), 
to_sfixed(-1631.0/65536.0,1,-nbitq), 
to_sfixed(-1964.0/65536.0,1,-nbitq), 
to_sfixed(505.0/65536.0,1,-nbitq), 
to_sfixed(-84.0/65536.0,1,-nbitq), 
to_sfixed(-817.0/65536.0,1,-nbitq), 
to_sfixed(-1475.0/65536.0,1,-nbitq), 
to_sfixed(-89.0/65536.0,1,-nbitq), 
to_sfixed(-2018.0/65536.0,1,-nbitq), 
to_sfixed(-3030.0/65536.0,1,-nbitq), 
to_sfixed(-3190.0/65536.0,1,-nbitq), 
to_sfixed(245.0/65536.0,1,-nbitq), 
to_sfixed(-264.0/65536.0,1,-nbitq), 
to_sfixed(-1495.0/65536.0,1,-nbitq), 
to_sfixed(4728.0/65536.0,1,-nbitq), 
to_sfixed(-2028.0/65536.0,1,-nbitq), 
to_sfixed(1412.0/65536.0,1,-nbitq), 
to_sfixed(3357.0/65536.0,1,-nbitq), 
to_sfixed(-1120.0/65536.0,1,-nbitq), 
to_sfixed(651.0/65536.0,1,-nbitq), 
to_sfixed(1064.0/65536.0,1,-nbitq), 
to_sfixed(2022.0/65536.0,1,-nbitq), 
to_sfixed(-298.0/65536.0,1,-nbitq), 
to_sfixed(3764.0/65536.0,1,-nbitq), 
to_sfixed(2824.0/65536.0,1,-nbitq), 
to_sfixed(909.0/65536.0,1,-nbitq), 
to_sfixed(2916.0/65536.0,1,-nbitq), 
to_sfixed(1047.0/65536.0,1,-nbitq), 
to_sfixed(-29.0/65536.0,1,-nbitq), 
to_sfixed(-3144.0/65536.0,1,-nbitq), 
to_sfixed(-525.0/65536.0,1,-nbitq), 
to_sfixed(-2621.0/65536.0,1,-nbitq), 
to_sfixed(-2551.0/65536.0,1,-nbitq), 
to_sfixed(1735.0/65536.0,1,-nbitq), 
to_sfixed(1582.0/65536.0,1,-nbitq), 
to_sfixed(401.0/65536.0,1,-nbitq), 
to_sfixed(245.0/65536.0,1,-nbitq), 
to_sfixed(-698.0/65536.0,1,-nbitq), 
to_sfixed(-693.0/65536.0,1,-nbitq), 
to_sfixed(1584.0/65536.0,1,-nbitq), 
to_sfixed(-2492.0/65536.0,1,-nbitq), 
to_sfixed(933.0/65536.0,1,-nbitq), 
to_sfixed(-957.0/65536.0,1,-nbitq), 
to_sfixed(1090.0/65536.0,1,-nbitq), 
to_sfixed(884.0/65536.0,1,-nbitq), 
to_sfixed(-879.0/65536.0,1,-nbitq), 
to_sfixed(3336.0/65536.0,1,-nbitq), 
to_sfixed(-3134.0/65536.0,1,-nbitq), 
to_sfixed(1371.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-737.0/65536.0,1,-nbitq), 
to_sfixed(1484.0/65536.0,1,-nbitq), 
to_sfixed(574.0/65536.0,1,-nbitq), 
to_sfixed(1847.0/65536.0,1,-nbitq), 
to_sfixed(-1398.0/65536.0,1,-nbitq), 
to_sfixed(-4849.0/65536.0,1,-nbitq), 
to_sfixed(-808.0/65536.0,1,-nbitq), 
to_sfixed(735.0/65536.0,1,-nbitq), 
to_sfixed(-2713.0/65536.0,1,-nbitq), 
to_sfixed(-1530.0/65536.0,1,-nbitq), 
to_sfixed(1204.0/65536.0,1,-nbitq), 
to_sfixed(-1603.0/65536.0,1,-nbitq), 
to_sfixed(-1817.0/65536.0,1,-nbitq), 
to_sfixed(17.0/65536.0,1,-nbitq), 
to_sfixed(1249.0/65536.0,1,-nbitq), 
to_sfixed(2633.0/65536.0,1,-nbitq), 
to_sfixed(756.0/65536.0,1,-nbitq), 
to_sfixed(1146.0/65536.0,1,-nbitq), 
to_sfixed(-996.0/65536.0,1,-nbitq), 
to_sfixed(-1756.0/65536.0,1,-nbitq), 
to_sfixed(-3790.0/65536.0,1,-nbitq), 
to_sfixed(2318.0/65536.0,1,-nbitq), 
to_sfixed(1187.0/65536.0,1,-nbitq), 
to_sfixed(1829.0/65536.0,1,-nbitq), 
to_sfixed(454.0/65536.0,1,-nbitq), 
to_sfixed(-780.0/65536.0,1,-nbitq), 
to_sfixed(1265.0/65536.0,1,-nbitq), 
to_sfixed(557.0/65536.0,1,-nbitq), 
to_sfixed(-836.0/65536.0,1,-nbitq), 
to_sfixed(-3022.0/65536.0,1,-nbitq), 
to_sfixed(2555.0/65536.0,1,-nbitq), 
to_sfixed(-2667.0/65536.0,1,-nbitq), 
to_sfixed(-4884.0/65536.0,1,-nbitq), 
to_sfixed(-1852.0/65536.0,1,-nbitq), 
to_sfixed(-2473.0/65536.0,1,-nbitq), 
to_sfixed(-2054.0/65536.0,1,-nbitq), 
to_sfixed(-2989.0/65536.0,1,-nbitq), 
to_sfixed(955.0/65536.0,1,-nbitq), 
to_sfixed(461.0/65536.0,1,-nbitq), 
to_sfixed(2154.0/65536.0,1,-nbitq), 
to_sfixed(-1172.0/65536.0,1,-nbitq), 
to_sfixed(889.0/65536.0,1,-nbitq), 
to_sfixed(-3648.0/65536.0,1,-nbitq), 
to_sfixed(2369.0/65536.0,1,-nbitq), 
to_sfixed(2626.0/65536.0,1,-nbitq), 
to_sfixed(3603.0/65536.0,1,-nbitq), 
to_sfixed(-398.0/65536.0,1,-nbitq), 
to_sfixed(105.0/65536.0,1,-nbitq), 
to_sfixed(-2219.0/65536.0,1,-nbitq), 
to_sfixed(-929.0/65536.0,1,-nbitq), 
to_sfixed(-1946.0/65536.0,1,-nbitq), 
to_sfixed(1302.0/65536.0,1,-nbitq), 
to_sfixed(1849.0/65536.0,1,-nbitq), 
to_sfixed(-2323.0/65536.0,1,-nbitq), 
to_sfixed(-1560.0/65536.0,1,-nbitq), 
to_sfixed(653.0/65536.0,1,-nbitq), 
to_sfixed(685.0/65536.0,1,-nbitq), 
to_sfixed(3146.0/65536.0,1,-nbitq), 
to_sfixed(-2636.0/65536.0,1,-nbitq), 
to_sfixed(1232.0/65536.0,1,-nbitq), 
to_sfixed(1320.0/65536.0,1,-nbitq), 
to_sfixed(2553.0/65536.0,1,-nbitq), 
to_sfixed(1110.0/65536.0,1,-nbitq), 
to_sfixed(-841.0/65536.0,1,-nbitq), 
to_sfixed(2697.0/65536.0,1,-nbitq), 
to_sfixed(252.0/65536.0,1,-nbitq), 
to_sfixed(-985.0/65536.0,1,-nbitq), 
to_sfixed(-3528.0/65536.0,1,-nbitq), 
to_sfixed(3701.0/65536.0,1,-nbitq), 
to_sfixed(-827.0/65536.0,1,-nbitq), 
to_sfixed(951.0/65536.0,1,-nbitq), 
to_sfixed(-715.0/65536.0,1,-nbitq), 
to_sfixed(1954.0/65536.0,1,-nbitq), 
to_sfixed(-156.0/65536.0,1,-nbitq), 
to_sfixed(-502.0/65536.0,1,-nbitq), 
to_sfixed(-1445.0/65536.0,1,-nbitq), 
to_sfixed(2072.0/65536.0,1,-nbitq), 
to_sfixed(1985.0/65536.0,1,-nbitq), 
to_sfixed(-2898.0/65536.0,1,-nbitq), 
to_sfixed(2732.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2852.0/65536.0,1,-nbitq), 
to_sfixed(-2302.0/65536.0,1,-nbitq), 
to_sfixed(1743.0/65536.0,1,-nbitq), 
to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(794.0/65536.0,1,-nbitq), 
to_sfixed(635.0/65536.0,1,-nbitq), 
to_sfixed(-2106.0/65536.0,1,-nbitq), 
to_sfixed(-601.0/65536.0,1,-nbitq), 
to_sfixed(-2363.0/65536.0,1,-nbitq), 
to_sfixed(-1505.0/65536.0,1,-nbitq), 
to_sfixed(-1754.0/65536.0,1,-nbitq), 
to_sfixed(-2475.0/65536.0,1,-nbitq), 
to_sfixed(317.0/65536.0,1,-nbitq), 
to_sfixed(-413.0/65536.0,1,-nbitq), 
to_sfixed(-687.0/65536.0,1,-nbitq), 
to_sfixed(-1449.0/65536.0,1,-nbitq), 
to_sfixed(-503.0/65536.0,1,-nbitq), 
to_sfixed(-1325.0/65536.0,1,-nbitq), 
to_sfixed(1071.0/65536.0,1,-nbitq), 
to_sfixed(1213.0/65536.0,1,-nbitq), 
to_sfixed(-3401.0/65536.0,1,-nbitq), 
to_sfixed(2689.0/65536.0,1,-nbitq), 
to_sfixed(-469.0/65536.0,1,-nbitq), 
to_sfixed(3894.0/65536.0,1,-nbitq), 
to_sfixed(1208.0/65536.0,1,-nbitq), 
to_sfixed(3997.0/65536.0,1,-nbitq), 
to_sfixed(1203.0/65536.0,1,-nbitq), 
to_sfixed(-1148.0/65536.0,1,-nbitq), 
to_sfixed(-2367.0/65536.0,1,-nbitq), 
to_sfixed(937.0/65536.0,1,-nbitq), 
to_sfixed(1066.0/65536.0,1,-nbitq), 
to_sfixed(-2440.0/65536.0,1,-nbitq), 
to_sfixed(-4142.0/65536.0,1,-nbitq), 
to_sfixed(-5434.0/65536.0,1,-nbitq), 
to_sfixed(-1651.0/65536.0,1,-nbitq), 
to_sfixed(-1765.0/65536.0,1,-nbitq), 
to_sfixed(2356.0/65536.0,1,-nbitq), 
to_sfixed(-3903.0/65536.0,1,-nbitq), 
to_sfixed(613.0/65536.0,1,-nbitq), 
to_sfixed(2149.0/65536.0,1,-nbitq), 
to_sfixed(-2119.0/65536.0,1,-nbitq), 
to_sfixed(-1177.0/65536.0,1,-nbitq), 
to_sfixed(-2594.0/65536.0,1,-nbitq), 
to_sfixed(3031.0/65536.0,1,-nbitq), 
to_sfixed(1323.0/65536.0,1,-nbitq), 
to_sfixed(775.0/65536.0,1,-nbitq), 
to_sfixed(2121.0/65536.0,1,-nbitq), 
to_sfixed(2663.0/65536.0,1,-nbitq), 
to_sfixed(-1608.0/65536.0,1,-nbitq), 
to_sfixed(-655.0/65536.0,1,-nbitq), 
to_sfixed(1533.0/65536.0,1,-nbitq), 
to_sfixed(-2500.0/65536.0,1,-nbitq), 
to_sfixed(-457.0/65536.0,1,-nbitq), 
to_sfixed(-1755.0/65536.0,1,-nbitq), 
to_sfixed(975.0/65536.0,1,-nbitq), 
to_sfixed(2884.0/65536.0,1,-nbitq), 
to_sfixed(173.0/65536.0,1,-nbitq), 
to_sfixed(1730.0/65536.0,1,-nbitq), 
to_sfixed(1601.0/65536.0,1,-nbitq), 
to_sfixed(652.0/65536.0,1,-nbitq), 
to_sfixed(-2183.0/65536.0,1,-nbitq), 
to_sfixed(2287.0/65536.0,1,-nbitq), 
to_sfixed(1547.0/65536.0,1,-nbitq), 
to_sfixed(1862.0/65536.0,1,-nbitq), 
to_sfixed(-1824.0/65536.0,1,-nbitq), 
to_sfixed(-81.0/65536.0,1,-nbitq), 
to_sfixed(-1382.0/65536.0,1,-nbitq), 
to_sfixed(-1626.0/65536.0,1,-nbitq), 
to_sfixed(-1046.0/65536.0,1,-nbitq), 
to_sfixed(-1716.0/65536.0,1,-nbitq), 
to_sfixed(2089.0/65536.0,1,-nbitq), 
to_sfixed(155.0/65536.0,1,-nbitq), 
to_sfixed(4158.0/65536.0,1,-nbitq), 
to_sfixed(2117.0/65536.0,1,-nbitq), 
to_sfixed(-1183.0/65536.0,1,-nbitq), 
to_sfixed(680.0/65536.0,1,-nbitq), 
to_sfixed(2366.0/65536.0,1,-nbitq), 
to_sfixed(653.0/65536.0,1,-nbitq), 
to_sfixed(988.0/65536.0,1,-nbitq), 
to_sfixed(1123.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1102.0/65536.0,1,-nbitq), 
to_sfixed(-689.0/65536.0,1,-nbitq), 
to_sfixed(3129.0/65536.0,1,-nbitq), 
to_sfixed(-3763.0/65536.0,1,-nbitq), 
to_sfixed(274.0/65536.0,1,-nbitq), 
to_sfixed(-2201.0/65536.0,1,-nbitq), 
to_sfixed(-316.0/65536.0,1,-nbitq), 
to_sfixed(1635.0/65536.0,1,-nbitq), 
to_sfixed(2685.0/65536.0,1,-nbitq), 
to_sfixed(46.0/65536.0,1,-nbitq), 
to_sfixed(-329.0/65536.0,1,-nbitq), 
to_sfixed(-1133.0/65536.0,1,-nbitq), 
to_sfixed(-544.0/65536.0,1,-nbitq), 
to_sfixed(-1806.0/65536.0,1,-nbitq), 
to_sfixed(1172.0/65536.0,1,-nbitq), 
to_sfixed(1166.0/65536.0,1,-nbitq), 
to_sfixed(-30.0/65536.0,1,-nbitq), 
to_sfixed(602.0/65536.0,1,-nbitq), 
to_sfixed(1519.0/65536.0,1,-nbitq), 
to_sfixed(386.0/65536.0,1,-nbitq), 
to_sfixed(1696.0/65536.0,1,-nbitq), 
to_sfixed(2723.0/65536.0,1,-nbitq), 
to_sfixed(-980.0/65536.0,1,-nbitq), 
to_sfixed(3187.0/65536.0,1,-nbitq), 
to_sfixed(2586.0/65536.0,1,-nbitq), 
to_sfixed(-1239.0/65536.0,1,-nbitq), 
to_sfixed(1547.0/65536.0,1,-nbitq), 
to_sfixed(1850.0/65536.0,1,-nbitq), 
to_sfixed(-880.0/65536.0,1,-nbitq), 
to_sfixed(346.0/65536.0,1,-nbitq), 
to_sfixed(-2315.0/65536.0,1,-nbitq), 
to_sfixed(-2540.0/65536.0,1,-nbitq), 
to_sfixed(-1057.0/65536.0,1,-nbitq), 
to_sfixed(-2326.0/65536.0,1,-nbitq), 
to_sfixed(2205.0/65536.0,1,-nbitq), 
to_sfixed(-2379.0/65536.0,1,-nbitq), 
to_sfixed(-2868.0/65536.0,1,-nbitq), 
to_sfixed(-3250.0/65536.0,1,-nbitq), 
to_sfixed(-2954.0/65536.0,1,-nbitq), 
to_sfixed(719.0/65536.0,1,-nbitq), 
to_sfixed(1098.0/65536.0,1,-nbitq), 
to_sfixed(-3079.0/65536.0,1,-nbitq), 
to_sfixed(-3283.0/65536.0,1,-nbitq), 
to_sfixed(1029.0/65536.0,1,-nbitq), 
to_sfixed(628.0/65536.0,1,-nbitq), 
to_sfixed(5313.0/65536.0,1,-nbitq), 
to_sfixed(3115.0/65536.0,1,-nbitq), 
to_sfixed(-1487.0/65536.0,1,-nbitq), 
to_sfixed(-545.0/65536.0,1,-nbitq), 
to_sfixed(665.0/65536.0,1,-nbitq), 
to_sfixed(1184.0/65536.0,1,-nbitq), 
to_sfixed(-1310.0/65536.0,1,-nbitq), 
to_sfixed(186.0/65536.0,1,-nbitq), 
to_sfixed(-1475.0/65536.0,1,-nbitq), 
to_sfixed(-1636.0/65536.0,1,-nbitq), 
to_sfixed(-368.0/65536.0,1,-nbitq), 
to_sfixed(827.0/65536.0,1,-nbitq), 
to_sfixed(1478.0/65536.0,1,-nbitq), 
to_sfixed(-1941.0/65536.0,1,-nbitq), 
to_sfixed(4347.0/65536.0,1,-nbitq), 
to_sfixed(-2256.0/65536.0,1,-nbitq), 
to_sfixed(-240.0/65536.0,1,-nbitq), 
to_sfixed(-1990.0/65536.0,1,-nbitq), 
to_sfixed(-549.0/65536.0,1,-nbitq), 
to_sfixed(3476.0/65536.0,1,-nbitq), 
to_sfixed(-689.0/65536.0,1,-nbitq), 
to_sfixed(159.0/65536.0,1,-nbitq), 
to_sfixed(-906.0/65536.0,1,-nbitq), 
to_sfixed(-124.0/65536.0,1,-nbitq), 
to_sfixed(-512.0/65536.0,1,-nbitq), 
to_sfixed(2320.0/65536.0,1,-nbitq), 
to_sfixed(515.0/65536.0,1,-nbitq), 
to_sfixed(4190.0/65536.0,1,-nbitq), 
to_sfixed(2513.0/65536.0,1,-nbitq), 
to_sfixed(-2515.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(2156.0/65536.0,1,-nbitq), 
to_sfixed(4674.0/65536.0,1,-nbitq), 
to_sfixed(-334.0/65536.0,1,-nbitq), 
to_sfixed(640.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2387.0/65536.0,1,-nbitq), 
to_sfixed(-1221.0/65536.0,1,-nbitq), 
to_sfixed(1339.0/65536.0,1,-nbitq), 
to_sfixed(-2275.0/65536.0,1,-nbitq), 
to_sfixed(-2061.0/65536.0,1,-nbitq), 
to_sfixed(-1942.0/65536.0,1,-nbitq), 
to_sfixed(-818.0/65536.0,1,-nbitq), 
to_sfixed(-1322.0/65536.0,1,-nbitq), 
to_sfixed(2322.0/65536.0,1,-nbitq), 
to_sfixed(-257.0/65536.0,1,-nbitq), 
to_sfixed(-240.0/65536.0,1,-nbitq), 
to_sfixed(-3357.0/65536.0,1,-nbitq), 
to_sfixed(-2847.0/65536.0,1,-nbitq), 
to_sfixed(441.0/65536.0,1,-nbitq), 
to_sfixed(2672.0/65536.0,1,-nbitq), 
to_sfixed(-888.0/65536.0,1,-nbitq), 
to_sfixed(1673.0/65536.0,1,-nbitq), 
to_sfixed(5.0/65536.0,1,-nbitq), 
to_sfixed(677.0/65536.0,1,-nbitq), 
to_sfixed(3215.0/65536.0,1,-nbitq), 
to_sfixed(-819.0/65536.0,1,-nbitq), 
to_sfixed(-2466.0/65536.0,1,-nbitq), 
to_sfixed(3683.0/65536.0,1,-nbitq), 
to_sfixed(3871.0/65536.0,1,-nbitq), 
to_sfixed(1348.0/65536.0,1,-nbitq), 
to_sfixed(-2694.0/65536.0,1,-nbitq), 
to_sfixed(1037.0/65536.0,1,-nbitq), 
to_sfixed(1655.0/65536.0,1,-nbitq), 
to_sfixed(-1198.0/65536.0,1,-nbitq), 
to_sfixed(-2274.0/65536.0,1,-nbitq), 
to_sfixed(-1677.0/65536.0,1,-nbitq), 
to_sfixed(-1058.0/65536.0,1,-nbitq), 
to_sfixed(-3627.0/65536.0,1,-nbitq), 
to_sfixed(-4328.0/65536.0,1,-nbitq), 
to_sfixed(-1383.0/65536.0,1,-nbitq), 
to_sfixed(-1879.0/65536.0,1,-nbitq), 
to_sfixed(-2729.0/65536.0,1,-nbitq), 
to_sfixed(-4270.0/65536.0,1,-nbitq), 
to_sfixed(-3437.0/65536.0,1,-nbitq), 
to_sfixed(2858.0/65536.0,1,-nbitq), 
to_sfixed(-379.0/65536.0,1,-nbitq), 
to_sfixed(714.0/65536.0,1,-nbitq), 
to_sfixed(738.0/65536.0,1,-nbitq), 
to_sfixed(1513.0/65536.0,1,-nbitq), 
to_sfixed(845.0/65536.0,1,-nbitq), 
to_sfixed(1058.0/65536.0,1,-nbitq), 
to_sfixed(-1378.0/65536.0,1,-nbitq), 
to_sfixed(-298.0/65536.0,1,-nbitq), 
to_sfixed(36.0/65536.0,1,-nbitq), 
to_sfixed(354.0/65536.0,1,-nbitq), 
to_sfixed(-2523.0/65536.0,1,-nbitq), 
to_sfixed(3628.0/65536.0,1,-nbitq), 
to_sfixed(944.0/65536.0,1,-nbitq), 
to_sfixed(20.0/65536.0,1,-nbitq), 
to_sfixed(264.0/65536.0,1,-nbitq), 
to_sfixed(-517.0/65536.0,1,-nbitq), 
to_sfixed(2536.0/65536.0,1,-nbitq), 
to_sfixed(1356.0/65536.0,1,-nbitq), 
to_sfixed(-2876.0/65536.0,1,-nbitq), 
to_sfixed(3092.0/65536.0,1,-nbitq), 
to_sfixed(2253.0/65536.0,1,-nbitq), 
to_sfixed(-2253.0/65536.0,1,-nbitq), 
to_sfixed(1088.0/65536.0,1,-nbitq), 
to_sfixed(-850.0/65536.0,1,-nbitq), 
to_sfixed(228.0/65536.0,1,-nbitq), 
to_sfixed(2924.0/65536.0,1,-nbitq), 
to_sfixed(437.0/65536.0,1,-nbitq), 
to_sfixed(-55.0/65536.0,1,-nbitq), 
to_sfixed(-1242.0/65536.0,1,-nbitq), 
to_sfixed(1696.0/65536.0,1,-nbitq), 
to_sfixed(-1599.0/65536.0,1,-nbitq), 
to_sfixed(-39.0/65536.0,1,-nbitq), 
to_sfixed(1817.0/65536.0,1,-nbitq), 
to_sfixed(-1913.0/65536.0,1,-nbitq), 
to_sfixed(-186.0/65536.0,1,-nbitq), 
to_sfixed(1482.0/65536.0,1,-nbitq), 
to_sfixed(-2426.0/65536.0,1,-nbitq), 
to_sfixed(1136.0/65536.0,1,-nbitq), 
to_sfixed(1031.0/65536.0,1,-nbitq), 
to_sfixed(1748.0/65536.0,1,-nbitq)  ), 
( to_sfixed(379.0/65536.0,1,-nbitq), 
to_sfixed(1984.0/65536.0,1,-nbitq), 
to_sfixed(-2121.0/65536.0,1,-nbitq), 
to_sfixed(180.0/65536.0,1,-nbitq), 
to_sfixed(3558.0/65536.0,1,-nbitq), 
to_sfixed(-1839.0/65536.0,1,-nbitq), 
to_sfixed(-1227.0/65536.0,1,-nbitq), 
to_sfixed(-3987.0/65536.0,1,-nbitq), 
to_sfixed(3837.0/65536.0,1,-nbitq), 
to_sfixed(-759.0/65536.0,1,-nbitq), 
to_sfixed(-2796.0/65536.0,1,-nbitq), 
to_sfixed(4718.0/65536.0,1,-nbitq), 
to_sfixed(-24.0/65536.0,1,-nbitq), 
to_sfixed(-911.0/65536.0,1,-nbitq), 
to_sfixed(2468.0/65536.0,1,-nbitq), 
to_sfixed(-1953.0/65536.0,1,-nbitq), 
to_sfixed(-1065.0/65536.0,1,-nbitq), 
to_sfixed(-139.0/65536.0,1,-nbitq), 
to_sfixed(3808.0/65536.0,1,-nbitq), 
to_sfixed(3038.0/65536.0,1,-nbitq), 
to_sfixed(40.0/65536.0,1,-nbitq), 
to_sfixed(-631.0/65536.0,1,-nbitq), 
to_sfixed(1123.0/65536.0,1,-nbitq), 
to_sfixed(3566.0/65536.0,1,-nbitq), 
to_sfixed(-1182.0/65536.0,1,-nbitq), 
to_sfixed(-1169.0/65536.0,1,-nbitq), 
to_sfixed(-2132.0/65536.0,1,-nbitq), 
to_sfixed(-524.0/65536.0,1,-nbitq), 
to_sfixed(-4837.0/65536.0,1,-nbitq), 
to_sfixed(-1151.0/65536.0,1,-nbitq), 
to_sfixed(2519.0/65536.0,1,-nbitq), 
to_sfixed(-1613.0/65536.0,1,-nbitq), 
to_sfixed(-4402.0/65536.0,1,-nbitq), 
to_sfixed(2135.0/65536.0,1,-nbitq), 
to_sfixed(-2366.0/65536.0,1,-nbitq), 
to_sfixed(-1362.0/65536.0,1,-nbitq), 
to_sfixed(-2807.0/65536.0,1,-nbitq), 
to_sfixed(-1636.0/65536.0,1,-nbitq), 
to_sfixed(-676.0/65536.0,1,-nbitq), 
to_sfixed(455.0/65536.0,1,-nbitq), 
to_sfixed(-1087.0/65536.0,1,-nbitq), 
to_sfixed(2034.0/65536.0,1,-nbitq), 
to_sfixed(-3619.0/65536.0,1,-nbitq), 
to_sfixed(-3003.0/65536.0,1,-nbitq), 
to_sfixed(3316.0/65536.0,1,-nbitq), 
to_sfixed(2352.0/65536.0,1,-nbitq), 
to_sfixed(-1314.0/65536.0,1,-nbitq), 
to_sfixed(967.0/65536.0,1,-nbitq), 
to_sfixed(-1900.0/65536.0,1,-nbitq), 
to_sfixed(4568.0/65536.0,1,-nbitq), 
to_sfixed(1728.0/65536.0,1,-nbitq), 
to_sfixed(1608.0/65536.0,1,-nbitq), 
to_sfixed(691.0/65536.0,1,-nbitq), 
to_sfixed(213.0/65536.0,1,-nbitq), 
to_sfixed(396.0/65536.0,1,-nbitq), 
to_sfixed(-113.0/65536.0,1,-nbitq), 
to_sfixed(2842.0/65536.0,1,-nbitq), 
to_sfixed(-2855.0/65536.0,1,-nbitq), 
to_sfixed(-1398.0/65536.0,1,-nbitq), 
to_sfixed(3185.0/65536.0,1,-nbitq), 
to_sfixed(-610.0/65536.0,1,-nbitq), 
to_sfixed(1197.0/65536.0,1,-nbitq), 
to_sfixed(-2044.0/65536.0,1,-nbitq), 
to_sfixed(2624.0/65536.0,1,-nbitq), 
to_sfixed(1877.0/65536.0,1,-nbitq), 
to_sfixed(255.0/65536.0,1,-nbitq), 
to_sfixed(-49.0/65536.0,1,-nbitq), 
to_sfixed(-1056.0/65536.0,1,-nbitq), 
to_sfixed(-2257.0/65536.0,1,-nbitq), 
to_sfixed(4118.0/65536.0,1,-nbitq), 
to_sfixed(1080.0/65536.0,1,-nbitq), 
to_sfixed(-30.0/65536.0,1,-nbitq), 
to_sfixed(1883.0/65536.0,1,-nbitq), 
to_sfixed(1416.0/65536.0,1,-nbitq), 
to_sfixed(-2661.0/65536.0,1,-nbitq), 
to_sfixed(1548.0/65536.0,1,-nbitq), 
to_sfixed(2447.0/65536.0,1,-nbitq), 
to_sfixed(1639.0/65536.0,1,-nbitq), 
to_sfixed(308.0/65536.0,1,-nbitq), 
to_sfixed(-1585.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-994.0/65536.0,1,-nbitq), 
to_sfixed(-2343.0/65536.0,1,-nbitq), 
to_sfixed(-5535.0/65536.0,1,-nbitq), 
to_sfixed(-2374.0/65536.0,1,-nbitq), 
to_sfixed(2395.0/65536.0,1,-nbitq), 
to_sfixed(-1128.0/65536.0,1,-nbitq), 
to_sfixed(3781.0/65536.0,1,-nbitq), 
to_sfixed(-1291.0/65536.0,1,-nbitq), 
to_sfixed(1494.0/65536.0,1,-nbitq), 
to_sfixed(2804.0/65536.0,1,-nbitq), 
to_sfixed(1240.0/65536.0,1,-nbitq), 
to_sfixed(7664.0/65536.0,1,-nbitq), 
to_sfixed(2655.0/65536.0,1,-nbitq), 
to_sfixed(3690.0/65536.0,1,-nbitq), 
to_sfixed(1482.0/65536.0,1,-nbitq), 
to_sfixed(2158.0/65536.0,1,-nbitq), 
to_sfixed(-1257.0/65536.0,1,-nbitq), 
to_sfixed(3128.0/65536.0,1,-nbitq), 
to_sfixed(1133.0/65536.0,1,-nbitq), 
to_sfixed(-1014.0/65536.0,1,-nbitq), 
to_sfixed(-2518.0/65536.0,1,-nbitq), 
to_sfixed(-1905.0/65536.0,1,-nbitq), 
to_sfixed(2912.0/65536.0,1,-nbitq), 
to_sfixed(845.0/65536.0,1,-nbitq), 
to_sfixed(1222.0/65536.0,1,-nbitq), 
to_sfixed(-530.0/65536.0,1,-nbitq), 
to_sfixed(-4381.0/65536.0,1,-nbitq), 
to_sfixed(-950.0/65536.0,1,-nbitq), 
to_sfixed(-6910.0/65536.0,1,-nbitq), 
to_sfixed(239.0/65536.0,1,-nbitq), 
to_sfixed(-1846.0/65536.0,1,-nbitq), 
to_sfixed(-71.0/65536.0,1,-nbitq), 
to_sfixed(-2032.0/65536.0,1,-nbitq), 
to_sfixed(1489.0/65536.0,1,-nbitq), 
to_sfixed(-3628.0/65536.0,1,-nbitq), 
to_sfixed(2588.0/65536.0,1,-nbitq), 
to_sfixed(-143.0/65536.0,1,-nbitq), 
to_sfixed(3382.0/65536.0,1,-nbitq), 
to_sfixed(4761.0/65536.0,1,-nbitq), 
to_sfixed(-2470.0/65536.0,1,-nbitq), 
to_sfixed(-4870.0/65536.0,1,-nbitq), 
to_sfixed(1865.0/65536.0,1,-nbitq), 
to_sfixed(-6398.0/65536.0,1,-nbitq), 
to_sfixed(1749.0/65536.0,1,-nbitq), 
to_sfixed(-126.0/65536.0,1,-nbitq), 
to_sfixed(-5506.0/65536.0,1,-nbitq), 
to_sfixed(-3088.0/65536.0,1,-nbitq), 
to_sfixed(2904.0/65536.0,1,-nbitq), 
to_sfixed(323.0/65536.0,1,-nbitq), 
to_sfixed(3799.0/65536.0,1,-nbitq), 
to_sfixed(2544.0/65536.0,1,-nbitq), 
to_sfixed(-2573.0/65536.0,1,-nbitq), 
to_sfixed(-113.0/65536.0,1,-nbitq), 
to_sfixed(17.0/65536.0,1,-nbitq), 
to_sfixed(-1147.0/65536.0,1,-nbitq), 
to_sfixed(-5089.0/65536.0,1,-nbitq), 
to_sfixed(3675.0/65536.0,1,-nbitq), 
to_sfixed(-2574.0/65536.0,1,-nbitq), 
to_sfixed(-2371.0/65536.0,1,-nbitq), 
to_sfixed(2349.0/65536.0,1,-nbitq), 
to_sfixed(1164.0/65536.0,1,-nbitq), 
to_sfixed(2178.0/65536.0,1,-nbitq), 
to_sfixed(1009.0/65536.0,1,-nbitq), 
to_sfixed(-163.0/65536.0,1,-nbitq), 
to_sfixed(4718.0/65536.0,1,-nbitq), 
to_sfixed(-2995.0/65536.0,1,-nbitq), 
to_sfixed(621.0/65536.0,1,-nbitq), 
to_sfixed(1684.0/65536.0,1,-nbitq), 
to_sfixed(-691.0/65536.0,1,-nbitq), 
to_sfixed(6633.0/65536.0,1,-nbitq), 
to_sfixed(-393.0/65536.0,1,-nbitq), 
to_sfixed(3473.0/65536.0,1,-nbitq), 
to_sfixed(202.0/65536.0,1,-nbitq), 
to_sfixed(1883.0/65536.0,1,-nbitq), 
to_sfixed(1710.0/65536.0,1,-nbitq), 
to_sfixed(2034.0/65536.0,1,-nbitq), 
to_sfixed(7408.0/65536.0,1,-nbitq), 
to_sfixed(-1897.0/65536.0,1,-nbitq), 
to_sfixed(75.0/65536.0,1,-nbitq), 
to_sfixed(-2210.0/65536.0,1,-nbitq)  ), 
( to_sfixed(203.0/65536.0,1,-nbitq), 
to_sfixed(-5405.0/65536.0,1,-nbitq), 
to_sfixed(-4213.0/65536.0,1,-nbitq), 
to_sfixed(-4561.0/65536.0,1,-nbitq), 
to_sfixed(-2316.0/65536.0,1,-nbitq), 
to_sfixed(-3624.0/65536.0,1,-nbitq), 
to_sfixed(755.0/65536.0,1,-nbitq), 
to_sfixed(2302.0/65536.0,1,-nbitq), 
to_sfixed(4030.0/65536.0,1,-nbitq), 
to_sfixed(-2488.0/65536.0,1,-nbitq), 
to_sfixed(614.0/65536.0,1,-nbitq), 
to_sfixed(6564.0/65536.0,1,-nbitq), 
to_sfixed(-1571.0/65536.0,1,-nbitq), 
to_sfixed(6033.0/65536.0,1,-nbitq), 
to_sfixed(-338.0/65536.0,1,-nbitq), 
to_sfixed(1045.0/65536.0,1,-nbitq), 
to_sfixed(-692.0/65536.0,1,-nbitq), 
to_sfixed(2097.0/65536.0,1,-nbitq), 
to_sfixed(-388.0/65536.0,1,-nbitq), 
to_sfixed(2125.0/65536.0,1,-nbitq), 
to_sfixed(544.0/65536.0,1,-nbitq), 
to_sfixed(1070.0/65536.0,1,-nbitq), 
to_sfixed(6520.0/65536.0,1,-nbitq), 
to_sfixed(1228.0/65536.0,1,-nbitq), 
to_sfixed(-2083.0/65536.0,1,-nbitq), 
to_sfixed(-3921.0/65536.0,1,-nbitq), 
to_sfixed(647.0/65536.0,1,-nbitq), 
to_sfixed(2885.0/65536.0,1,-nbitq), 
to_sfixed(-7733.0/65536.0,1,-nbitq), 
to_sfixed(1757.0/65536.0,1,-nbitq), 
to_sfixed(3645.0/65536.0,1,-nbitq), 
to_sfixed(-6120.0/65536.0,1,-nbitq), 
to_sfixed(-947.0/65536.0,1,-nbitq), 
to_sfixed(6716.0/65536.0,1,-nbitq), 
to_sfixed(-1290.0/65536.0,1,-nbitq), 
to_sfixed(1677.0/65536.0,1,-nbitq), 
to_sfixed(3351.0/65536.0,1,-nbitq), 
to_sfixed(5112.0/65536.0,1,-nbitq), 
to_sfixed(12102.0/65536.0,1,-nbitq), 
to_sfixed(-6944.0/65536.0,1,-nbitq), 
to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(-2101.0/65536.0,1,-nbitq), 
to_sfixed(-3955.0/65536.0,1,-nbitq), 
to_sfixed(5089.0/65536.0,1,-nbitq), 
to_sfixed(1392.0/65536.0,1,-nbitq), 
to_sfixed(-10540.0/65536.0,1,-nbitq), 
to_sfixed(1456.0/65536.0,1,-nbitq), 
to_sfixed(369.0/65536.0,1,-nbitq), 
to_sfixed(307.0/65536.0,1,-nbitq), 
to_sfixed(2804.0/65536.0,1,-nbitq), 
to_sfixed(383.0/65536.0,1,-nbitq), 
to_sfixed(-3980.0/65536.0,1,-nbitq), 
to_sfixed(1114.0/65536.0,1,-nbitq), 
to_sfixed(-2907.0/65536.0,1,-nbitq), 
to_sfixed(-2416.0/65536.0,1,-nbitq), 
to_sfixed(-2976.0/65536.0,1,-nbitq), 
to_sfixed(-228.0/65536.0,1,-nbitq), 
to_sfixed(-1746.0/65536.0,1,-nbitq), 
to_sfixed(-196.0/65536.0,1,-nbitq), 
to_sfixed(-5526.0/65536.0,1,-nbitq), 
to_sfixed(-2339.0/65536.0,1,-nbitq), 
to_sfixed(2469.0/65536.0,1,-nbitq), 
to_sfixed(2515.0/65536.0,1,-nbitq), 
to_sfixed(1708.0/65536.0,1,-nbitq), 
to_sfixed(4273.0/65536.0,1,-nbitq), 
to_sfixed(-4506.0/65536.0,1,-nbitq), 
to_sfixed(2936.0/65536.0,1,-nbitq), 
to_sfixed(8105.0/65536.0,1,-nbitq), 
to_sfixed(-1992.0/65536.0,1,-nbitq), 
to_sfixed(4925.0/65536.0,1,-nbitq), 
to_sfixed(-2065.0/65536.0,1,-nbitq), 
to_sfixed(8773.0/65536.0,1,-nbitq), 
to_sfixed(-151.0/65536.0,1,-nbitq), 
to_sfixed(1959.0/65536.0,1,-nbitq), 
to_sfixed(-902.0/65536.0,1,-nbitq), 
to_sfixed(2005.0/65536.0,1,-nbitq), 
to_sfixed(6979.0/65536.0,1,-nbitq), 
to_sfixed(-5283.0/65536.0,1,-nbitq), 
to_sfixed(1205.0/65536.0,1,-nbitq), 
to_sfixed(-1603.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2157.0/65536.0,1,-nbitq), 
to_sfixed(-1246.0/65536.0,1,-nbitq), 
to_sfixed(-2866.0/65536.0,1,-nbitq), 
to_sfixed(-4150.0/65536.0,1,-nbitq), 
to_sfixed(-6170.0/65536.0,1,-nbitq), 
to_sfixed(-5308.0/65536.0,1,-nbitq), 
to_sfixed(52.0/65536.0,1,-nbitq), 
to_sfixed(2992.0/65536.0,1,-nbitq), 
to_sfixed(-755.0/65536.0,1,-nbitq), 
to_sfixed(-457.0/65536.0,1,-nbitq), 
to_sfixed(-1343.0/65536.0,1,-nbitq), 
to_sfixed(9027.0/65536.0,1,-nbitq), 
to_sfixed(2354.0/65536.0,1,-nbitq), 
to_sfixed(13.0/65536.0,1,-nbitq), 
to_sfixed(1593.0/65536.0,1,-nbitq), 
to_sfixed(-548.0/65536.0,1,-nbitq), 
to_sfixed(-98.0/65536.0,1,-nbitq), 
to_sfixed(-3207.0/65536.0,1,-nbitq), 
to_sfixed(1516.0/65536.0,1,-nbitq), 
to_sfixed(3084.0/65536.0,1,-nbitq), 
to_sfixed(-2826.0/65536.0,1,-nbitq), 
to_sfixed(-2222.0/65536.0,1,-nbitq), 
to_sfixed(-1075.0/65536.0,1,-nbitq), 
to_sfixed(-3385.0/65536.0,1,-nbitq), 
to_sfixed(1683.0/65536.0,1,-nbitq), 
to_sfixed(-4649.0/65536.0,1,-nbitq), 
to_sfixed(3517.0/65536.0,1,-nbitq), 
to_sfixed(1059.0/65536.0,1,-nbitq), 
to_sfixed(-7906.0/65536.0,1,-nbitq), 
to_sfixed(-1574.0/65536.0,1,-nbitq), 
to_sfixed(-240.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(2056.0/65536.0,1,-nbitq), 
to_sfixed(3852.0/65536.0,1,-nbitq), 
to_sfixed(1360.0/65536.0,1,-nbitq), 
to_sfixed(-1484.0/65536.0,1,-nbitq), 
to_sfixed(1227.0/65536.0,1,-nbitq), 
to_sfixed(5303.0/65536.0,1,-nbitq), 
to_sfixed(10802.0/65536.0,1,-nbitq), 
to_sfixed(-3896.0/65536.0,1,-nbitq), 
to_sfixed(1419.0/65536.0,1,-nbitq), 
to_sfixed(569.0/65536.0,1,-nbitq), 
to_sfixed(3640.0/65536.0,1,-nbitq), 
to_sfixed(4907.0/65536.0,1,-nbitq), 
to_sfixed(738.0/65536.0,1,-nbitq), 
to_sfixed(-2413.0/65536.0,1,-nbitq), 
to_sfixed(724.0/65536.0,1,-nbitq), 
to_sfixed(-155.0/65536.0,1,-nbitq), 
to_sfixed(3397.0/65536.0,1,-nbitq), 
to_sfixed(3460.0/65536.0,1,-nbitq), 
to_sfixed(-1385.0/65536.0,1,-nbitq), 
to_sfixed(-3002.0/65536.0,1,-nbitq), 
to_sfixed(-2429.0/65536.0,1,-nbitq), 
to_sfixed(-9555.0/65536.0,1,-nbitq), 
to_sfixed(2205.0/65536.0,1,-nbitq), 
to_sfixed(-2293.0/65536.0,1,-nbitq), 
to_sfixed(1945.0/65536.0,1,-nbitq), 
to_sfixed(1073.0/65536.0,1,-nbitq), 
to_sfixed(2485.0/65536.0,1,-nbitq), 
to_sfixed(-5728.0/65536.0,1,-nbitq), 
to_sfixed(-1499.0/65536.0,1,-nbitq), 
to_sfixed(1332.0/65536.0,1,-nbitq), 
to_sfixed(498.0/65536.0,1,-nbitq), 
to_sfixed(-1887.0/65536.0,1,-nbitq), 
to_sfixed(458.0/65536.0,1,-nbitq), 
to_sfixed(-2919.0/65536.0,1,-nbitq), 
to_sfixed(7379.0/65536.0,1,-nbitq), 
to_sfixed(7426.0/65536.0,1,-nbitq), 
to_sfixed(2583.0/65536.0,1,-nbitq), 
to_sfixed(6577.0/65536.0,1,-nbitq), 
to_sfixed(-2664.0/65536.0,1,-nbitq), 
to_sfixed(7844.0/65536.0,1,-nbitq), 
to_sfixed(-826.0/65536.0,1,-nbitq), 
to_sfixed(755.0/65536.0,1,-nbitq), 
to_sfixed(1214.0/65536.0,1,-nbitq), 
to_sfixed(-2104.0/65536.0,1,-nbitq), 
to_sfixed(4291.0/65536.0,1,-nbitq), 
to_sfixed(-3803.0/65536.0,1,-nbitq), 
to_sfixed(1816.0/65536.0,1,-nbitq), 
to_sfixed(-934.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4024.0/65536.0,1,-nbitq), 
to_sfixed(2579.0/65536.0,1,-nbitq), 
to_sfixed(-2591.0/65536.0,1,-nbitq), 
to_sfixed(-7653.0/65536.0,1,-nbitq), 
to_sfixed(-6435.0/65536.0,1,-nbitq), 
to_sfixed(-2359.0/65536.0,1,-nbitq), 
to_sfixed(-43.0/65536.0,1,-nbitq), 
to_sfixed(1031.0/65536.0,1,-nbitq), 
to_sfixed(1847.0/65536.0,1,-nbitq), 
to_sfixed(-719.0/65536.0,1,-nbitq), 
to_sfixed(-3025.0/65536.0,1,-nbitq), 
to_sfixed(7189.0/65536.0,1,-nbitq), 
to_sfixed(-2193.0/65536.0,1,-nbitq), 
to_sfixed(-3527.0/65536.0,1,-nbitq), 
to_sfixed(2490.0/65536.0,1,-nbitq), 
to_sfixed(-1881.0/65536.0,1,-nbitq), 
to_sfixed(-2389.0/65536.0,1,-nbitq), 
to_sfixed(-8902.0/65536.0,1,-nbitq), 
to_sfixed(4888.0/65536.0,1,-nbitq), 
to_sfixed(-885.0/65536.0,1,-nbitq), 
to_sfixed(-1805.0/65536.0,1,-nbitq), 
to_sfixed(-5425.0/65536.0,1,-nbitq), 
to_sfixed(5864.0/65536.0,1,-nbitq), 
to_sfixed(460.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(-3530.0/65536.0,1,-nbitq), 
to_sfixed(3918.0/65536.0,1,-nbitq), 
to_sfixed(2925.0/65536.0,1,-nbitq), 
to_sfixed(-6634.0/65536.0,1,-nbitq), 
to_sfixed(-40.0/65536.0,1,-nbitq), 
to_sfixed(-913.0/65536.0,1,-nbitq), 
to_sfixed(-2766.0/65536.0,1,-nbitq), 
to_sfixed(2547.0/65536.0,1,-nbitq), 
to_sfixed(4742.0/65536.0,1,-nbitq), 
to_sfixed(-1645.0/65536.0,1,-nbitq), 
to_sfixed(3265.0/65536.0,1,-nbitq), 
to_sfixed(4228.0/65536.0,1,-nbitq), 
to_sfixed(10661.0/65536.0,1,-nbitq), 
to_sfixed(7505.0/65536.0,1,-nbitq), 
to_sfixed(-181.0/65536.0,1,-nbitq), 
to_sfixed(3492.0/65536.0,1,-nbitq), 
to_sfixed(-1284.0/65536.0,1,-nbitq), 
to_sfixed(5077.0/65536.0,1,-nbitq), 
to_sfixed(5352.0/65536.0,1,-nbitq), 
to_sfixed(-128.0/65536.0,1,-nbitq), 
to_sfixed(-1542.0/65536.0,1,-nbitq), 
to_sfixed(1370.0/65536.0,1,-nbitq), 
to_sfixed(-5517.0/65536.0,1,-nbitq), 
to_sfixed(1068.0/65536.0,1,-nbitq), 
to_sfixed(2283.0/65536.0,1,-nbitq), 
to_sfixed(1017.0/65536.0,1,-nbitq), 
to_sfixed(-1264.0/65536.0,1,-nbitq), 
to_sfixed(2165.0/65536.0,1,-nbitq), 
to_sfixed(-13657.0/65536.0,1,-nbitq), 
to_sfixed(-1964.0/65536.0,1,-nbitq), 
to_sfixed(-6673.0/65536.0,1,-nbitq), 
to_sfixed(3118.0/65536.0,1,-nbitq), 
to_sfixed(198.0/65536.0,1,-nbitq), 
to_sfixed(462.0/65536.0,1,-nbitq), 
to_sfixed(-11593.0/65536.0,1,-nbitq), 
to_sfixed(-2115.0/65536.0,1,-nbitq), 
to_sfixed(1861.0/65536.0,1,-nbitq), 
to_sfixed(-264.0/65536.0,1,-nbitq), 
to_sfixed(1099.0/65536.0,1,-nbitq), 
to_sfixed(2944.0/65536.0,1,-nbitq), 
to_sfixed(220.0/65536.0,1,-nbitq), 
to_sfixed(5598.0/65536.0,1,-nbitq), 
to_sfixed(10237.0/65536.0,1,-nbitq), 
to_sfixed(1216.0/65536.0,1,-nbitq), 
to_sfixed(6253.0/65536.0,1,-nbitq), 
to_sfixed(-67.0/65536.0,1,-nbitq), 
to_sfixed(6277.0/65536.0,1,-nbitq), 
to_sfixed(-2582.0/65536.0,1,-nbitq), 
to_sfixed(-2379.0/65536.0,1,-nbitq), 
to_sfixed(-2922.0/65536.0,1,-nbitq), 
to_sfixed(859.0/65536.0,1,-nbitq), 
to_sfixed(7560.0/65536.0,1,-nbitq), 
to_sfixed(1793.0/65536.0,1,-nbitq), 
to_sfixed(872.0/65536.0,1,-nbitq), 
to_sfixed(-5150.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2547.0/65536.0,1,-nbitq), 
to_sfixed(191.0/65536.0,1,-nbitq), 
to_sfixed(-8637.0/65536.0,1,-nbitq), 
to_sfixed(-9830.0/65536.0,1,-nbitq), 
to_sfixed(-5878.0/65536.0,1,-nbitq), 
to_sfixed(-182.0/65536.0,1,-nbitq), 
to_sfixed(-494.0/65536.0,1,-nbitq), 
to_sfixed(-4138.0/65536.0,1,-nbitq), 
to_sfixed(2797.0/65536.0,1,-nbitq), 
to_sfixed(-302.0/65536.0,1,-nbitq), 
to_sfixed(-176.0/65536.0,1,-nbitq), 
to_sfixed(-872.0/65536.0,1,-nbitq), 
to_sfixed(1414.0/65536.0,1,-nbitq), 
to_sfixed(-6500.0/65536.0,1,-nbitq), 
to_sfixed(-541.0/65536.0,1,-nbitq), 
to_sfixed(-1049.0/65536.0,1,-nbitq), 
to_sfixed(-2957.0/65536.0,1,-nbitq), 
to_sfixed(-3830.0/65536.0,1,-nbitq), 
to_sfixed(1261.0/65536.0,1,-nbitq), 
to_sfixed(-1724.0/65536.0,1,-nbitq), 
to_sfixed(-2808.0/65536.0,1,-nbitq), 
to_sfixed(-3821.0/65536.0,1,-nbitq), 
to_sfixed(1578.0/65536.0,1,-nbitq), 
to_sfixed(5775.0/65536.0,1,-nbitq), 
to_sfixed(-3173.0/65536.0,1,-nbitq), 
to_sfixed(-7576.0/65536.0,1,-nbitq), 
to_sfixed(3802.0/65536.0,1,-nbitq), 
to_sfixed(-627.0/65536.0,1,-nbitq), 
to_sfixed(-430.0/65536.0,1,-nbitq), 
to_sfixed(-1620.0/65536.0,1,-nbitq), 
to_sfixed(769.0/65536.0,1,-nbitq), 
to_sfixed(-2763.0/65536.0,1,-nbitq), 
to_sfixed(3288.0/65536.0,1,-nbitq), 
to_sfixed(326.0/65536.0,1,-nbitq), 
to_sfixed(2032.0/65536.0,1,-nbitq), 
to_sfixed(-1179.0/65536.0,1,-nbitq), 
to_sfixed(3301.0/65536.0,1,-nbitq), 
to_sfixed(7330.0/65536.0,1,-nbitq), 
to_sfixed(10481.0/65536.0,1,-nbitq), 
to_sfixed(-282.0/65536.0,1,-nbitq), 
to_sfixed(1211.0/65536.0,1,-nbitq), 
to_sfixed(-2148.0/65536.0,1,-nbitq), 
to_sfixed(784.0/65536.0,1,-nbitq), 
to_sfixed(1714.0/65536.0,1,-nbitq), 
to_sfixed(-471.0/65536.0,1,-nbitq), 
to_sfixed(-786.0/65536.0,1,-nbitq), 
to_sfixed(2089.0/65536.0,1,-nbitq), 
to_sfixed(-2282.0/65536.0,1,-nbitq), 
to_sfixed(902.0/65536.0,1,-nbitq), 
to_sfixed(3158.0/65536.0,1,-nbitq), 
to_sfixed(-1943.0/65536.0,1,-nbitq), 
to_sfixed(-1437.0/65536.0,1,-nbitq), 
to_sfixed(-1699.0/65536.0,1,-nbitq), 
to_sfixed(-9806.0/65536.0,1,-nbitq), 
to_sfixed(-240.0/65536.0,1,-nbitq), 
to_sfixed(-3726.0/65536.0,1,-nbitq), 
to_sfixed(196.0/65536.0,1,-nbitq), 
to_sfixed(-606.0/65536.0,1,-nbitq), 
to_sfixed(570.0/65536.0,1,-nbitq), 
to_sfixed(-13168.0/65536.0,1,-nbitq), 
to_sfixed(195.0/65536.0,1,-nbitq), 
to_sfixed(916.0/65536.0,1,-nbitq), 
to_sfixed(1894.0/65536.0,1,-nbitq), 
to_sfixed(1765.0/65536.0,1,-nbitq), 
to_sfixed(5189.0/65536.0,1,-nbitq), 
to_sfixed(-3987.0/65536.0,1,-nbitq), 
to_sfixed(130.0/65536.0,1,-nbitq), 
to_sfixed(9952.0/65536.0,1,-nbitq), 
to_sfixed(4538.0/65536.0,1,-nbitq), 
to_sfixed(13469.0/65536.0,1,-nbitq), 
to_sfixed(-3575.0/65536.0,1,-nbitq), 
to_sfixed(3643.0/65536.0,1,-nbitq), 
to_sfixed(-5818.0/65536.0,1,-nbitq), 
to_sfixed(-523.0/65536.0,1,-nbitq), 
to_sfixed(-1005.0/65536.0,1,-nbitq), 
to_sfixed(-1658.0/65536.0,1,-nbitq), 
to_sfixed(1719.0/65536.0,1,-nbitq), 
to_sfixed(2461.0/65536.0,1,-nbitq), 
to_sfixed(-571.0/65536.0,1,-nbitq), 
to_sfixed(-1488.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3765.0/65536.0,1,-nbitq), 
to_sfixed(3097.0/65536.0,1,-nbitq), 
to_sfixed(-8518.0/65536.0,1,-nbitq), 
to_sfixed(-13807.0/65536.0,1,-nbitq), 
to_sfixed(-5736.0/65536.0,1,-nbitq), 
to_sfixed(2289.0/65536.0,1,-nbitq), 
to_sfixed(1760.0/65536.0,1,-nbitq), 
to_sfixed(-279.0/65536.0,1,-nbitq), 
to_sfixed(6597.0/65536.0,1,-nbitq), 
to_sfixed(1675.0/65536.0,1,-nbitq), 
to_sfixed(2845.0/65536.0,1,-nbitq), 
to_sfixed(1487.0/65536.0,1,-nbitq), 
to_sfixed(-3389.0/65536.0,1,-nbitq), 
to_sfixed(-3416.0/65536.0,1,-nbitq), 
to_sfixed(695.0/65536.0,1,-nbitq), 
to_sfixed(-720.0/65536.0,1,-nbitq), 
to_sfixed(1360.0/65536.0,1,-nbitq), 
to_sfixed(-3410.0/65536.0,1,-nbitq), 
to_sfixed(3655.0/65536.0,1,-nbitq), 
to_sfixed(-2436.0/65536.0,1,-nbitq), 
to_sfixed(-3871.0/65536.0,1,-nbitq), 
to_sfixed(714.0/65536.0,1,-nbitq), 
to_sfixed(5173.0/65536.0,1,-nbitq), 
to_sfixed(5589.0/65536.0,1,-nbitq), 
to_sfixed(-5042.0/65536.0,1,-nbitq), 
to_sfixed(-9441.0/65536.0,1,-nbitq), 
to_sfixed(687.0/65536.0,1,-nbitq), 
to_sfixed(-337.0/65536.0,1,-nbitq), 
to_sfixed(233.0/65536.0,1,-nbitq), 
to_sfixed(292.0/65536.0,1,-nbitq), 
to_sfixed(-1586.0/65536.0,1,-nbitq), 
to_sfixed(-10897.0/65536.0,1,-nbitq), 
to_sfixed(1597.0/65536.0,1,-nbitq), 
to_sfixed(-1045.0/65536.0,1,-nbitq), 
to_sfixed(-1812.0/65536.0,1,-nbitq), 
to_sfixed(-3235.0/65536.0,1,-nbitq), 
to_sfixed(6581.0/65536.0,1,-nbitq), 
to_sfixed(5487.0/65536.0,1,-nbitq), 
to_sfixed(7696.0/65536.0,1,-nbitq), 
to_sfixed(2865.0/65536.0,1,-nbitq), 
to_sfixed(-4783.0/65536.0,1,-nbitq), 
to_sfixed(-593.0/65536.0,1,-nbitq), 
to_sfixed(1868.0/65536.0,1,-nbitq), 
to_sfixed(851.0/65536.0,1,-nbitq), 
to_sfixed(-1041.0/65536.0,1,-nbitq), 
to_sfixed(-6738.0/65536.0,1,-nbitq), 
to_sfixed(124.0/65536.0,1,-nbitq), 
to_sfixed(4635.0/65536.0,1,-nbitq), 
to_sfixed(2477.0/65536.0,1,-nbitq), 
to_sfixed(1067.0/65536.0,1,-nbitq), 
to_sfixed(2280.0/65536.0,1,-nbitq), 
to_sfixed(-1573.0/65536.0,1,-nbitq), 
to_sfixed(-6339.0/65536.0,1,-nbitq), 
to_sfixed(-9252.0/65536.0,1,-nbitq), 
to_sfixed(-2446.0/65536.0,1,-nbitq), 
to_sfixed(-5985.0/65536.0,1,-nbitq), 
to_sfixed(1406.0/65536.0,1,-nbitq), 
to_sfixed(775.0/65536.0,1,-nbitq), 
to_sfixed(-1013.0/65536.0,1,-nbitq), 
to_sfixed(-12906.0/65536.0,1,-nbitq), 
to_sfixed(1659.0/65536.0,1,-nbitq), 
to_sfixed(-705.0/65536.0,1,-nbitq), 
to_sfixed(999.0/65536.0,1,-nbitq), 
to_sfixed(-1460.0/65536.0,1,-nbitq), 
to_sfixed(1113.0/65536.0,1,-nbitq), 
to_sfixed(-5316.0/65536.0,1,-nbitq), 
to_sfixed(1901.0/65536.0,1,-nbitq), 
to_sfixed(13381.0/65536.0,1,-nbitq), 
to_sfixed(4072.0/65536.0,1,-nbitq), 
to_sfixed(12540.0/65536.0,1,-nbitq), 
to_sfixed(-1154.0/65536.0,1,-nbitq), 
to_sfixed(-4482.0/65536.0,1,-nbitq), 
to_sfixed(-4055.0/65536.0,1,-nbitq), 
to_sfixed(851.0/65536.0,1,-nbitq), 
to_sfixed(-136.0/65536.0,1,-nbitq), 
to_sfixed(2134.0/65536.0,1,-nbitq), 
to_sfixed(3020.0/65536.0,1,-nbitq), 
to_sfixed(3878.0/65536.0,1,-nbitq), 
to_sfixed(2147.0/65536.0,1,-nbitq), 
to_sfixed(-2597.0/65536.0,1,-nbitq)  ), 
( to_sfixed(6086.0/65536.0,1,-nbitq), 
to_sfixed(27.0/65536.0,1,-nbitq), 
to_sfixed(-7780.0/65536.0,1,-nbitq), 
to_sfixed(-9585.0/65536.0,1,-nbitq), 
to_sfixed(-3117.0/65536.0,1,-nbitq), 
to_sfixed(-2870.0/65536.0,1,-nbitq), 
to_sfixed(-1833.0/65536.0,1,-nbitq), 
to_sfixed(-4440.0/65536.0,1,-nbitq), 
to_sfixed(7076.0/65536.0,1,-nbitq), 
to_sfixed(804.0/65536.0,1,-nbitq), 
to_sfixed(-1872.0/65536.0,1,-nbitq), 
to_sfixed(-8892.0/65536.0,1,-nbitq), 
to_sfixed(1319.0/65536.0,1,-nbitq), 
to_sfixed(-276.0/65536.0,1,-nbitq), 
to_sfixed(1762.0/65536.0,1,-nbitq), 
to_sfixed(1431.0/65536.0,1,-nbitq), 
to_sfixed(1712.0/65536.0,1,-nbitq), 
to_sfixed(-5436.0/65536.0,1,-nbitq), 
to_sfixed(5446.0/65536.0,1,-nbitq), 
to_sfixed(-1174.0/65536.0,1,-nbitq), 
to_sfixed(-6171.0/65536.0,1,-nbitq), 
to_sfixed(443.0/65536.0,1,-nbitq), 
to_sfixed(3467.0/65536.0,1,-nbitq), 
to_sfixed(6156.0/65536.0,1,-nbitq), 
to_sfixed(-2321.0/65536.0,1,-nbitq), 
to_sfixed(-4361.0/65536.0,1,-nbitq), 
to_sfixed(-246.0/65536.0,1,-nbitq), 
to_sfixed(833.0/65536.0,1,-nbitq), 
to_sfixed(1019.0/65536.0,1,-nbitq), 
to_sfixed(-990.0/65536.0,1,-nbitq), 
to_sfixed(789.0/65536.0,1,-nbitq), 
to_sfixed(-5514.0/65536.0,1,-nbitq), 
to_sfixed(2395.0/65536.0,1,-nbitq), 
to_sfixed(-1649.0/65536.0,1,-nbitq), 
to_sfixed(1774.0/65536.0,1,-nbitq), 
to_sfixed(-2836.0/65536.0,1,-nbitq), 
to_sfixed(3568.0/65536.0,1,-nbitq), 
to_sfixed(6829.0/65536.0,1,-nbitq), 
to_sfixed(1810.0/65536.0,1,-nbitq), 
to_sfixed(2157.0/65536.0,1,-nbitq), 
to_sfixed(-890.0/65536.0,1,-nbitq), 
to_sfixed(-2058.0/65536.0,1,-nbitq), 
to_sfixed(-3308.0/65536.0,1,-nbitq), 
to_sfixed(-1254.0/65536.0,1,-nbitq), 
to_sfixed(36.0/65536.0,1,-nbitq), 
to_sfixed(-2533.0/65536.0,1,-nbitq), 
to_sfixed(-1110.0/65536.0,1,-nbitq), 
to_sfixed(5833.0/65536.0,1,-nbitq), 
to_sfixed(652.0/65536.0,1,-nbitq), 
to_sfixed(-1359.0/65536.0,1,-nbitq), 
to_sfixed(-1101.0/65536.0,1,-nbitq), 
to_sfixed(-728.0/65536.0,1,-nbitq), 
to_sfixed(-9388.0/65536.0,1,-nbitq), 
to_sfixed(-7508.0/65536.0,1,-nbitq), 
to_sfixed(131.0/65536.0,1,-nbitq), 
to_sfixed(-7159.0/65536.0,1,-nbitq), 
to_sfixed(-906.0/65536.0,1,-nbitq), 
to_sfixed(-2344.0/65536.0,1,-nbitq), 
to_sfixed(-2023.0/65536.0,1,-nbitq), 
to_sfixed(-14268.0/65536.0,1,-nbitq), 
to_sfixed(3538.0/65536.0,1,-nbitq), 
to_sfixed(1066.0/65536.0,1,-nbitq), 
to_sfixed(3196.0/65536.0,1,-nbitq), 
to_sfixed(-3152.0/65536.0,1,-nbitq), 
to_sfixed(3699.0/65536.0,1,-nbitq), 
to_sfixed(-4932.0/65536.0,1,-nbitq), 
to_sfixed(2373.0/65536.0,1,-nbitq), 
to_sfixed(8911.0/65536.0,1,-nbitq), 
to_sfixed(11258.0/65536.0,1,-nbitq), 
to_sfixed(8955.0/65536.0,1,-nbitq), 
to_sfixed(417.0/65536.0,1,-nbitq), 
to_sfixed(68.0/65536.0,1,-nbitq), 
to_sfixed(-4578.0/65536.0,1,-nbitq), 
to_sfixed(-2557.0/65536.0,1,-nbitq), 
to_sfixed(2755.0/65536.0,1,-nbitq), 
to_sfixed(2108.0/65536.0,1,-nbitq), 
to_sfixed(3351.0/65536.0,1,-nbitq), 
to_sfixed(294.0/65536.0,1,-nbitq), 
to_sfixed(1585.0/65536.0,1,-nbitq), 
to_sfixed(-214.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3155.0/65536.0,1,-nbitq), 
to_sfixed(-1514.0/65536.0,1,-nbitq), 
to_sfixed(-1192.0/65536.0,1,-nbitq), 
to_sfixed(-4007.0/65536.0,1,-nbitq), 
to_sfixed(1371.0/65536.0,1,-nbitq), 
to_sfixed(3036.0/65536.0,1,-nbitq), 
to_sfixed(1473.0/65536.0,1,-nbitq), 
to_sfixed(-1753.0/65536.0,1,-nbitq), 
to_sfixed(6890.0/65536.0,1,-nbitq), 
to_sfixed(-2325.0/65536.0,1,-nbitq), 
to_sfixed(-187.0/65536.0,1,-nbitq), 
to_sfixed(-14575.0/65536.0,1,-nbitq), 
to_sfixed(-894.0/65536.0,1,-nbitq), 
to_sfixed(7857.0/65536.0,1,-nbitq), 
to_sfixed(719.0/65536.0,1,-nbitq), 
to_sfixed(-2156.0/65536.0,1,-nbitq), 
to_sfixed(276.0/65536.0,1,-nbitq), 
to_sfixed(-4266.0/65536.0,1,-nbitq), 
to_sfixed(1651.0/65536.0,1,-nbitq), 
to_sfixed(2217.0/65536.0,1,-nbitq), 
to_sfixed(-10967.0/65536.0,1,-nbitq), 
to_sfixed(-2414.0/65536.0,1,-nbitq), 
to_sfixed(-2716.0/65536.0,1,-nbitq), 
to_sfixed(8173.0/65536.0,1,-nbitq), 
to_sfixed(-4924.0/65536.0,1,-nbitq), 
to_sfixed(6205.0/65536.0,1,-nbitq), 
to_sfixed(6215.0/65536.0,1,-nbitq), 
to_sfixed(-196.0/65536.0,1,-nbitq), 
to_sfixed(1914.0/65536.0,1,-nbitq), 
to_sfixed(1115.0/65536.0,1,-nbitq), 
to_sfixed(3082.0/65536.0,1,-nbitq), 
to_sfixed(-8616.0/65536.0,1,-nbitq), 
to_sfixed(-314.0/65536.0,1,-nbitq), 
to_sfixed(-1831.0/65536.0,1,-nbitq), 
to_sfixed(-56.0/65536.0,1,-nbitq), 
to_sfixed(-1863.0/65536.0,1,-nbitq), 
to_sfixed(5430.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(-1134.0/65536.0,1,-nbitq), 
to_sfixed(1.0/65536.0,1,-nbitq), 
to_sfixed(-736.0/65536.0,1,-nbitq), 
to_sfixed(-2328.0/65536.0,1,-nbitq), 
to_sfixed(-5020.0/65536.0,1,-nbitq), 
to_sfixed(-5678.0/65536.0,1,-nbitq), 
to_sfixed(-292.0/65536.0,1,-nbitq), 
to_sfixed(-931.0/65536.0,1,-nbitq), 
to_sfixed(-3022.0/65536.0,1,-nbitq), 
to_sfixed(4187.0/65536.0,1,-nbitq), 
to_sfixed(1122.0/65536.0,1,-nbitq), 
to_sfixed(-1208.0/65536.0,1,-nbitq), 
to_sfixed(2081.0/65536.0,1,-nbitq), 
to_sfixed(2810.0/65536.0,1,-nbitq), 
to_sfixed(-5396.0/65536.0,1,-nbitq), 
to_sfixed(-3307.0/65536.0,1,-nbitq), 
to_sfixed(-21.0/65536.0,1,-nbitq), 
to_sfixed(-5751.0/65536.0,1,-nbitq), 
to_sfixed(-2673.0/65536.0,1,-nbitq), 
to_sfixed(-2096.0/65536.0,1,-nbitq), 
to_sfixed(-1253.0/65536.0,1,-nbitq), 
to_sfixed(-4831.0/65536.0,1,-nbitq), 
to_sfixed(274.0/65536.0,1,-nbitq), 
to_sfixed(-1781.0/65536.0,1,-nbitq), 
to_sfixed(-457.0/65536.0,1,-nbitq), 
to_sfixed(417.0/65536.0,1,-nbitq), 
to_sfixed(2480.0/65536.0,1,-nbitq), 
to_sfixed(-4943.0/65536.0,1,-nbitq), 
to_sfixed(-981.0/65536.0,1,-nbitq), 
to_sfixed(5784.0/65536.0,1,-nbitq), 
to_sfixed(8727.0/65536.0,1,-nbitq), 
to_sfixed(-1638.0/65536.0,1,-nbitq), 
to_sfixed(-3174.0/65536.0,1,-nbitq), 
to_sfixed(-1339.0/65536.0,1,-nbitq), 
to_sfixed(-271.0/65536.0,1,-nbitq), 
to_sfixed(-1405.0/65536.0,1,-nbitq), 
to_sfixed(-826.0/65536.0,1,-nbitq), 
to_sfixed(1788.0/65536.0,1,-nbitq), 
to_sfixed(3812.0/65536.0,1,-nbitq), 
to_sfixed(-5933.0/65536.0,1,-nbitq), 
to_sfixed(87.0/65536.0,1,-nbitq), 
to_sfixed(154.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2496.0/65536.0,1,-nbitq), 
to_sfixed(2065.0/65536.0,1,-nbitq), 
to_sfixed(-31.0/65536.0,1,-nbitq), 
to_sfixed(-4358.0/65536.0,1,-nbitq), 
to_sfixed(-12.0/65536.0,1,-nbitq), 
to_sfixed(2386.0/65536.0,1,-nbitq), 
to_sfixed(1724.0/65536.0,1,-nbitq), 
to_sfixed(-3030.0/65536.0,1,-nbitq), 
to_sfixed(3908.0/65536.0,1,-nbitq), 
to_sfixed(-1691.0/65536.0,1,-nbitq), 
to_sfixed(-1748.0/65536.0,1,-nbitq), 
to_sfixed(-14786.0/65536.0,1,-nbitq), 
to_sfixed(382.0/65536.0,1,-nbitq), 
to_sfixed(7309.0/65536.0,1,-nbitq), 
to_sfixed(-1319.0/65536.0,1,-nbitq), 
to_sfixed(1832.0/65536.0,1,-nbitq), 
to_sfixed(1988.0/65536.0,1,-nbitq), 
to_sfixed(-337.0/65536.0,1,-nbitq), 
to_sfixed(3685.0/65536.0,1,-nbitq), 
to_sfixed(786.0/65536.0,1,-nbitq), 
to_sfixed(-10375.0/65536.0,1,-nbitq), 
to_sfixed(-3224.0/65536.0,1,-nbitq), 
to_sfixed(-7655.0/65536.0,1,-nbitq), 
to_sfixed(5201.0/65536.0,1,-nbitq), 
to_sfixed(-3083.0/65536.0,1,-nbitq), 
to_sfixed(6495.0/65536.0,1,-nbitq), 
to_sfixed(2902.0/65536.0,1,-nbitq), 
to_sfixed(3193.0/65536.0,1,-nbitq), 
to_sfixed(-2882.0/65536.0,1,-nbitq), 
to_sfixed(3306.0/65536.0,1,-nbitq), 
to_sfixed(6294.0/65536.0,1,-nbitq), 
to_sfixed(-3360.0/65536.0,1,-nbitq), 
to_sfixed(4869.0/65536.0,1,-nbitq), 
to_sfixed(-748.0/65536.0,1,-nbitq), 
to_sfixed(-1205.0/65536.0,1,-nbitq), 
to_sfixed(-3351.0/65536.0,1,-nbitq), 
to_sfixed(5138.0/65536.0,1,-nbitq), 
to_sfixed(-4806.0/65536.0,1,-nbitq), 
to_sfixed(5091.0/65536.0,1,-nbitq), 
to_sfixed(3156.0/65536.0,1,-nbitq), 
to_sfixed(-2029.0/65536.0,1,-nbitq), 
to_sfixed(1821.0/65536.0,1,-nbitq), 
to_sfixed(-10051.0/65536.0,1,-nbitq), 
to_sfixed(-5700.0/65536.0,1,-nbitq), 
to_sfixed(-1108.0/65536.0,1,-nbitq), 
to_sfixed(-4807.0/65536.0,1,-nbitq), 
to_sfixed(577.0/65536.0,1,-nbitq), 
to_sfixed(-198.0/65536.0,1,-nbitq), 
to_sfixed(-1780.0/65536.0,1,-nbitq), 
to_sfixed(-1131.0/65536.0,1,-nbitq), 
to_sfixed(-1463.0/65536.0,1,-nbitq), 
to_sfixed(501.0/65536.0,1,-nbitq), 
to_sfixed(701.0/65536.0,1,-nbitq), 
to_sfixed(-3002.0/65536.0,1,-nbitq), 
to_sfixed(362.0/65536.0,1,-nbitq), 
to_sfixed(-7587.0/65536.0,1,-nbitq), 
to_sfixed(-2806.0/65536.0,1,-nbitq), 
to_sfixed(879.0/65536.0,1,-nbitq), 
to_sfixed(-96.0/65536.0,1,-nbitq), 
to_sfixed(-4291.0/65536.0,1,-nbitq), 
to_sfixed(418.0/65536.0,1,-nbitq), 
to_sfixed(-884.0/65536.0,1,-nbitq), 
to_sfixed(823.0/65536.0,1,-nbitq), 
to_sfixed(-1991.0/65536.0,1,-nbitq), 
to_sfixed(3429.0/65536.0,1,-nbitq), 
to_sfixed(71.0/65536.0,1,-nbitq), 
to_sfixed(5169.0/65536.0,1,-nbitq), 
to_sfixed(6924.0/65536.0,1,-nbitq), 
to_sfixed(4263.0/65536.0,1,-nbitq), 
to_sfixed(-2133.0/65536.0,1,-nbitq), 
to_sfixed(1017.0/65536.0,1,-nbitq), 
to_sfixed(3647.0/65536.0,1,-nbitq), 
to_sfixed(819.0/65536.0,1,-nbitq), 
to_sfixed(900.0/65536.0,1,-nbitq), 
to_sfixed(-2824.0/65536.0,1,-nbitq), 
to_sfixed(2530.0/65536.0,1,-nbitq), 
to_sfixed(7615.0/65536.0,1,-nbitq), 
to_sfixed(-6210.0/65536.0,1,-nbitq), 
to_sfixed(-3022.0/65536.0,1,-nbitq), 
to_sfixed(1703.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2057.0/65536.0,1,-nbitq), 
to_sfixed(3244.0/65536.0,1,-nbitq), 
to_sfixed(5161.0/65536.0,1,-nbitq), 
to_sfixed(-664.0/65536.0,1,-nbitq), 
to_sfixed(1810.0/65536.0,1,-nbitq), 
to_sfixed(7660.0/65536.0,1,-nbitq), 
to_sfixed(3862.0/65536.0,1,-nbitq), 
to_sfixed(-7608.0/65536.0,1,-nbitq), 
to_sfixed(3551.0/65536.0,1,-nbitq), 
to_sfixed(-1988.0/65536.0,1,-nbitq), 
to_sfixed(-1002.0/65536.0,1,-nbitq), 
to_sfixed(-10472.0/65536.0,1,-nbitq), 
to_sfixed(325.0/65536.0,1,-nbitq), 
to_sfixed(667.0/65536.0,1,-nbitq), 
to_sfixed(-3848.0/65536.0,1,-nbitq), 
to_sfixed(-1310.0/65536.0,1,-nbitq), 
to_sfixed(2030.0/65536.0,1,-nbitq), 
to_sfixed(478.0/65536.0,1,-nbitq), 
to_sfixed(1719.0/65536.0,1,-nbitq), 
to_sfixed(-715.0/65536.0,1,-nbitq), 
to_sfixed(-5407.0/65536.0,1,-nbitq), 
to_sfixed(-2543.0/65536.0,1,-nbitq), 
to_sfixed(-10246.0/65536.0,1,-nbitq), 
to_sfixed(560.0/65536.0,1,-nbitq), 
to_sfixed(-2139.0/65536.0,1,-nbitq), 
to_sfixed(9946.0/65536.0,1,-nbitq), 
to_sfixed(3569.0/65536.0,1,-nbitq), 
to_sfixed(1744.0/65536.0,1,-nbitq), 
to_sfixed(260.0/65536.0,1,-nbitq), 
to_sfixed(-903.0/65536.0,1,-nbitq), 
to_sfixed(5075.0/65536.0,1,-nbitq), 
to_sfixed(-517.0/65536.0,1,-nbitq), 
to_sfixed(990.0/65536.0,1,-nbitq), 
to_sfixed(1651.0/65536.0,1,-nbitq), 
to_sfixed(1102.0/65536.0,1,-nbitq), 
to_sfixed(-1473.0/65536.0,1,-nbitq), 
to_sfixed(6234.0/65536.0,1,-nbitq), 
to_sfixed(-3409.0/65536.0,1,-nbitq), 
to_sfixed(1741.0/65536.0,1,-nbitq), 
to_sfixed(-2289.0/65536.0,1,-nbitq), 
to_sfixed(-4863.0/65536.0,1,-nbitq), 
to_sfixed(-457.0/65536.0,1,-nbitq), 
to_sfixed(-4679.0/65536.0,1,-nbitq), 
to_sfixed(-6223.0/65536.0,1,-nbitq), 
to_sfixed(2498.0/65536.0,1,-nbitq), 
to_sfixed(-4196.0/65536.0,1,-nbitq), 
to_sfixed(1260.0/65536.0,1,-nbitq), 
to_sfixed(-2009.0/65536.0,1,-nbitq), 
to_sfixed(-272.0/65536.0,1,-nbitq), 
to_sfixed(3620.0/65536.0,1,-nbitq), 
to_sfixed(-2479.0/65536.0,1,-nbitq), 
to_sfixed(-7605.0/65536.0,1,-nbitq), 
to_sfixed(692.0/65536.0,1,-nbitq), 
to_sfixed(3893.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(1540.0/65536.0,1,-nbitq), 
to_sfixed(1190.0/65536.0,1,-nbitq), 
to_sfixed(2016.0/65536.0,1,-nbitq), 
to_sfixed(-629.0/65536.0,1,-nbitq), 
to_sfixed(-4161.0/65536.0,1,-nbitq), 
to_sfixed(-636.0/65536.0,1,-nbitq), 
to_sfixed(2364.0/65536.0,1,-nbitq), 
to_sfixed(1476.0/65536.0,1,-nbitq), 
to_sfixed(-847.0/65536.0,1,-nbitq), 
to_sfixed(3820.0/65536.0,1,-nbitq), 
to_sfixed(-4486.0/65536.0,1,-nbitq), 
to_sfixed(2666.0/65536.0,1,-nbitq), 
to_sfixed(7462.0/65536.0,1,-nbitq), 
to_sfixed(7089.0/65536.0,1,-nbitq), 
to_sfixed(-6997.0/65536.0,1,-nbitq), 
to_sfixed(827.0/65536.0,1,-nbitq), 
to_sfixed(1691.0/65536.0,1,-nbitq), 
to_sfixed(-2532.0/65536.0,1,-nbitq), 
to_sfixed(1013.0/65536.0,1,-nbitq), 
to_sfixed(-1942.0/65536.0,1,-nbitq), 
to_sfixed(-2767.0/65536.0,1,-nbitq), 
to_sfixed(1894.0/65536.0,1,-nbitq), 
to_sfixed(-5903.0/65536.0,1,-nbitq), 
to_sfixed(-1346.0/65536.0,1,-nbitq), 
to_sfixed(624.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1623.0/65536.0,1,-nbitq), 
to_sfixed(3001.0/65536.0,1,-nbitq), 
to_sfixed(2119.0/65536.0,1,-nbitq), 
to_sfixed(6535.0/65536.0,1,-nbitq), 
to_sfixed(8595.0/65536.0,1,-nbitq), 
to_sfixed(5425.0/65536.0,1,-nbitq), 
to_sfixed(2008.0/65536.0,1,-nbitq), 
to_sfixed(-7744.0/65536.0,1,-nbitq), 
to_sfixed(313.0/65536.0,1,-nbitq), 
to_sfixed(-1181.0/65536.0,1,-nbitq), 
to_sfixed(-89.0/65536.0,1,-nbitq), 
to_sfixed(-10264.0/65536.0,1,-nbitq), 
to_sfixed(1395.0/65536.0,1,-nbitq), 
to_sfixed(5678.0/65536.0,1,-nbitq), 
to_sfixed(-304.0/65536.0,1,-nbitq), 
to_sfixed(69.0/65536.0,1,-nbitq), 
to_sfixed(1590.0/65536.0,1,-nbitq), 
to_sfixed(1563.0/65536.0,1,-nbitq), 
to_sfixed(-1837.0/65536.0,1,-nbitq), 
to_sfixed(434.0/65536.0,1,-nbitq), 
to_sfixed(-4309.0/65536.0,1,-nbitq), 
to_sfixed(-7059.0/65536.0,1,-nbitq), 
to_sfixed(-4602.0/65536.0,1,-nbitq), 
to_sfixed(-3059.0/65536.0,1,-nbitq), 
to_sfixed(-1895.0/65536.0,1,-nbitq), 
to_sfixed(7315.0/65536.0,1,-nbitq), 
to_sfixed(4137.0/65536.0,1,-nbitq), 
to_sfixed(1526.0/65536.0,1,-nbitq), 
to_sfixed(4047.0/65536.0,1,-nbitq), 
to_sfixed(-1368.0/65536.0,1,-nbitq), 
to_sfixed(1764.0/65536.0,1,-nbitq), 
to_sfixed(71.0/65536.0,1,-nbitq), 
to_sfixed(2091.0/65536.0,1,-nbitq), 
to_sfixed(3893.0/65536.0,1,-nbitq), 
to_sfixed(836.0/65536.0,1,-nbitq), 
to_sfixed(273.0/65536.0,1,-nbitq), 
to_sfixed(8354.0/65536.0,1,-nbitq), 
to_sfixed(1493.0/65536.0,1,-nbitq), 
to_sfixed(285.0/65536.0,1,-nbitq), 
to_sfixed(1408.0/65536.0,1,-nbitq), 
to_sfixed(-6032.0/65536.0,1,-nbitq), 
to_sfixed(1387.0/65536.0,1,-nbitq), 
to_sfixed(-3710.0/65536.0,1,-nbitq), 
to_sfixed(-4220.0/65536.0,1,-nbitq), 
to_sfixed(465.0/65536.0,1,-nbitq), 
to_sfixed(-4354.0/65536.0,1,-nbitq), 
to_sfixed(-4719.0/65536.0,1,-nbitq), 
to_sfixed(-1075.0/65536.0,1,-nbitq), 
to_sfixed(-2432.0/65536.0,1,-nbitq), 
to_sfixed(-941.0/65536.0,1,-nbitq), 
to_sfixed(1689.0/65536.0,1,-nbitq), 
to_sfixed(-5372.0/65536.0,1,-nbitq), 
to_sfixed(-2130.0/65536.0,1,-nbitq), 
to_sfixed(-2272.0/65536.0,1,-nbitq), 
to_sfixed(338.0/65536.0,1,-nbitq), 
to_sfixed(697.0/65536.0,1,-nbitq), 
to_sfixed(993.0/65536.0,1,-nbitq), 
to_sfixed(1253.0/65536.0,1,-nbitq), 
to_sfixed(1048.0/65536.0,1,-nbitq), 
to_sfixed(495.0/65536.0,1,-nbitq), 
to_sfixed(1510.0/65536.0,1,-nbitq), 
to_sfixed(-3086.0/65536.0,1,-nbitq), 
to_sfixed(2075.0/65536.0,1,-nbitq), 
to_sfixed(371.0/65536.0,1,-nbitq), 
to_sfixed(1980.0/65536.0,1,-nbitq), 
to_sfixed(-4748.0/65536.0,1,-nbitq), 
to_sfixed(2611.0/65536.0,1,-nbitq), 
to_sfixed(4711.0/65536.0,1,-nbitq), 
to_sfixed(5616.0/65536.0,1,-nbitq), 
to_sfixed(-7357.0/65536.0,1,-nbitq), 
to_sfixed(-2760.0/65536.0,1,-nbitq), 
to_sfixed(314.0/65536.0,1,-nbitq), 
to_sfixed(1903.0/65536.0,1,-nbitq), 
to_sfixed(-258.0/65536.0,1,-nbitq), 
to_sfixed(-2824.0/65536.0,1,-nbitq), 
to_sfixed(5174.0/65536.0,1,-nbitq), 
to_sfixed(2089.0/65536.0,1,-nbitq), 
to_sfixed(-6719.0/65536.0,1,-nbitq), 
to_sfixed(-1126.0/65536.0,1,-nbitq), 
to_sfixed(-1705.0/65536.0,1,-nbitq)  ), 
( to_sfixed(938.0/65536.0,1,-nbitq), 
to_sfixed(2065.0/65536.0,1,-nbitq), 
to_sfixed(5225.0/65536.0,1,-nbitq), 
to_sfixed(-146.0/65536.0,1,-nbitq), 
to_sfixed(6787.0/65536.0,1,-nbitq), 
to_sfixed(5544.0/65536.0,1,-nbitq), 
to_sfixed(249.0/65536.0,1,-nbitq), 
to_sfixed(-3490.0/65536.0,1,-nbitq), 
to_sfixed(-1677.0/65536.0,1,-nbitq), 
to_sfixed(1666.0/65536.0,1,-nbitq), 
to_sfixed(-1243.0/65536.0,1,-nbitq), 
to_sfixed(-2766.0/65536.0,1,-nbitq), 
to_sfixed(-4111.0/65536.0,1,-nbitq), 
to_sfixed(4063.0/65536.0,1,-nbitq), 
to_sfixed(2182.0/65536.0,1,-nbitq), 
to_sfixed(-2940.0/65536.0,1,-nbitq), 
to_sfixed(-2715.0/65536.0,1,-nbitq), 
to_sfixed(2448.0/65536.0,1,-nbitq), 
to_sfixed(21.0/65536.0,1,-nbitq), 
to_sfixed(-1288.0/65536.0,1,-nbitq), 
to_sfixed(-3277.0/65536.0,1,-nbitq), 
to_sfixed(-427.0/65536.0,1,-nbitq), 
to_sfixed(-2390.0/65536.0,1,-nbitq), 
to_sfixed(1572.0/65536.0,1,-nbitq), 
to_sfixed(143.0/65536.0,1,-nbitq), 
to_sfixed(6866.0/65536.0,1,-nbitq), 
to_sfixed(3740.0/65536.0,1,-nbitq), 
to_sfixed(1312.0/65536.0,1,-nbitq), 
to_sfixed(4627.0/65536.0,1,-nbitq), 
to_sfixed(-1151.0/65536.0,1,-nbitq), 
to_sfixed(3774.0/65536.0,1,-nbitq), 
to_sfixed(3327.0/65536.0,1,-nbitq), 
to_sfixed(2786.0/65536.0,1,-nbitq), 
to_sfixed(6521.0/65536.0,1,-nbitq), 
to_sfixed(-4308.0/65536.0,1,-nbitq), 
to_sfixed(1064.0/65536.0,1,-nbitq), 
to_sfixed(6971.0/65536.0,1,-nbitq), 
to_sfixed(7748.0/65536.0,1,-nbitq), 
to_sfixed(-1926.0/65536.0,1,-nbitq), 
to_sfixed(-799.0/65536.0,1,-nbitq), 
to_sfixed(-1647.0/65536.0,1,-nbitq), 
to_sfixed(1440.0/65536.0,1,-nbitq), 
to_sfixed(-1360.0/65536.0,1,-nbitq), 
to_sfixed(-3813.0/65536.0,1,-nbitq), 
to_sfixed(-980.0/65536.0,1,-nbitq), 
to_sfixed(-4094.0/65536.0,1,-nbitq), 
to_sfixed(-4681.0/65536.0,1,-nbitq), 
to_sfixed(-3741.0/65536.0,1,-nbitq), 
to_sfixed(1098.0/65536.0,1,-nbitq), 
to_sfixed(4081.0/65536.0,1,-nbitq), 
to_sfixed(2029.0/65536.0,1,-nbitq), 
to_sfixed(-6798.0/65536.0,1,-nbitq), 
to_sfixed(-4610.0/65536.0,1,-nbitq), 
to_sfixed(-3796.0/65536.0,1,-nbitq), 
to_sfixed(303.0/65536.0,1,-nbitq), 
to_sfixed(-1894.0/65536.0,1,-nbitq), 
to_sfixed(-744.0/65536.0,1,-nbitq), 
to_sfixed(-550.0/65536.0,1,-nbitq), 
to_sfixed(-3122.0/65536.0,1,-nbitq), 
to_sfixed(-3441.0/65536.0,1,-nbitq), 
to_sfixed(-3339.0/65536.0,1,-nbitq), 
to_sfixed(-2748.0/65536.0,1,-nbitq), 
to_sfixed(466.0/65536.0,1,-nbitq), 
to_sfixed(2024.0/65536.0,1,-nbitq), 
to_sfixed(-821.0/65536.0,1,-nbitq), 
to_sfixed(929.0/65536.0,1,-nbitq), 
to_sfixed(-707.0/65536.0,1,-nbitq), 
to_sfixed(4352.0/65536.0,1,-nbitq), 
to_sfixed(6276.0/65536.0,1,-nbitq), 
to_sfixed(-7278.0/65536.0,1,-nbitq), 
to_sfixed(-2449.0/65536.0,1,-nbitq), 
to_sfixed(-3816.0/65536.0,1,-nbitq), 
to_sfixed(837.0/65536.0,1,-nbitq), 
to_sfixed(-2140.0/65536.0,1,-nbitq), 
to_sfixed(2465.0/65536.0,1,-nbitq), 
to_sfixed(7423.0/65536.0,1,-nbitq), 
to_sfixed(6558.0/65536.0,1,-nbitq), 
to_sfixed(-2949.0/65536.0,1,-nbitq), 
to_sfixed(1162.0/65536.0,1,-nbitq), 
to_sfixed(1791.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3060.0/65536.0,1,-nbitq), 
to_sfixed(2360.0/65536.0,1,-nbitq), 
to_sfixed(1767.0/65536.0,1,-nbitq), 
to_sfixed(3310.0/65536.0,1,-nbitq), 
to_sfixed(7868.0/65536.0,1,-nbitq), 
to_sfixed(5525.0/65536.0,1,-nbitq), 
to_sfixed(4091.0/65536.0,1,-nbitq), 
to_sfixed(-2052.0/65536.0,1,-nbitq), 
to_sfixed(-865.0/65536.0,1,-nbitq), 
to_sfixed(-279.0/65536.0,1,-nbitq), 
to_sfixed(2004.0/65536.0,1,-nbitq), 
to_sfixed(-9874.0/65536.0,1,-nbitq), 
to_sfixed(-3165.0/65536.0,1,-nbitq), 
to_sfixed(5734.0/65536.0,1,-nbitq), 
to_sfixed(2314.0/65536.0,1,-nbitq), 
to_sfixed(16.0/65536.0,1,-nbitq), 
to_sfixed(-3055.0/65536.0,1,-nbitq), 
to_sfixed(1053.0/65536.0,1,-nbitq), 
to_sfixed(4.0/65536.0,1,-nbitq), 
to_sfixed(-1197.0/65536.0,1,-nbitq), 
to_sfixed(-4032.0/65536.0,1,-nbitq), 
to_sfixed(3873.0/65536.0,1,-nbitq), 
to_sfixed(315.0/65536.0,1,-nbitq), 
to_sfixed(6162.0/65536.0,1,-nbitq), 
to_sfixed(2137.0/65536.0,1,-nbitq), 
to_sfixed(7769.0/65536.0,1,-nbitq), 
to_sfixed(1791.0/65536.0,1,-nbitq), 
to_sfixed(-2061.0/65536.0,1,-nbitq), 
to_sfixed(-885.0/65536.0,1,-nbitq), 
to_sfixed(-1666.0/65536.0,1,-nbitq), 
to_sfixed(4099.0/65536.0,1,-nbitq), 
to_sfixed(-1652.0/65536.0,1,-nbitq), 
to_sfixed(3977.0/65536.0,1,-nbitq), 
to_sfixed(4429.0/65536.0,1,-nbitq), 
to_sfixed(-3366.0/65536.0,1,-nbitq), 
to_sfixed(-4378.0/65536.0,1,-nbitq), 
to_sfixed(5813.0/65536.0,1,-nbitq), 
to_sfixed(1276.0/65536.0,1,-nbitq), 
to_sfixed(-2448.0/65536.0,1,-nbitq), 
to_sfixed(424.0/65536.0,1,-nbitq), 
to_sfixed(2734.0/65536.0,1,-nbitq), 
to_sfixed(-2379.0/65536.0,1,-nbitq), 
to_sfixed(-2083.0/65536.0,1,-nbitq), 
to_sfixed(-8895.0/65536.0,1,-nbitq), 
to_sfixed(3084.0/65536.0,1,-nbitq), 
to_sfixed(3938.0/65536.0,1,-nbitq), 
to_sfixed(-3248.0/65536.0,1,-nbitq), 
to_sfixed(-4133.0/65536.0,1,-nbitq), 
to_sfixed(945.0/65536.0,1,-nbitq), 
to_sfixed(1654.0/65536.0,1,-nbitq), 
to_sfixed(491.0/65536.0,1,-nbitq), 
to_sfixed(-10119.0/65536.0,1,-nbitq), 
to_sfixed(-9424.0/65536.0,1,-nbitq), 
to_sfixed(872.0/65536.0,1,-nbitq), 
to_sfixed(3879.0/65536.0,1,-nbitq), 
to_sfixed(-1020.0/65536.0,1,-nbitq), 
to_sfixed(726.0/65536.0,1,-nbitq), 
to_sfixed(1097.0/65536.0,1,-nbitq), 
to_sfixed(-191.0/65536.0,1,-nbitq), 
to_sfixed(-7734.0/65536.0,1,-nbitq), 
to_sfixed(-4474.0/65536.0,1,-nbitq), 
to_sfixed(-1432.0/65536.0,1,-nbitq), 
to_sfixed(2879.0/65536.0,1,-nbitq), 
to_sfixed(-2700.0/65536.0,1,-nbitq), 
to_sfixed(-4194.0/65536.0,1,-nbitq), 
to_sfixed(1013.0/65536.0,1,-nbitq), 
to_sfixed(-4043.0/65536.0,1,-nbitq), 
to_sfixed(2388.0/65536.0,1,-nbitq), 
to_sfixed(4643.0/65536.0,1,-nbitq), 
to_sfixed(-9084.0/65536.0,1,-nbitq), 
to_sfixed(-180.0/65536.0,1,-nbitq), 
to_sfixed(-2717.0/65536.0,1,-nbitq), 
to_sfixed(2662.0/65536.0,1,-nbitq), 
to_sfixed(-2638.0/65536.0,1,-nbitq), 
to_sfixed(614.0/65536.0,1,-nbitq), 
to_sfixed(3787.0/65536.0,1,-nbitq), 
to_sfixed(10264.0/65536.0,1,-nbitq), 
to_sfixed(-1923.0/65536.0,1,-nbitq), 
to_sfixed(943.0/65536.0,1,-nbitq), 
to_sfixed(-2619.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2512.0/65536.0,1,-nbitq), 
to_sfixed(-2179.0/65536.0,1,-nbitq), 
to_sfixed(3881.0/65536.0,1,-nbitq), 
to_sfixed(-2346.0/65536.0,1,-nbitq), 
to_sfixed(6417.0/65536.0,1,-nbitq), 
to_sfixed(-94.0/65536.0,1,-nbitq), 
to_sfixed(849.0/65536.0,1,-nbitq), 
to_sfixed(-1974.0/65536.0,1,-nbitq), 
to_sfixed(-1849.0/65536.0,1,-nbitq), 
to_sfixed(921.0/65536.0,1,-nbitq), 
to_sfixed(-1191.0/65536.0,1,-nbitq), 
to_sfixed(-4826.0/65536.0,1,-nbitq), 
to_sfixed(-367.0/65536.0,1,-nbitq), 
to_sfixed(3526.0/65536.0,1,-nbitq), 
to_sfixed(1385.0/65536.0,1,-nbitq), 
to_sfixed(-2912.0/65536.0,1,-nbitq), 
to_sfixed(-3175.0/65536.0,1,-nbitq), 
to_sfixed(-1512.0/65536.0,1,-nbitq), 
to_sfixed(-754.0/65536.0,1,-nbitq), 
to_sfixed(833.0/65536.0,1,-nbitq), 
to_sfixed(-3834.0/65536.0,1,-nbitq), 
to_sfixed(2878.0/65536.0,1,-nbitq), 
to_sfixed(7554.0/65536.0,1,-nbitq), 
to_sfixed(11458.0/65536.0,1,-nbitq), 
to_sfixed(2018.0/65536.0,1,-nbitq), 
to_sfixed(1594.0/65536.0,1,-nbitq), 
to_sfixed(1097.0/65536.0,1,-nbitq), 
to_sfixed(2111.0/65536.0,1,-nbitq), 
to_sfixed(-847.0/65536.0,1,-nbitq), 
to_sfixed(3153.0/65536.0,1,-nbitq), 
to_sfixed(3200.0/65536.0,1,-nbitq), 
to_sfixed(-1267.0/65536.0,1,-nbitq), 
to_sfixed(3582.0/65536.0,1,-nbitq), 
to_sfixed(4345.0/65536.0,1,-nbitq), 
to_sfixed(-2895.0/65536.0,1,-nbitq), 
to_sfixed(-2162.0/65536.0,1,-nbitq), 
to_sfixed(5994.0/65536.0,1,-nbitq), 
to_sfixed(1580.0/65536.0,1,-nbitq), 
to_sfixed(2400.0/65536.0,1,-nbitq), 
to_sfixed(3053.0/65536.0,1,-nbitq), 
to_sfixed(2061.0/65536.0,1,-nbitq), 
to_sfixed(426.0/65536.0,1,-nbitq), 
to_sfixed(-6902.0/65536.0,1,-nbitq), 
to_sfixed(-4428.0/65536.0,1,-nbitq), 
to_sfixed(2395.0/65536.0,1,-nbitq), 
to_sfixed(4734.0/65536.0,1,-nbitq), 
to_sfixed(1363.0/65536.0,1,-nbitq), 
to_sfixed(1282.0/65536.0,1,-nbitq), 
to_sfixed(-2437.0/65536.0,1,-nbitq), 
to_sfixed(-277.0/65536.0,1,-nbitq), 
to_sfixed(1873.0/65536.0,1,-nbitq), 
to_sfixed(-8651.0/65536.0,1,-nbitq), 
to_sfixed(-4827.0/65536.0,1,-nbitq), 
to_sfixed(-1313.0/65536.0,1,-nbitq), 
to_sfixed(2387.0/65536.0,1,-nbitq), 
to_sfixed(2202.0/65536.0,1,-nbitq), 
to_sfixed(-1899.0/65536.0,1,-nbitq), 
to_sfixed(1462.0/65536.0,1,-nbitq), 
to_sfixed(59.0/65536.0,1,-nbitq), 
to_sfixed(116.0/65536.0,1,-nbitq), 
to_sfixed(-2433.0/65536.0,1,-nbitq), 
to_sfixed(1800.0/65536.0,1,-nbitq), 
to_sfixed(-2224.0/65536.0,1,-nbitq), 
to_sfixed(-1296.0/65536.0,1,-nbitq), 
to_sfixed(-3618.0/65536.0,1,-nbitq), 
to_sfixed(-910.0/65536.0,1,-nbitq), 
to_sfixed(-4718.0/65536.0,1,-nbitq), 
to_sfixed(2878.0/65536.0,1,-nbitq), 
to_sfixed(684.0/65536.0,1,-nbitq), 
to_sfixed(-4992.0/65536.0,1,-nbitq), 
to_sfixed(-3272.0/65536.0,1,-nbitq), 
to_sfixed(1343.0/65536.0,1,-nbitq), 
to_sfixed(2331.0/65536.0,1,-nbitq), 
to_sfixed(2683.0/65536.0,1,-nbitq), 
to_sfixed(-262.0/65536.0,1,-nbitq), 
to_sfixed(600.0/65536.0,1,-nbitq), 
to_sfixed(8757.0/65536.0,1,-nbitq), 
to_sfixed(697.0/65536.0,1,-nbitq), 
to_sfixed(-2589.0/65536.0,1,-nbitq), 
to_sfixed(1379.0/65536.0,1,-nbitq)  ), 
( to_sfixed(996.0/65536.0,1,-nbitq), 
to_sfixed(-996.0/65536.0,1,-nbitq), 
to_sfixed(63.0/65536.0,1,-nbitq), 
to_sfixed(-1490.0/65536.0,1,-nbitq), 
to_sfixed(5868.0/65536.0,1,-nbitq), 
to_sfixed(1426.0/65536.0,1,-nbitq), 
to_sfixed(2791.0/65536.0,1,-nbitq), 
to_sfixed(-2603.0/65536.0,1,-nbitq), 
to_sfixed(3159.0/65536.0,1,-nbitq), 
to_sfixed(2237.0/65536.0,1,-nbitq), 
to_sfixed(-3669.0/65536.0,1,-nbitq), 
to_sfixed(2211.0/65536.0,1,-nbitq), 
to_sfixed(-3321.0/65536.0,1,-nbitq), 
to_sfixed(5129.0/65536.0,1,-nbitq), 
to_sfixed(-767.0/65536.0,1,-nbitq), 
to_sfixed(-2409.0/65536.0,1,-nbitq), 
to_sfixed(-1478.0/65536.0,1,-nbitq), 
to_sfixed(-775.0/65536.0,1,-nbitq), 
to_sfixed(-214.0/65536.0,1,-nbitq), 
to_sfixed(-1835.0/65536.0,1,-nbitq), 
to_sfixed(-6665.0/65536.0,1,-nbitq), 
to_sfixed(3495.0/65536.0,1,-nbitq), 
to_sfixed(816.0/65536.0,1,-nbitq), 
to_sfixed(9765.0/65536.0,1,-nbitq), 
to_sfixed(-612.0/65536.0,1,-nbitq), 
to_sfixed(1829.0/65536.0,1,-nbitq), 
to_sfixed(-3481.0/65536.0,1,-nbitq), 
to_sfixed(101.0/65536.0,1,-nbitq), 
to_sfixed(-4376.0/65536.0,1,-nbitq), 
to_sfixed(-1388.0/65536.0,1,-nbitq), 
to_sfixed(-438.0/65536.0,1,-nbitq), 
to_sfixed(-2530.0/65536.0,1,-nbitq), 
to_sfixed(2292.0/65536.0,1,-nbitq), 
to_sfixed(1205.0/65536.0,1,-nbitq), 
to_sfixed(-2079.0/65536.0,1,-nbitq), 
to_sfixed(-564.0/65536.0,1,-nbitq), 
to_sfixed(1631.0/65536.0,1,-nbitq), 
to_sfixed(-2061.0/65536.0,1,-nbitq), 
to_sfixed(1881.0/65536.0,1,-nbitq), 
to_sfixed(-1074.0/65536.0,1,-nbitq), 
to_sfixed(-599.0/65536.0,1,-nbitq), 
to_sfixed(-1781.0/65536.0,1,-nbitq), 
to_sfixed(-7244.0/65536.0,1,-nbitq), 
to_sfixed(-5956.0/65536.0,1,-nbitq), 
to_sfixed(2529.0/65536.0,1,-nbitq), 
to_sfixed(2096.0/65536.0,1,-nbitq), 
to_sfixed(263.0/65536.0,1,-nbitq), 
to_sfixed(3655.0/65536.0,1,-nbitq), 
to_sfixed(-937.0/65536.0,1,-nbitq), 
to_sfixed(2711.0/65536.0,1,-nbitq), 
to_sfixed(30.0/65536.0,1,-nbitq), 
to_sfixed(-4072.0/65536.0,1,-nbitq), 
to_sfixed(-2374.0/65536.0,1,-nbitq), 
to_sfixed(-1737.0/65536.0,1,-nbitq), 
to_sfixed(3477.0/65536.0,1,-nbitq), 
to_sfixed(4199.0/65536.0,1,-nbitq), 
to_sfixed(-125.0/65536.0,1,-nbitq), 
to_sfixed(-164.0/65536.0,1,-nbitq), 
to_sfixed(-1250.0/65536.0,1,-nbitq), 
to_sfixed(31.0/65536.0,1,-nbitq), 
to_sfixed(-832.0/65536.0,1,-nbitq), 
to_sfixed(-2565.0/65536.0,1,-nbitq), 
to_sfixed(-1599.0/65536.0,1,-nbitq), 
to_sfixed(-582.0/65536.0,1,-nbitq), 
to_sfixed(-2608.0/65536.0,1,-nbitq), 
to_sfixed(1681.0/65536.0,1,-nbitq), 
to_sfixed(-4942.0/65536.0,1,-nbitq), 
to_sfixed(-130.0/65536.0,1,-nbitq), 
to_sfixed(-3716.0/65536.0,1,-nbitq), 
to_sfixed(-6595.0/65536.0,1,-nbitq), 
to_sfixed(76.0/65536.0,1,-nbitq), 
to_sfixed(-734.0/65536.0,1,-nbitq), 
to_sfixed(1400.0/65536.0,1,-nbitq), 
to_sfixed(-832.0/65536.0,1,-nbitq), 
to_sfixed(711.0/65536.0,1,-nbitq), 
to_sfixed(-274.0/65536.0,1,-nbitq), 
to_sfixed(6586.0/65536.0,1,-nbitq), 
to_sfixed(3144.0/65536.0,1,-nbitq), 
to_sfixed(-658.0/65536.0,1,-nbitq), 
to_sfixed(3815.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-115.0/65536.0,1,-nbitq), 
to_sfixed(449.0/65536.0,1,-nbitq), 
to_sfixed(2938.0/65536.0,1,-nbitq), 
to_sfixed(-4480.0/65536.0,1,-nbitq), 
to_sfixed(1630.0/65536.0,1,-nbitq), 
to_sfixed(-1738.0/65536.0,1,-nbitq), 
to_sfixed(-1563.0/65536.0,1,-nbitq), 
to_sfixed(-5261.0/65536.0,1,-nbitq), 
to_sfixed(-3838.0/65536.0,1,-nbitq), 
to_sfixed(-1566.0/65536.0,1,-nbitq), 
to_sfixed(724.0/65536.0,1,-nbitq), 
to_sfixed(241.0/65536.0,1,-nbitq), 
to_sfixed(1020.0/65536.0,1,-nbitq), 
to_sfixed(1179.0/65536.0,1,-nbitq), 
to_sfixed(310.0/65536.0,1,-nbitq), 
to_sfixed(-1182.0/65536.0,1,-nbitq), 
to_sfixed(-1697.0/65536.0,1,-nbitq), 
to_sfixed(-3459.0/65536.0,1,-nbitq), 
to_sfixed(987.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(-4901.0/65536.0,1,-nbitq), 
to_sfixed(730.0/65536.0,1,-nbitq), 
to_sfixed(86.0/65536.0,1,-nbitq), 
to_sfixed(6757.0/65536.0,1,-nbitq), 
to_sfixed(269.0/65536.0,1,-nbitq), 
to_sfixed(3622.0/65536.0,1,-nbitq), 
to_sfixed(-2318.0/65536.0,1,-nbitq), 
to_sfixed(1523.0/65536.0,1,-nbitq), 
to_sfixed(-2475.0/65536.0,1,-nbitq), 
to_sfixed(2577.0/65536.0,1,-nbitq), 
to_sfixed(-3064.0/65536.0,1,-nbitq), 
to_sfixed(1127.0/65536.0,1,-nbitq), 
to_sfixed(443.0/65536.0,1,-nbitq), 
to_sfixed(1258.0/65536.0,1,-nbitq), 
to_sfixed(-1946.0/65536.0,1,-nbitq), 
to_sfixed(1276.0/65536.0,1,-nbitq), 
to_sfixed(4705.0/65536.0,1,-nbitq), 
to_sfixed(-387.0/65536.0,1,-nbitq), 
to_sfixed(835.0/65536.0,1,-nbitq), 
to_sfixed(1439.0/65536.0,1,-nbitq), 
to_sfixed(-3959.0/65536.0,1,-nbitq), 
to_sfixed(-1310.0/65536.0,1,-nbitq), 
to_sfixed(-5302.0/65536.0,1,-nbitq), 
to_sfixed(-871.0/65536.0,1,-nbitq), 
to_sfixed(-2020.0/65536.0,1,-nbitq), 
to_sfixed(2432.0/65536.0,1,-nbitq), 
to_sfixed(597.0/65536.0,1,-nbitq), 
to_sfixed(3547.0/65536.0,1,-nbitq), 
to_sfixed(3354.0/65536.0,1,-nbitq), 
to_sfixed(4006.0/65536.0,1,-nbitq), 
to_sfixed(857.0/65536.0,1,-nbitq), 
to_sfixed(-2928.0/65536.0,1,-nbitq), 
to_sfixed(-1036.0/65536.0,1,-nbitq), 
to_sfixed(-1499.0/65536.0,1,-nbitq), 
to_sfixed(2159.0/65536.0,1,-nbitq), 
to_sfixed(2569.0/65536.0,1,-nbitq), 
to_sfixed(-640.0/65536.0,1,-nbitq), 
to_sfixed(-1186.0/65536.0,1,-nbitq), 
to_sfixed(512.0/65536.0,1,-nbitq), 
to_sfixed(1266.0/65536.0,1,-nbitq), 
to_sfixed(2564.0/65536.0,1,-nbitq), 
to_sfixed(-2855.0/65536.0,1,-nbitq), 
to_sfixed(-2150.0/65536.0,1,-nbitq), 
to_sfixed(-2516.0/65536.0,1,-nbitq), 
to_sfixed(-39.0/65536.0,1,-nbitq), 
to_sfixed(-1537.0/65536.0,1,-nbitq), 
to_sfixed(-6026.0/65536.0,1,-nbitq), 
to_sfixed(-6442.0/65536.0,1,-nbitq), 
to_sfixed(-1260.0/65536.0,1,-nbitq), 
to_sfixed(-6465.0/65536.0,1,-nbitq), 
to_sfixed(1586.0/65536.0,1,-nbitq), 
to_sfixed(76.0/65536.0,1,-nbitq), 
to_sfixed(41.0/65536.0,1,-nbitq), 
to_sfixed(1981.0/65536.0,1,-nbitq), 
to_sfixed(2067.0/65536.0,1,-nbitq), 
to_sfixed(-3585.0/65536.0,1,-nbitq), 
to_sfixed(222.0/65536.0,1,-nbitq), 
to_sfixed(-2850.0/65536.0,1,-nbitq), 
to_sfixed(-529.0/65536.0,1,-nbitq), 
to_sfixed(270.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2661.0/65536.0,1,-nbitq), 
to_sfixed(-1292.0/65536.0,1,-nbitq), 
to_sfixed(4602.0/65536.0,1,-nbitq), 
to_sfixed(-1254.0/65536.0,1,-nbitq), 
to_sfixed(85.0/65536.0,1,-nbitq), 
to_sfixed(302.0/65536.0,1,-nbitq), 
to_sfixed(49.0/65536.0,1,-nbitq), 
to_sfixed(-3299.0/65536.0,1,-nbitq), 
to_sfixed(-3537.0/65536.0,1,-nbitq), 
to_sfixed(984.0/65536.0,1,-nbitq), 
to_sfixed(-227.0/65536.0,1,-nbitq), 
to_sfixed(3966.0/65536.0,1,-nbitq), 
to_sfixed(2336.0/65536.0,1,-nbitq), 
to_sfixed(-872.0/65536.0,1,-nbitq), 
to_sfixed(691.0/65536.0,1,-nbitq), 
to_sfixed(196.0/65536.0,1,-nbitq), 
to_sfixed(-1197.0/65536.0,1,-nbitq), 
to_sfixed(109.0/65536.0,1,-nbitq), 
to_sfixed(1341.0/65536.0,1,-nbitq), 
to_sfixed(-1957.0/65536.0,1,-nbitq), 
to_sfixed(-757.0/65536.0,1,-nbitq), 
to_sfixed(395.0/65536.0,1,-nbitq), 
to_sfixed(604.0/65536.0,1,-nbitq), 
to_sfixed(1519.0/65536.0,1,-nbitq), 
to_sfixed(-2473.0/65536.0,1,-nbitq), 
to_sfixed(-1088.0/65536.0,1,-nbitq), 
to_sfixed(-3655.0/65536.0,1,-nbitq), 
to_sfixed(-2066.0/65536.0,1,-nbitq), 
to_sfixed(-1784.0/65536.0,1,-nbitq), 
to_sfixed(-2280.0/65536.0,1,-nbitq), 
to_sfixed(786.0/65536.0,1,-nbitq), 
to_sfixed(-791.0/65536.0,1,-nbitq), 
to_sfixed(-338.0/65536.0,1,-nbitq), 
to_sfixed(1642.0/65536.0,1,-nbitq), 
to_sfixed(1700.0/65536.0,1,-nbitq), 
to_sfixed(-1930.0/65536.0,1,-nbitq), 
to_sfixed(-427.0/65536.0,1,-nbitq), 
to_sfixed(1525.0/65536.0,1,-nbitq), 
to_sfixed(-1473.0/65536.0,1,-nbitq), 
to_sfixed(-1154.0/65536.0,1,-nbitq), 
to_sfixed(-4117.0/65536.0,1,-nbitq), 
to_sfixed(-2739.0/65536.0,1,-nbitq), 
to_sfixed(-3369.0/65536.0,1,-nbitq), 
to_sfixed(-494.0/65536.0,1,-nbitq), 
to_sfixed(-419.0/65536.0,1,-nbitq), 
to_sfixed(4067.0/65536.0,1,-nbitq), 
to_sfixed(-192.0/65536.0,1,-nbitq), 
to_sfixed(-82.0/65536.0,1,-nbitq), 
to_sfixed(-2021.0/65536.0,1,-nbitq), 
to_sfixed(3820.0/65536.0,1,-nbitq), 
to_sfixed(-2056.0/65536.0,1,-nbitq), 
to_sfixed(-2561.0/65536.0,1,-nbitq), 
to_sfixed(-1122.0/65536.0,1,-nbitq), 
to_sfixed(-2344.0/65536.0,1,-nbitq), 
to_sfixed(4987.0/65536.0,1,-nbitq), 
to_sfixed(2254.0/65536.0,1,-nbitq), 
to_sfixed(-757.0/65536.0,1,-nbitq), 
to_sfixed(-2890.0/65536.0,1,-nbitq), 
to_sfixed(-1851.0/65536.0,1,-nbitq), 
to_sfixed(779.0/65536.0,1,-nbitq), 
to_sfixed(2056.0/65536.0,1,-nbitq), 
to_sfixed(-2695.0/65536.0,1,-nbitq), 
to_sfixed(-519.0/65536.0,1,-nbitq), 
to_sfixed(2363.0/65536.0,1,-nbitq), 
to_sfixed(1178.0/65536.0,1,-nbitq), 
to_sfixed(1191.0/65536.0,1,-nbitq), 
to_sfixed(-1755.0/65536.0,1,-nbitq), 
to_sfixed(-5468.0/65536.0,1,-nbitq), 
to_sfixed(245.0/65536.0,1,-nbitq), 
to_sfixed(-3258.0/65536.0,1,-nbitq), 
to_sfixed(294.0/65536.0,1,-nbitq), 
to_sfixed(-5752.0/65536.0,1,-nbitq), 
to_sfixed(-2620.0/65536.0,1,-nbitq), 
to_sfixed(1090.0/65536.0,1,-nbitq), 
to_sfixed(1154.0/65536.0,1,-nbitq), 
to_sfixed(2548.0/65536.0,1,-nbitq), 
to_sfixed(-1489.0/65536.0,1,-nbitq), 
to_sfixed(262.0/65536.0,1,-nbitq), 
to_sfixed(-2073.0/65536.0,1,-nbitq), 
to_sfixed(782.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1937.0/65536.0,1,-nbitq), 
to_sfixed(641.0/65536.0,1,-nbitq), 
to_sfixed(623.0/65536.0,1,-nbitq), 
to_sfixed(-4006.0/65536.0,1,-nbitq), 
to_sfixed(-1871.0/65536.0,1,-nbitq), 
to_sfixed(749.0/65536.0,1,-nbitq), 
to_sfixed(-1196.0/65536.0,1,-nbitq), 
to_sfixed(-410.0/65536.0,1,-nbitq), 
to_sfixed(1270.0/65536.0,1,-nbitq), 
to_sfixed(2863.0/65536.0,1,-nbitq), 
to_sfixed(1882.0/65536.0,1,-nbitq), 
to_sfixed(423.0/65536.0,1,-nbitq), 
to_sfixed(1785.0/65536.0,1,-nbitq), 
to_sfixed(527.0/65536.0,1,-nbitq), 
to_sfixed(-64.0/65536.0,1,-nbitq), 
to_sfixed(78.0/65536.0,1,-nbitq), 
to_sfixed(-593.0/65536.0,1,-nbitq), 
to_sfixed(2299.0/65536.0,1,-nbitq), 
to_sfixed(2862.0/65536.0,1,-nbitq), 
to_sfixed(1658.0/65536.0,1,-nbitq), 
to_sfixed(-2675.0/65536.0,1,-nbitq), 
to_sfixed(-1442.0/65536.0,1,-nbitq), 
to_sfixed(1192.0/65536.0,1,-nbitq), 
to_sfixed(-541.0/65536.0,1,-nbitq), 
to_sfixed(1838.0/65536.0,1,-nbitq), 
to_sfixed(-1703.0/65536.0,1,-nbitq), 
to_sfixed(-3636.0/65536.0,1,-nbitq), 
to_sfixed(-743.0/65536.0,1,-nbitq), 
to_sfixed(1548.0/65536.0,1,-nbitq), 
to_sfixed(87.0/65536.0,1,-nbitq), 
to_sfixed(1161.0/65536.0,1,-nbitq), 
to_sfixed(-1437.0/65536.0,1,-nbitq), 
to_sfixed(176.0/65536.0,1,-nbitq), 
to_sfixed(1461.0/65536.0,1,-nbitq), 
to_sfixed(1948.0/65536.0,1,-nbitq), 
to_sfixed(330.0/65536.0,1,-nbitq), 
to_sfixed(343.0/65536.0,1,-nbitq), 
to_sfixed(-1819.0/65536.0,1,-nbitq), 
to_sfixed(353.0/65536.0,1,-nbitq), 
to_sfixed(-652.0/65536.0,1,-nbitq), 
to_sfixed(-5587.0/65536.0,1,-nbitq), 
to_sfixed(-993.0/65536.0,1,-nbitq), 
to_sfixed(-340.0/65536.0,1,-nbitq), 
to_sfixed(2781.0/65536.0,1,-nbitq), 
to_sfixed(-902.0/65536.0,1,-nbitq), 
to_sfixed(3704.0/65536.0,1,-nbitq), 
to_sfixed(3556.0/65536.0,1,-nbitq), 
to_sfixed(923.0/65536.0,1,-nbitq), 
to_sfixed(-2303.0/65536.0,1,-nbitq), 
to_sfixed(521.0/65536.0,1,-nbitq), 
to_sfixed(-97.0/65536.0,1,-nbitq), 
to_sfixed(-2037.0/65536.0,1,-nbitq), 
to_sfixed(3582.0/65536.0,1,-nbitq), 
to_sfixed(601.0/65536.0,1,-nbitq), 
to_sfixed(592.0/65536.0,1,-nbitq), 
to_sfixed(371.0/65536.0,1,-nbitq), 
to_sfixed(-1655.0/65536.0,1,-nbitq), 
to_sfixed(684.0/65536.0,1,-nbitq), 
to_sfixed(-264.0/65536.0,1,-nbitq), 
to_sfixed(677.0/65536.0,1,-nbitq), 
to_sfixed(-3253.0/65536.0,1,-nbitq), 
to_sfixed(-920.0/65536.0,1,-nbitq), 
to_sfixed(-2717.0/65536.0,1,-nbitq), 
to_sfixed(736.0/65536.0,1,-nbitq), 
to_sfixed(691.0/65536.0,1,-nbitq), 
to_sfixed(994.0/65536.0,1,-nbitq), 
to_sfixed(-330.0/65536.0,1,-nbitq), 
to_sfixed(-85.0/65536.0,1,-nbitq), 
to_sfixed(-3226.0/65536.0,1,-nbitq), 
to_sfixed(-1736.0/65536.0,1,-nbitq), 
to_sfixed(-980.0/65536.0,1,-nbitq), 
to_sfixed(11.0/65536.0,1,-nbitq), 
to_sfixed(-988.0/65536.0,1,-nbitq), 
to_sfixed(-2592.0/65536.0,1,-nbitq), 
to_sfixed(981.0/65536.0,1,-nbitq), 
to_sfixed(2613.0/65536.0,1,-nbitq), 
to_sfixed(1712.0/65536.0,1,-nbitq), 
to_sfixed(3910.0/65536.0,1,-nbitq), 
to_sfixed(262.0/65536.0,1,-nbitq), 
to_sfixed(527.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1187.0/65536.0,1,-nbitq), 
to_sfixed(-1641.0/65536.0,1,-nbitq), 
to_sfixed(1104.0/65536.0,1,-nbitq), 
to_sfixed(-1902.0/65536.0,1,-nbitq), 
to_sfixed(-605.0/65536.0,1,-nbitq), 
to_sfixed(115.0/65536.0,1,-nbitq), 
to_sfixed(-1159.0/65536.0,1,-nbitq), 
to_sfixed(-2272.0/65536.0,1,-nbitq), 
to_sfixed(-3122.0/65536.0,1,-nbitq), 
to_sfixed(1380.0/65536.0,1,-nbitq), 
to_sfixed(-357.0/65536.0,1,-nbitq), 
to_sfixed(1382.0/65536.0,1,-nbitq), 
to_sfixed(59.0/65536.0,1,-nbitq), 
to_sfixed(138.0/65536.0,1,-nbitq), 
to_sfixed(1890.0/65536.0,1,-nbitq), 
to_sfixed(-2114.0/65536.0,1,-nbitq), 
to_sfixed(510.0/65536.0,1,-nbitq), 
to_sfixed(1108.0/65536.0,1,-nbitq), 
to_sfixed(1813.0/65536.0,1,-nbitq), 
to_sfixed(160.0/65536.0,1,-nbitq), 
to_sfixed(-1451.0/65536.0,1,-nbitq), 
to_sfixed(-2479.0/65536.0,1,-nbitq), 
to_sfixed(35.0/65536.0,1,-nbitq), 
to_sfixed(80.0/65536.0,1,-nbitq), 
to_sfixed(1726.0/65536.0,1,-nbitq), 
to_sfixed(-1179.0/65536.0,1,-nbitq), 
to_sfixed(-2708.0/65536.0,1,-nbitq), 
to_sfixed(-1270.0/65536.0,1,-nbitq), 
to_sfixed(1167.0/65536.0,1,-nbitq), 
to_sfixed(-2105.0/65536.0,1,-nbitq), 
to_sfixed(2480.0/65536.0,1,-nbitq), 
to_sfixed(-816.0/65536.0,1,-nbitq), 
to_sfixed(-884.0/65536.0,1,-nbitq), 
to_sfixed(-124.0/65536.0,1,-nbitq), 
to_sfixed(-583.0/65536.0,1,-nbitq), 
to_sfixed(763.0/65536.0,1,-nbitq), 
to_sfixed(519.0/65536.0,1,-nbitq), 
to_sfixed(-438.0/65536.0,1,-nbitq), 
to_sfixed(-1898.0/65536.0,1,-nbitq), 
to_sfixed(3042.0/65536.0,1,-nbitq), 
to_sfixed(-1265.0/65536.0,1,-nbitq), 
to_sfixed(-3291.0/65536.0,1,-nbitq), 
to_sfixed(-4408.0/65536.0,1,-nbitq), 
to_sfixed(-720.0/65536.0,1,-nbitq), 
to_sfixed(2821.0/65536.0,1,-nbitq), 
to_sfixed(3757.0/65536.0,1,-nbitq), 
to_sfixed(-237.0/65536.0,1,-nbitq), 
to_sfixed(-984.0/65536.0,1,-nbitq), 
to_sfixed(2318.0/65536.0,1,-nbitq), 
to_sfixed(644.0/65536.0,1,-nbitq), 
to_sfixed(1783.0/65536.0,1,-nbitq), 
to_sfixed(774.0/65536.0,1,-nbitq), 
to_sfixed(874.0/65536.0,1,-nbitq), 
to_sfixed(-3004.0/65536.0,1,-nbitq), 
to_sfixed(1299.0/65536.0,1,-nbitq), 
to_sfixed(3946.0/65536.0,1,-nbitq), 
to_sfixed(3060.0/65536.0,1,-nbitq), 
to_sfixed(1278.0/65536.0,1,-nbitq), 
to_sfixed(2400.0/65536.0,1,-nbitq), 
to_sfixed(5838.0/65536.0,1,-nbitq), 
to_sfixed(1274.0/65536.0,1,-nbitq), 
to_sfixed(-2922.0/65536.0,1,-nbitq), 
to_sfixed(1919.0/65536.0,1,-nbitq), 
to_sfixed(2490.0/65536.0,1,-nbitq), 
to_sfixed(-1289.0/65536.0,1,-nbitq), 
to_sfixed(-1335.0/65536.0,1,-nbitq), 
to_sfixed(-2247.0/65536.0,1,-nbitq), 
to_sfixed(-1714.0/65536.0,1,-nbitq), 
to_sfixed(1318.0/65536.0,1,-nbitq), 
to_sfixed(2681.0/65536.0,1,-nbitq), 
to_sfixed(3246.0/65536.0,1,-nbitq), 
to_sfixed(-1625.0/65536.0,1,-nbitq), 
to_sfixed(1456.0/65536.0,1,-nbitq), 
to_sfixed(1602.0/65536.0,1,-nbitq), 
to_sfixed(492.0/65536.0,1,-nbitq), 
to_sfixed(614.0/65536.0,1,-nbitq), 
to_sfixed(1207.0/65536.0,1,-nbitq), 
to_sfixed(2997.0/65536.0,1,-nbitq), 
to_sfixed(-2294.0/65536.0,1,-nbitq), 
to_sfixed(467.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1475.0/65536.0,1,-nbitq), 
to_sfixed(-767.0/65536.0,1,-nbitq), 
to_sfixed(827.0/65536.0,1,-nbitq), 
to_sfixed(-2692.0/65536.0,1,-nbitq), 
to_sfixed(-1342.0/65536.0,1,-nbitq), 
to_sfixed(-328.0/65536.0,1,-nbitq), 
to_sfixed(-1056.0/65536.0,1,-nbitq), 
to_sfixed(28.0/65536.0,1,-nbitq), 
to_sfixed(1077.0/65536.0,1,-nbitq), 
to_sfixed(3042.0/65536.0,1,-nbitq), 
to_sfixed(-2458.0/65536.0,1,-nbitq), 
to_sfixed(1192.0/65536.0,1,-nbitq), 
to_sfixed(952.0/65536.0,1,-nbitq), 
to_sfixed(1322.0/65536.0,1,-nbitq), 
to_sfixed(3399.0/65536.0,1,-nbitq), 
to_sfixed(1067.0/65536.0,1,-nbitq), 
to_sfixed(2719.0/65536.0,1,-nbitq), 
to_sfixed(-204.0/65536.0,1,-nbitq), 
to_sfixed(2785.0/65536.0,1,-nbitq), 
to_sfixed(3344.0/65536.0,1,-nbitq), 
to_sfixed(-3344.0/65536.0,1,-nbitq), 
to_sfixed(-2518.0/65536.0,1,-nbitq), 
to_sfixed(2036.0/65536.0,1,-nbitq), 
to_sfixed(2787.0/65536.0,1,-nbitq), 
to_sfixed(-1811.0/65536.0,1,-nbitq), 
to_sfixed(-891.0/65536.0,1,-nbitq), 
to_sfixed(-1096.0/65536.0,1,-nbitq), 
to_sfixed(-2564.0/65536.0,1,-nbitq), 
to_sfixed(-831.0/65536.0,1,-nbitq), 
to_sfixed(-1746.0/65536.0,1,-nbitq), 
to_sfixed(-2403.0/65536.0,1,-nbitq), 
to_sfixed(2458.0/65536.0,1,-nbitq), 
to_sfixed(-2190.0/65536.0,1,-nbitq), 
to_sfixed(-4534.0/65536.0,1,-nbitq), 
to_sfixed(1052.0/65536.0,1,-nbitq), 
to_sfixed(-1953.0/65536.0,1,-nbitq), 
to_sfixed(2643.0/65536.0,1,-nbitq), 
to_sfixed(-411.0/65536.0,1,-nbitq), 
to_sfixed(-1308.0/65536.0,1,-nbitq), 
to_sfixed(2626.0/65536.0,1,-nbitq), 
to_sfixed(-3828.0/65536.0,1,-nbitq), 
to_sfixed(-51.0/65536.0,1,-nbitq), 
to_sfixed(-1738.0/65536.0,1,-nbitq), 
to_sfixed(63.0/65536.0,1,-nbitq), 
to_sfixed(-753.0/65536.0,1,-nbitq), 
to_sfixed(4131.0/65536.0,1,-nbitq), 
to_sfixed(-1367.0/65536.0,1,-nbitq), 
to_sfixed(-317.0/65536.0,1,-nbitq), 
to_sfixed(3148.0/65536.0,1,-nbitq), 
to_sfixed(1923.0/65536.0,1,-nbitq), 
to_sfixed(-1829.0/65536.0,1,-nbitq), 
to_sfixed(196.0/65536.0,1,-nbitq), 
to_sfixed(3106.0/65536.0,1,-nbitq), 
to_sfixed(-1432.0/65536.0,1,-nbitq), 
to_sfixed(626.0/65536.0,1,-nbitq), 
to_sfixed(-1759.0/65536.0,1,-nbitq), 
to_sfixed(2535.0/65536.0,1,-nbitq), 
to_sfixed(-2282.0/65536.0,1,-nbitq), 
to_sfixed(1582.0/65536.0,1,-nbitq), 
to_sfixed(5025.0/65536.0,1,-nbitq), 
to_sfixed(-875.0/65536.0,1,-nbitq), 
to_sfixed(-774.0/65536.0,1,-nbitq), 
to_sfixed(159.0/65536.0,1,-nbitq), 
to_sfixed(-1135.0/65536.0,1,-nbitq), 
to_sfixed(3339.0/65536.0,1,-nbitq), 
to_sfixed(-461.0/65536.0,1,-nbitq), 
to_sfixed(328.0/65536.0,1,-nbitq), 
to_sfixed(-1392.0/65536.0,1,-nbitq), 
to_sfixed(-1650.0/65536.0,1,-nbitq), 
to_sfixed(434.0/65536.0,1,-nbitq), 
to_sfixed(-1071.0/65536.0,1,-nbitq), 
to_sfixed(643.0/65536.0,1,-nbitq), 
to_sfixed(2600.0/65536.0,1,-nbitq), 
to_sfixed(-2374.0/65536.0,1,-nbitq), 
to_sfixed(-2924.0/65536.0,1,-nbitq), 
to_sfixed(-720.0/65536.0,1,-nbitq), 
to_sfixed(-2868.0/65536.0,1,-nbitq), 
to_sfixed(401.0/65536.0,1,-nbitq), 
to_sfixed(-89.0/65536.0,1,-nbitq), 
to_sfixed(3262.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2079.0/65536.0,1,-nbitq), 
to_sfixed(2607.0/65536.0,1,-nbitq), 
to_sfixed(-540.0/65536.0,1,-nbitq), 
to_sfixed(-26.0/65536.0,1,-nbitq), 
to_sfixed(-3418.0/65536.0,1,-nbitq), 
to_sfixed(-2296.0/65536.0,1,-nbitq), 
to_sfixed(-465.0/65536.0,1,-nbitq), 
to_sfixed(-2890.0/65536.0,1,-nbitq), 
to_sfixed(-3314.0/65536.0,1,-nbitq), 
to_sfixed(-2388.0/65536.0,1,-nbitq), 
to_sfixed(-2003.0/65536.0,1,-nbitq), 
to_sfixed(-2875.0/65536.0,1,-nbitq), 
to_sfixed(-1095.0/65536.0,1,-nbitq), 
to_sfixed(-1896.0/65536.0,1,-nbitq), 
to_sfixed(2215.0/65536.0,1,-nbitq), 
to_sfixed(3019.0/65536.0,1,-nbitq), 
to_sfixed(-948.0/65536.0,1,-nbitq), 
to_sfixed(3382.0/65536.0,1,-nbitq), 
to_sfixed(-310.0/65536.0,1,-nbitq), 
to_sfixed(-2150.0/65536.0,1,-nbitq), 
to_sfixed(-560.0/65536.0,1,-nbitq), 
to_sfixed(-2857.0/65536.0,1,-nbitq), 
to_sfixed(836.0/65536.0,1,-nbitq), 
to_sfixed(2423.0/65536.0,1,-nbitq), 
to_sfixed(800.0/65536.0,1,-nbitq), 
to_sfixed(1293.0/65536.0,1,-nbitq), 
to_sfixed(-2977.0/65536.0,1,-nbitq), 
to_sfixed(1921.0/65536.0,1,-nbitq), 
to_sfixed(-3607.0/65536.0,1,-nbitq), 
to_sfixed(-2642.0/65536.0,1,-nbitq), 
to_sfixed(372.0/65536.0,1,-nbitq), 
to_sfixed(-1569.0/65536.0,1,-nbitq), 
to_sfixed(-4036.0/65536.0,1,-nbitq), 
to_sfixed(-3832.0/65536.0,1,-nbitq), 
to_sfixed(-930.0/65536.0,1,-nbitq), 
to_sfixed(-1990.0/65536.0,1,-nbitq), 
to_sfixed(-1715.0/65536.0,1,-nbitq), 
to_sfixed(-2924.0/65536.0,1,-nbitq), 
to_sfixed(-2160.0/65536.0,1,-nbitq), 
to_sfixed(715.0/65536.0,1,-nbitq), 
to_sfixed(-87.0/65536.0,1,-nbitq), 
to_sfixed(-1991.0/65536.0,1,-nbitq), 
to_sfixed(-4017.0/65536.0,1,-nbitq), 
to_sfixed(3135.0/65536.0,1,-nbitq), 
to_sfixed(1950.0/65536.0,1,-nbitq), 
to_sfixed(1609.0/65536.0,1,-nbitq), 
to_sfixed(-2335.0/65536.0,1,-nbitq), 
to_sfixed(-2196.0/65536.0,1,-nbitq), 
to_sfixed(1526.0/65536.0,1,-nbitq), 
to_sfixed(1468.0/65536.0,1,-nbitq), 
to_sfixed(2099.0/65536.0,1,-nbitq), 
to_sfixed(1759.0/65536.0,1,-nbitq), 
to_sfixed(-1223.0/65536.0,1,-nbitq), 
to_sfixed(1701.0/65536.0,1,-nbitq), 
to_sfixed(352.0/65536.0,1,-nbitq), 
to_sfixed(649.0/65536.0,1,-nbitq), 
to_sfixed(-1225.0/65536.0,1,-nbitq), 
to_sfixed(-995.0/65536.0,1,-nbitq), 
to_sfixed(-550.0/65536.0,1,-nbitq), 
to_sfixed(4892.0/65536.0,1,-nbitq), 
to_sfixed(-57.0/65536.0,1,-nbitq), 
to_sfixed(-2656.0/65536.0,1,-nbitq), 
to_sfixed(3154.0/65536.0,1,-nbitq), 
to_sfixed(1278.0/65536.0,1,-nbitq), 
to_sfixed(-522.0/65536.0,1,-nbitq), 
to_sfixed(-491.0/65536.0,1,-nbitq), 
to_sfixed(2899.0/65536.0,1,-nbitq), 
to_sfixed(-944.0/65536.0,1,-nbitq), 
to_sfixed(-1819.0/65536.0,1,-nbitq), 
to_sfixed(2793.0/65536.0,1,-nbitq), 
to_sfixed(1276.0/65536.0,1,-nbitq), 
to_sfixed(155.0/65536.0,1,-nbitq), 
to_sfixed(1385.0/65536.0,1,-nbitq), 
to_sfixed(1501.0/65536.0,1,-nbitq), 
to_sfixed(1122.0/65536.0,1,-nbitq), 
to_sfixed(1855.0/65536.0,1,-nbitq), 
to_sfixed(2108.0/65536.0,1,-nbitq), 
to_sfixed(3257.0/65536.0,1,-nbitq), 
to_sfixed(-1400.0/65536.0,1,-nbitq), 
to_sfixed(228.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-607.0/65536.0,1,-nbitq), 
to_sfixed(1292.0/65536.0,1,-nbitq), 
to_sfixed(2110.0/65536.0,1,-nbitq), 
to_sfixed(-494.0/65536.0,1,-nbitq), 
to_sfixed(878.0/65536.0,1,-nbitq), 
to_sfixed(-2555.0/65536.0,1,-nbitq), 
to_sfixed(2111.0/65536.0,1,-nbitq), 
to_sfixed(-283.0/65536.0,1,-nbitq), 
to_sfixed(-374.0/65536.0,1,-nbitq), 
to_sfixed(2986.0/65536.0,1,-nbitq), 
to_sfixed(2048.0/65536.0,1,-nbitq), 
to_sfixed(2554.0/65536.0,1,-nbitq), 
to_sfixed(1388.0/65536.0,1,-nbitq), 
to_sfixed(-2207.0/65536.0,1,-nbitq), 
to_sfixed(1051.0/65536.0,1,-nbitq), 
to_sfixed(-2482.0/65536.0,1,-nbitq), 
to_sfixed(-2347.0/65536.0,1,-nbitq), 
to_sfixed(2444.0/65536.0,1,-nbitq), 
to_sfixed(3616.0/65536.0,1,-nbitq), 
to_sfixed(3430.0/65536.0,1,-nbitq), 
to_sfixed(-179.0/65536.0,1,-nbitq), 
to_sfixed(-1754.0/65536.0,1,-nbitq), 
to_sfixed(-569.0/65536.0,1,-nbitq), 
to_sfixed(4313.0/65536.0,1,-nbitq), 
to_sfixed(-2021.0/65536.0,1,-nbitq), 
to_sfixed(2731.0/65536.0,1,-nbitq), 
to_sfixed(-3913.0/65536.0,1,-nbitq), 
to_sfixed(-1665.0/65536.0,1,-nbitq), 
to_sfixed(2126.0/65536.0,1,-nbitq), 
to_sfixed(-1017.0/65536.0,1,-nbitq), 
to_sfixed(-1099.0/65536.0,1,-nbitq), 
to_sfixed(-1302.0/65536.0,1,-nbitq), 
to_sfixed(-2487.0/65536.0,1,-nbitq), 
to_sfixed(-5711.0/65536.0,1,-nbitq), 
to_sfixed(-2202.0/65536.0,1,-nbitq), 
to_sfixed(-2941.0/65536.0,1,-nbitq), 
to_sfixed(-1694.0/65536.0,1,-nbitq), 
to_sfixed(-3173.0/65536.0,1,-nbitq), 
to_sfixed(-415.0/65536.0,1,-nbitq), 
to_sfixed(-2457.0/65536.0,1,-nbitq), 
to_sfixed(-1143.0/65536.0,1,-nbitq), 
to_sfixed(-310.0/65536.0,1,-nbitq), 
to_sfixed(-1390.0/65536.0,1,-nbitq), 
to_sfixed(82.0/65536.0,1,-nbitq), 
to_sfixed(-1665.0/65536.0,1,-nbitq), 
to_sfixed(-450.0/65536.0,1,-nbitq), 
to_sfixed(1520.0/65536.0,1,-nbitq), 
to_sfixed(-121.0/65536.0,1,-nbitq), 
to_sfixed(-765.0/65536.0,1,-nbitq), 
to_sfixed(1208.0/65536.0,1,-nbitq), 
to_sfixed(-1577.0/65536.0,1,-nbitq), 
to_sfixed(-1056.0/65536.0,1,-nbitq), 
to_sfixed(1942.0/65536.0,1,-nbitq), 
to_sfixed(-2083.0/65536.0,1,-nbitq), 
to_sfixed(869.0/65536.0,1,-nbitq), 
to_sfixed(-1016.0/65536.0,1,-nbitq), 
to_sfixed(1668.0/65536.0,1,-nbitq), 
to_sfixed(2068.0/65536.0,1,-nbitq), 
to_sfixed(-2784.0/65536.0,1,-nbitq), 
to_sfixed(5538.0/65536.0,1,-nbitq), 
to_sfixed(-3436.0/65536.0,1,-nbitq), 
to_sfixed(1425.0/65536.0,1,-nbitq), 
to_sfixed(3040.0/65536.0,1,-nbitq), 
to_sfixed(-920.0/65536.0,1,-nbitq), 
to_sfixed(-172.0/65536.0,1,-nbitq), 
to_sfixed(144.0/65536.0,1,-nbitq), 
to_sfixed(-1770.0/65536.0,1,-nbitq), 
to_sfixed(-3763.0/65536.0,1,-nbitq), 
to_sfixed(-926.0/65536.0,1,-nbitq), 
to_sfixed(379.0/65536.0,1,-nbitq), 
to_sfixed(324.0/65536.0,1,-nbitq), 
to_sfixed(-2676.0/65536.0,1,-nbitq), 
to_sfixed(-1593.0/65536.0,1,-nbitq), 
to_sfixed(-2753.0/65536.0,1,-nbitq), 
to_sfixed(1229.0/65536.0,1,-nbitq), 
to_sfixed(2842.0/65536.0,1,-nbitq), 
to_sfixed(-2230.0/65536.0,1,-nbitq), 
to_sfixed(4932.0/65536.0,1,-nbitq), 
to_sfixed(2208.0/65536.0,1,-nbitq), 
to_sfixed(2920.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1353.0/65536.0,1,-nbitq), 
to_sfixed(4036.0/65536.0,1,-nbitq), 
to_sfixed(3338.0/65536.0,1,-nbitq), 
to_sfixed(-745.0/65536.0,1,-nbitq), 
to_sfixed(-708.0/65536.0,1,-nbitq), 
to_sfixed(-4618.0/65536.0,1,-nbitq), 
to_sfixed(-2503.0/65536.0,1,-nbitq), 
to_sfixed(-2232.0/65536.0,1,-nbitq), 
to_sfixed(508.0/65536.0,1,-nbitq), 
to_sfixed(-1045.0/65536.0,1,-nbitq), 
to_sfixed(-1968.0/65536.0,1,-nbitq), 
to_sfixed(2694.0/65536.0,1,-nbitq), 
to_sfixed(-1999.0/65536.0,1,-nbitq), 
to_sfixed(-265.0/65536.0,1,-nbitq), 
to_sfixed(-1365.0/65536.0,1,-nbitq), 
to_sfixed(1994.0/65536.0,1,-nbitq), 
to_sfixed(-955.0/65536.0,1,-nbitq), 
to_sfixed(-783.0/65536.0,1,-nbitq), 
to_sfixed(1808.0/65536.0,1,-nbitq), 
to_sfixed(1231.0/65536.0,1,-nbitq), 
to_sfixed(-427.0/65536.0,1,-nbitq), 
to_sfixed(-819.0/65536.0,1,-nbitq), 
to_sfixed(873.0/65536.0,1,-nbitq), 
to_sfixed(3547.0/65536.0,1,-nbitq), 
to_sfixed(-1934.0/65536.0,1,-nbitq), 
to_sfixed(-518.0/65536.0,1,-nbitq), 
to_sfixed(-1007.0/65536.0,1,-nbitq), 
to_sfixed(1964.0/65536.0,1,-nbitq), 
to_sfixed(4371.0/65536.0,1,-nbitq), 
to_sfixed(-2296.0/65536.0,1,-nbitq), 
to_sfixed(-1815.0/65536.0,1,-nbitq), 
to_sfixed(-2404.0/65536.0,1,-nbitq), 
to_sfixed(-1965.0/65536.0,1,-nbitq), 
to_sfixed(-1455.0/65536.0,1,-nbitq), 
to_sfixed(1934.0/65536.0,1,-nbitq), 
to_sfixed(228.0/65536.0,1,-nbitq), 
to_sfixed(-193.0/65536.0,1,-nbitq), 
to_sfixed(-1980.0/65536.0,1,-nbitq), 
to_sfixed(-589.0/65536.0,1,-nbitq), 
to_sfixed(-210.0/65536.0,1,-nbitq), 
to_sfixed(-1693.0/65536.0,1,-nbitq), 
to_sfixed(-3306.0/65536.0,1,-nbitq), 
to_sfixed(914.0/65536.0,1,-nbitq), 
to_sfixed(2834.0/65536.0,1,-nbitq), 
to_sfixed(3312.0/65536.0,1,-nbitq), 
to_sfixed(585.0/65536.0,1,-nbitq), 
to_sfixed(2522.0/65536.0,1,-nbitq), 
to_sfixed(682.0/65536.0,1,-nbitq), 
to_sfixed(-1806.0/65536.0,1,-nbitq), 
to_sfixed(-967.0/65536.0,1,-nbitq), 
to_sfixed(2580.0/65536.0,1,-nbitq), 
to_sfixed(3442.0/65536.0,1,-nbitq), 
to_sfixed(3156.0/65536.0,1,-nbitq), 
to_sfixed(-6339.0/65536.0,1,-nbitq), 
to_sfixed(2147.0/65536.0,1,-nbitq), 
to_sfixed(3003.0/65536.0,1,-nbitq), 
to_sfixed(-673.0/65536.0,1,-nbitq), 
to_sfixed(703.0/65536.0,1,-nbitq), 
to_sfixed(-1252.0/65536.0,1,-nbitq), 
to_sfixed(31.0/65536.0,1,-nbitq), 
to_sfixed(1256.0/65536.0,1,-nbitq), 
to_sfixed(1237.0/65536.0,1,-nbitq), 
to_sfixed(759.0/65536.0,1,-nbitq), 
to_sfixed(58.0/65536.0,1,-nbitq), 
to_sfixed(-477.0/65536.0,1,-nbitq), 
to_sfixed(-3284.0/65536.0,1,-nbitq), 
to_sfixed(40.0/65536.0,1,-nbitq), 
to_sfixed(-1352.0/65536.0,1,-nbitq), 
to_sfixed(279.0/65536.0,1,-nbitq), 
to_sfixed(1066.0/65536.0,1,-nbitq), 
to_sfixed(-51.0/65536.0,1,-nbitq), 
to_sfixed(-2435.0/65536.0,1,-nbitq), 
to_sfixed(-891.0/65536.0,1,-nbitq), 
to_sfixed(1380.0/65536.0,1,-nbitq), 
to_sfixed(-2288.0/65536.0,1,-nbitq), 
to_sfixed(3730.0/65536.0,1,-nbitq), 
to_sfixed(451.0/65536.0,1,-nbitq), 
to_sfixed(4880.0/65536.0,1,-nbitq), 
to_sfixed(-2872.0/65536.0,1,-nbitq), 
to_sfixed(2191.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2093.0/65536.0,1,-nbitq), 
to_sfixed(4350.0/65536.0,1,-nbitq), 
to_sfixed(2623.0/65536.0,1,-nbitq), 
to_sfixed(-68.0/65536.0,1,-nbitq), 
to_sfixed(-1024.0/65536.0,1,-nbitq), 
to_sfixed(-3484.0/65536.0,1,-nbitq), 
to_sfixed(-1326.0/65536.0,1,-nbitq), 
to_sfixed(1074.0/65536.0,1,-nbitq), 
to_sfixed(2993.0/65536.0,1,-nbitq), 
to_sfixed(-706.0/65536.0,1,-nbitq), 
to_sfixed(-941.0/65536.0,1,-nbitq), 
to_sfixed(-206.0/65536.0,1,-nbitq), 
to_sfixed(-1810.0/65536.0,1,-nbitq), 
to_sfixed(1283.0/65536.0,1,-nbitq), 
to_sfixed(3550.0/65536.0,1,-nbitq), 
to_sfixed(551.0/65536.0,1,-nbitq), 
to_sfixed(1988.0/65536.0,1,-nbitq), 
to_sfixed(4331.0/65536.0,1,-nbitq), 
to_sfixed(325.0/65536.0,1,-nbitq), 
to_sfixed(-2318.0/65536.0,1,-nbitq), 
to_sfixed(1696.0/65536.0,1,-nbitq), 
to_sfixed(-3331.0/65536.0,1,-nbitq), 
to_sfixed(1728.0/65536.0,1,-nbitq), 
to_sfixed(-1464.0/65536.0,1,-nbitq), 
to_sfixed(2683.0/65536.0,1,-nbitq), 
to_sfixed(-1789.0/65536.0,1,-nbitq), 
to_sfixed(-19.0/65536.0,1,-nbitq), 
to_sfixed(-2187.0/65536.0,1,-nbitq), 
to_sfixed(-737.0/65536.0,1,-nbitq), 
to_sfixed(-381.0/65536.0,1,-nbitq), 
to_sfixed(1523.0/65536.0,1,-nbitq), 
to_sfixed(980.0/65536.0,1,-nbitq), 
to_sfixed(-2693.0/65536.0,1,-nbitq), 
to_sfixed(-3086.0/65536.0,1,-nbitq), 
to_sfixed(-415.0/65536.0,1,-nbitq), 
to_sfixed(-501.0/65536.0,1,-nbitq), 
to_sfixed(-1467.0/65536.0,1,-nbitq), 
to_sfixed(-2656.0/65536.0,1,-nbitq), 
to_sfixed(7.0/65536.0,1,-nbitq), 
to_sfixed(2147.0/65536.0,1,-nbitq), 
to_sfixed(967.0/65536.0,1,-nbitq), 
to_sfixed(257.0/65536.0,1,-nbitq), 
to_sfixed(1804.0/65536.0,1,-nbitq), 
to_sfixed(-1479.0/65536.0,1,-nbitq), 
to_sfixed(-29.0/65536.0,1,-nbitq), 
to_sfixed(975.0/65536.0,1,-nbitq), 
to_sfixed(26.0/65536.0,1,-nbitq), 
to_sfixed(-943.0/65536.0,1,-nbitq), 
to_sfixed(3603.0/65536.0,1,-nbitq), 
to_sfixed(4293.0/65536.0,1,-nbitq), 
to_sfixed(-1849.0/65536.0,1,-nbitq), 
to_sfixed(-1479.0/65536.0,1,-nbitq), 
to_sfixed(133.0/65536.0,1,-nbitq), 
to_sfixed(-4046.0/65536.0,1,-nbitq), 
to_sfixed(-1381.0/65536.0,1,-nbitq), 
to_sfixed(-498.0/65536.0,1,-nbitq), 
to_sfixed(1781.0/65536.0,1,-nbitq), 
to_sfixed(1887.0/65536.0,1,-nbitq), 
to_sfixed(-2591.0/65536.0,1,-nbitq), 
to_sfixed(201.0/65536.0,1,-nbitq), 
to_sfixed(-1354.0/65536.0,1,-nbitq), 
to_sfixed(-1649.0/65536.0,1,-nbitq), 
to_sfixed(809.0/65536.0,1,-nbitq), 
to_sfixed(2061.0/65536.0,1,-nbitq), 
to_sfixed(1472.0/65536.0,1,-nbitq), 
to_sfixed(1588.0/65536.0,1,-nbitq), 
to_sfixed(2527.0/65536.0,1,-nbitq), 
to_sfixed(-3053.0/65536.0,1,-nbitq), 
to_sfixed(2075.0/65536.0,1,-nbitq), 
to_sfixed(610.0/65536.0,1,-nbitq), 
to_sfixed(514.0/65536.0,1,-nbitq), 
to_sfixed(-1633.0/65536.0,1,-nbitq), 
to_sfixed(-831.0/65536.0,1,-nbitq), 
to_sfixed(-518.0/65536.0,1,-nbitq), 
to_sfixed(2087.0/65536.0,1,-nbitq), 
to_sfixed(3992.0/65536.0,1,-nbitq), 
to_sfixed(113.0/65536.0,1,-nbitq), 
to_sfixed(4924.0/65536.0,1,-nbitq), 
to_sfixed(-2862.0/65536.0,1,-nbitq), 
to_sfixed(700.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2275.0/65536.0,1,-nbitq), 
to_sfixed(3779.0/65536.0,1,-nbitq), 
to_sfixed(-3739.0/65536.0,1,-nbitq), 
to_sfixed(-4624.0/65536.0,1,-nbitq), 
to_sfixed(514.0/65536.0,1,-nbitq), 
to_sfixed(2.0/65536.0,1,-nbitq), 
to_sfixed(2383.0/65536.0,1,-nbitq), 
to_sfixed(1550.0/65536.0,1,-nbitq), 
to_sfixed(1898.0/65536.0,1,-nbitq), 
to_sfixed(-1837.0/65536.0,1,-nbitq), 
to_sfixed(-602.0/65536.0,1,-nbitq), 
to_sfixed(5303.0/65536.0,1,-nbitq), 
to_sfixed(-2436.0/65536.0,1,-nbitq), 
to_sfixed(5321.0/65536.0,1,-nbitq), 
to_sfixed(1394.0/65536.0,1,-nbitq), 
to_sfixed(395.0/65536.0,1,-nbitq), 
to_sfixed(1514.0/65536.0,1,-nbitq), 
to_sfixed(5940.0/65536.0,1,-nbitq), 
to_sfixed(2331.0/65536.0,1,-nbitq), 
to_sfixed(495.0/65536.0,1,-nbitq), 
to_sfixed(-2407.0/65536.0,1,-nbitq), 
to_sfixed(-1264.0/65536.0,1,-nbitq), 
to_sfixed(8221.0/65536.0,1,-nbitq), 
to_sfixed(3232.0/65536.0,1,-nbitq), 
to_sfixed(1215.0/65536.0,1,-nbitq), 
to_sfixed(-6200.0/65536.0,1,-nbitq), 
to_sfixed(-3448.0/65536.0,1,-nbitq), 
to_sfixed(-16.0/65536.0,1,-nbitq), 
to_sfixed(-1610.0/65536.0,1,-nbitq), 
to_sfixed(3133.0/65536.0,1,-nbitq), 
to_sfixed(2172.0/65536.0,1,-nbitq), 
to_sfixed(-1309.0/65536.0,1,-nbitq), 
to_sfixed(-3199.0/65536.0,1,-nbitq), 
to_sfixed(-3715.0/65536.0,1,-nbitq), 
to_sfixed(2132.0/65536.0,1,-nbitq), 
to_sfixed(2361.0/65536.0,1,-nbitq), 
to_sfixed(-2114.0/65536.0,1,-nbitq), 
to_sfixed(-2399.0/65536.0,1,-nbitq), 
to_sfixed(-455.0/65536.0,1,-nbitq), 
to_sfixed(-2920.0/65536.0,1,-nbitq), 
to_sfixed(-3043.0/65536.0,1,-nbitq), 
to_sfixed(-134.0/65536.0,1,-nbitq), 
to_sfixed(-3376.0/65536.0,1,-nbitq), 
to_sfixed(-2517.0/65536.0,1,-nbitq), 
to_sfixed(1805.0/65536.0,1,-nbitq), 
to_sfixed(-1205.0/65536.0,1,-nbitq), 
to_sfixed(-3636.0/65536.0,1,-nbitq), 
to_sfixed(-2963.0/65536.0,1,-nbitq), 
to_sfixed(-1779.0/65536.0,1,-nbitq), 
to_sfixed(4539.0/65536.0,1,-nbitq), 
to_sfixed(2383.0/65536.0,1,-nbitq), 
to_sfixed(-1929.0/65536.0,1,-nbitq), 
to_sfixed(1677.0/65536.0,1,-nbitq), 
to_sfixed(-584.0/65536.0,1,-nbitq), 
to_sfixed(1669.0/65536.0,1,-nbitq), 
to_sfixed(-1697.0/65536.0,1,-nbitq), 
to_sfixed(2712.0/65536.0,1,-nbitq), 
to_sfixed(-1122.0/65536.0,1,-nbitq), 
to_sfixed(-911.0/65536.0,1,-nbitq), 
to_sfixed(785.0/65536.0,1,-nbitq), 
to_sfixed(-1592.0/65536.0,1,-nbitq), 
to_sfixed(88.0/65536.0,1,-nbitq), 
to_sfixed(1186.0/65536.0,1,-nbitq), 
to_sfixed(-282.0/65536.0,1,-nbitq), 
to_sfixed(2661.0/65536.0,1,-nbitq), 
to_sfixed(32.0/65536.0,1,-nbitq), 
to_sfixed(3451.0/65536.0,1,-nbitq), 
to_sfixed(-3868.0/65536.0,1,-nbitq), 
to_sfixed(-950.0/65536.0,1,-nbitq), 
to_sfixed(4545.0/65536.0,1,-nbitq), 
to_sfixed(-1354.0/65536.0,1,-nbitq), 
to_sfixed(75.0/65536.0,1,-nbitq), 
to_sfixed(-2172.0/65536.0,1,-nbitq), 
to_sfixed(-2355.0/65536.0,1,-nbitq), 
to_sfixed(-660.0/65536.0,1,-nbitq), 
to_sfixed(-528.0/65536.0,1,-nbitq), 
to_sfixed(4831.0/65536.0,1,-nbitq), 
to_sfixed(-428.0/65536.0,1,-nbitq), 
to_sfixed(-2387.0/65536.0,1,-nbitq), 
to_sfixed(2870.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2596.0/65536.0,1,-nbitq), 
to_sfixed(-1007.0/65536.0,1,-nbitq), 
to_sfixed(-8153.0/65536.0,1,-nbitq), 
to_sfixed(-318.0/65536.0,1,-nbitq), 
to_sfixed(-289.0/65536.0,1,-nbitq), 
to_sfixed(-1969.0/65536.0,1,-nbitq), 
to_sfixed(2836.0/65536.0,1,-nbitq), 
to_sfixed(-153.0/65536.0,1,-nbitq), 
to_sfixed(3673.0/65536.0,1,-nbitq), 
to_sfixed(2475.0/65536.0,1,-nbitq), 
to_sfixed(2513.0/65536.0,1,-nbitq), 
to_sfixed(4480.0/65536.0,1,-nbitq), 
to_sfixed(-2010.0/65536.0,1,-nbitq), 
to_sfixed(-1187.0/65536.0,1,-nbitq), 
to_sfixed(-1843.0/65536.0,1,-nbitq), 
to_sfixed(1624.0/65536.0,1,-nbitq), 
to_sfixed(-2683.0/65536.0,1,-nbitq), 
to_sfixed(2605.0/65536.0,1,-nbitq), 
to_sfixed(1013.0/65536.0,1,-nbitq), 
to_sfixed(447.0/65536.0,1,-nbitq), 
to_sfixed(-3177.0/65536.0,1,-nbitq), 
to_sfixed(-772.0/65536.0,1,-nbitq), 
to_sfixed(9308.0/65536.0,1,-nbitq), 
to_sfixed(-2577.0/65536.0,1,-nbitq), 
to_sfixed(840.0/65536.0,1,-nbitq), 
to_sfixed(-7992.0/65536.0,1,-nbitq), 
to_sfixed(-197.0/65536.0,1,-nbitq), 
to_sfixed(-1642.0/65536.0,1,-nbitq), 
to_sfixed(-5420.0/65536.0,1,-nbitq), 
to_sfixed(2176.0/65536.0,1,-nbitq), 
to_sfixed(-424.0/65536.0,1,-nbitq), 
to_sfixed(-3867.0/65536.0,1,-nbitq), 
to_sfixed(-62.0/65536.0,1,-nbitq), 
to_sfixed(-989.0/65536.0,1,-nbitq), 
to_sfixed(-1697.0/65536.0,1,-nbitq), 
to_sfixed(-1808.0/65536.0,1,-nbitq), 
to_sfixed(-1535.0/65536.0,1,-nbitq), 
to_sfixed(1679.0/65536.0,1,-nbitq), 
to_sfixed(9784.0/65536.0,1,-nbitq), 
to_sfixed(169.0/65536.0,1,-nbitq), 
to_sfixed(-1919.0/65536.0,1,-nbitq), 
to_sfixed(138.0/65536.0,1,-nbitq), 
to_sfixed(-2333.0/65536.0,1,-nbitq), 
to_sfixed(1842.0/65536.0,1,-nbitq), 
to_sfixed(2786.0/65536.0,1,-nbitq), 
to_sfixed(-21.0/65536.0,1,-nbitq), 
to_sfixed(158.0/65536.0,1,-nbitq), 
to_sfixed(-4684.0/65536.0,1,-nbitq), 
to_sfixed(3180.0/65536.0,1,-nbitq), 
to_sfixed(-553.0/65536.0,1,-nbitq), 
to_sfixed(770.0/65536.0,1,-nbitq), 
to_sfixed(-3666.0/65536.0,1,-nbitq), 
to_sfixed(1059.0/65536.0,1,-nbitq), 
to_sfixed(-805.0/65536.0,1,-nbitq), 
to_sfixed(2253.0/65536.0,1,-nbitq), 
to_sfixed(-2659.0/65536.0,1,-nbitq), 
to_sfixed(3947.0/65536.0,1,-nbitq), 
to_sfixed(-2138.0/65536.0,1,-nbitq), 
to_sfixed(1084.0/65536.0,1,-nbitq), 
to_sfixed(-2835.0/65536.0,1,-nbitq), 
to_sfixed(-3451.0/65536.0,1,-nbitq), 
to_sfixed(-1408.0/65536.0,1,-nbitq), 
to_sfixed(2708.0/65536.0,1,-nbitq), 
to_sfixed(-2738.0/65536.0,1,-nbitq), 
to_sfixed(1770.0/65536.0,1,-nbitq), 
to_sfixed(-3182.0/65536.0,1,-nbitq), 
to_sfixed(5285.0/65536.0,1,-nbitq), 
to_sfixed(5267.0/65536.0,1,-nbitq), 
to_sfixed(1875.0/65536.0,1,-nbitq), 
to_sfixed(4042.0/65536.0,1,-nbitq), 
to_sfixed(2033.0/65536.0,1,-nbitq), 
to_sfixed(4158.0/65536.0,1,-nbitq), 
to_sfixed(-715.0/65536.0,1,-nbitq), 
to_sfixed(-131.0/65536.0,1,-nbitq), 
to_sfixed(-2219.0/65536.0,1,-nbitq), 
to_sfixed(1808.0/65536.0,1,-nbitq), 
to_sfixed(2743.0/65536.0,1,-nbitq), 
to_sfixed(2977.0/65536.0,1,-nbitq), 
to_sfixed(2956.0/65536.0,1,-nbitq), 
to_sfixed(2424.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-168.0/65536.0,1,-nbitq), 
to_sfixed(-88.0/65536.0,1,-nbitq), 
to_sfixed(-8556.0/65536.0,1,-nbitq), 
to_sfixed(-5937.0/65536.0,1,-nbitq), 
to_sfixed(-5003.0/65536.0,1,-nbitq), 
to_sfixed(-1134.0/65536.0,1,-nbitq), 
to_sfixed(449.0/65536.0,1,-nbitq), 
to_sfixed(3632.0/65536.0,1,-nbitq), 
to_sfixed(-871.0/65536.0,1,-nbitq), 
to_sfixed(446.0/65536.0,1,-nbitq), 
to_sfixed(2326.0/65536.0,1,-nbitq), 
to_sfixed(6901.0/65536.0,1,-nbitq), 
to_sfixed(2039.0/65536.0,1,-nbitq), 
to_sfixed(-3092.0/65536.0,1,-nbitq), 
to_sfixed(-4301.0/65536.0,1,-nbitq), 
to_sfixed(-1757.0/65536.0,1,-nbitq), 
to_sfixed(-536.0/65536.0,1,-nbitq), 
to_sfixed(1707.0/65536.0,1,-nbitq), 
to_sfixed(-4866.0/65536.0,1,-nbitq), 
to_sfixed(182.0/65536.0,1,-nbitq), 
to_sfixed(75.0/65536.0,1,-nbitq), 
to_sfixed(-625.0/65536.0,1,-nbitq), 
to_sfixed(9550.0/65536.0,1,-nbitq), 
to_sfixed(-269.0/65536.0,1,-nbitq), 
to_sfixed(-799.0/65536.0,1,-nbitq), 
to_sfixed(-7024.0/65536.0,1,-nbitq), 
to_sfixed(165.0/65536.0,1,-nbitq), 
to_sfixed(-1199.0/65536.0,1,-nbitq), 
to_sfixed(-4313.0/65536.0,1,-nbitq), 
to_sfixed(1436.0/65536.0,1,-nbitq), 
to_sfixed(-2055.0/65536.0,1,-nbitq), 
to_sfixed(-7324.0/65536.0,1,-nbitq), 
to_sfixed(-757.0/65536.0,1,-nbitq), 
to_sfixed(-1418.0/65536.0,1,-nbitq), 
to_sfixed(-2864.0/65536.0,1,-nbitq), 
to_sfixed(-940.0/65536.0,1,-nbitq), 
to_sfixed(260.0/65536.0,1,-nbitq), 
to_sfixed(4108.0/65536.0,1,-nbitq), 
to_sfixed(12527.0/65536.0,1,-nbitq), 
to_sfixed(-2917.0/65536.0,1,-nbitq), 
to_sfixed(-1336.0/65536.0,1,-nbitq), 
to_sfixed(-3257.0/65536.0,1,-nbitq), 
to_sfixed(1276.0/65536.0,1,-nbitq), 
to_sfixed(-790.0/65536.0,1,-nbitq), 
to_sfixed(-1812.0/65536.0,1,-nbitq), 
to_sfixed(1117.0/65536.0,1,-nbitq), 
to_sfixed(-3431.0/65536.0,1,-nbitq), 
to_sfixed(-6758.0/65536.0,1,-nbitq), 
to_sfixed(786.0/65536.0,1,-nbitq), 
to_sfixed(2676.0/65536.0,1,-nbitq), 
to_sfixed(2555.0/65536.0,1,-nbitq), 
to_sfixed(-5535.0/65536.0,1,-nbitq), 
to_sfixed(-490.0/65536.0,1,-nbitq), 
to_sfixed(-5920.0/65536.0,1,-nbitq), 
to_sfixed(4583.0/65536.0,1,-nbitq), 
to_sfixed(-6002.0/65536.0,1,-nbitq), 
to_sfixed(1928.0/65536.0,1,-nbitq), 
to_sfixed(-1563.0/65536.0,1,-nbitq), 
to_sfixed(2892.0/65536.0,1,-nbitq), 
to_sfixed(-3387.0/65536.0,1,-nbitq), 
to_sfixed(-2427.0/65536.0,1,-nbitq), 
to_sfixed(124.0/65536.0,1,-nbitq), 
to_sfixed(-2324.0/65536.0,1,-nbitq), 
to_sfixed(262.0/65536.0,1,-nbitq), 
to_sfixed(-150.0/65536.0,1,-nbitq), 
to_sfixed(-7129.0/65536.0,1,-nbitq), 
to_sfixed(5479.0/65536.0,1,-nbitq), 
to_sfixed(6356.0/65536.0,1,-nbitq), 
to_sfixed(-2570.0/65536.0,1,-nbitq), 
to_sfixed(2842.0/65536.0,1,-nbitq), 
to_sfixed(1541.0/65536.0,1,-nbitq), 
to_sfixed(2627.0/65536.0,1,-nbitq), 
to_sfixed(-1629.0/65536.0,1,-nbitq), 
to_sfixed(1598.0/65536.0,1,-nbitq), 
to_sfixed(1657.0/65536.0,1,-nbitq), 
to_sfixed(1290.0/65536.0,1,-nbitq), 
to_sfixed(5839.0/65536.0,1,-nbitq), 
to_sfixed(-1423.0/65536.0,1,-nbitq), 
to_sfixed(-435.0/65536.0,1,-nbitq), 
to_sfixed(1287.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1026.0/65536.0,1,-nbitq), 
to_sfixed(3260.0/65536.0,1,-nbitq), 
to_sfixed(-10880.0/65536.0,1,-nbitq), 
to_sfixed(-1717.0/65536.0,1,-nbitq), 
to_sfixed(-519.0/65536.0,1,-nbitq), 
to_sfixed(-1067.0/65536.0,1,-nbitq), 
to_sfixed(2966.0/65536.0,1,-nbitq), 
to_sfixed(547.0/65536.0,1,-nbitq), 
to_sfixed(2019.0/65536.0,1,-nbitq), 
to_sfixed(2799.0/65536.0,1,-nbitq), 
to_sfixed(-315.0/65536.0,1,-nbitq), 
to_sfixed(9729.0/65536.0,1,-nbitq), 
to_sfixed(-618.0/65536.0,1,-nbitq), 
to_sfixed(-5586.0/65536.0,1,-nbitq), 
to_sfixed(-108.0/65536.0,1,-nbitq), 
to_sfixed(-1814.0/65536.0,1,-nbitq), 
to_sfixed(46.0/65536.0,1,-nbitq), 
to_sfixed(-981.0/65536.0,1,-nbitq), 
to_sfixed(-3014.0/65536.0,1,-nbitq), 
to_sfixed(12.0/65536.0,1,-nbitq), 
to_sfixed(3926.0/65536.0,1,-nbitq), 
to_sfixed(-627.0/65536.0,1,-nbitq), 
to_sfixed(8663.0/65536.0,1,-nbitq), 
to_sfixed(-1086.0/65536.0,1,-nbitq), 
to_sfixed(4103.0/65536.0,1,-nbitq), 
to_sfixed(-4110.0/65536.0,1,-nbitq), 
to_sfixed(-1597.0/65536.0,1,-nbitq), 
to_sfixed(-753.0/65536.0,1,-nbitq), 
to_sfixed(-5375.0/65536.0,1,-nbitq), 
to_sfixed(2523.0/65536.0,1,-nbitq), 
to_sfixed(-2359.0/65536.0,1,-nbitq), 
to_sfixed(-4505.0/65536.0,1,-nbitq), 
to_sfixed(2163.0/65536.0,1,-nbitq), 
to_sfixed(-2887.0/65536.0,1,-nbitq), 
to_sfixed(-2561.0/65536.0,1,-nbitq), 
to_sfixed(1490.0/65536.0,1,-nbitq), 
to_sfixed(4486.0/65536.0,1,-nbitq), 
to_sfixed(9330.0/65536.0,1,-nbitq), 
to_sfixed(9693.0/65536.0,1,-nbitq), 
to_sfixed(2864.0/65536.0,1,-nbitq), 
to_sfixed(1679.0/65536.0,1,-nbitq), 
to_sfixed(409.0/65536.0,1,-nbitq), 
to_sfixed(1903.0/65536.0,1,-nbitq), 
to_sfixed(471.0/65536.0,1,-nbitq), 
to_sfixed(-2313.0/65536.0,1,-nbitq), 
to_sfixed(1089.0/65536.0,1,-nbitq), 
to_sfixed(-1259.0/65536.0,1,-nbitq), 
to_sfixed(-6114.0/65536.0,1,-nbitq), 
to_sfixed(3195.0/65536.0,1,-nbitq), 
to_sfixed(3186.0/65536.0,1,-nbitq), 
to_sfixed(2859.0/65536.0,1,-nbitq), 
to_sfixed(-2356.0/65536.0,1,-nbitq), 
to_sfixed(-3443.0/65536.0,1,-nbitq), 
to_sfixed(-6463.0/65536.0,1,-nbitq), 
to_sfixed(3528.0/65536.0,1,-nbitq), 
to_sfixed(-6011.0/65536.0,1,-nbitq), 
to_sfixed(1490.0/65536.0,1,-nbitq), 
to_sfixed(1658.0/65536.0,1,-nbitq), 
to_sfixed(1495.0/65536.0,1,-nbitq), 
to_sfixed(-5190.0/65536.0,1,-nbitq), 
to_sfixed(-5526.0/65536.0,1,-nbitq), 
to_sfixed(-2739.0/65536.0,1,-nbitq), 
to_sfixed(1624.0/65536.0,1,-nbitq), 
to_sfixed(1704.0/65536.0,1,-nbitq), 
to_sfixed(-64.0/65536.0,1,-nbitq), 
to_sfixed(-7138.0/65536.0,1,-nbitq), 
to_sfixed(5834.0/65536.0,1,-nbitq), 
to_sfixed(11972.0/65536.0,1,-nbitq), 
to_sfixed(-3026.0/65536.0,1,-nbitq), 
to_sfixed(8603.0/65536.0,1,-nbitq), 
to_sfixed(1916.0/65536.0,1,-nbitq), 
to_sfixed(-1254.0/65536.0,1,-nbitq), 
to_sfixed(-3727.0/65536.0,1,-nbitq), 
to_sfixed(2408.0/65536.0,1,-nbitq), 
to_sfixed(2070.0/65536.0,1,-nbitq), 
to_sfixed(-1032.0/65536.0,1,-nbitq), 
to_sfixed(5856.0/65536.0,1,-nbitq), 
to_sfixed(1382.0/65536.0,1,-nbitq), 
to_sfixed(-627.0/65536.0,1,-nbitq), 
to_sfixed(-751.0/65536.0,1,-nbitq)  ), 
( to_sfixed(159.0/65536.0,1,-nbitq), 
to_sfixed(3041.0/65536.0,1,-nbitq), 
to_sfixed(-9331.0/65536.0,1,-nbitq), 
to_sfixed(-2795.0/65536.0,1,-nbitq), 
to_sfixed(-1448.0/65536.0,1,-nbitq), 
to_sfixed(816.0/65536.0,1,-nbitq), 
to_sfixed(2029.0/65536.0,1,-nbitq), 
to_sfixed(942.0/65536.0,1,-nbitq), 
to_sfixed(3495.0/65536.0,1,-nbitq), 
to_sfixed(693.0/65536.0,1,-nbitq), 
to_sfixed(3090.0/65536.0,1,-nbitq), 
to_sfixed(8389.0/65536.0,1,-nbitq), 
to_sfixed(-1628.0/65536.0,1,-nbitq), 
to_sfixed(-7458.0/65536.0,1,-nbitq), 
to_sfixed(-2818.0/65536.0,1,-nbitq), 
to_sfixed(206.0/65536.0,1,-nbitq), 
to_sfixed(-1813.0/65536.0,1,-nbitq), 
to_sfixed(-6173.0/65536.0,1,-nbitq), 
to_sfixed(1470.0/65536.0,1,-nbitq), 
to_sfixed(469.0/65536.0,1,-nbitq), 
to_sfixed(1460.0/65536.0,1,-nbitq), 
to_sfixed(-2368.0/65536.0,1,-nbitq), 
to_sfixed(5519.0/65536.0,1,-nbitq), 
to_sfixed(981.0/65536.0,1,-nbitq), 
to_sfixed(-1192.0/65536.0,1,-nbitq), 
to_sfixed(-8329.0/65536.0,1,-nbitq), 
to_sfixed(-72.0/65536.0,1,-nbitq), 
to_sfixed(-3.0/65536.0,1,-nbitq), 
to_sfixed(2797.0/65536.0,1,-nbitq), 
to_sfixed(-1386.0/65536.0,1,-nbitq), 
to_sfixed(2993.0/65536.0,1,-nbitq), 
to_sfixed(-6756.0/65536.0,1,-nbitq), 
to_sfixed(1457.0/65536.0,1,-nbitq), 
to_sfixed(-1428.0/65536.0,1,-nbitq), 
to_sfixed(-3550.0/65536.0,1,-nbitq), 
to_sfixed(-2714.0/65536.0,1,-nbitq), 
to_sfixed(1306.0/65536.0,1,-nbitq), 
to_sfixed(9069.0/65536.0,1,-nbitq), 
to_sfixed(2596.0/65536.0,1,-nbitq), 
to_sfixed(697.0/65536.0,1,-nbitq), 
to_sfixed(-992.0/65536.0,1,-nbitq), 
to_sfixed(-2191.0/65536.0,1,-nbitq), 
to_sfixed(444.0/65536.0,1,-nbitq), 
to_sfixed(199.0/65536.0,1,-nbitq), 
to_sfixed(-1953.0/65536.0,1,-nbitq), 
to_sfixed(1352.0/65536.0,1,-nbitq), 
to_sfixed(782.0/65536.0,1,-nbitq), 
to_sfixed(-8498.0/65536.0,1,-nbitq), 
to_sfixed(3039.0/65536.0,1,-nbitq), 
to_sfixed(853.0/65536.0,1,-nbitq), 
to_sfixed(-374.0/65536.0,1,-nbitq), 
to_sfixed(1161.0/65536.0,1,-nbitq), 
to_sfixed(-4380.0/65536.0,1,-nbitq), 
to_sfixed(-5757.0/65536.0,1,-nbitq), 
to_sfixed(1253.0/65536.0,1,-nbitq), 
to_sfixed(-6098.0/65536.0,1,-nbitq), 
to_sfixed(2501.0/65536.0,1,-nbitq), 
to_sfixed(1338.0/65536.0,1,-nbitq), 
to_sfixed(-1288.0/65536.0,1,-nbitq), 
to_sfixed(-7313.0/65536.0,1,-nbitq), 
to_sfixed(-5672.0/65536.0,1,-nbitq), 
to_sfixed(-1509.0/65536.0,1,-nbitq), 
to_sfixed(-715.0/65536.0,1,-nbitq), 
to_sfixed(-3068.0/65536.0,1,-nbitq), 
to_sfixed(553.0/65536.0,1,-nbitq), 
to_sfixed(-7389.0/65536.0,1,-nbitq), 
to_sfixed(4308.0/65536.0,1,-nbitq), 
to_sfixed(11420.0/65536.0,1,-nbitq), 
to_sfixed(3866.0/65536.0,1,-nbitq), 
to_sfixed(9867.0/65536.0,1,-nbitq), 
to_sfixed(1897.0/65536.0,1,-nbitq), 
to_sfixed(-1943.0/65536.0,1,-nbitq), 
to_sfixed(-4522.0/65536.0,1,-nbitq), 
to_sfixed(-2185.0/65536.0,1,-nbitq), 
to_sfixed(-1989.0/65536.0,1,-nbitq), 
to_sfixed(-2672.0/65536.0,1,-nbitq), 
to_sfixed(7224.0/65536.0,1,-nbitq), 
to_sfixed(3776.0/65536.0,1,-nbitq), 
to_sfixed(2317.0/65536.0,1,-nbitq), 
to_sfixed(-2839.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2984.0/65536.0,1,-nbitq), 
to_sfixed(6141.0/65536.0,1,-nbitq), 
to_sfixed(-7120.0/65536.0,1,-nbitq), 
to_sfixed(-2050.0/65536.0,1,-nbitq), 
to_sfixed(-3464.0/65536.0,1,-nbitq), 
to_sfixed(1581.0/65536.0,1,-nbitq), 
to_sfixed(3441.0/65536.0,1,-nbitq), 
to_sfixed(1047.0/65536.0,1,-nbitq), 
to_sfixed(1182.0/65536.0,1,-nbitq), 
to_sfixed(-2671.0/65536.0,1,-nbitq), 
to_sfixed(3490.0/65536.0,1,-nbitq), 
to_sfixed(1155.0/65536.0,1,-nbitq), 
to_sfixed(-1262.0/65536.0,1,-nbitq), 
to_sfixed(-7319.0/65536.0,1,-nbitq), 
to_sfixed(-1986.0/65536.0,1,-nbitq), 
to_sfixed(-1929.0/65536.0,1,-nbitq), 
to_sfixed(-1008.0/65536.0,1,-nbitq), 
to_sfixed(-3726.0/65536.0,1,-nbitq), 
to_sfixed(1326.0/65536.0,1,-nbitq), 
to_sfixed(1389.0/65536.0,1,-nbitq), 
to_sfixed(-1568.0/65536.0,1,-nbitq), 
to_sfixed(1159.0/65536.0,1,-nbitq), 
to_sfixed(-1718.0/65536.0,1,-nbitq), 
to_sfixed(1236.0/65536.0,1,-nbitq), 
to_sfixed(896.0/65536.0,1,-nbitq), 
to_sfixed(-5563.0/65536.0,1,-nbitq), 
to_sfixed(-2288.0/65536.0,1,-nbitq), 
to_sfixed(2081.0/65536.0,1,-nbitq), 
to_sfixed(137.0/65536.0,1,-nbitq), 
to_sfixed(-630.0/65536.0,1,-nbitq), 
to_sfixed(999.0/65536.0,1,-nbitq), 
to_sfixed(-5981.0/65536.0,1,-nbitq), 
to_sfixed(2811.0/65536.0,1,-nbitq), 
to_sfixed(-773.0/65536.0,1,-nbitq), 
to_sfixed(-246.0/65536.0,1,-nbitq), 
to_sfixed(2453.0/65536.0,1,-nbitq), 
to_sfixed(3163.0/65536.0,1,-nbitq), 
to_sfixed(4857.0/65536.0,1,-nbitq), 
to_sfixed(5620.0/65536.0,1,-nbitq), 
to_sfixed(3435.0/65536.0,1,-nbitq), 
to_sfixed(490.0/65536.0,1,-nbitq), 
to_sfixed(-1979.0/65536.0,1,-nbitq), 
to_sfixed(-1060.0/65536.0,1,-nbitq), 
to_sfixed(1642.0/65536.0,1,-nbitq), 
to_sfixed(2051.0/65536.0,1,-nbitq), 
to_sfixed(-1258.0/65536.0,1,-nbitq), 
to_sfixed(-2179.0/65536.0,1,-nbitq), 
to_sfixed(-3618.0/65536.0,1,-nbitq), 
to_sfixed(244.0/65536.0,1,-nbitq), 
to_sfixed(1739.0/65536.0,1,-nbitq), 
to_sfixed(1073.0/65536.0,1,-nbitq), 
to_sfixed(3471.0/65536.0,1,-nbitq), 
to_sfixed(-7042.0/65536.0,1,-nbitq), 
to_sfixed(-1858.0/65536.0,1,-nbitq), 
to_sfixed(1509.0/65536.0,1,-nbitq), 
to_sfixed(-4520.0/65536.0,1,-nbitq), 
to_sfixed(627.0/65536.0,1,-nbitq), 
to_sfixed(308.0/65536.0,1,-nbitq), 
to_sfixed(366.0/65536.0,1,-nbitq), 
to_sfixed(-7322.0/65536.0,1,-nbitq), 
to_sfixed(-3578.0/65536.0,1,-nbitq), 
to_sfixed(-74.0/65536.0,1,-nbitq), 
to_sfixed(-2386.0/65536.0,1,-nbitq), 
to_sfixed(2546.0/65536.0,1,-nbitq), 
to_sfixed(-771.0/65536.0,1,-nbitq), 
to_sfixed(-4179.0/65536.0,1,-nbitq), 
to_sfixed(7112.0/65536.0,1,-nbitq), 
to_sfixed(10583.0/65536.0,1,-nbitq), 
to_sfixed(8667.0/65536.0,1,-nbitq), 
to_sfixed(8765.0/65536.0,1,-nbitq), 
to_sfixed(-2420.0/65536.0,1,-nbitq), 
to_sfixed(259.0/65536.0,1,-nbitq), 
to_sfixed(-1063.0/65536.0,1,-nbitq), 
to_sfixed(-1544.0/65536.0,1,-nbitq), 
to_sfixed(351.0/65536.0,1,-nbitq), 
to_sfixed(-302.0/65536.0,1,-nbitq), 
to_sfixed(1441.0/65536.0,1,-nbitq), 
to_sfixed(6383.0/65536.0,1,-nbitq), 
to_sfixed(-416.0/65536.0,1,-nbitq), 
to_sfixed(1205.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3162.0/65536.0,1,-nbitq), 
to_sfixed(3225.0/65536.0,1,-nbitq), 
to_sfixed(-4661.0/65536.0,1,-nbitq), 
to_sfixed(-4020.0/65536.0,1,-nbitq), 
to_sfixed(-5290.0/65536.0,1,-nbitq), 
to_sfixed(3460.0/65536.0,1,-nbitq), 
to_sfixed(-163.0/65536.0,1,-nbitq), 
to_sfixed(-1397.0/65536.0,1,-nbitq), 
to_sfixed(2824.0/65536.0,1,-nbitq), 
to_sfixed(1595.0/65536.0,1,-nbitq), 
to_sfixed(1493.0/65536.0,1,-nbitq), 
to_sfixed(-2805.0/65536.0,1,-nbitq), 
to_sfixed(-1316.0/65536.0,1,-nbitq), 
to_sfixed(-5113.0/65536.0,1,-nbitq), 
to_sfixed(-2623.0/65536.0,1,-nbitq), 
to_sfixed(-69.0/65536.0,1,-nbitq), 
to_sfixed(1382.0/65536.0,1,-nbitq), 
to_sfixed(1024.0/65536.0,1,-nbitq), 
to_sfixed(3130.0/65536.0,1,-nbitq), 
to_sfixed(-488.0/65536.0,1,-nbitq), 
to_sfixed(-3353.0/65536.0,1,-nbitq), 
to_sfixed(-5403.0/65536.0,1,-nbitq), 
to_sfixed(-5664.0/65536.0,1,-nbitq), 
to_sfixed(3705.0/65536.0,1,-nbitq), 
to_sfixed(1645.0/65536.0,1,-nbitq), 
to_sfixed(-2125.0/65536.0,1,-nbitq), 
to_sfixed(1858.0/65536.0,1,-nbitq), 
to_sfixed(-1864.0/65536.0,1,-nbitq), 
to_sfixed(2147.0/65536.0,1,-nbitq), 
to_sfixed(-2606.0/65536.0,1,-nbitq), 
to_sfixed(-74.0/65536.0,1,-nbitq), 
to_sfixed(-4972.0/65536.0,1,-nbitq), 
to_sfixed(3898.0/65536.0,1,-nbitq), 
to_sfixed(474.0/65536.0,1,-nbitq), 
to_sfixed(-2365.0/65536.0,1,-nbitq), 
to_sfixed(1927.0/65536.0,1,-nbitq), 
to_sfixed(5491.0/65536.0,1,-nbitq), 
to_sfixed(2911.0/65536.0,1,-nbitq), 
to_sfixed(3088.0/65536.0,1,-nbitq), 
to_sfixed(-764.0/65536.0,1,-nbitq), 
to_sfixed(-212.0/65536.0,1,-nbitq), 
to_sfixed(-2135.0/65536.0,1,-nbitq), 
to_sfixed(467.0/65536.0,1,-nbitq), 
to_sfixed(-542.0/65536.0,1,-nbitq), 
to_sfixed(3318.0/65536.0,1,-nbitq), 
to_sfixed(-1625.0/65536.0,1,-nbitq), 
to_sfixed(-2027.0/65536.0,1,-nbitq), 
to_sfixed(-3935.0/65536.0,1,-nbitq), 
to_sfixed(-1632.0/65536.0,1,-nbitq), 
to_sfixed(353.0/65536.0,1,-nbitq), 
to_sfixed(1534.0/65536.0,1,-nbitq), 
to_sfixed(160.0/65536.0,1,-nbitq), 
to_sfixed(-7142.0/65536.0,1,-nbitq), 
to_sfixed(3359.0/65536.0,1,-nbitq), 
to_sfixed(242.0/65536.0,1,-nbitq), 
to_sfixed(-1645.0/65536.0,1,-nbitq), 
to_sfixed(928.0/65536.0,1,-nbitq), 
to_sfixed(1480.0/65536.0,1,-nbitq), 
to_sfixed(877.0/65536.0,1,-nbitq), 
to_sfixed(-6618.0/65536.0,1,-nbitq), 
to_sfixed(-5038.0/65536.0,1,-nbitq), 
to_sfixed(-1292.0/65536.0,1,-nbitq), 
to_sfixed(-1994.0/65536.0,1,-nbitq), 
to_sfixed(-564.0/65536.0,1,-nbitq), 
to_sfixed(2175.0/65536.0,1,-nbitq), 
to_sfixed(-4808.0/65536.0,1,-nbitq), 
to_sfixed(3754.0/65536.0,1,-nbitq), 
to_sfixed(6299.0/65536.0,1,-nbitq), 
to_sfixed(8631.0/65536.0,1,-nbitq), 
to_sfixed(1791.0/65536.0,1,-nbitq), 
to_sfixed(-3246.0/65536.0,1,-nbitq), 
to_sfixed(377.0/65536.0,1,-nbitq), 
to_sfixed(-2311.0/65536.0,1,-nbitq), 
to_sfixed(-382.0/65536.0,1,-nbitq), 
to_sfixed(-1943.0/65536.0,1,-nbitq), 
to_sfixed(976.0/65536.0,1,-nbitq), 
to_sfixed(1726.0/65536.0,1,-nbitq), 
to_sfixed(8529.0/65536.0,1,-nbitq), 
to_sfixed(-1944.0/65536.0,1,-nbitq), 
to_sfixed(-900.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1059.0/65536.0,1,-nbitq), 
to_sfixed(4108.0/65536.0,1,-nbitq), 
to_sfixed(-1338.0/65536.0,1,-nbitq), 
to_sfixed(-782.0/65536.0,1,-nbitq), 
to_sfixed(349.0/65536.0,1,-nbitq), 
to_sfixed(1532.0/65536.0,1,-nbitq), 
to_sfixed(2726.0/65536.0,1,-nbitq), 
to_sfixed(-1582.0/65536.0,1,-nbitq), 
to_sfixed(4227.0/65536.0,1,-nbitq), 
to_sfixed(-1342.0/65536.0,1,-nbitq), 
to_sfixed(3040.0/65536.0,1,-nbitq), 
to_sfixed(-7582.0/65536.0,1,-nbitq), 
to_sfixed(2239.0/65536.0,1,-nbitq), 
to_sfixed(-1451.0/65536.0,1,-nbitq), 
to_sfixed(-1933.0/65536.0,1,-nbitq), 
to_sfixed(1062.0/65536.0,1,-nbitq), 
to_sfixed(517.0/65536.0,1,-nbitq), 
to_sfixed(-261.0/65536.0,1,-nbitq), 
to_sfixed(1257.0/65536.0,1,-nbitq), 
to_sfixed(3471.0/65536.0,1,-nbitq), 
to_sfixed(-4194.0/65536.0,1,-nbitq), 
to_sfixed(-3776.0/65536.0,1,-nbitq), 
to_sfixed(-3694.0/65536.0,1,-nbitq), 
to_sfixed(1932.0/65536.0,1,-nbitq), 
to_sfixed(2087.0/65536.0,1,-nbitq), 
to_sfixed(1050.0/65536.0,1,-nbitq), 
to_sfixed(3058.0/65536.0,1,-nbitq), 
to_sfixed(-2067.0/65536.0,1,-nbitq), 
to_sfixed(39.0/65536.0,1,-nbitq), 
to_sfixed(1566.0/65536.0,1,-nbitq), 
to_sfixed(3137.0/65536.0,1,-nbitq), 
to_sfixed(-3664.0/65536.0,1,-nbitq), 
to_sfixed(2661.0/65536.0,1,-nbitq), 
to_sfixed(-3414.0/65536.0,1,-nbitq), 
to_sfixed(-300.0/65536.0,1,-nbitq), 
to_sfixed(665.0/65536.0,1,-nbitq), 
to_sfixed(3542.0/65536.0,1,-nbitq), 
to_sfixed(4125.0/65536.0,1,-nbitq), 
to_sfixed(-742.0/65536.0,1,-nbitq), 
to_sfixed(648.0/65536.0,1,-nbitq), 
to_sfixed(1537.0/65536.0,1,-nbitq), 
to_sfixed(-1710.0/65536.0,1,-nbitq), 
to_sfixed(-3046.0/65536.0,1,-nbitq), 
to_sfixed(849.0/65536.0,1,-nbitq), 
to_sfixed(1983.0/65536.0,1,-nbitq), 
to_sfixed(5020.0/65536.0,1,-nbitq), 
to_sfixed(1400.0/65536.0,1,-nbitq), 
to_sfixed(3963.0/65536.0,1,-nbitq), 
to_sfixed(2698.0/65536.0,1,-nbitq), 
to_sfixed(4139.0/65536.0,1,-nbitq), 
to_sfixed(118.0/65536.0,1,-nbitq), 
to_sfixed(2474.0/65536.0,1,-nbitq), 
to_sfixed(-1229.0/65536.0,1,-nbitq), 
to_sfixed(-701.0/65536.0,1,-nbitq), 
to_sfixed(541.0/65536.0,1,-nbitq), 
to_sfixed(-6101.0/65536.0,1,-nbitq), 
to_sfixed(3086.0/65536.0,1,-nbitq), 
to_sfixed(-2020.0/65536.0,1,-nbitq), 
to_sfixed(2019.0/65536.0,1,-nbitq), 
to_sfixed(-8225.0/65536.0,1,-nbitq), 
to_sfixed(-3284.0/65536.0,1,-nbitq), 
to_sfixed(-2573.0/65536.0,1,-nbitq), 
to_sfixed(1918.0/65536.0,1,-nbitq), 
to_sfixed(-2554.0/65536.0,1,-nbitq), 
to_sfixed(2428.0/65536.0,1,-nbitq), 
to_sfixed(-2449.0/65536.0,1,-nbitq), 
to_sfixed(1894.0/65536.0,1,-nbitq), 
to_sfixed(3560.0/65536.0,1,-nbitq), 
to_sfixed(5166.0/65536.0,1,-nbitq), 
to_sfixed(1558.0/65536.0,1,-nbitq), 
to_sfixed(-2390.0/65536.0,1,-nbitq), 
to_sfixed(-139.0/65536.0,1,-nbitq), 
to_sfixed(-1485.0/65536.0,1,-nbitq), 
to_sfixed(-1269.0/65536.0,1,-nbitq), 
to_sfixed(-1380.0/65536.0,1,-nbitq), 
to_sfixed(-898.0/65536.0,1,-nbitq), 
to_sfixed(3157.0/65536.0,1,-nbitq), 
to_sfixed(2532.0/65536.0,1,-nbitq), 
to_sfixed(-1908.0/65536.0,1,-nbitq), 
to_sfixed(4219.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3877.0/65536.0,1,-nbitq), 
to_sfixed(-1311.0/65536.0,1,-nbitq), 
to_sfixed(-1589.0/65536.0,1,-nbitq), 
to_sfixed(2871.0/65536.0,1,-nbitq), 
to_sfixed(-227.0/65536.0,1,-nbitq), 
to_sfixed(-2040.0/65536.0,1,-nbitq), 
to_sfixed(-86.0/65536.0,1,-nbitq), 
to_sfixed(-526.0/65536.0,1,-nbitq), 
to_sfixed(6961.0/65536.0,1,-nbitq), 
to_sfixed(1956.0/65536.0,1,-nbitq), 
to_sfixed(-814.0/65536.0,1,-nbitq), 
to_sfixed(-10277.0/65536.0,1,-nbitq), 
to_sfixed(1657.0/65536.0,1,-nbitq), 
to_sfixed(3441.0/65536.0,1,-nbitq), 
to_sfixed(317.0/65536.0,1,-nbitq), 
to_sfixed(-50.0/65536.0,1,-nbitq), 
to_sfixed(1110.0/65536.0,1,-nbitq), 
to_sfixed(-2125.0/65536.0,1,-nbitq), 
to_sfixed(-1770.0/65536.0,1,-nbitq), 
to_sfixed(3534.0/65536.0,1,-nbitq), 
to_sfixed(-1158.0/65536.0,1,-nbitq), 
to_sfixed(-640.0/65536.0,1,-nbitq), 
to_sfixed(-8224.0/65536.0,1,-nbitq), 
to_sfixed(3125.0/65536.0,1,-nbitq), 
to_sfixed(-2046.0/65536.0,1,-nbitq), 
to_sfixed(3949.0/65536.0,1,-nbitq), 
to_sfixed(3215.0/65536.0,1,-nbitq), 
to_sfixed(1762.0/65536.0,1,-nbitq), 
to_sfixed(1015.0/65536.0,1,-nbitq), 
to_sfixed(727.0/65536.0,1,-nbitq), 
to_sfixed(-237.0/65536.0,1,-nbitq), 
to_sfixed(-1770.0/65536.0,1,-nbitq), 
to_sfixed(-395.0/65536.0,1,-nbitq), 
to_sfixed(679.0/65536.0,1,-nbitq), 
to_sfixed(184.0/65536.0,1,-nbitq), 
to_sfixed(-1132.0/65536.0,1,-nbitq), 
to_sfixed(4259.0/65536.0,1,-nbitq), 
to_sfixed(2530.0/65536.0,1,-nbitq), 
to_sfixed(143.0/65536.0,1,-nbitq), 
to_sfixed(2550.0/65536.0,1,-nbitq), 
to_sfixed(-43.0/65536.0,1,-nbitq), 
to_sfixed(-1275.0/65536.0,1,-nbitq), 
to_sfixed(-3997.0/65536.0,1,-nbitq), 
to_sfixed(-1979.0/65536.0,1,-nbitq), 
to_sfixed(830.0/65536.0,1,-nbitq), 
to_sfixed(2562.0/65536.0,1,-nbitq), 
to_sfixed(-2860.0/65536.0,1,-nbitq), 
to_sfixed(3819.0/65536.0,1,-nbitq), 
to_sfixed(2214.0/65536.0,1,-nbitq), 
to_sfixed(2864.0/65536.0,1,-nbitq), 
to_sfixed(1651.0/65536.0,1,-nbitq), 
to_sfixed(-3933.0/65536.0,1,-nbitq), 
to_sfixed(-3329.0/65536.0,1,-nbitq), 
to_sfixed(3230.0/65536.0,1,-nbitq), 
to_sfixed(-1239.0/65536.0,1,-nbitq), 
to_sfixed(-2981.0/65536.0,1,-nbitq), 
to_sfixed(3454.0/65536.0,1,-nbitq), 
to_sfixed(510.0/65536.0,1,-nbitq), 
to_sfixed(2752.0/65536.0,1,-nbitq), 
to_sfixed(-7314.0/65536.0,1,-nbitq), 
to_sfixed(1627.0/65536.0,1,-nbitq), 
to_sfixed(-1427.0/65536.0,1,-nbitq), 
to_sfixed(1820.0/65536.0,1,-nbitq), 
to_sfixed(-2802.0/65536.0,1,-nbitq), 
to_sfixed(1305.0/65536.0,1,-nbitq), 
to_sfixed(-1090.0/65536.0,1,-nbitq), 
to_sfixed(5029.0/65536.0,1,-nbitq), 
to_sfixed(4226.0/65536.0,1,-nbitq), 
to_sfixed(9353.0/65536.0,1,-nbitq), 
to_sfixed(-948.0/65536.0,1,-nbitq), 
to_sfixed(-4089.0/65536.0,1,-nbitq), 
to_sfixed(-154.0/65536.0,1,-nbitq), 
to_sfixed(-2550.0/65536.0,1,-nbitq), 
to_sfixed(274.0/65536.0,1,-nbitq), 
to_sfixed(44.0/65536.0,1,-nbitq), 
to_sfixed(-119.0/65536.0,1,-nbitq), 
to_sfixed(2278.0/65536.0,1,-nbitq), 
to_sfixed(689.0/65536.0,1,-nbitq), 
to_sfixed(1238.0/65536.0,1,-nbitq), 
to_sfixed(2453.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4080.0/65536.0,1,-nbitq), 
to_sfixed(1254.0/65536.0,1,-nbitq), 
to_sfixed(-2562.0/65536.0,1,-nbitq), 
to_sfixed(1950.0/65536.0,1,-nbitq), 
to_sfixed(5328.0/65536.0,1,-nbitq), 
to_sfixed(-880.0/65536.0,1,-nbitq), 
to_sfixed(3949.0/65536.0,1,-nbitq), 
to_sfixed(-4578.0/65536.0,1,-nbitq), 
to_sfixed(2747.0/65536.0,1,-nbitq), 
to_sfixed(-630.0/65536.0,1,-nbitq), 
to_sfixed(2434.0/65536.0,1,-nbitq), 
to_sfixed(-10489.0/65536.0,1,-nbitq), 
to_sfixed(576.0/65536.0,1,-nbitq), 
to_sfixed(1048.0/65536.0,1,-nbitq), 
to_sfixed(-1807.0/65536.0,1,-nbitq), 
to_sfixed(135.0/65536.0,1,-nbitq), 
to_sfixed(207.0/65536.0,1,-nbitq), 
to_sfixed(-2659.0/65536.0,1,-nbitq), 
to_sfixed(3744.0/65536.0,1,-nbitq), 
to_sfixed(-1775.0/65536.0,1,-nbitq), 
to_sfixed(-656.0/65536.0,1,-nbitq), 
to_sfixed(-4732.0/65536.0,1,-nbitq), 
to_sfixed(-6164.0/65536.0,1,-nbitq), 
to_sfixed(2010.0/65536.0,1,-nbitq), 
to_sfixed(1723.0/65536.0,1,-nbitq), 
to_sfixed(8753.0/65536.0,1,-nbitq), 
to_sfixed(5238.0/65536.0,1,-nbitq), 
to_sfixed(738.0/65536.0,1,-nbitq), 
to_sfixed(275.0/65536.0,1,-nbitq), 
to_sfixed(-1268.0/65536.0,1,-nbitq), 
to_sfixed(-85.0/65536.0,1,-nbitq), 
to_sfixed(-1658.0/65536.0,1,-nbitq), 
to_sfixed(1677.0/65536.0,1,-nbitq), 
to_sfixed(-2688.0/65536.0,1,-nbitq), 
to_sfixed(-752.0/65536.0,1,-nbitq), 
to_sfixed(-1468.0/65536.0,1,-nbitq), 
to_sfixed(2646.0/65536.0,1,-nbitq), 
to_sfixed(-55.0/65536.0,1,-nbitq), 
to_sfixed(-785.0/65536.0,1,-nbitq), 
to_sfixed(-54.0/65536.0,1,-nbitq), 
to_sfixed(-1500.0/65536.0,1,-nbitq), 
to_sfixed(-1593.0/65536.0,1,-nbitq), 
to_sfixed(-1959.0/65536.0,1,-nbitq), 
to_sfixed(-6144.0/65536.0,1,-nbitq), 
to_sfixed(-2344.0/65536.0,1,-nbitq), 
to_sfixed(717.0/65536.0,1,-nbitq), 
to_sfixed(-3736.0/65536.0,1,-nbitq), 
to_sfixed(2211.0/65536.0,1,-nbitq), 
to_sfixed(2155.0/65536.0,1,-nbitq), 
to_sfixed(-355.0/65536.0,1,-nbitq), 
to_sfixed(866.0/65536.0,1,-nbitq), 
to_sfixed(-3955.0/65536.0,1,-nbitq), 
to_sfixed(-4554.0/65536.0,1,-nbitq), 
to_sfixed(5825.0/65536.0,1,-nbitq), 
to_sfixed(-1250.0/65536.0,1,-nbitq), 
to_sfixed(-167.0/65536.0,1,-nbitq), 
to_sfixed(2858.0/65536.0,1,-nbitq), 
to_sfixed(781.0/65536.0,1,-nbitq), 
to_sfixed(2333.0/65536.0,1,-nbitq), 
to_sfixed(-3919.0/65536.0,1,-nbitq), 
to_sfixed(1664.0/65536.0,1,-nbitq), 
to_sfixed(-1635.0/65536.0,1,-nbitq), 
to_sfixed(2726.0/65536.0,1,-nbitq), 
to_sfixed(-1309.0/65536.0,1,-nbitq), 
to_sfixed(529.0/65536.0,1,-nbitq), 
to_sfixed(-3107.0/65536.0,1,-nbitq), 
to_sfixed(1435.0/65536.0,1,-nbitq), 
to_sfixed(2660.0/65536.0,1,-nbitq), 
to_sfixed(10560.0/65536.0,1,-nbitq), 
to_sfixed(-4273.0/65536.0,1,-nbitq), 
to_sfixed(-645.0/65536.0,1,-nbitq), 
to_sfixed(1582.0/65536.0,1,-nbitq), 
to_sfixed(1170.0/65536.0,1,-nbitq), 
to_sfixed(-1603.0/65536.0,1,-nbitq), 
to_sfixed(-2339.0/65536.0,1,-nbitq), 
to_sfixed(-68.0/65536.0,1,-nbitq), 
to_sfixed(4266.0/65536.0,1,-nbitq), 
to_sfixed(2554.0/65536.0,1,-nbitq), 
to_sfixed(-1168.0/65536.0,1,-nbitq), 
to_sfixed(532.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1708.0/65536.0,1,-nbitq), 
to_sfixed(-3400.0/65536.0,1,-nbitq), 
to_sfixed(2256.0/65536.0,1,-nbitq), 
to_sfixed(6195.0/65536.0,1,-nbitq), 
to_sfixed(10209.0/65536.0,1,-nbitq), 
to_sfixed(2857.0/65536.0,1,-nbitq), 
to_sfixed(5257.0/65536.0,1,-nbitq), 
to_sfixed(-5774.0/65536.0,1,-nbitq), 
to_sfixed(-2305.0/65536.0,1,-nbitq), 
to_sfixed(738.0/65536.0,1,-nbitq), 
to_sfixed(-527.0/65536.0,1,-nbitq), 
to_sfixed(-6417.0/65536.0,1,-nbitq), 
to_sfixed(-905.0/65536.0,1,-nbitq), 
to_sfixed(5433.0/65536.0,1,-nbitq), 
to_sfixed(-1230.0/65536.0,1,-nbitq), 
to_sfixed(-1422.0/65536.0,1,-nbitq), 
to_sfixed(2217.0/65536.0,1,-nbitq), 
to_sfixed(799.0/65536.0,1,-nbitq), 
to_sfixed(2727.0/65536.0,1,-nbitq), 
to_sfixed(3256.0/65536.0,1,-nbitq), 
to_sfixed(-1691.0/65536.0,1,-nbitq), 
to_sfixed(-682.0/65536.0,1,-nbitq), 
to_sfixed(-5207.0/65536.0,1,-nbitq), 
to_sfixed(4244.0/65536.0,1,-nbitq), 
to_sfixed(1091.0/65536.0,1,-nbitq), 
to_sfixed(9359.0/65536.0,1,-nbitq), 
to_sfixed(3378.0/65536.0,1,-nbitq), 
to_sfixed(-696.0/65536.0,1,-nbitq), 
to_sfixed(2594.0/65536.0,1,-nbitq), 
to_sfixed(-1876.0/65536.0,1,-nbitq), 
to_sfixed(3733.0/65536.0,1,-nbitq), 
to_sfixed(-1332.0/65536.0,1,-nbitq), 
to_sfixed(738.0/65536.0,1,-nbitq), 
to_sfixed(-1641.0/65536.0,1,-nbitq), 
to_sfixed(-2869.0/65536.0,1,-nbitq), 
to_sfixed(-3005.0/65536.0,1,-nbitq), 
to_sfixed(3022.0/65536.0,1,-nbitq), 
to_sfixed(1220.0/65536.0,1,-nbitq), 
to_sfixed(-6059.0/65536.0,1,-nbitq), 
to_sfixed(2065.0/65536.0,1,-nbitq), 
to_sfixed(-326.0/65536.0,1,-nbitq), 
to_sfixed(-1949.0/65536.0,1,-nbitq), 
to_sfixed(-2591.0/65536.0,1,-nbitq), 
to_sfixed(-7762.0/65536.0,1,-nbitq), 
to_sfixed(1805.0/65536.0,1,-nbitq), 
to_sfixed(-621.0/65536.0,1,-nbitq), 
to_sfixed(-131.0/65536.0,1,-nbitq), 
to_sfixed(-2725.0/65536.0,1,-nbitq), 
to_sfixed(1921.0/65536.0,1,-nbitq), 
to_sfixed(-1455.0/65536.0,1,-nbitq), 
to_sfixed(-1852.0/65536.0,1,-nbitq), 
to_sfixed(-1647.0/65536.0,1,-nbitq), 
to_sfixed(-3786.0/65536.0,1,-nbitq), 
to_sfixed(2608.0/65536.0,1,-nbitq), 
to_sfixed(-2734.0/65536.0,1,-nbitq), 
to_sfixed(-1554.0/65536.0,1,-nbitq), 
to_sfixed(1437.0/65536.0,1,-nbitq), 
to_sfixed(-2379.0/65536.0,1,-nbitq), 
to_sfixed(74.0/65536.0,1,-nbitq), 
to_sfixed(-2696.0/65536.0,1,-nbitq), 
to_sfixed(-1305.0/65536.0,1,-nbitq), 
to_sfixed(-1650.0/65536.0,1,-nbitq), 
to_sfixed(-1217.0/65536.0,1,-nbitq), 
to_sfixed(471.0/65536.0,1,-nbitq), 
to_sfixed(1103.0/65536.0,1,-nbitq), 
to_sfixed(-2511.0/65536.0,1,-nbitq), 
to_sfixed(5314.0/65536.0,1,-nbitq), 
to_sfixed(6025.0/65536.0,1,-nbitq), 
to_sfixed(3721.0/65536.0,1,-nbitq), 
to_sfixed(-3958.0/65536.0,1,-nbitq), 
to_sfixed(-3171.0/65536.0,1,-nbitq), 
to_sfixed(2216.0/65536.0,1,-nbitq), 
to_sfixed(952.0/65536.0,1,-nbitq), 
to_sfixed(-1325.0/65536.0,1,-nbitq), 
to_sfixed(11.0/65536.0,1,-nbitq), 
to_sfixed(4323.0/65536.0,1,-nbitq), 
to_sfixed(4398.0/65536.0,1,-nbitq), 
to_sfixed(-2027.0/65536.0,1,-nbitq), 
to_sfixed(-1867.0/65536.0,1,-nbitq), 
to_sfixed(3.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3195.0/65536.0,1,-nbitq), 
to_sfixed(-1373.0/65536.0,1,-nbitq), 
to_sfixed(2639.0/65536.0,1,-nbitq), 
to_sfixed(3771.0/65536.0,1,-nbitq), 
to_sfixed(6335.0/65536.0,1,-nbitq), 
to_sfixed(1429.0/65536.0,1,-nbitq), 
to_sfixed(54.0/65536.0,1,-nbitq), 
to_sfixed(-357.0/65536.0,1,-nbitq), 
to_sfixed(-3136.0/65536.0,1,-nbitq), 
to_sfixed(1928.0/65536.0,1,-nbitq), 
to_sfixed(-1154.0/65536.0,1,-nbitq), 
to_sfixed(-1120.0/65536.0,1,-nbitq), 
to_sfixed(-764.0/65536.0,1,-nbitq), 
to_sfixed(6302.0/65536.0,1,-nbitq), 
to_sfixed(-124.0/65536.0,1,-nbitq), 
to_sfixed(-1235.0/65536.0,1,-nbitq), 
to_sfixed(-1372.0/65536.0,1,-nbitq), 
to_sfixed(2179.0/65536.0,1,-nbitq), 
to_sfixed(6887.0/65536.0,1,-nbitq), 
to_sfixed(-2135.0/65536.0,1,-nbitq), 
to_sfixed(-3858.0/65536.0,1,-nbitq), 
to_sfixed(368.0/65536.0,1,-nbitq), 
to_sfixed(-1963.0/65536.0,1,-nbitq), 
to_sfixed(1864.0/65536.0,1,-nbitq), 
to_sfixed(639.0/65536.0,1,-nbitq), 
to_sfixed(10768.0/65536.0,1,-nbitq), 
to_sfixed(1241.0/65536.0,1,-nbitq), 
to_sfixed(-2828.0/65536.0,1,-nbitq), 
to_sfixed(98.0/65536.0,1,-nbitq), 
to_sfixed(-14.0/65536.0,1,-nbitq), 
to_sfixed(682.0/65536.0,1,-nbitq), 
to_sfixed(2512.0/65536.0,1,-nbitq), 
to_sfixed(-1035.0/65536.0,1,-nbitq), 
to_sfixed(2482.0/65536.0,1,-nbitq), 
to_sfixed(-2419.0/65536.0,1,-nbitq), 
to_sfixed(-1935.0/65536.0,1,-nbitq), 
to_sfixed(6407.0/65536.0,1,-nbitq), 
to_sfixed(6675.0/65536.0,1,-nbitq), 
to_sfixed(-6646.0/65536.0,1,-nbitq), 
to_sfixed(3568.0/65536.0,1,-nbitq), 
to_sfixed(4122.0/65536.0,1,-nbitq), 
to_sfixed(563.0/65536.0,1,-nbitq), 
to_sfixed(-2366.0/65536.0,1,-nbitq), 
to_sfixed(-4636.0/65536.0,1,-nbitq), 
to_sfixed(2478.0/65536.0,1,-nbitq), 
to_sfixed(1831.0/65536.0,1,-nbitq), 
to_sfixed(-468.0/65536.0,1,-nbitq), 
to_sfixed(-3537.0/65536.0,1,-nbitq), 
to_sfixed(2355.0/65536.0,1,-nbitq), 
to_sfixed(1073.0/65536.0,1,-nbitq), 
to_sfixed(274.0/65536.0,1,-nbitq), 
to_sfixed(-1939.0/65536.0,1,-nbitq), 
to_sfixed(-426.0/65536.0,1,-nbitq), 
to_sfixed(-2013.0/65536.0,1,-nbitq), 
to_sfixed(60.0/65536.0,1,-nbitq), 
to_sfixed(2477.0/65536.0,1,-nbitq), 
to_sfixed(1420.0/65536.0,1,-nbitq), 
to_sfixed(316.0/65536.0,1,-nbitq), 
to_sfixed(978.0/65536.0,1,-nbitq), 
to_sfixed(-2637.0/65536.0,1,-nbitq), 
to_sfixed(-3754.0/65536.0,1,-nbitq), 
to_sfixed(-2261.0/65536.0,1,-nbitq), 
to_sfixed(-741.0/65536.0,1,-nbitq), 
to_sfixed(-1899.0/65536.0,1,-nbitq), 
to_sfixed(-1691.0/65536.0,1,-nbitq), 
to_sfixed(805.0/65536.0,1,-nbitq), 
to_sfixed(650.0/65536.0,1,-nbitq), 
to_sfixed(1926.0/65536.0,1,-nbitq), 
to_sfixed(4610.0/65536.0,1,-nbitq), 
to_sfixed(-3575.0/65536.0,1,-nbitq), 
to_sfixed(986.0/65536.0,1,-nbitq), 
to_sfixed(1333.0/65536.0,1,-nbitq), 
to_sfixed(-4944.0/65536.0,1,-nbitq), 
to_sfixed(2201.0/65536.0,1,-nbitq), 
to_sfixed(1090.0/65536.0,1,-nbitq), 
to_sfixed(6522.0/65536.0,1,-nbitq), 
to_sfixed(5213.0/65536.0,1,-nbitq), 
to_sfixed(3088.0/65536.0,1,-nbitq), 
to_sfixed(-2932.0/65536.0,1,-nbitq), 
to_sfixed(3544.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-965.0/65536.0,1,-nbitq), 
to_sfixed(-1490.0/65536.0,1,-nbitq), 
to_sfixed(952.0/65536.0,1,-nbitq), 
to_sfixed(784.0/65536.0,1,-nbitq), 
to_sfixed(7174.0/65536.0,1,-nbitq), 
to_sfixed(646.0/65536.0,1,-nbitq), 
to_sfixed(2100.0/65536.0,1,-nbitq), 
to_sfixed(-2432.0/65536.0,1,-nbitq), 
to_sfixed(-2639.0/65536.0,1,-nbitq), 
to_sfixed(-2231.0/65536.0,1,-nbitq), 
to_sfixed(-1175.0/65536.0,1,-nbitq), 
to_sfixed(-6027.0/65536.0,1,-nbitq), 
to_sfixed(1828.0/65536.0,1,-nbitq), 
to_sfixed(3855.0/65536.0,1,-nbitq), 
to_sfixed(412.0/65536.0,1,-nbitq), 
to_sfixed(2289.0/65536.0,1,-nbitq), 
to_sfixed(-1429.0/65536.0,1,-nbitq), 
to_sfixed(-4107.0/65536.0,1,-nbitq), 
to_sfixed(1795.0/65536.0,1,-nbitq), 
to_sfixed(-266.0/65536.0,1,-nbitq), 
to_sfixed(-3650.0/65536.0,1,-nbitq), 
to_sfixed(3256.0/65536.0,1,-nbitq), 
to_sfixed(4326.0/65536.0,1,-nbitq), 
to_sfixed(2260.0/65536.0,1,-nbitq), 
to_sfixed(1920.0/65536.0,1,-nbitq), 
to_sfixed(5048.0/65536.0,1,-nbitq), 
to_sfixed(1233.0/65536.0,1,-nbitq), 
to_sfixed(2546.0/65536.0,1,-nbitq), 
to_sfixed(-1515.0/65536.0,1,-nbitq), 
to_sfixed(2574.0/65536.0,1,-nbitq), 
to_sfixed(1162.0/65536.0,1,-nbitq), 
to_sfixed(-1031.0/65536.0,1,-nbitq), 
to_sfixed(70.0/65536.0,1,-nbitq), 
to_sfixed(-951.0/65536.0,1,-nbitq), 
to_sfixed(-483.0/65536.0,1,-nbitq), 
to_sfixed(-1971.0/65536.0,1,-nbitq), 
to_sfixed(1342.0/65536.0,1,-nbitq), 
to_sfixed(822.0/65536.0,1,-nbitq), 
to_sfixed(-2031.0/65536.0,1,-nbitq), 
to_sfixed(-1202.0/65536.0,1,-nbitq), 
to_sfixed(2191.0/65536.0,1,-nbitq), 
to_sfixed(-68.0/65536.0,1,-nbitq), 
to_sfixed(-6668.0/65536.0,1,-nbitq), 
to_sfixed(-4051.0/65536.0,1,-nbitq), 
to_sfixed(-1792.0/65536.0,1,-nbitq), 
to_sfixed(5402.0/65536.0,1,-nbitq), 
to_sfixed(2669.0/65536.0,1,-nbitq), 
to_sfixed(-735.0/65536.0,1,-nbitq), 
to_sfixed(-1213.0/65536.0,1,-nbitq), 
to_sfixed(1640.0/65536.0,1,-nbitq), 
to_sfixed(2925.0/65536.0,1,-nbitq), 
to_sfixed(-6480.0/65536.0,1,-nbitq), 
to_sfixed(-5503.0/65536.0,1,-nbitq), 
to_sfixed(-2151.0/65536.0,1,-nbitq), 
to_sfixed(1637.0/65536.0,1,-nbitq), 
to_sfixed(-2828.0/65536.0,1,-nbitq), 
to_sfixed(2633.0/65536.0,1,-nbitq), 
to_sfixed(-2118.0/65536.0,1,-nbitq), 
to_sfixed(594.0/65536.0,1,-nbitq), 
to_sfixed(-58.0/65536.0,1,-nbitq), 
to_sfixed(-6562.0/65536.0,1,-nbitq), 
to_sfixed(-767.0/65536.0,1,-nbitq), 
to_sfixed(2518.0/65536.0,1,-nbitq), 
to_sfixed(2111.0/65536.0,1,-nbitq), 
to_sfixed(2996.0/65536.0,1,-nbitq), 
to_sfixed(652.0/65536.0,1,-nbitq), 
to_sfixed(537.0/65536.0,1,-nbitq), 
to_sfixed(2536.0/65536.0,1,-nbitq), 
to_sfixed(-955.0/65536.0,1,-nbitq), 
to_sfixed(-8863.0/65536.0,1,-nbitq), 
to_sfixed(-3531.0/65536.0,1,-nbitq), 
to_sfixed(3325.0/65536.0,1,-nbitq), 
to_sfixed(-703.0/65536.0,1,-nbitq), 
to_sfixed(634.0/65536.0,1,-nbitq), 
to_sfixed(348.0/65536.0,1,-nbitq), 
to_sfixed(2936.0/65536.0,1,-nbitq), 
to_sfixed(2825.0/65536.0,1,-nbitq), 
to_sfixed(-557.0/65536.0,1,-nbitq), 
to_sfixed(-1577.0/65536.0,1,-nbitq), 
to_sfixed(-286.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2503.0/65536.0,1,-nbitq), 
to_sfixed(456.0/65536.0,1,-nbitq), 
to_sfixed(2101.0/65536.0,1,-nbitq), 
to_sfixed(-2952.0/65536.0,1,-nbitq), 
to_sfixed(5053.0/65536.0,1,-nbitq), 
to_sfixed(-3014.0/65536.0,1,-nbitq), 
to_sfixed(2579.0/65536.0,1,-nbitq), 
to_sfixed(-3177.0/65536.0,1,-nbitq), 
to_sfixed(372.0/65536.0,1,-nbitq), 
to_sfixed(2128.0/65536.0,1,-nbitq), 
to_sfixed(-1328.0/65536.0,1,-nbitq), 
to_sfixed(-2039.0/65536.0,1,-nbitq), 
to_sfixed(-1840.0/65536.0,1,-nbitq), 
to_sfixed(2773.0/65536.0,1,-nbitq), 
to_sfixed(1661.0/65536.0,1,-nbitq), 
to_sfixed(-1166.0/65536.0,1,-nbitq), 
to_sfixed(2348.0/65536.0,1,-nbitq), 
to_sfixed(-3744.0/65536.0,1,-nbitq), 
to_sfixed(2586.0/65536.0,1,-nbitq), 
to_sfixed(-2053.0/65536.0,1,-nbitq), 
to_sfixed(-5354.0/65536.0,1,-nbitq), 
to_sfixed(2214.0/65536.0,1,-nbitq), 
to_sfixed(394.0/65536.0,1,-nbitq), 
to_sfixed(6757.0/65536.0,1,-nbitq), 
to_sfixed(175.0/65536.0,1,-nbitq), 
to_sfixed(2723.0/65536.0,1,-nbitq), 
to_sfixed(-582.0/65536.0,1,-nbitq), 
to_sfixed(2160.0/65536.0,1,-nbitq), 
to_sfixed(-5402.0/65536.0,1,-nbitq), 
to_sfixed(2098.0/65536.0,1,-nbitq), 
to_sfixed(-2392.0/65536.0,1,-nbitq), 
to_sfixed(-2183.0/65536.0,1,-nbitq), 
to_sfixed(-2014.0/65536.0,1,-nbitq), 
to_sfixed(-1719.0/65536.0,1,-nbitq), 
to_sfixed(-3458.0/65536.0,1,-nbitq), 
to_sfixed(-606.0/65536.0,1,-nbitq), 
to_sfixed(3272.0/65536.0,1,-nbitq), 
to_sfixed(-1629.0/65536.0,1,-nbitq), 
to_sfixed(511.0/65536.0,1,-nbitq), 
to_sfixed(843.0/65536.0,1,-nbitq), 
to_sfixed(-2250.0/65536.0,1,-nbitq), 
to_sfixed(279.0/65536.0,1,-nbitq), 
to_sfixed(-4974.0/65536.0,1,-nbitq), 
to_sfixed(-3287.0/65536.0,1,-nbitq), 
to_sfixed(-122.0/65536.0,1,-nbitq), 
to_sfixed(2362.0/65536.0,1,-nbitq), 
to_sfixed(-1979.0/65536.0,1,-nbitq), 
to_sfixed(967.0/65536.0,1,-nbitq), 
to_sfixed(-273.0/65536.0,1,-nbitq), 
to_sfixed(4492.0/65536.0,1,-nbitq), 
to_sfixed(-1315.0/65536.0,1,-nbitq), 
to_sfixed(-5646.0/65536.0,1,-nbitq), 
to_sfixed(-4354.0/65536.0,1,-nbitq), 
to_sfixed(-2135.0/65536.0,1,-nbitq), 
to_sfixed(3717.0/65536.0,1,-nbitq), 
to_sfixed(542.0/65536.0,1,-nbitq), 
to_sfixed(782.0/65536.0,1,-nbitq), 
to_sfixed(1497.0/65536.0,1,-nbitq), 
to_sfixed(-602.0/65536.0,1,-nbitq), 
to_sfixed(-2760.0/65536.0,1,-nbitq), 
to_sfixed(-689.0/65536.0,1,-nbitq), 
to_sfixed(-2102.0/65536.0,1,-nbitq), 
to_sfixed(969.0/65536.0,1,-nbitq), 
to_sfixed(-1377.0/65536.0,1,-nbitq), 
to_sfixed(-2095.0/65536.0,1,-nbitq), 
to_sfixed(-1139.0/65536.0,1,-nbitq), 
to_sfixed(-2937.0/65536.0,1,-nbitq), 
to_sfixed(-949.0/65536.0,1,-nbitq), 
to_sfixed(410.0/65536.0,1,-nbitq), 
to_sfixed(-5543.0/65536.0,1,-nbitq), 
to_sfixed(1513.0/65536.0,1,-nbitq), 
to_sfixed(2033.0/65536.0,1,-nbitq), 
to_sfixed(-653.0/65536.0,1,-nbitq), 
to_sfixed(274.0/65536.0,1,-nbitq), 
to_sfixed(656.0/65536.0,1,-nbitq), 
to_sfixed(-1664.0/65536.0,1,-nbitq), 
to_sfixed(1532.0/65536.0,1,-nbitq), 
to_sfixed(1101.0/65536.0,1,-nbitq), 
to_sfixed(-3552.0/65536.0,1,-nbitq), 
to_sfixed(2242.0/65536.0,1,-nbitq)  ), 
( to_sfixed(918.0/65536.0,1,-nbitq), 
to_sfixed(-3207.0/65536.0,1,-nbitq), 
to_sfixed(932.0/65536.0,1,-nbitq), 
to_sfixed(-1017.0/65536.0,1,-nbitq), 
to_sfixed(4794.0/65536.0,1,-nbitq), 
to_sfixed(-4502.0/65536.0,1,-nbitq), 
to_sfixed(2349.0/65536.0,1,-nbitq), 
to_sfixed(-1716.0/65536.0,1,-nbitq), 
to_sfixed(-462.0/65536.0,1,-nbitq), 
to_sfixed(-2939.0/65536.0,1,-nbitq), 
to_sfixed(1798.0/65536.0,1,-nbitq), 
to_sfixed(3797.0/65536.0,1,-nbitq), 
to_sfixed(-2476.0/65536.0,1,-nbitq), 
to_sfixed(5204.0/65536.0,1,-nbitq), 
to_sfixed(-1749.0/65536.0,1,-nbitq), 
to_sfixed(-1407.0/65536.0,1,-nbitq), 
to_sfixed(-1674.0/65536.0,1,-nbitq), 
to_sfixed(-4267.0/65536.0,1,-nbitq), 
to_sfixed(4023.0/65536.0,1,-nbitq), 
to_sfixed(610.0/65536.0,1,-nbitq), 
to_sfixed(-3618.0/65536.0,1,-nbitq), 
to_sfixed(-465.0/65536.0,1,-nbitq), 
to_sfixed(3772.0/65536.0,1,-nbitq), 
to_sfixed(4148.0/65536.0,1,-nbitq), 
to_sfixed(-3733.0/65536.0,1,-nbitq), 
to_sfixed(-957.0/65536.0,1,-nbitq), 
to_sfixed(1582.0/65536.0,1,-nbitq), 
to_sfixed(-1838.0/65536.0,1,-nbitq), 
to_sfixed(-237.0/65536.0,1,-nbitq), 
to_sfixed(-1568.0/65536.0,1,-nbitq), 
to_sfixed(-1190.0/65536.0,1,-nbitq), 
to_sfixed(755.0/65536.0,1,-nbitq), 
to_sfixed(2031.0/65536.0,1,-nbitq), 
to_sfixed(915.0/65536.0,1,-nbitq), 
to_sfixed(2269.0/65536.0,1,-nbitq), 
to_sfixed(-2736.0/65536.0,1,-nbitq), 
to_sfixed(2484.0/65536.0,1,-nbitq), 
to_sfixed(-4502.0/65536.0,1,-nbitq), 
to_sfixed(2697.0/65536.0,1,-nbitq), 
to_sfixed(236.0/65536.0,1,-nbitq), 
to_sfixed(-269.0/65536.0,1,-nbitq), 
to_sfixed(-2528.0/65536.0,1,-nbitq), 
to_sfixed(-7761.0/65536.0,1,-nbitq), 
to_sfixed(-286.0/65536.0,1,-nbitq), 
to_sfixed(-2648.0/65536.0,1,-nbitq), 
to_sfixed(5945.0/65536.0,1,-nbitq), 
to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(497.0/65536.0,1,-nbitq), 
to_sfixed(1903.0/65536.0,1,-nbitq), 
to_sfixed(3000.0/65536.0,1,-nbitq), 
to_sfixed(-2158.0/65536.0,1,-nbitq), 
to_sfixed(-4377.0/65536.0,1,-nbitq), 
to_sfixed(-4658.0/65536.0,1,-nbitq), 
to_sfixed(-1150.0/65536.0,1,-nbitq), 
to_sfixed(4398.0/65536.0,1,-nbitq), 
to_sfixed(438.0/65536.0,1,-nbitq), 
to_sfixed(2442.0/65536.0,1,-nbitq), 
to_sfixed(941.0/65536.0,1,-nbitq), 
to_sfixed(-1945.0/65536.0,1,-nbitq), 
to_sfixed(2209.0/65536.0,1,-nbitq), 
to_sfixed(128.0/65536.0,1,-nbitq), 
to_sfixed(-3148.0/65536.0,1,-nbitq), 
to_sfixed(-675.0/65536.0,1,-nbitq), 
to_sfixed(-1078.0/65536.0,1,-nbitq), 
to_sfixed(998.0/65536.0,1,-nbitq), 
to_sfixed(-1557.0/65536.0,1,-nbitq), 
to_sfixed(365.0/65536.0,1,-nbitq), 
to_sfixed(1403.0/65536.0,1,-nbitq), 
to_sfixed(-212.0/65536.0,1,-nbitq), 
to_sfixed(-3353.0/65536.0,1,-nbitq), 
to_sfixed(2272.0/65536.0,1,-nbitq), 
to_sfixed(1941.0/65536.0,1,-nbitq), 
to_sfixed(-2516.0/65536.0,1,-nbitq), 
to_sfixed(896.0/65536.0,1,-nbitq), 
to_sfixed(-2214.0/65536.0,1,-nbitq), 
to_sfixed(-2275.0/65536.0,1,-nbitq), 
to_sfixed(1285.0/65536.0,1,-nbitq), 
to_sfixed(-1401.0/65536.0,1,-nbitq), 
to_sfixed(-372.0/65536.0,1,-nbitq), 
to_sfixed(1085.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-39.0/65536.0,1,-nbitq), 
to_sfixed(-289.0/65536.0,1,-nbitq), 
to_sfixed(5980.0/65536.0,1,-nbitq), 
to_sfixed(-4146.0/65536.0,1,-nbitq), 
to_sfixed(5008.0/65536.0,1,-nbitq), 
to_sfixed(-1380.0/65536.0,1,-nbitq), 
to_sfixed(-2376.0/65536.0,1,-nbitq), 
to_sfixed(-655.0/65536.0,1,-nbitq), 
to_sfixed(81.0/65536.0,1,-nbitq), 
to_sfixed(1655.0/65536.0,1,-nbitq), 
to_sfixed(2926.0/65536.0,1,-nbitq), 
to_sfixed(2959.0/65536.0,1,-nbitq), 
to_sfixed(-3235.0/65536.0,1,-nbitq), 
to_sfixed(1547.0/65536.0,1,-nbitq), 
to_sfixed(-3329.0/65536.0,1,-nbitq), 
to_sfixed(586.0/65536.0,1,-nbitq), 
to_sfixed(-2187.0/65536.0,1,-nbitq), 
to_sfixed(-1089.0/65536.0,1,-nbitq), 
to_sfixed(833.0/65536.0,1,-nbitq), 
to_sfixed(-1319.0/65536.0,1,-nbitq), 
to_sfixed(-675.0/65536.0,1,-nbitq), 
to_sfixed(-26.0/65536.0,1,-nbitq), 
to_sfixed(-1518.0/65536.0,1,-nbitq), 
to_sfixed(4874.0/65536.0,1,-nbitq), 
to_sfixed(1101.0/65536.0,1,-nbitq), 
to_sfixed(-1059.0/65536.0,1,-nbitq), 
to_sfixed(50.0/65536.0,1,-nbitq), 
to_sfixed(1327.0/65536.0,1,-nbitq), 
to_sfixed(-939.0/65536.0,1,-nbitq), 
to_sfixed(2746.0/65536.0,1,-nbitq), 
to_sfixed(-3816.0/65536.0,1,-nbitq), 
to_sfixed(-2024.0/65536.0,1,-nbitq), 
to_sfixed(956.0/65536.0,1,-nbitq), 
to_sfixed(1872.0/65536.0,1,-nbitq), 
to_sfixed(1613.0/65536.0,1,-nbitq), 
to_sfixed(691.0/65536.0,1,-nbitq), 
to_sfixed(487.0/65536.0,1,-nbitq), 
to_sfixed(-2559.0/65536.0,1,-nbitq), 
to_sfixed(1875.0/65536.0,1,-nbitq), 
to_sfixed(597.0/65536.0,1,-nbitq), 
to_sfixed(-4498.0/65536.0,1,-nbitq), 
to_sfixed(1934.0/65536.0,1,-nbitq), 
to_sfixed(-2072.0/65536.0,1,-nbitq), 
to_sfixed(2514.0/65536.0,1,-nbitq), 
to_sfixed(322.0/65536.0,1,-nbitq), 
to_sfixed(4714.0/65536.0,1,-nbitq), 
to_sfixed(-848.0/65536.0,1,-nbitq), 
to_sfixed(-518.0/65536.0,1,-nbitq), 
to_sfixed(-697.0/65536.0,1,-nbitq), 
to_sfixed(1063.0/65536.0,1,-nbitq), 
to_sfixed(-938.0/65536.0,1,-nbitq), 
to_sfixed(-5014.0/65536.0,1,-nbitq), 
to_sfixed(-188.0/65536.0,1,-nbitq), 
to_sfixed(2563.0/65536.0,1,-nbitq), 
to_sfixed(5000.0/65536.0,1,-nbitq), 
to_sfixed(320.0/65536.0,1,-nbitq), 
to_sfixed(-1969.0/65536.0,1,-nbitq), 
to_sfixed(2003.0/65536.0,1,-nbitq), 
to_sfixed(-2410.0/65536.0,1,-nbitq), 
to_sfixed(2901.0/65536.0,1,-nbitq), 
to_sfixed(1570.0/65536.0,1,-nbitq), 
to_sfixed(-1859.0/65536.0,1,-nbitq), 
to_sfixed(-937.0/65536.0,1,-nbitq), 
to_sfixed(2090.0/65536.0,1,-nbitq), 
to_sfixed(8.0/65536.0,1,-nbitq), 
to_sfixed(2933.0/65536.0,1,-nbitq), 
to_sfixed(-1957.0/65536.0,1,-nbitq), 
to_sfixed(-3893.0/65536.0,1,-nbitq), 
to_sfixed(-3038.0/65536.0,1,-nbitq), 
to_sfixed(-3214.0/65536.0,1,-nbitq), 
to_sfixed(1883.0/65536.0,1,-nbitq), 
to_sfixed(-1062.0/65536.0,1,-nbitq), 
to_sfixed(492.0/65536.0,1,-nbitq), 
to_sfixed(176.0/65536.0,1,-nbitq), 
to_sfixed(1261.0/65536.0,1,-nbitq), 
to_sfixed(2820.0/65536.0,1,-nbitq), 
to_sfixed(-1460.0/65536.0,1,-nbitq), 
to_sfixed(3040.0/65536.0,1,-nbitq), 
to_sfixed(1036.0/65536.0,1,-nbitq), 
to_sfixed(4657.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1737.0/65536.0,1,-nbitq), 
to_sfixed(718.0/65536.0,1,-nbitq), 
to_sfixed(4583.0/65536.0,1,-nbitq), 
to_sfixed(-555.0/65536.0,1,-nbitq), 
to_sfixed(2171.0/65536.0,1,-nbitq), 
to_sfixed(-3584.0/65536.0,1,-nbitq), 
to_sfixed(-1758.0/65536.0,1,-nbitq), 
to_sfixed(-2880.0/65536.0,1,-nbitq), 
to_sfixed(521.0/65536.0,1,-nbitq), 
to_sfixed(355.0/65536.0,1,-nbitq), 
to_sfixed(-2367.0/65536.0,1,-nbitq), 
to_sfixed(-347.0/65536.0,1,-nbitq), 
to_sfixed(-2691.0/65536.0,1,-nbitq), 
to_sfixed(2214.0/65536.0,1,-nbitq), 
to_sfixed(-2046.0/65536.0,1,-nbitq), 
to_sfixed(2538.0/65536.0,1,-nbitq), 
to_sfixed(1685.0/65536.0,1,-nbitq), 
to_sfixed(390.0/65536.0,1,-nbitq), 
to_sfixed(-1107.0/65536.0,1,-nbitq), 
to_sfixed(-120.0/65536.0,1,-nbitq), 
to_sfixed(-544.0/65536.0,1,-nbitq), 
to_sfixed(3001.0/65536.0,1,-nbitq), 
to_sfixed(3739.0/65536.0,1,-nbitq), 
to_sfixed(-1397.0/65536.0,1,-nbitq), 
to_sfixed(-708.0/65536.0,1,-nbitq), 
to_sfixed(-1927.0/65536.0,1,-nbitq), 
to_sfixed(355.0/65536.0,1,-nbitq), 
to_sfixed(2341.0/65536.0,1,-nbitq), 
to_sfixed(2108.0/65536.0,1,-nbitq), 
to_sfixed(-557.0/65536.0,1,-nbitq), 
to_sfixed(-3267.0/65536.0,1,-nbitq), 
to_sfixed(-2937.0/65536.0,1,-nbitq), 
to_sfixed(-2841.0/65536.0,1,-nbitq), 
to_sfixed(-2738.0/65536.0,1,-nbitq), 
to_sfixed(-2565.0/65536.0,1,-nbitq), 
to_sfixed(2351.0/65536.0,1,-nbitq), 
to_sfixed(2374.0/65536.0,1,-nbitq), 
to_sfixed(-1756.0/65536.0,1,-nbitq), 
to_sfixed(1162.0/65536.0,1,-nbitq), 
to_sfixed(2130.0/65536.0,1,-nbitq), 
to_sfixed(-6471.0/65536.0,1,-nbitq), 
to_sfixed(-3130.0/65536.0,1,-nbitq), 
to_sfixed(-1446.0/65536.0,1,-nbitq), 
to_sfixed(-447.0/65536.0,1,-nbitq), 
to_sfixed(-1739.0/65536.0,1,-nbitq), 
to_sfixed(1228.0/65536.0,1,-nbitq), 
to_sfixed(1482.0/65536.0,1,-nbitq), 
to_sfixed(2800.0/65536.0,1,-nbitq), 
to_sfixed(1446.0/65536.0,1,-nbitq), 
to_sfixed(1004.0/65536.0,1,-nbitq), 
to_sfixed(880.0/65536.0,1,-nbitq), 
to_sfixed(-4883.0/65536.0,1,-nbitq), 
to_sfixed(497.0/65536.0,1,-nbitq), 
to_sfixed(-3135.0/65536.0,1,-nbitq), 
to_sfixed(881.0/65536.0,1,-nbitq), 
to_sfixed(13.0/65536.0,1,-nbitq), 
to_sfixed(2194.0/65536.0,1,-nbitq), 
to_sfixed(-1705.0/65536.0,1,-nbitq), 
to_sfixed(1797.0/65536.0,1,-nbitq), 
to_sfixed(4451.0/65536.0,1,-nbitq), 
to_sfixed(1466.0/65536.0,1,-nbitq), 
to_sfixed(2350.0/65536.0,1,-nbitq), 
to_sfixed(1762.0/65536.0,1,-nbitq), 
to_sfixed(517.0/65536.0,1,-nbitq), 
to_sfixed(975.0/65536.0,1,-nbitq), 
to_sfixed(-184.0/65536.0,1,-nbitq), 
to_sfixed(-3705.0/65536.0,1,-nbitq), 
to_sfixed(-3847.0/65536.0,1,-nbitq), 
to_sfixed(-194.0/65536.0,1,-nbitq), 
to_sfixed(-1714.0/65536.0,1,-nbitq), 
to_sfixed(-30.0/65536.0,1,-nbitq), 
to_sfixed(-4075.0/65536.0,1,-nbitq), 
to_sfixed(392.0/65536.0,1,-nbitq), 
to_sfixed(1784.0/65536.0,1,-nbitq), 
to_sfixed(-979.0/65536.0,1,-nbitq), 
to_sfixed(-487.0/65536.0,1,-nbitq), 
to_sfixed(273.0/65536.0,1,-nbitq), 
to_sfixed(3677.0/65536.0,1,-nbitq), 
to_sfixed(-842.0/65536.0,1,-nbitq), 
to_sfixed(-712.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-834.0/65536.0,1,-nbitq), 
to_sfixed(2604.0/65536.0,1,-nbitq), 
to_sfixed(2470.0/65536.0,1,-nbitq), 
to_sfixed(917.0/65536.0,1,-nbitq), 
to_sfixed(-1413.0/65536.0,1,-nbitq), 
to_sfixed(-4068.0/65536.0,1,-nbitq), 
to_sfixed(132.0/65536.0,1,-nbitq), 
to_sfixed(-1421.0/65536.0,1,-nbitq), 
to_sfixed(-2266.0/65536.0,1,-nbitq), 
to_sfixed(-610.0/65536.0,1,-nbitq), 
to_sfixed(441.0/65536.0,1,-nbitq), 
to_sfixed(-2423.0/65536.0,1,-nbitq), 
to_sfixed(-36.0/65536.0,1,-nbitq), 
to_sfixed(-3097.0/65536.0,1,-nbitq), 
to_sfixed(-2828.0/65536.0,1,-nbitq), 
to_sfixed(226.0/65536.0,1,-nbitq), 
to_sfixed(1185.0/65536.0,1,-nbitq), 
to_sfixed(224.0/65536.0,1,-nbitq), 
to_sfixed(2841.0/65536.0,1,-nbitq), 
to_sfixed(3048.0/65536.0,1,-nbitq), 
to_sfixed(1037.0/65536.0,1,-nbitq), 
to_sfixed(1289.0/65536.0,1,-nbitq), 
to_sfixed(3164.0/65536.0,1,-nbitq), 
to_sfixed(1393.0/65536.0,1,-nbitq), 
to_sfixed(231.0/65536.0,1,-nbitq), 
to_sfixed(-442.0/65536.0,1,-nbitq), 
to_sfixed(943.0/65536.0,1,-nbitq), 
to_sfixed(236.0/65536.0,1,-nbitq), 
to_sfixed(-1439.0/65536.0,1,-nbitq), 
to_sfixed(835.0/65536.0,1,-nbitq), 
to_sfixed(-2726.0/65536.0,1,-nbitq), 
to_sfixed(248.0/65536.0,1,-nbitq), 
to_sfixed(229.0/65536.0,1,-nbitq), 
to_sfixed(326.0/65536.0,1,-nbitq), 
to_sfixed(1822.0/65536.0,1,-nbitq), 
to_sfixed(1142.0/65536.0,1,-nbitq), 
to_sfixed(-2110.0/65536.0,1,-nbitq), 
to_sfixed(824.0/65536.0,1,-nbitq), 
to_sfixed(1444.0/65536.0,1,-nbitq), 
to_sfixed(-1626.0/65536.0,1,-nbitq), 
to_sfixed(-1350.0/65536.0,1,-nbitq), 
to_sfixed(2267.0/65536.0,1,-nbitq), 
to_sfixed(-3247.0/65536.0,1,-nbitq), 
to_sfixed(-1867.0/65536.0,1,-nbitq), 
to_sfixed(142.0/65536.0,1,-nbitq), 
to_sfixed(3836.0/65536.0,1,-nbitq), 
to_sfixed(3181.0/65536.0,1,-nbitq), 
to_sfixed(-917.0/65536.0,1,-nbitq), 
to_sfixed(-897.0/65536.0,1,-nbitq), 
to_sfixed(298.0/65536.0,1,-nbitq), 
to_sfixed(-1483.0/65536.0,1,-nbitq), 
to_sfixed(-1140.0/65536.0,1,-nbitq), 
to_sfixed(-1966.0/65536.0,1,-nbitq), 
to_sfixed(-3128.0/65536.0,1,-nbitq), 
to_sfixed(3972.0/65536.0,1,-nbitq), 
to_sfixed(-14.0/65536.0,1,-nbitq), 
to_sfixed(2431.0/65536.0,1,-nbitq), 
to_sfixed(-890.0/65536.0,1,-nbitq), 
to_sfixed(1775.0/65536.0,1,-nbitq), 
to_sfixed(5465.0/65536.0,1,-nbitq), 
to_sfixed(-3340.0/65536.0,1,-nbitq), 
to_sfixed(1079.0/65536.0,1,-nbitq), 
to_sfixed(3113.0/65536.0,1,-nbitq), 
to_sfixed(-1437.0/65536.0,1,-nbitq), 
to_sfixed(129.0/65536.0,1,-nbitq), 
to_sfixed(3506.0/65536.0,1,-nbitq), 
to_sfixed(-553.0/65536.0,1,-nbitq), 
to_sfixed(-3813.0/65536.0,1,-nbitq), 
to_sfixed(-1072.0/65536.0,1,-nbitq), 
to_sfixed(266.0/65536.0,1,-nbitq), 
to_sfixed(160.0/65536.0,1,-nbitq), 
to_sfixed(-1676.0/65536.0,1,-nbitq), 
to_sfixed(270.0/65536.0,1,-nbitq), 
to_sfixed(-2817.0/65536.0,1,-nbitq), 
to_sfixed(-1104.0/65536.0,1,-nbitq), 
to_sfixed(4744.0/65536.0,1,-nbitq), 
to_sfixed(-554.0/65536.0,1,-nbitq), 
to_sfixed(1737.0/65536.0,1,-nbitq), 
to_sfixed(-515.0/65536.0,1,-nbitq), 
to_sfixed(4129.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-450.0/65536.0,1,-nbitq), 
to_sfixed(2606.0/65536.0,1,-nbitq), 
to_sfixed(4324.0/65536.0,1,-nbitq), 
to_sfixed(441.0/65536.0,1,-nbitq), 
to_sfixed(-2256.0/65536.0,1,-nbitq), 
to_sfixed(-4431.0/65536.0,1,-nbitq), 
to_sfixed(1998.0/65536.0,1,-nbitq), 
to_sfixed(196.0/65536.0,1,-nbitq), 
to_sfixed(-2151.0/65536.0,1,-nbitq), 
to_sfixed(-1525.0/65536.0,1,-nbitq), 
to_sfixed(807.0/65536.0,1,-nbitq), 
to_sfixed(-960.0/65536.0,1,-nbitq), 
to_sfixed(1459.0/65536.0,1,-nbitq), 
to_sfixed(-2142.0/65536.0,1,-nbitq), 
to_sfixed(2054.0/65536.0,1,-nbitq), 
to_sfixed(-20.0/65536.0,1,-nbitq), 
to_sfixed(-2515.0/65536.0,1,-nbitq), 
to_sfixed(3023.0/65536.0,1,-nbitq), 
to_sfixed(1653.0/65536.0,1,-nbitq), 
to_sfixed(2759.0/65536.0,1,-nbitq), 
to_sfixed(-3352.0/65536.0,1,-nbitq), 
to_sfixed(2420.0/65536.0,1,-nbitq), 
to_sfixed(1014.0/65536.0,1,-nbitq), 
to_sfixed(-897.0/65536.0,1,-nbitq), 
to_sfixed(-2108.0/65536.0,1,-nbitq), 
to_sfixed(439.0/65536.0,1,-nbitq), 
to_sfixed(-840.0/65536.0,1,-nbitq), 
to_sfixed(2006.0/65536.0,1,-nbitq), 
to_sfixed(-2240.0/65536.0,1,-nbitq), 
to_sfixed(-492.0/65536.0,1,-nbitq), 
to_sfixed(-1698.0/65536.0,1,-nbitq), 
to_sfixed(1997.0/65536.0,1,-nbitq), 
to_sfixed(94.0/65536.0,1,-nbitq), 
to_sfixed(-1821.0/65536.0,1,-nbitq), 
to_sfixed(2798.0/65536.0,1,-nbitq), 
to_sfixed(-941.0/65536.0,1,-nbitq), 
to_sfixed(1693.0/65536.0,1,-nbitq), 
to_sfixed(-3867.0/65536.0,1,-nbitq), 
to_sfixed(-2592.0/65536.0,1,-nbitq), 
to_sfixed(-785.0/65536.0,1,-nbitq), 
to_sfixed(-4015.0/65536.0,1,-nbitq), 
to_sfixed(-2461.0/65536.0,1,-nbitq), 
to_sfixed(-4297.0/65536.0,1,-nbitq), 
to_sfixed(3671.0/65536.0,1,-nbitq), 
to_sfixed(1896.0/65536.0,1,-nbitq), 
to_sfixed(4724.0/65536.0,1,-nbitq), 
to_sfixed(1442.0/65536.0,1,-nbitq), 
to_sfixed(2079.0/65536.0,1,-nbitq), 
to_sfixed(3258.0/65536.0,1,-nbitq), 
to_sfixed(2523.0/65536.0,1,-nbitq), 
to_sfixed(-1520.0/65536.0,1,-nbitq), 
to_sfixed(2199.0/65536.0,1,-nbitq), 
to_sfixed(1482.0/65536.0,1,-nbitq), 
to_sfixed(-2107.0/65536.0,1,-nbitq), 
to_sfixed(2815.0/65536.0,1,-nbitq), 
to_sfixed(2009.0/65536.0,1,-nbitq), 
to_sfixed(-1281.0/65536.0,1,-nbitq), 
to_sfixed(-1444.0/65536.0,1,-nbitq), 
to_sfixed(-1595.0/65536.0,1,-nbitq), 
to_sfixed(4123.0/65536.0,1,-nbitq), 
to_sfixed(1144.0/65536.0,1,-nbitq), 
to_sfixed(-2417.0/65536.0,1,-nbitq), 
to_sfixed(1409.0/65536.0,1,-nbitq), 
to_sfixed(-2494.0/65536.0,1,-nbitq), 
to_sfixed(1756.0/65536.0,1,-nbitq), 
to_sfixed(-1833.0/65536.0,1,-nbitq), 
to_sfixed(2294.0/65536.0,1,-nbitq), 
to_sfixed(-2723.0/65536.0,1,-nbitq), 
to_sfixed(785.0/65536.0,1,-nbitq), 
to_sfixed(2197.0/65536.0,1,-nbitq), 
to_sfixed(2872.0/65536.0,1,-nbitq), 
to_sfixed(2281.0/65536.0,1,-nbitq), 
to_sfixed(1350.0/65536.0,1,-nbitq), 
to_sfixed(-1412.0/65536.0,1,-nbitq), 
to_sfixed(-2888.0/65536.0,1,-nbitq), 
to_sfixed(1023.0/65536.0,1,-nbitq), 
to_sfixed(-2337.0/65536.0,1,-nbitq), 
to_sfixed(247.0/65536.0,1,-nbitq), 
to_sfixed(1603.0/65536.0,1,-nbitq), 
to_sfixed(-1093.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3178.0/65536.0,1,-nbitq), 
to_sfixed(1420.0/65536.0,1,-nbitq), 
to_sfixed(250.0/65536.0,1,-nbitq), 
to_sfixed(89.0/65536.0,1,-nbitq), 
to_sfixed(-2973.0/65536.0,1,-nbitq), 
to_sfixed(642.0/65536.0,1,-nbitq), 
to_sfixed(1891.0/65536.0,1,-nbitq), 
to_sfixed(-1135.0/65536.0,1,-nbitq), 
to_sfixed(-1041.0/65536.0,1,-nbitq), 
to_sfixed(1068.0/65536.0,1,-nbitq), 
to_sfixed(-3242.0/65536.0,1,-nbitq), 
to_sfixed(2103.0/65536.0,1,-nbitq), 
to_sfixed(-1318.0/65536.0,1,-nbitq), 
to_sfixed(-560.0/65536.0,1,-nbitq), 
to_sfixed(-2551.0/65536.0,1,-nbitq), 
to_sfixed(2302.0/65536.0,1,-nbitq), 
to_sfixed(-826.0/65536.0,1,-nbitq), 
to_sfixed(1324.0/65536.0,1,-nbitq), 
to_sfixed(-1030.0/65536.0,1,-nbitq), 
to_sfixed(2432.0/65536.0,1,-nbitq), 
to_sfixed(924.0/65536.0,1,-nbitq), 
to_sfixed(1819.0/65536.0,1,-nbitq), 
to_sfixed(560.0/65536.0,1,-nbitq), 
to_sfixed(495.0/65536.0,1,-nbitq), 
to_sfixed(2919.0/65536.0,1,-nbitq), 
to_sfixed(1468.0/65536.0,1,-nbitq), 
to_sfixed(69.0/65536.0,1,-nbitq), 
to_sfixed(3076.0/65536.0,1,-nbitq), 
to_sfixed(-401.0/65536.0,1,-nbitq), 
to_sfixed(-1329.0/65536.0,1,-nbitq), 
to_sfixed(-2983.0/65536.0,1,-nbitq), 
to_sfixed(2867.0/65536.0,1,-nbitq), 
to_sfixed(-2385.0/65536.0,1,-nbitq), 
to_sfixed(-3704.0/65536.0,1,-nbitq), 
to_sfixed(1411.0/65536.0,1,-nbitq), 
to_sfixed(-2091.0/65536.0,1,-nbitq), 
to_sfixed(-1849.0/65536.0,1,-nbitq), 
to_sfixed(-2217.0/65536.0,1,-nbitq), 
to_sfixed(-324.0/65536.0,1,-nbitq), 
to_sfixed(1762.0/65536.0,1,-nbitq), 
to_sfixed(-62.0/65536.0,1,-nbitq), 
to_sfixed(-2722.0/65536.0,1,-nbitq), 
to_sfixed(-1102.0/65536.0,1,-nbitq), 
to_sfixed(216.0/65536.0,1,-nbitq), 
to_sfixed(2116.0/65536.0,1,-nbitq), 
to_sfixed(2093.0/65536.0,1,-nbitq), 
to_sfixed(-1231.0/65536.0,1,-nbitq), 
to_sfixed(2660.0/65536.0,1,-nbitq), 
to_sfixed(3470.0/65536.0,1,-nbitq), 
to_sfixed(4467.0/65536.0,1,-nbitq), 
to_sfixed(1713.0/65536.0,1,-nbitq), 
to_sfixed(756.0/65536.0,1,-nbitq), 
to_sfixed(576.0/65536.0,1,-nbitq), 
to_sfixed(-633.0/65536.0,1,-nbitq), 
to_sfixed(578.0/65536.0,1,-nbitq), 
to_sfixed(-1731.0/65536.0,1,-nbitq), 
to_sfixed(2293.0/65536.0,1,-nbitq), 
to_sfixed(-2738.0/65536.0,1,-nbitq), 
to_sfixed(263.0/65536.0,1,-nbitq), 
to_sfixed(4590.0/65536.0,1,-nbitq), 
to_sfixed(-3872.0/65536.0,1,-nbitq), 
to_sfixed(-941.0/65536.0,1,-nbitq), 
to_sfixed(1147.0/65536.0,1,-nbitq), 
to_sfixed(-1067.0/65536.0,1,-nbitq), 
to_sfixed(1057.0/65536.0,1,-nbitq), 
to_sfixed(-225.0/65536.0,1,-nbitq), 
to_sfixed(1777.0/65536.0,1,-nbitq), 
to_sfixed(1324.0/65536.0,1,-nbitq), 
to_sfixed(3498.0/65536.0,1,-nbitq), 
to_sfixed(-2601.0/65536.0,1,-nbitq), 
to_sfixed(2777.0/65536.0,1,-nbitq), 
to_sfixed(-208.0/65536.0,1,-nbitq), 
to_sfixed(2217.0/65536.0,1,-nbitq), 
to_sfixed(1588.0/65536.0,1,-nbitq), 
to_sfixed(-47.0/65536.0,1,-nbitq), 
to_sfixed(-1875.0/65536.0,1,-nbitq), 
to_sfixed(2855.0/65536.0,1,-nbitq), 
to_sfixed(4288.0/65536.0,1,-nbitq), 
to_sfixed(1074.0/65536.0,1,-nbitq), 
to_sfixed(3189.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-247.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(3178.0/65536.0,1,-nbitq), 
to_sfixed(1852.0/65536.0,1,-nbitq), 
to_sfixed(1035.0/65536.0,1,-nbitq), 
to_sfixed(342.0/65536.0,1,-nbitq), 
to_sfixed(2702.0/65536.0,1,-nbitq), 
to_sfixed(2405.0/65536.0,1,-nbitq), 
to_sfixed(-255.0/65536.0,1,-nbitq), 
to_sfixed(2665.0/65536.0,1,-nbitq), 
to_sfixed(1579.0/65536.0,1,-nbitq), 
to_sfixed(-460.0/65536.0,1,-nbitq), 
to_sfixed(50.0/65536.0,1,-nbitq), 
to_sfixed(6.0/65536.0,1,-nbitq), 
to_sfixed(1574.0/65536.0,1,-nbitq), 
to_sfixed(-2817.0/65536.0,1,-nbitq), 
to_sfixed(-3124.0/65536.0,1,-nbitq), 
to_sfixed(2600.0/65536.0,1,-nbitq), 
to_sfixed(993.0/65536.0,1,-nbitq), 
to_sfixed(1335.0/65536.0,1,-nbitq), 
to_sfixed(-2796.0/65536.0,1,-nbitq), 
to_sfixed(3606.0/65536.0,1,-nbitq), 
to_sfixed(-277.0/65536.0,1,-nbitq), 
to_sfixed(-760.0/65536.0,1,-nbitq), 
to_sfixed(178.0/65536.0,1,-nbitq), 
to_sfixed(90.0/65536.0,1,-nbitq), 
to_sfixed(-2382.0/65536.0,1,-nbitq), 
to_sfixed(1705.0/65536.0,1,-nbitq), 
to_sfixed(-2100.0/65536.0,1,-nbitq), 
to_sfixed(-2449.0/65536.0,1,-nbitq), 
to_sfixed(-1118.0/65536.0,1,-nbitq), 
to_sfixed(1276.0/65536.0,1,-nbitq), 
to_sfixed(-5268.0/65536.0,1,-nbitq), 
to_sfixed(-3497.0/65536.0,1,-nbitq), 
to_sfixed(1780.0/65536.0,1,-nbitq), 
to_sfixed(-1409.0/65536.0,1,-nbitq), 
to_sfixed(-1510.0/65536.0,1,-nbitq), 
to_sfixed(1388.0/65536.0,1,-nbitq), 
to_sfixed(-1006.0/65536.0,1,-nbitq), 
to_sfixed(-1258.0/65536.0,1,-nbitq), 
to_sfixed(-2751.0/65536.0,1,-nbitq), 
to_sfixed(-1404.0/65536.0,1,-nbitq), 
to_sfixed(-515.0/65536.0,1,-nbitq), 
to_sfixed(1816.0/65536.0,1,-nbitq), 
to_sfixed(511.0/65536.0,1,-nbitq), 
to_sfixed(187.0/65536.0,1,-nbitq), 
to_sfixed(-2439.0/65536.0,1,-nbitq), 
to_sfixed(118.0/65536.0,1,-nbitq), 
to_sfixed(909.0/65536.0,1,-nbitq), 
to_sfixed(-1095.0/65536.0,1,-nbitq), 
to_sfixed(1425.0/65536.0,1,-nbitq), 
to_sfixed(1611.0/65536.0,1,-nbitq), 
to_sfixed(2969.0/65536.0,1,-nbitq), 
to_sfixed(75.0/65536.0,1,-nbitq), 
to_sfixed(426.0/65536.0,1,-nbitq), 
to_sfixed(-1185.0/65536.0,1,-nbitq), 
to_sfixed(127.0/65536.0,1,-nbitq), 
to_sfixed(2895.0/65536.0,1,-nbitq), 
to_sfixed(771.0/65536.0,1,-nbitq), 
to_sfixed(5522.0/65536.0,1,-nbitq), 
to_sfixed(296.0/65536.0,1,-nbitq), 
to_sfixed(1491.0/65536.0,1,-nbitq), 
to_sfixed(-407.0/65536.0,1,-nbitq), 
to_sfixed(-1310.0/65536.0,1,-nbitq), 
to_sfixed(-579.0/65536.0,1,-nbitq), 
to_sfixed(2402.0/65536.0,1,-nbitq), 
to_sfixed(424.0/65536.0,1,-nbitq), 
to_sfixed(-3064.0/65536.0,1,-nbitq), 
to_sfixed(641.0/65536.0,1,-nbitq), 
to_sfixed(-1320.0/65536.0,1,-nbitq), 
to_sfixed(-349.0/65536.0,1,-nbitq), 
to_sfixed(1591.0/65536.0,1,-nbitq), 
to_sfixed(818.0/65536.0,1,-nbitq), 
to_sfixed(390.0/65536.0,1,-nbitq), 
to_sfixed(-1971.0/65536.0,1,-nbitq), 
to_sfixed(-1773.0/65536.0,1,-nbitq), 
to_sfixed(559.0/65536.0,1,-nbitq), 
to_sfixed(-1004.0/65536.0,1,-nbitq), 
to_sfixed(-600.0/65536.0,1,-nbitq), 
to_sfixed(2010.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-189.0/65536.0,1,-nbitq), 
to_sfixed(-2247.0/65536.0,1,-nbitq), 
to_sfixed(3861.0/65536.0,1,-nbitq), 
to_sfixed(-2298.0/65536.0,1,-nbitq), 
to_sfixed(-577.0/65536.0,1,-nbitq), 
to_sfixed(-4325.0/65536.0,1,-nbitq), 
to_sfixed(-964.0/65536.0,1,-nbitq), 
to_sfixed(-1793.0/65536.0,1,-nbitq), 
to_sfixed(-463.0/65536.0,1,-nbitq), 
to_sfixed(4.0/65536.0,1,-nbitq), 
to_sfixed(-865.0/65536.0,1,-nbitq), 
to_sfixed(2748.0/65536.0,1,-nbitq), 
to_sfixed(1449.0/65536.0,1,-nbitq), 
to_sfixed(-2099.0/65536.0,1,-nbitq), 
to_sfixed(730.0/65536.0,1,-nbitq), 
to_sfixed(1555.0/65536.0,1,-nbitq), 
to_sfixed(-2670.0/65536.0,1,-nbitq), 
to_sfixed(-1200.0/65536.0,1,-nbitq), 
to_sfixed(1688.0/65536.0,1,-nbitq), 
to_sfixed(1722.0/65536.0,1,-nbitq), 
to_sfixed(-2579.0/65536.0,1,-nbitq), 
to_sfixed(-1943.0/65536.0,1,-nbitq), 
to_sfixed(1052.0/65536.0,1,-nbitq), 
to_sfixed(1652.0/65536.0,1,-nbitq), 
to_sfixed(-2094.0/65536.0,1,-nbitq), 
to_sfixed(2140.0/65536.0,1,-nbitq), 
to_sfixed(-2351.0/65536.0,1,-nbitq), 
to_sfixed(-2227.0/65536.0,1,-nbitq), 
to_sfixed(1616.0/65536.0,1,-nbitq), 
to_sfixed(1421.0/65536.0,1,-nbitq), 
to_sfixed(-923.0/65536.0,1,-nbitq), 
to_sfixed(-739.0/65536.0,1,-nbitq), 
to_sfixed(-4691.0/65536.0,1,-nbitq), 
to_sfixed(-517.0/65536.0,1,-nbitq), 
to_sfixed(2542.0/65536.0,1,-nbitq), 
to_sfixed(2421.0/65536.0,1,-nbitq), 
to_sfixed(2215.0/65536.0,1,-nbitq), 
to_sfixed(645.0/65536.0,1,-nbitq), 
to_sfixed(-4392.0/65536.0,1,-nbitq), 
to_sfixed(697.0/65536.0,1,-nbitq), 
to_sfixed(-2732.0/65536.0,1,-nbitq), 
to_sfixed(-3316.0/65536.0,1,-nbitq), 
to_sfixed(-3313.0/65536.0,1,-nbitq), 
to_sfixed(-2041.0/65536.0,1,-nbitq), 
to_sfixed(419.0/65536.0,1,-nbitq), 
to_sfixed(2952.0/65536.0,1,-nbitq), 
to_sfixed(2602.0/65536.0,1,-nbitq), 
to_sfixed(45.0/65536.0,1,-nbitq), 
to_sfixed(884.0/65536.0,1,-nbitq), 
to_sfixed(2226.0/65536.0,1,-nbitq), 
to_sfixed(2944.0/65536.0,1,-nbitq), 
to_sfixed(-2062.0/65536.0,1,-nbitq), 
to_sfixed(-2502.0/65536.0,1,-nbitq), 
to_sfixed(-3253.0/65536.0,1,-nbitq), 
to_sfixed(3385.0/65536.0,1,-nbitq), 
to_sfixed(3107.0/65536.0,1,-nbitq), 
to_sfixed(-1313.0/65536.0,1,-nbitq), 
to_sfixed(3334.0/65536.0,1,-nbitq), 
to_sfixed(1197.0/65536.0,1,-nbitq), 
to_sfixed(5312.0/65536.0,1,-nbitq), 
to_sfixed(-2280.0/65536.0,1,-nbitq), 
to_sfixed(590.0/65536.0,1,-nbitq), 
to_sfixed(851.0/65536.0,1,-nbitq), 
to_sfixed(124.0/65536.0,1,-nbitq), 
to_sfixed(3024.0/65536.0,1,-nbitq), 
to_sfixed(838.0/65536.0,1,-nbitq), 
to_sfixed(543.0/65536.0,1,-nbitq), 
to_sfixed(834.0/65536.0,1,-nbitq), 
to_sfixed(552.0/65536.0,1,-nbitq), 
to_sfixed(-2272.0/65536.0,1,-nbitq), 
to_sfixed(-170.0/65536.0,1,-nbitq), 
to_sfixed(564.0/65536.0,1,-nbitq), 
to_sfixed(2693.0/65536.0,1,-nbitq), 
to_sfixed(571.0/65536.0,1,-nbitq), 
to_sfixed(-1448.0/65536.0,1,-nbitq), 
to_sfixed(-360.0/65536.0,1,-nbitq), 
to_sfixed(1195.0/65536.0,1,-nbitq), 
to_sfixed(-1286.0/65536.0,1,-nbitq), 
to_sfixed(-2330.0/65536.0,1,-nbitq), 
to_sfixed(3920.0/65536.0,1,-nbitq)  ), 
( to_sfixed(195.0/65536.0,1,-nbitq), 
to_sfixed(-951.0/65536.0,1,-nbitq), 
to_sfixed(1648.0/65536.0,1,-nbitq), 
to_sfixed(-1648.0/65536.0,1,-nbitq), 
to_sfixed(1138.0/65536.0,1,-nbitq), 
to_sfixed(426.0/65536.0,1,-nbitq), 
to_sfixed(1929.0/65536.0,1,-nbitq), 
to_sfixed(1249.0/65536.0,1,-nbitq), 
to_sfixed(-1730.0/65536.0,1,-nbitq), 
to_sfixed(-1728.0/65536.0,1,-nbitq), 
to_sfixed(622.0/65536.0,1,-nbitq), 
to_sfixed(904.0/65536.0,1,-nbitq), 
to_sfixed(-650.0/65536.0,1,-nbitq), 
to_sfixed(370.0/65536.0,1,-nbitq), 
to_sfixed(3064.0/65536.0,1,-nbitq), 
to_sfixed(1438.0/65536.0,1,-nbitq), 
to_sfixed(-2850.0/65536.0,1,-nbitq), 
to_sfixed(1681.0/65536.0,1,-nbitq), 
to_sfixed(3974.0/65536.0,1,-nbitq), 
to_sfixed(3201.0/65536.0,1,-nbitq), 
to_sfixed(1104.0/65536.0,1,-nbitq), 
to_sfixed(3634.0/65536.0,1,-nbitq), 
to_sfixed(-684.0/65536.0,1,-nbitq), 
to_sfixed(-256.0/65536.0,1,-nbitq), 
to_sfixed(-1221.0/65536.0,1,-nbitq), 
to_sfixed(-1714.0/65536.0,1,-nbitq), 
to_sfixed(-2455.0/65536.0,1,-nbitq), 
to_sfixed(-2280.0/65536.0,1,-nbitq), 
to_sfixed(-2028.0/65536.0,1,-nbitq), 
to_sfixed(2748.0/65536.0,1,-nbitq), 
to_sfixed(955.0/65536.0,1,-nbitq), 
to_sfixed(-3417.0/65536.0,1,-nbitq), 
to_sfixed(-3309.0/65536.0,1,-nbitq), 
to_sfixed(-466.0/65536.0,1,-nbitq), 
to_sfixed(2420.0/65536.0,1,-nbitq), 
to_sfixed(2729.0/65536.0,1,-nbitq), 
to_sfixed(-214.0/65536.0,1,-nbitq), 
to_sfixed(-3565.0/65536.0,1,-nbitq), 
to_sfixed(1608.0/65536.0,1,-nbitq), 
to_sfixed(-26.0/65536.0,1,-nbitq), 
to_sfixed(-4168.0/65536.0,1,-nbitq), 
to_sfixed(-543.0/65536.0,1,-nbitq), 
to_sfixed(-4921.0/65536.0,1,-nbitq), 
to_sfixed(-1146.0/65536.0,1,-nbitq), 
to_sfixed(2601.0/65536.0,1,-nbitq), 
to_sfixed(903.0/65536.0,1,-nbitq), 
to_sfixed(-2547.0/65536.0,1,-nbitq), 
to_sfixed(-172.0/65536.0,1,-nbitq), 
to_sfixed(-2124.0/65536.0,1,-nbitq), 
to_sfixed(835.0/65536.0,1,-nbitq), 
to_sfixed(-608.0/65536.0,1,-nbitq), 
to_sfixed(-3098.0/65536.0,1,-nbitq), 
to_sfixed(2317.0/65536.0,1,-nbitq), 
to_sfixed(1829.0/65536.0,1,-nbitq), 
to_sfixed(1869.0/65536.0,1,-nbitq), 
to_sfixed(1485.0/65536.0,1,-nbitq), 
to_sfixed(-2442.0/65536.0,1,-nbitq), 
to_sfixed(2214.0/65536.0,1,-nbitq), 
to_sfixed(2922.0/65536.0,1,-nbitq), 
to_sfixed(397.0/65536.0,1,-nbitq), 
to_sfixed(-3288.0/65536.0,1,-nbitq), 
to_sfixed(280.0/65536.0,1,-nbitq), 
to_sfixed(2926.0/65536.0,1,-nbitq), 
to_sfixed(2545.0/65536.0,1,-nbitq), 
to_sfixed(-1532.0/65536.0,1,-nbitq), 
to_sfixed(-611.0/65536.0,1,-nbitq), 
to_sfixed(317.0/65536.0,1,-nbitq), 
to_sfixed(728.0/65536.0,1,-nbitq), 
to_sfixed(929.0/65536.0,1,-nbitq), 
to_sfixed(3883.0/65536.0,1,-nbitq), 
to_sfixed(-2584.0/65536.0,1,-nbitq), 
to_sfixed(-2615.0/65536.0,1,-nbitq), 
to_sfixed(-1466.0/65536.0,1,-nbitq), 
to_sfixed(-2501.0/65536.0,1,-nbitq), 
to_sfixed(-2125.0/65536.0,1,-nbitq), 
to_sfixed(404.0/65536.0,1,-nbitq), 
to_sfixed(929.0/65536.0,1,-nbitq), 
to_sfixed(3542.0/65536.0,1,-nbitq), 
to_sfixed(1863.0/65536.0,1,-nbitq), 
to_sfixed(26.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2013.0/65536.0,1,-nbitq), 
to_sfixed(1934.0/65536.0,1,-nbitq), 
to_sfixed(1132.0/65536.0,1,-nbitq), 
to_sfixed(441.0/65536.0,1,-nbitq), 
to_sfixed(-1002.0/65536.0,1,-nbitq), 
to_sfixed(-2174.0/65536.0,1,-nbitq), 
to_sfixed(691.0/65536.0,1,-nbitq), 
to_sfixed(-568.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(2484.0/65536.0,1,-nbitq), 
to_sfixed(-2023.0/65536.0,1,-nbitq), 
to_sfixed(5636.0/65536.0,1,-nbitq), 
to_sfixed(1924.0/65536.0,1,-nbitq), 
to_sfixed(3077.0/65536.0,1,-nbitq), 
to_sfixed(590.0/65536.0,1,-nbitq), 
to_sfixed(1729.0/65536.0,1,-nbitq), 
to_sfixed(-2847.0/65536.0,1,-nbitq), 
to_sfixed(-650.0/65536.0,1,-nbitq), 
to_sfixed(2398.0/65536.0,1,-nbitq), 
to_sfixed(-352.0/65536.0,1,-nbitq), 
to_sfixed(-3668.0/65536.0,1,-nbitq), 
to_sfixed(585.0/65536.0,1,-nbitq), 
to_sfixed(2755.0/65536.0,1,-nbitq), 
to_sfixed(-705.0/65536.0,1,-nbitq), 
to_sfixed(-4363.0/65536.0,1,-nbitq), 
to_sfixed(-2087.0/65536.0,1,-nbitq), 
to_sfixed(-1334.0/65536.0,1,-nbitq), 
to_sfixed(1539.0/65536.0,1,-nbitq), 
to_sfixed(-3614.0/65536.0,1,-nbitq), 
to_sfixed(491.0/65536.0,1,-nbitq), 
to_sfixed(-3135.0/65536.0,1,-nbitq), 
to_sfixed(833.0/65536.0,1,-nbitq), 
to_sfixed(-5618.0/65536.0,1,-nbitq), 
to_sfixed(-3995.0/65536.0,1,-nbitq), 
to_sfixed(1006.0/65536.0,1,-nbitq), 
to_sfixed(-339.0/65536.0,1,-nbitq), 
to_sfixed(3964.0/65536.0,1,-nbitq), 
to_sfixed(-2531.0/65536.0,1,-nbitq), 
to_sfixed(2476.0/65536.0,1,-nbitq), 
to_sfixed(-1301.0/65536.0,1,-nbitq), 
to_sfixed(-513.0/65536.0,1,-nbitq), 
to_sfixed(-1618.0/65536.0,1,-nbitq), 
to_sfixed(-2699.0/65536.0,1,-nbitq), 
to_sfixed(-535.0/65536.0,1,-nbitq), 
to_sfixed(2604.0/65536.0,1,-nbitq), 
to_sfixed(1942.0/65536.0,1,-nbitq), 
to_sfixed(-1839.0/65536.0,1,-nbitq), 
to_sfixed(-781.0/65536.0,1,-nbitq), 
to_sfixed(834.0/65536.0,1,-nbitq), 
to_sfixed(2651.0/65536.0,1,-nbitq), 
to_sfixed(803.0/65536.0,1,-nbitq), 
to_sfixed(-793.0/65536.0,1,-nbitq), 
to_sfixed(-2977.0/65536.0,1,-nbitq), 
to_sfixed(2264.0/65536.0,1,-nbitq), 
to_sfixed(2659.0/65536.0,1,-nbitq), 
to_sfixed(-56.0/65536.0,1,-nbitq), 
to_sfixed(1829.0/65536.0,1,-nbitq), 
to_sfixed(3510.0/65536.0,1,-nbitq), 
to_sfixed(2318.0/65536.0,1,-nbitq), 
to_sfixed(-471.0/65536.0,1,-nbitq), 
to_sfixed(2515.0/65536.0,1,-nbitq), 
to_sfixed(-1234.0/65536.0,1,-nbitq), 
to_sfixed(2057.0/65536.0,1,-nbitq), 
to_sfixed(1039.0/65536.0,1,-nbitq), 
to_sfixed(2597.0/65536.0,1,-nbitq), 
to_sfixed(-2509.0/65536.0,1,-nbitq), 
to_sfixed(1339.0/65536.0,1,-nbitq), 
to_sfixed(-2328.0/65536.0,1,-nbitq), 
to_sfixed(2434.0/65536.0,1,-nbitq), 
to_sfixed(778.0/65536.0,1,-nbitq), 
to_sfixed(2455.0/65536.0,1,-nbitq), 
to_sfixed(-3543.0/65536.0,1,-nbitq), 
to_sfixed(689.0/65536.0,1,-nbitq), 
to_sfixed(138.0/65536.0,1,-nbitq), 
to_sfixed(30.0/65536.0,1,-nbitq), 
to_sfixed(1318.0/65536.0,1,-nbitq), 
to_sfixed(3746.0/65536.0,1,-nbitq), 
to_sfixed(3069.0/65536.0,1,-nbitq), 
to_sfixed(2018.0/65536.0,1,-nbitq), 
to_sfixed(-104.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-888.0/65536.0,1,-nbitq), 
to_sfixed(3342.0/65536.0,1,-nbitq), 
to_sfixed(-6127.0/65536.0,1,-nbitq), 
to_sfixed(-173.0/65536.0,1,-nbitq), 
to_sfixed(-1494.0/65536.0,1,-nbitq), 
to_sfixed(-4820.0/65536.0,1,-nbitq), 
to_sfixed(-647.0/65536.0,1,-nbitq), 
to_sfixed(-753.0/65536.0,1,-nbitq), 
to_sfixed(125.0/65536.0,1,-nbitq), 
to_sfixed(1125.0/65536.0,1,-nbitq), 
to_sfixed(-4998.0/65536.0,1,-nbitq), 
to_sfixed(4244.0/65536.0,1,-nbitq), 
to_sfixed(317.0/65536.0,1,-nbitq), 
to_sfixed(-1440.0/65536.0,1,-nbitq), 
to_sfixed(1913.0/65536.0,1,-nbitq), 
to_sfixed(-1732.0/65536.0,1,-nbitq), 
to_sfixed(-634.0/65536.0,1,-nbitq), 
to_sfixed(2921.0/65536.0,1,-nbitq), 
to_sfixed(-1673.0/65536.0,1,-nbitq), 
to_sfixed(2007.0/65536.0,1,-nbitq), 
to_sfixed(166.0/65536.0,1,-nbitq), 
to_sfixed(-468.0/65536.0,1,-nbitq), 
to_sfixed(8396.0/65536.0,1,-nbitq), 
to_sfixed(3354.0/65536.0,1,-nbitq), 
to_sfixed(-1021.0/65536.0,1,-nbitq), 
to_sfixed(-1967.0/65536.0,1,-nbitq), 
to_sfixed(-2752.0/65536.0,1,-nbitq), 
to_sfixed(-2623.0/65536.0,1,-nbitq), 
to_sfixed(-3082.0/65536.0,1,-nbitq), 
to_sfixed(2412.0/65536.0,1,-nbitq), 
to_sfixed(-3522.0/65536.0,1,-nbitq), 
to_sfixed(443.0/65536.0,1,-nbitq), 
to_sfixed(-1592.0/65536.0,1,-nbitq), 
to_sfixed(-2440.0/65536.0,1,-nbitq), 
to_sfixed(-1809.0/65536.0,1,-nbitq), 
to_sfixed(-547.0/65536.0,1,-nbitq), 
to_sfixed(2464.0/65536.0,1,-nbitq), 
to_sfixed(12.0/65536.0,1,-nbitq), 
to_sfixed(6029.0/65536.0,1,-nbitq), 
to_sfixed(156.0/65536.0,1,-nbitq), 
to_sfixed(-1105.0/65536.0,1,-nbitq), 
to_sfixed(-3230.0/65536.0,1,-nbitq), 
to_sfixed(422.0/65536.0,1,-nbitq), 
to_sfixed(-4562.0/65536.0,1,-nbitq), 
to_sfixed(-1469.0/65536.0,1,-nbitq), 
to_sfixed(3668.0/65536.0,1,-nbitq), 
to_sfixed(-2320.0/65536.0,1,-nbitq), 
to_sfixed(-1116.0/65536.0,1,-nbitq), 
to_sfixed(1267.0/65536.0,1,-nbitq), 
to_sfixed(3436.0/65536.0,1,-nbitq), 
to_sfixed(-1966.0/65536.0,1,-nbitq), 
to_sfixed(-2763.0/65536.0,1,-nbitq), 
to_sfixed(1835.0/65536.0,1,-nbitq), 
to_sfixed(4105.0/65536.0,1,-nbitq), 
to_sfixed(2929.0/65536.0,1,-nbitq), 
to_sfixed(-4857.0/65536.0,1,-nbitq), 
to_sfixed(-1691.0/65536.0,1,-nbitq), 
to_sfixed(-479.0/65536.0,1,-nbitq), 
to_sfixed(1698.0/65536.0,1,-nbitq), 
to_sfixed(272.0/65536.0,1,-nbitq), 
to_sfixed(-2613.0/65536.0,1,-nbitq), 
to_sfixed(-633.0/65536.0,1,-nbitq), 
to_sfixed(1885.0/65536.0,1,-nbitq), 
to_sfixed(-2679.0/65536.0,1,-nbitq), 
to_sfixed(939.0/65536.0,1,-nbitq), 
to_sfixed(190.0/65536.0,1,-nbitq), 
to_sfixed(2406.0/65536.0,1,-nbitq), 
to_sfixed(-1491.0/65536.0,1,-nbitq), 
to_sfixed(-874.0/65536.0,1,-nbitq), 
to_sfixed(777.0/65536.0,1,-nbitq), 
to_sfixed(-2341.0/65536.0,1,-nbitq), 
to_sfixed(-2101.0/65536.0,1,-nbitq), 
to_sfixed(-221.0/65536.0,1,-nbitq), 
to_sfixed(632.0/65536.0,1,-nbitq), 
to_sfixed(-2376.0/65536.0,1,-nbitq), 
to_sfixed(1323.0/65536.0,1,-nbitq), 
to_sfixed(5278.0/65536.0,1,-nbitq), 
to_sfixed(-166.0/65536.0,1,-nbitq), 
to_sfixed(-2510.0/65536.0,1,-nbitq), 
to_sfixed(-197.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3401.0/65536.0,1,-nbitq), 
to_sfixed(3162.0/65536.0,1,-nbitq), 
to_sfixed(-4896.0/65536.0,1,-nbitq), 
to_sfixed(-2468.0/65536.0,1,-nbitq), 
to_sfixed(-1879.0/65536.0,1,-nbitq), 
to_sfixed(-633.0/65536.0,1,-nbitq), 
to_sfixed(4547.0/65536.0,1,-nbitq), 
to_sfixed(1036.0/65536.0,1,-nbitq), 
to_sfixed(-1200.0/65536.0,1,-nbitq), 
to_sfixed(1835.0/65536.0,1,-nbitq), 
to_sfixed(2146.0/65536.0,1,-nbitq), 
to_sfixed(4520.0/65536.0,1,-nbitq), 
to_sfixed(-1733.0/65536.0,1,-nbitq), 
to_sfixed(-2948.0/65536.0,1,-nbitq), 
to_sfixed(-4191.0/65536.0,1,-nbitq), 
to_sfixed(-1155.0/65536.0,1,-nbitq), 
to_sfixed(-1735.0/65536.0,1,-nbitq), 
to_sfixed(-537.0/65536.0,1,-nbitq), 
to_sfixed(-2336.0/65536.0,1,-nbitq), 
to_sfixed(-1278.0/65536.0,1,-nbitq), 
to_sfixed(750.0/65536.0,1,-nbitq), 
to_sfixed(4874.0/65536.0,1,-nbitq), 
to_sfixed(5629.0/65536.0,1,-nbitq), 
to_sfixed(-1658.0/65536.0,1,-nbitq), 
to_sfixed(1811.0/65536.0,1,-nbitq), 
to_sfixed(-4477.0/65536.0,1,-nbitq), 
to_sfixed(-2680.0/65536.0,1,-nbitq), 
to_sfixed(-468.0/65536.0,1,-nbitq), 
to_sfixed(-5101.0/65536.0,1,-nbitq), 
to_sfixed(-1499.0/65536.0,1,-nbitq), 
to_sfixed(1907.0/65536.0,1,-nbitq), 
to_sfixed(-2717.0/65536.0,1,-nbitq), 
to_sfixed(-4237.0/65536.0,1,-nbitq), 
to_sfixed(-4289.0/65536.0,1,-nbitq), 
to_sfixed(-2701.0/65536.0,1,-nbitq), 
to_sfixed(2960.0/65536.0,1,-nbitq), 
to_sfixed(2085.0/65536.0,1,-nbitq), 
to_sfixed(-1078.0/65536.0,1,-nbitq), 
to_sfixed(5194.0/65536.0,1,-nbitq), 
to_sfixed(980.0/65536.0,1,-nbitq), 
to_sfixed(-2060.0/65536.0,1,-nbitq), 
to_sfixed(1084.0/65536.0,1,-nbitq), 
to_sfixed(-218.0/65536.0,1,-nbitq), 
to_sfixed(1661.0/65536.0,1,-nbitq), 
to_sfixed(-719.0/65536.0,1,-nbitq), 
to_sfixed(3356.0/65536.0,1,-nbitq), 
to_sfixed(-3142.0/65536.0,1,-nbitq), 
to_sfixed(-2738.0/65536.0,1,-nbitq), 
to_sfixed(224.0/65536.0,1,-nbitq), 
to_sfixed(191.0/65536.0,1,-nbitq), 
to_sfixed(63.0/65536.0,1,-nbitq), 
to_sfixed(-4786.0/65536.0,1,-nbitq), 
to_sfixed(1201.0/65536.0,1,-nbitq), 
to_sfixed(1250.0/65536.0,1,-nbitq), 
to_sfixed(5028.0/65536.0,1,-nbitq), 
to_sfixed(-4052.0/65536.0,1,-nbitq), 
to_sfixed(-108.0/65536.0,1,-nbitq), 
to_sfixed(4118.0/65536.0,1,-nbitq), 
to_sfixed(3493.0/65536.0,1,-nbitq), 
to_sfixed(-4410.0/65536.0,1,-nbitq), 
to_sfixed(1111.0/65536.0,1,-nbitq), 
to_sfixed(2727.0/65536.0,1,-nbitq), 
to_sfixed(1911.0/65536.0,1,-nbitq), 
to_sfixed(1668.0/65536.0,1,-nbitq), 
to_sfixed(1426.0/65536.0,1,-nbitq), 
to_sfixed(-1878.0/65536.0,1,-nbitq), 
to_sfixed(5625.0/65536.0,1,-nbitq), 
to_sfixed(3637.0/65536.0,1,-nbitq), 
to_sfixed(4902.0/65536.0,1,-nbitq), 
to_sfixed(7146.0/65536.0,1,-nbitq), 
to_sfixed(2146.0/65536.0,1,-nbitq), 
to_sfixed(1223.0/65536.0,1,-nbitq), 
to_sfixed(-1341.0/65536.0,1,-nbitq), 
to_sfixed(348.0/65536.0,1,-nbitq), 
to_sfixed(-1985.0/65536.0,1,-nbitq), 
to_sfixed(677.0/65536.0,1,-nbitq), 
to_sfixed(130.0/65536.0,1,-nbitq), 
to_sfixed(3794.0/65536.0,1,-nbitq), 
to_sfixed(1365.0/65536.0,1,-nbitq), 
to_sfixed(1415.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3058.0/65536.0,1,-nbitq), 
to_sfixed(199.0/65536.0,1,-nbitq), 
to_sfixed(-9285.0/65536.0,1,-nbitq), 
to_sfixed(-3520.0/65536.0,1,-nbitq), 
to_sfixed(314.0/65536.0,1,-nbitq), 
to_sfixed(-591.0/65536.0,1,-nbitq), 
to_sfixed(5031.0/65536.0,1,-nbitq), 
to_sfixed(2472.0/65536.0,1,-nbitq), 
to_sfixed(-730.0/65536.0,1,-nbitq), 
to_sfixed(2639.0/65536.0,1,-nbitq), 
to_sfixed(233.0/65536.0,1,-nbitq), 
to_sfixed(3638.0/65536.0,1,-nbitq), 
to_sfixed(1892.0/65536.0,1,-nbitq), 
to_sfixed(-6165.0/65536.0,1,-nbitq), 
to_sfixed(528.0/65536.0,1,-nbitq), 
to_sfixed(-1923.0/65536.0,1,-nbitq), 
to_sfixed(661.0/65536.0,1,-nbitq), 
to_sfixed(761.0/65536.0,1,-nbitq), 
to_sfixed(-3602.0/65536.0,1,-nbitq), 
to_sfixed(2908.0/65536.0,1,-nbitq), 
to_sfixed(4053.0/65536.0,1,-nbitq), 
to_sfixed(1286.0/65536.0,1,-nbitq), 
to_sfixed(3122.0/65536.0,1,-nbitq), 
to_sfixed(-2738.0/65536.0,1,-nbitq), 
to_sfixed(2024.0/65536.0,1,-nbitq), 
to_sfixed(-2021.0/65536.0,1,-nbitq), 
to_sfixed(-4602.0/65536.0,1,-nbitq), 
to_sfixed(1487.0/65536.0,1,-nbitq), 
to_sfixed(-5959.0/65536.0,1,-nbitq), 
to_sfixed(-2939.0/65536.0,1,-nbitq), 
to_sfixed(-74.0/65536.0,1,-nbitq), 
to_sfixed(-2228.0/65536.0,1,-nbitq), 
to_sfixed(-1124.0/65536.0,1,-nbitq), 
to_sfixed(917.0/65536.0,1,-nbitq), 
to_sfixed(-1575.0/65536.0,1,-nbitq), 
to_sfixed(1998.0/65536.0,1,-nbitq), 
to_sfixed(-774.0/65536.0,1,-nbitq), 
to_sfixed(2644.0/65536.0,1,-nbitq), 
to_sfixed(10699.0/65536.0,1,-nbitq), 
to_sfixed(1476.0/65536.0,1,-nbitq), 
to_sfixed(-2570.0/65536.0,1,-nbitq), 
to_sfixed(-1077.0/65536.0,1,-nbitq), 
to_sfixed(9.0/65536.0,1,-nbitq), 
to_sfixed(-1668.0/65536.0,1,-nbitq), 
to_sfixed(-343.0/65536.0,1,-nbitq), 
to_sfixed(973.0/65536.0,1,-nbitq), 
to_sfixed(-4356.0/65536.0,1,-nbitq), 
to_sfixed(-6840.0/65536.0,1,-nbitq), 
to_sfixed(993.0/65536.0,1,-nbitq), 
to_sfixed(3149.0/65536.0,1,-nbitq), 
to_sfixed(510.0/65536.0,1,-nbitq), 
to_sfixed(-4720.0/65536.0,1,-nbitq), 
to_sfixed(-1294.0/65536.0,1,-nbitq), 
to_sfixed(-2210.0/65536.0,1,-nbitq), 
to_sfixed(1554.0/65536.0,1,-nbitq), 
to_sfixed(-4873.0/65536.0,1,-nbitq), 
to_sfixed(-1541.0/65536.0,1,-nbitq), 
to_sfixed(3849.0/65536.0,1,-nbitq), 
to_sfixed(-1426.0/65536.0,1,-nbitq), 
to_sfixed(-6831.0/65536.0,1,-nbitq), 
to_sfixed(-2112.0/65536.0,1,-nbitq), 
to_sfixed(227.0/65536.0,1,-nbitq), 
to_sfixed(-1021.0/65536.0,1,-nbitq), 
to_sfixed(-442.0/65536.0,1,-nbitq), 
to_sfixed(1508.0/65536.0,1,-nbitq), 
to_sfixed(-6697.0/65536.0,1,-nbitq), 
to_sfixed(4876.0/65536.0,1,-nbitq), 
to_sfixed(2304.0/65536.0,1,-nbitq), 
to_sfixed(2990.0/65536.0,1,-nbitq), 
to_sfixed(9937.0/65536.0,1,-nbitq), 
to_sfixed(1730.0/65536.0,1,-nbitq), 
to_sfixed(-3537.0/65536.0,1,-nbitq), 
to_sfixed(-3078.0/65536.0,1,-nbitq), 
to_sfixed(2150.0/65536.0,1,-nbitq), 
to_sfixed(-1663.0/65536.0,1,-nbitq), 
to_sfixed(1295.0/65536.0,1,-nbitq), 
to_sfixed(125.0/65536.0,1,-nbitq), 
to_sfixed(1645.0/65536.0,1,-nbitq), 
to_sfixed(-2551.0/65536.0,1,-nbitq), 
to_sfixed(-60.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-615.0/65536.0,1,-nbitq), 
to_sfixed(2572.0/65536.0,1,-nbitq), 
to_sfixed(-6189.0/65536.0,1,-nbitq), 
to_sfixed(-4960.0/65536.0,1,-nbitq), 
to_sfixed(-476.0/65536.0,1,-nbitq), 
to_sfixed(588.0/65536.0,1,-nbitq), 
to_sfixed(2422.0/65536.0,1,-nbitq), 
to_sfixed(271.0/65536.0,1,-nbitq), 
to_sfixed(-15.0/65536.0,1,-nbitq), 
to_sfixed(-1793.0/65536.0,1,-nbitq), 
to_sfixed(-873.0/65536.0,1,-nbitq), 
to_sfixed(5086.0/65536.0,1,-nbitq), 
to_sfixed(1503.0/65536.0,1,-nbitq), 
to_sfixed(-5736.0/65536.0,1,-nbitq), 
to_sfixed(-4848.0/65536.0,1,-nbitq), 
to_sfixed(961.0/65536.0,1,-nbitq), 
to_sfixed(1593.0/65536.0,1,-nbitq), 
to_sfixed(-475.0/65536.0,1,-nbitq), 
to_sfixed(-844.0/65536.0,1,-nbitq), 
to_sfixed(2738.0/65536.0,1,-nbitq), 
to_sfixed(2337.0/65536.0,1,-nbitq), 
to_sfixed(2691.0/65536.0,1,-nbitq), 
to_sfixed(3395.0/65536.0,1,-nbitq), 
to_sfixed(-2572.0/65536.0,1,-nbitq), 
to_sfixed(4210.0/65536.0,1,-nbitq), 
to_sfixed(-5277.0/65536.0,1,-nbitq), 
to_sfixed(-477.0/65536.0,1,-nbitq), 
to_sfixed(2230.0/65536.0,1,-nbitq), 
to_sfixed(-1191.0/65536.0,1,-nbitq), 
to_sfixed(562.0/65536.0,1,-nbitq), 
to_sfixed(2741.0/65536.0,1,-nbitq), 
to_sfixed(-7158.0/65536.0,1,-nbitq), 
to_sfixed(784.0/65536.0,1,-nbitq), 
to_sfixed(-178.0/65536.0,1,-nbitq), 
to_sfixed(-290.0/65536.0,1,-nbitq), 
to_sfixed(1346.0/65536.0,1,-nbitq), 
to_sfixed(-561.0/65536.0,1,-nbitq), 
to_sfixed(4699.0/65536.0,1,-nbitq), 
to_sfixed(5210.0/65536.0,1,-nbitq), 
to_sfixed(229.0/65536.0,1,-nbitq), 
to_sfixed(-2717.0/65536.0,1,-nbitq), 
to_sfixed(1606.0/65536.0,1,-nbitq), 
to_sfixed(54.0/65536.0,1,-nbitq), 
to_sfixed(347.0/65536.0,1,-nbitq), 
to_sfixed(152.0/65536.0,1,-nbitq), 
to_sfixed(-1857.0/65536.0,1,-nbitq), 
to_sfixed(481.0/65536.0,1,-nbitq), 
to_sfixed(-5327.0/65536.0,1,-nbitq), 
to_sfixed(-2426.0/65536.0,1,-nbitq), 
to_sfixed(2041.0/65536.0,1,-nbitq), 
to_sfixed(2139.0/65536.0,1,-nbitq), 
to_sfixed(-6199.0/65536.0,1,-nbitq), 
to_sfixed(1553.0/65536.0,1,-nbitq), 
to_sfixed(-873.0/65536.0,1,-nbitq), 
to_sfixed(326.0/65536.0,1,-nbitq), 
to_sfixed(-5559.0/65536.0,1,-nbitq), 
to_sfixed(3134.0/65536.0,1,-nbitq), 
to_sfixed(3757.0/65536.0,1,-nbitq), 
to_sfixed(-735.0/65536.0,1,-nbitq), 
to_sfixed(-5715.0/65536.0,1,-nbitq), 
to_sfixed(-837.0/65536.0,1,-nbitq), 
to_sfixed(-2477.0/65536.0,1,-nbitq), 
to_sfixed(1576.0/65536.0,1,-nbitq), 
to_sfixed(-3194.0/65536.0,1,-nbitq), 
to_sfixed(3561.0/65536.0,1,-nbitq), 
to_sfixed(-6012.0/65536.0,1,-nbitq), 
to_sfixed(8290.0/65536.0,1,-nbitq), 
to_sfixed(6474.0/65536.0,1,-nbitq), 
to_sfixed(2466.0/65536.0,1,-nbitq), 
to_sfixed(6295.0/65536.0,1,-nbitq), 
to_sfixed(2173.0/65536.0,1,-nbitq), 
to_sfixed(-3288.0/65536.0,1,-nbitq), 
to_sfixed(-4085.0/65536.0,1,-nbitq), 
to_sfixed(-2154.0/65536.0,1,-nbitq), 
to_sfixed(-130.0/65536.0,1,-nbitq), 
to_sfixed(3587.0/65536.0,1,-nbitq), 
to_sfixed(3611.0/65536.0,1,-nbitq), 
to_sfixed(5936.0/65536.0,1,-nbitq), 
to_sfixed(1894.0/65536.0,1,-nbitq), 
to_sfixed(1436.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2217.0/65536.0,1,-nbitq), 
to_sfixed(3533.0/65536.0,1,-nbitq), 
to_sfixed(-8627.0/65536.0,1,-nbitq), 
to_sfixed(-5038.0/65536.0,1,-nbitq), 
to_sfixed(-344.0/65536.0,1,-nbitq), 
to_sfixed(3125.0/65536.0,1,-nbitq), 
to_sfixed(294.0/65536.0,1,-nbitq), 
to_sfixed(1255.0/65536.0,1,-nbitq), 
to_sfixed(3576.0/65536.0,1,-nbitq), 
to_sfixed(2521.0/65536.0,1,-nbitq), 
to_sfixed(895.0/65536.0,1,-nbitq), 
to_sfixed(5045.0/65536.0,1,-nbitq), 
to_sfixed(-2593.0/65536.0,1,-nbitq), 
to_sfixed(-4489.0/65536.0,1,-nbitq), 
to_sfixed(-1242.0/65536.0,1,-nbitq), 
to_sfixed(-126.0/65536.0,1,-nbitq), 
to_sfixed(353.0/65536.0,1,-nbitq), 
to_sfixed(1395.0/65536.0,1,-nbitq), 
to_sfixed(1041.0/65536.0,1,-nbitq), 
to_sfixed(-1754.0/65536.0,1,-nbitq), 
to_sfixed(3850.0/65536.0,1,-nbitq), 
to_sfixed(-918.0/65536.0,1,-nbitq), 
to_sfixed(1861.0/65536.0,1,-nbitq), 
to_sfixed(-1291.0/65536.0,1,-nbitq), 
to_sfixed(3918.0/65536.0,1,-nbitq), 
to_sfixed(660.0/65536.0,1,-nbitq), 
to_sfixed(-4220.0/65536.0,1,-nbitq), 
to_sfixed(2676.0/65536.0,1,-nbitq), 
to_sfixed(2522.0/65536.0,1,-nbitq), 
to_sfixed(-3173.0/65536.0,1,-nbitq), 
to_sfixed(1908.0/65536.0,1,-nbitq), 
to_sfixed(-4375.0/65536.0,1,-nbitq), 
to_sfixed(3140.0/65536.0,1,-nbitq), 
to_sfixed(-2172.0/65536.0,1,-nbitq), 
to_sfixed(-225.0/65536.0,1,-nbitq), 
to_sfixed(1048.0/65536.0,1,-nbitq), 
to_sfixed(4346.0/65536.0,1,-nbitq), 
to_sfixed(1669.0/65536.0,1,-nbitq), 
to_sfixed(3723.0/65536.0,1,-nbitq), 
to_sfixed(-1025.0/65536.0,1,-nbitq), 
to_sfixed(-3562.0/65536.0,1,-nbitq), 
to_sfixed(-2667.0/65536.0,1,-nbitq), 
to_sfixed(6173.0/65536.0,1,-nbitq), 
to_sfixed(-457.0/65536.0,1,-nbitq), 
to_sfixed(3132.0/65536.0,1,-nbitq), 
to_sfixed(969.0/65536.0,1,-nbitq), 
to_sfixed(-2691.0/65536.0,1,-nbitq), 
to_sfixed(-10434.0/65536.0,1,-nbitq), 
to_sfixed(1838.0/65536.0,1,-nbitq), 
to_sfixed(619.0/65536.0,1,-nbitq), 
to_sfixed(-2537.0/65536.0,1,-nbitq), 
to_sfixed(119.0/65536.0,1,-nbitq), 
to_sfixed(-2123.0/65536.0,1,-nbitq), 
to_sfixed(-4566.0/65536.0,1,-nbitq), 
to_sfixed(-1522.0/65536.0,1,-nbitq), 
to_sfixed(-5967.0/65536.0,1,-nbitq), 
to_sfixed(1562.0/65536.0,1,-nbitq), 
to_sfixed(2090.0/65536.0,1,-nbitq), 
to_sfixed(-1803.0/65536.0,1,-nbitq), 
to_sfixed(-6996.0/65536.0,1,-nbitq), 
to_sfixed(-3801.0/65536.0,1,-nbitq), 
to_sfixed(-1714.0/65536.0,1,-nbitq), 
to_sfixed(-548.0/65536.0,1,-nbitq), 
to_sfixed(1764.0/65536.0,1,-nbitq), 
to_sfixed(2576.0/65536.0,1,-nbitq), 
to_sfixed(-4619.0/65536.0,1,-nbitq), 
to_sfixed(7451.0/65536.0,1,-nbitq), 
to_sfixed(5959.0/65536.0,1,-nbitq), 
to_sfixed(-926.0/65536.0,1,-nbitq), 
to_sfixed(10441.0/65536.0,1,-nbitq), 
to_sfixed(-436.0/65536.0,1,-nbitq), 
to_sfixed(-3521.0/65536.0,1,-nbitq), 
to_sfixed(-5318.0/65536.0,1,-nbitq), 
to_sfixed(-1646.0/65536.0,1,-nbitq), 
to_sfixed(629.0/65536.0,1,-nbitq), 
to_sfixed(4346.0/65536.0,1,-nbitq), 
to_sfixed(1062.0/65536.0,1,-nbitq), 
to_sfixed(3644.0/65536.0,1,-nbitq), 
to_sfixed(1063.0/65536.0,1,-nbitq), 
to_sfixed(243.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1436.0/65536.0,1,-nbitq), 
to_sfixed(1871.0/65536.0,1,-nbitq), 
to_sfixed(-7207.0/65536.0,1,-nbitq), 
to_sfixed(-953.0/65536.0,1,-nbitq), 
to_sfixed(4002.0/65536.0,1,-nbitq), 
to_sfixed(3234.0/65536.0,1,-nbitq), 
to_sfixed(2788.0/65536.0,1,-nbitq), 
to_sfixed(299.0/65536.0,1,-nbitq), 
to_sfixed(2164.0/65536.0,1,-nbitq), 
to_sfixed(-2425.0/65536.0,1,-nbitq), 
to_sfixed(1426.0/65536.0,1,-nbitq), 
to_sfixed(9751.0/65536.0,1,-nbitq), 
to_sfixed(-53.0/65536.0,1,-nbitq), 
to_sfixed(-6226.0/65536.0,1,-nbitq), 
to_sfixed(-2804.0/65536.0,1,-nbitq), 
to_sfixed(-428.0/65536.0,1,-nbitq), 
to_sfixed(-1899.0/65536.0,1,-nbitq), 
to_sfixed(521.0/65536.0,1,-nbitq), 
to_sfixed(-2314.0/65536.0,1,-nbitq), 
to_sfixed(1714.0/65536.0,1,-nbitq), 
to_sfixed(5616.0/65536.0,1,-nbitq), 
to_sfixed(-42.0/65536.0,1,-nbitq), 
to_sfixed(2875.0/65536.0,1,-nbitq), 
to_sfixed(-1036.0/65536.0,1,-nbitq), 
to_sfixed(4033.0/65536.0,1,-nbitq), 
to_sfixed(-2211.0/65536.0,1,-nbitq), 
to_sfixed(-2064.0/65536.0,1,-nbitq), 
to_sfixed(542.0/65536.0,1,-nbitq), 
to_sfixed(959.0/65536.0,1,-nbitq), 
to_sfixed(-706.0/65536.0,1,-nbitq), 
to_sfixed(-1773.0/65536.0,1,-nbitq), 
to_sfixed(-6404.0/65536.0,1,-nbitq), 
to_sfixed(767.0/65536.0,1,-nbitq), 
to_sfixed(-2444.0/65536.0,1,-nbitq), 
to_sfixed(-983.0/65536.0,1,-nbitq), 
to_sfixed(-2632.0/65536.0,1,-nbitq), 
to_sfixed(3614.0/65536.0,1,-nbitq), 
to_sfixed(1871.0/65536.0,1,-nbitq), 
to_sfixed(-322.0/65536.0,1,-nbitq), 
to_sfixed(-1868.0/65536.0,1,-nbitq), 
to_sfixed(-1064.0/65536.0,1,-nbitq), 
to_sfixed(2045.0/65536.0,1,-nbitq), 
to_sfixed(5867.0/65536.0,1,-nbitq), 
to_sfixed(420.0/65536.0,1,-nbitq), 
to_sfixed(-1410.0/65536.0,1,-nbitq), 
to_sfixed(407.0/65536.0,1,-nbitq), 
to_sfixed(-1214.0/65536.0,1,-nbitq), 
to_sfixed(-5287.0/65536.0,1,-nbitq), 
to_sfixed(-1722.0/65536.0,1,-nbitq), 
to_sfixed(-1182.0/65536.0,1,-nbitq), 
to_sfixed(606.0/65536.0,1,-nbitq), 
to_sfixed(1583.0/65536.0,1,-nbitq), 
to_sfixed(-1036.0/65536.0,1,-nbitq), 
to_sfixed(-3197.0/65536.0,1,-nbitq), 
to_sfixed(-2106.0/65536.0,1,-nbitq), 
to_sfixed(-5505.0/65536.0,1,-nbitq), 
to_sfixed(3409.0/65536.0,1,-nbitq), 
to_sfixed(2616.0/65536.0,1,-nbitq), 
to_sfixed(2356.0/65536.0,1,-nbitq), 
to_sfixed(-7188.0/65536.0,1,-nbitq), 
to_sfixed(-2735.0/65536.0,1,-nbitq), 
to_sfixed(1656.0/65536.0,1,-nbitq), 
to_sfixed(-1129.0/65536.0,1,-nbitq), 
to_sfixed(-2180.0/65536.0,1,-nbitq), 
to_sfixed(98.0/65536.0,1,-nbitq), 
to_sfixed(-3744.0/65536.0,1,-nbitq), 
to_sfixed(4350.0/65536.0,1,-nbitq), 
to_sfixed(8077.0/65536.0,1,-nbitq), 
to_sfixed(-707.0/65536.0,1,-nbitq), 
to_sfixed(7561.0/65536.0,1,-nbitq), 
to_sfixed(-2858.0/65536.0,1,-nbitq), 
to_sfixed(-2150.0/65536.0,1,-nbitq), 
to_sfixed(-2774.0/65536.0,1,-nbitq), 
to_sfixed(-1284.0/65536.0,1,-nbitq), 
to_sfixed(-1486.0/65536.0,1,-nbitq), 
to_sfixed(2085.0/65536.0,1,-nbitq), 
to_sfixed(1039.0/65536.0,1,-nbitq), 
to_sfixed(6872.0/65536.0,1,-nbitq), 
to_sfixed(-1622.0/65536.0,1,-nbitq), 
to_sfixed(3602.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1751.0/65536.0,1,-nbitq), 
to_sfixed(2193.0/65536.0,1,-nbitq), 
to_sfixed(-2787.0/65536.0,1,-nbitq), 
to_sfixed(-1370.0/65536.0,1,-nbitq), 
to_sfixed(4510.0/65536.0,1,-nbitq), 
to_sfixed(1836.0/65536.0,1,-nbitq), 
to_sfixed(404.0/65536.0,1,-nbitq), 
to_sfixed(896.0/65536.0,1,-nbitq), 
to_sfixed(2448.0/65536.0,1,-nbitq), 
to_sfixed(451.0/65536.0,1,-nbitq), 
to_sfixed(3712.0/65536.0,1,-nbitq), 
to_sfixed(3450.0/65536.0,1,-nbitq), 
to_sfixed(2072.0/65536.0,1,-nbitq), 
to_sfixed(-1547.0/65536.0,1,-nbitq), 
to_sfixed(-2788.0/65536.0,1,-nbitq), 
to_sfixed(-1937.0/65536.0,1,-nbitq), 
to_sfixed(105.0/65536.0,1,-nbitq), 
to_sfixed(571.0/65536.0,1,-nbitq), 
to_sfixed(-2131.0/65536.0,1,-nbitq), 
to_sfixed(-1958.0/65536.0,1,-nbitq), 
to_sfixed(3790.0/65536.0,1,-nbitq), 
to_sfixed(-158.0/65536.0,1,-nbitq), 
to_sfixed(-3445.0/65536.0,1,-nbitq), 
to_sfixed(2801.0/65536.0,1,-nbitq), 
to_sfixed(2732.0/65536.0,1,-nbitq), 
to_sfixed(1754.0/65536.0,1,-nbitq), 
to_sfixed(1851.0/65536.0,1,-nbitq), 
to_sfixed(-1512.0/65536.0,1,-nbitq), 
to_sfixed(-578.0/65536.0,1,-nbitq), 
to_sfixed(139.0/65536.0,1,-nbitq), 
to_sfixed(2468.0/65536.0,1,-nbitq), 
to_sfixed(-3477.0/65536.0,1,-nbitq), 
to_sfixed(364.0/65536.0,1,-nbitq), 
to_sfixed(-982.0/65536.0,1,-nbitq), 
to_sfixed(-4219.0/65536.0,1,-nbitq), 
to_sfixed(986.0/65536.0,1,-nbitq), 
to_sfixed(1692.0/65536.0,1,-nbitq), 
to_sfixed(4825.0/65536.0,1,-nbitq), 
to_sfixed(-1012.0/65536.0,1,-nbitq), 
to_sfixed(-788.0/65536.0,1,-nbitq), 
to_sfixed(2555.0/65536.0,1,-nbitq), 
to_sfixed(-2690.0/65536.0,1,-nbitq), 
to_sfixed(307.0/65536.0,1,-nbitq), 
to_sfixed(-2461.0/65536.0,1,-nbitq), 
to_sfixed(825.0/65536.0,1,-nbitq), 
to_sfixed(2221.0/65536.0,1,-nbitq), 
to_sfixed(-3807.0/65536.0,1,-nbitq), 
to_sfixed(-6576.0/65536.0,1,-nbitq), 
to_sfixed(-1585.0/65536.0,1,-nbitq), 
to_sfixed(594.0/65536.0,1,-nbitq), 
to_sfixed(-764.0/65536.0,1,-nbitq), 
to_sfixed(1042.0/65536.0,1,-nbitq), 
to_sfixed(1616.0/65536.0,1,-nbitq), 
to_sfixed(-6776.0/65536.0,1,-nbitq), 
to_sfixed(-3046.0/65536.0,1,-nbitq), 
to_sfixed(-1362.0/65536.0,1,-nbitq), 
to_sfixed(3502.0/65536.0,1,-nbitq), 
to_sfixed(404.0/65536.0,1,-nbitq), 
to_sfixed(-2392.0/65536.0,1,-nbitq), 
to_sfixed(-3628.0/65536.0,1,-nbitq), 
to_sfixed(-2185.0/65536.0,1,-nbitq), 
to_sfixed(-1042.0/65536.0,1,-nbitq), 
to_sfixed(-1804.0/65536.0,1,-nbitq), 
to_sfixed(-2393.0/65536.0,1,-nbitq), 
to_sfixed(1228.0/65536.0,1,-nbitq), 
to_sfixed(-970.0/65536.0,1,-nbitq), 
to_sfixed(4614.0/65536.0,1,-nbitq), 
to_sfixed(7050.0/65536.0,1,-nbitq), 
to_sfixed(4169.0/65536.0,1,-nbitq), 
to_sfixed(5105.0/65536.0,1,-nbitq), 
to_sfixed(-1126.0/65536.0,1,-nbitq), 
to_sfixed(-4899.0/65536.0,1,-nbitq), 
to_sfixed(-1187.0/65536.0,1,-nbitq), 
to_sfixed(-3282.0/65536.0,1,-nbitq), 
to_sfixed(1322.0/65536.0,1,-nbitq), 
to_sfixed(77.0/65536.0,1,-nbitq), 
to_sfixed(2233.0/65536.0,1,-nbitq), 
to_sfixed(3245.0/65536.0,1,-nbitq), 
to_sfixed(-1403.0/65536.0,1,-nbitq), 
to_sfixed(2855.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3296.0/65536.0,1,-nbitq), 
to_sfixed(63.0/65536.0,1,-nbitq), 
to_sfixed(310.0/65536.0,1,-nbitq), 
to_sfixed(3443.0/65536.0,1,-nbitq), 
to_sfixed(782.0/65536.0,1,-nbitq), 
to_sfixed(2496.0/65536.0,1,-nbitq), 
to_sfixed(547.0/65536.0,1,-nbitq), 
to_sfixed(1488.0/65536.0,1,-nbitq), 
to_sfixed(501.0/65536.0,1,-nbitq), 
to_sfixed(1077.0/65536.0,1,-nbitq), 
to_sfixed(5043.0/65536.0,1,-nbitq), 
to_sfixed(3613.0/65536.0,1,-nbitq), 
to_sfixed(299.0/65536.0,1,-nbitq), 
to_sfixed(38.0/65536.0,1,-nbitq), 
to_sfixed(-1681.0/65536.0,1,-nbitq), 
to_sfixed(-1707.0/65536.0,1,-nbitq), 
to_sfixed(1581.0/65536.0,1,-nbitq), 
to_sfixed(-1579.0/65536.0,1,-nbitq), 
to_sfixed(852.0/65536.0,1,-nbitq), 
to_sfixed(1266.0/65536.0,1,-nbitq), 
to_sfixed(-752.0/65536.0,1,-nbitq), 
to_sfixed(-4438.0/65536.0,1,-nbitq), 
to_sfixed(-3598.0/65536.0,1,-nbitq), 
to_sfixed(2924.0/65536.0,1,-nbitq), 
to_sfixed(5651.0/65536.0,1,-nbitq), 
to_sfixed(7738.0/65536.0,1,-nbitq), 
to_sfixed(2926.0/65536.0,1,-nbitq), 
to_sfixed(233.0/65536.0,1,-nbitq), 
to_sfixed(3886.0/65536.0,1,-nbitq), 
to_sfixed(2778.0/65536.0,1,-nbitq), 
to_sfixed(1589.0/65536.0,1,-nbitq), 
to_sfixed(-1143.0/65536.0,1,-nbitq), 
to_sfixed(2418.0/65536.0,1,-nbitq), 
to_sfixed(1018.0/65536.0,1,-nbitq), 
to_sfixed(-2472.0/65536.0,1,-nbitq), 
to_sfixed(-1125.0/65536.0,1,-nbitq), 
to_sfixed(4793.0/65536.0,1,-nbitq), 
to_sfixed(2772.0/65536.0,1,-nbitq), 
to_sfixed(-2494.0/65536.0,1,-nbitq), 
to_sfixed(-881.0/65536.0,1,-nbitq), 
to_sfixed(-468.0/65536.0,1,-nbitq), 
to_sfixed(2460.0/65536.0,1,-nbitq), 
to_sfixed(-2950.0/65536.0,1,-nbitq), 
to_sfixed(-3121.0/65536.0,1,-nbitq), 
to_sfixed(3276.0/65536.0,1,-nbitq), 
to_sfixed(6871.0/65536.0,1,-nbitq), 
to_sfixed(-3040.0/65536.0,1,-nbitq), 
to_sfixed(267.0/65536.0,1,-nbitq), 
to_sfixed(3141.0/65536.0,1,-nbitq), 
to_sfixed(-1011.0/65536.0,1,-nbitq), 
to_sfixed(-1679.0/65536.0,1,-nbitq), 
to_sfixed(5145.0/65536.0,1,-nbitq), 
to_sfixed(2242.0/65536.0,1,-nbitq), 
to_sfixed(-3802.0/65536.0,1,-nbitq), 
to_sfixed(-1084.0/65536.0,1,-nbitq), 
to_sfixed(2209.0/65536.0,1,-nbitq), 
to_sfixed(-1282.0/65536.0,1,-nbitq), 
to_sfixed(-2808.0/65536.0,1,-nbitq), 
to_sfixed(-909.0/65536.0,1,-nbitq), 
to_sfixed(-4447.0/65536.0,1,-nbitq), 
to_sfixed(-1203.0/65536.0,1,-nbitq), 
to_sfixed(-380.0/65536.0,1,-nbitq), 
to_sfixed(-1009.0/65536.0,1,-nbitq), 
to_sfixed(-1851.0/65536.0,1,-nbitq), 
to_sfixed(-558.0/65536.0,1,-nbitq), 
to_sfixed(-5228.0/65536.0,1,-nbitq), 
to_sfixed(1317.0/65536.0,1,-nbitq), 
to_sfixed(3196.0/65536.0,1,-nbitq), 
to_sfixed(3303.0/65536.0,1,-nbitq), 
to_sfixed(-1885.0/65536.0,1,-nbitq), 
to_sfixed(608.0/65536.0,1,-nbitq), 
to_sfixed(1258.0/65536.0,1,-nbitq), 
to_sfixed(-4865.0/65536.0,1,-nbitq), 
to_sfixed(855.0/65536.0,1,-nbitq), 
to_sfixed(2332.0/65536.0,1,-nbitq), 
to_sfixed(2977.0/65536.0,1,-nbitq), 
to_sfixed(-488.0/65536.0,1,-nbitq), 
to_sfixed(-1966.0/65536.0,1,-nbitq), 
to_sfixed(-2767.0/65536.0,1,-nbitq), 
to_sfixed(1013.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1491.0/65536.0,1,-nbitq), 
to_sfixed(-2624.0/65536.0,1,-nbitq), 
to_sfixed(-832.0/65536.0,1,-nbitq), 
to_sfixed(5252.0/65536.0,1,-nbitq), 
to_sfixed(5629.0/65536.0,1,-nbitq), 
to_sfixed(1450.0/65536.0,1,-nbitq), 
to_sfixed(2184.0/65536.0,1,-nbitq), 
to_sfixed(-526.0/65536.0,1,-nbitq), 
to_sfixed(-1387.0/65536.0,1,-nbitq), 
to_sfixed(923.0/65536.0,1,-nbitq), 
to_sfixed(1469.0/65536.0,1,-nbitq), 
to_sfixed(-729.0/65536.0,1,-nbitq), 
to_sfixed(-1701.0/65536.0,1,-nbitq), 
to_sfixed(1278.0/65536.0,1,-nbitq), 
to_sfixed(-2522.0/65536.0,1,-nbitq), 
to_sfixed(-1805.0/65536.0,1,-nbitq), 
to_sfixed(-1684.0/65536.0,1,-nbitq), 
to_sfixed(996.0/65536.0,1,-nbitq), 
to_sfixed(3986.0/65536.0,1,-nbitq), 
to_sfixed(376.0/65536.0,1,-nbitq), 
to_sfixed(-14.0/65536.0,1,-nbitq), 
to_sfixed(-11195.0/65536.0,1,-nbitq), 
to_sfixed(-6755.0/65536.0,1,-nbitq), 
to_sfixed(-356.0/65536.0,1,-nbitq), 
to_sfixed(3832.0/65536.0,1,-nbitq), 
to_sfixed(8692.0/65536.0,1,-nbitq), 
to_sfixed(4019.0/65536.0,1,-nbitq), 
to_sfixed(2790.0/65536.0,1,-nbitq), 
to_sfixed(2393.0/65536.0,1,-nbitq), 
to_sfixed(904.0/65536.0,1,-nbitq), 
to_sfixed(-1719.0/65536.0,1,-nbitq), 
to_sfixed(-1365.0/65536.0,1,-nbitq), 
to_sfixed(553.0/65536.0,1,-nbitq), 
to_sfixed(-67.0/65536.0,1,-nbitq), 
to_sfixed(-3192.0/65536.0,1,-nbitq), 
to_sfixed(-2600.0/65536.0,1,-nbitq), 
to_sfixed(350.0/65536.0,1,-nbitq), 
to_sfixed(326.0/65536.0,1,-nbitq), 
to_sfixed(-1346.0/65536.0,1,-nbitq), 
to_sfixed(2199.0/65536.0,1,-nbitq), 
to_sfixed(2285.0/65536.0,1,-nbitq), 
to_sfixed(1116.0/65536.0,1,-nbitq), 
to_sfixed(-2056.0/65536.0,1,-nbitq), 
to_sfixed(-2088.0/65536.0,1,-nbitq), 
to_sfixed(1627.0/65536.0,1,-nbitq), 
to_sfixed(7007.0/65536.0,1,-nbitq), 
to_sfixed(16.0/65536.0,1,-nbitq), 
to_sfixed(-1137.0/65536.0,1,-nbitq), 
to_sfixed(-2223.0/65536.0,1,-nbitq), 
to_sfixed(4124.0/65536.0,1,-nbitq), 
to_sfixed(-442.0/65536.0,1,-nbitq), 
to_sfixed(3931.0/65536.0,1,-nbitq), 
to_sfixed(327.0/65536.0,1,-nbitq), 
to_sfixed(-3410.0/65536.0,1,-nbitq), 
to_sfixed(-3087.0/65536.0,1,-nbitq), 
to_sfixed(-560.0/65536.0,1,-nbitq), 
to_sfixed(-449.0/65536.0,1,-nbitq), 
to_sfixed(-1843.0/65536.0,1,-nbitq), 
to_sfixed(1244.0/65536.0,1,-nbitq), 
to_sfixed(1992.0/65536.0,1,-nbitq), 
to_sfixed(371.0/65536.0,1,-nbitq), 
to_sfixed(2176.0/65536.0,1,-nbitq), 
to_sfixed(1426.0/65536.0,1,-nbitq), 
to_sfixed(-302.0/65536.0,1,-nbitq), 
to_sfixed(1567.0/65536.0,1,-nbitq), 
to_sfixed(-640.0/65536.0,1,-nbitq), 
to_sfixed(2166.0/65536.0,1,-nbitq), 
to_sfixed(5500.0/65536.0,1,-nbitq), 
to_sfixed(3501.0/65536.0,1,-nbitq), 
to_sfixed(-2650.0/65536.0,1,-nbitq), 
to_sfixed(747.0/65536.0,1,-nbitq), 
to_sfixed(129.0/65536.0,1,-nbitq), 
to_sfixed(-2226.0/65536.0,1,-nbitq), 
to_sfixed(-860.0/65536.0,1,-nbitq), 
to_sfixed(1977.0/65536.0,1,-nbitq), 
to_sfixed(1053.0/65536.0,1,-nbitq), 
to_sfixed(-681.0/65536.0,1,-nbitq), 
to_sfixed(934.0/65536.0,1,-nbitq), 
to_sfixed(-3173.0/65536.0,1,-nbitq), 
to_sfixed(-518.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2169.0/65536.0,1,-nbitq), 
to_sfixed(-828.0/65536.0,1,-nbitq), 
to_sfixed(6499.0/65536.0,1,-nbitq), 
to_sfixed(811.0/65536.0,1,-nbitq), 
to_sfixed(4160.0/65536.0,1,-nbitq), 
to_sfixed(2281.0/65536.0,1,-nbitq), 
to_sfixed(-599.0/65536.0,1,-nbitq), 
to_sfixed(-827.0/65536.0,1,-nbitq), 
to_sfixed(1075.0/65536.0,1,-nbitq), 
to_sfixed(-269.0/65536.0,1,-nbitq), 
to_sfixed(1169.0/65536.0,1,-nbitq), 
to_sfixed(4660.0/65536.0,1,-nbitq), 
to_sfixed(-2190.0/65536.0,1,-nbitq), 
to_sfixed(-1259.0/65536.0,1,-nbitq), 
to_sfixed(1327.0/65536.0,1,-nbitq), 
to_sfixed(-1845.0/65536.0,1,-nbitq), 
to_sfixed(1354.0/65536.0,1,-nbitq), 
to_sfixed(1660.0/65536.0,1,-nbitq), 
to_sfixed(600.0/65536.0,1,-nbitq), 
to_sfixed(-819.0/65536.0,1,-nbitq), 
to_sfixed(-3941.0/65536.0,1,-nbitq), 
to_sfixed(-3406.0/65536.0,1,-nbitq), 
to_sfixed(-2043.0/65536.0,1,-nbitq), 
to_sfixed(110.0/65536.0,1,-nbitq), 
to_sfixed(137.0/65536.0,1,-nbitq), 
to_sfixed(6006.0/65536.0,1,-nbitq), 
to_sfixed(663.0/65536.0,1,-nbitq), 
to_sfixed(-2413.0/65536.0,1,-nbitq), 
to_sfixed(-854.0/65536.0,1,-nbitq), 
to_sfixed(-3427.0/65536.0,1,-nbitq), 
to_sfixed(2417.0/65536.0,1,-nbitq), 
to_sfixed(1867.0/65536.0,1,-nbitq), 
to_sfixed(4728.0/65536.0,1,-nbitq), 
to_sfixed(-1666.0/65536.0,1,-nbitq), 
to_sfixed(1650.0/65536.0,1,-nbitq), 
to_sfixed(933.0/65536.0,1,-nbitq), 
to_sfixed(5870.0/65536.0,1,-nbitq), 
to_sfixed(430.0/65536.0,1,-nbitq), 
to_sfixed(-590.0/65536.0,1,-nbitq), 
to_sfixed(2365.0/65536.0,1,-nbitq), 
to_sfixed(3955.0/65536.0,1,-nbitq), 
to_sfixed(2814.0/65536.0,1,-nbitq), 
to_sfixed(-3338.0/65536.0,1,-nbitq), 
to_sfixed(-665.0/65536.0,1,-nbitq), 
to_sfixed(1958.0/65536.0,1,-nbitq), 
to_sfixed(4182.0/65536.0,1,-nbitq), 
to_sfixed(61.0/65536.0,1,-nbitq), 
to_sfixed(-2461.0/65536.0,1,-nbitq), 
to_sfixed(1523.0/65536.0,1,-nbitq), 
to_sfixed(-571.0/65536.0,1,-nbitq), 
to_sfixed(-1006.0/65536.0,1,-nbitq), 
to_sfixed(1489.0/65536.0,1,-nbitq), 
to_sfixed(-3400.0/65536.0,1,-nbitq), 
to_sfixed(-2397.0/65536.0,1,-nbitq), 
to_sfixed(-527.0/65536.0,1,-nbitq), 
to_sfixed(537.0/65536.0,1,-nbitq), 
to_sfixed(-1730.0/65536.0,1,-nbitq), 
to_sfixed(-521.0/65536.0,1,-nbitq), 
to_sfixed(2790.0/65536.0,1,-nbitq), 
to_sfixed(1315.0/65536.0,1,-nbitq), 
to_sfixed(116.0/65536.0,1,-nbitq), 
to_sfixed(-2065.0/65536.0,1,-nbitq), 
to_sfixed(-1270.0/65536.0,1,-nbitq), 
to_sfixed(126.0/65536.0,1,-nbitq), 
to_sfixed(-214.0/65536.0,1,-nbitq), 
to_sfixed(2761.0/65536.0,1,-nbitq), 
to_sfixed(442.0/65536.0,1,-nbitq), 
to_sfixed(1952.0/65536.0,1,-nbitq), 
to_sfixed(3086.0/65536.0,1,-nbitq), 
to_sfixed(-3194.0/65536.0,1,-nbitq), 
to_sfixed(-2602.0/65536.0,1,-nbitq), 
to_sfixed(-1103.0/65536.0,1,-nbitq), 
to_sfixed(-5204.0/65536.0,1,-nbitq), 
to_sfixed(2466.0/65536.0,1,-nbitq), 
to_sfixed(317.0/65536.0,1,-nbitq), 
to_sfixed(-1064.0/65536.0,1,-nbitq), 
to_sfixed(-1135.0/65536.0,1,-nbitq), 
to_sfixed(-673.0/65536.0,1,-nbitq), 
to_sfixed(-1762.0/65536.0,1,-nbitq), 
to_sfixed(1239.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1465.0/65536.0,1,-nbitq), 
to_sfixed(824.0/65536.0,1,-nbitq), 
to_sfixed(2675.0/65536.0,1,-nbitq), 
to_sfixed(4.0/65536.0,1,-nbitq), 
to_sfixed(3522.0/65536.0,1,-nbitq), 
to_sfixed(-2782.0/65536.0,1,-nbitq), 
to_sfixed(-533.0/65536.0,1,-nbitq), 
to_sfixed(1174.0/65536.0,1,-nbitq), 
to_sfixed(1252.0/65536.0,1,-nbitq), 
to_sfixed(642.0/65536.0,1,-nbitq), 
to_sfixed(293.0/65536.0,1,-nbitq), 
to_sfixed(29.0/65536.0,1,-nbitq), 
to_sfixed(31.0/65536.0,1,-nbitq), 
to_sfixed(-682.0/65536.0,1,-nbitq), 
to_sfixed(1390.0/65536.0,1,-nbitq), 
to_sfixed(2496.0/65536.0,1,-nbitq), 
to_sfixed(1973.0/65536.0,1,-nbitq), 
to_sfixed(284.0/65536.0,1,-nbitq), 
to_sfixed(337.0/65536.0,1,-nbitq), 
to_sfixed(-35.0/65536.0,1,-nbitq), 
to_sfixed(-2890.0/65536.0,1,-nbitq), 
to_sfixed(329.0/65536.0,1,-nbitq), 
to_sfixed(549.0/65536.0,1,-nbitq), 
to_sfixed(1536.0/65536.0,1,-nbitq), 
to_sfixed(-867.0/65536.0,1,-nbitq), 
to_sfixed(5534.0/65536.0,1,-nbitq), 
to_sfixed(-2273.0/65536.0,1,-nbitq), 
to_sfixed(1208.0/65536.0,1,-nbitq), 
to_sfixed(-2882.0/65536.0,1,-nbitq), 
to_sfixed(-983.0/65536.0,1,-nbitq), 
to_sfixed(-469.0/65536.0,1,-nbitq), 
to_sfixed(1955.0/65536.0,1,-nbitq), 
to_sfixed(458.0/65536.0,1,-nbitq), 
to_sfixed(1616.0/65536.0,1,-nbitq), 
to_sfixed(-1223.0/65536.0,1,-nbitq), 
to_sfixed(-2042.0/65536.0,1,-nbitq), 
to_sfixed(3927.0/65536.0,1,-nbitq), 
to_sfixed(786.0/65536.0,1,-nbitq), 
to_sfixed(-252.0/65536.0,1,-nbitq), 
to_sfixed(1514.0/65536.0,1,-nbitq), 
to_sfixed(3151.0/65536.0,1,-nbitq), 
to_sfixed(-2156.0/65536.0,1,-nbitq), 
to_sfixed(-4854.0/65536.0,1,-nbitq), 
to_sfixed(-704.0/65536.0,1,-nbitq), 
to_sfixed(610.0/65536.0,1,-nbitq), 
to_sfixed(4675.0/65536.0,1,-nbitq), 
to_sfixed(132.0/65536.0,1,-nbitq), 
to_sfixed(-2285.0/65536.0,1,-nbitq), 
to_sfixed(477.0/65536.0,1,-nbitq), 
to_sfixed(2786.0/65536.0,1,-nbitq), 
to_sfixed(878.0/65536.0,1,-nbitq), 
to_sfixed(-2800.0/65536.0,1,-nbitq), 
to_sfixed(-3648.0/65536.0,1,-nbitq), 
to_sfixed(-219.0/65536.0,1,-nbitq), 
to_sfixed(834.0/65536.0,1,-nbitq), 
to_sfixed(4667.0/65536.0,1,-nbitq), 
to_sfixed(-2601.0/65536.0,1,-nbitq), 
to_sfixed(956.0/65536.0,1,-nbitq), 
to_sfixed(716.0/65536.0,1,-nbitq), 
to_sfixed(-133.0/65536.0,1,-nbitq), 
to_sfixed(-5867.0/65536.0,1,-nbitq), 
to_sfixed(-1823.0/65536.0,1,-nbitq), 
to_sfixed(2429.0/65536.0,1,-nbitq), 
to_sfixed(-1786.0/65536.0,1,-nbitq), 
to_sfixed(3064.0/65536.0,1,-nbitq), 
to_sfixed(170.0/65536.0,1,-nbitq), 
to_sfixed(1278.0/65536.0,1,-nbitq), 
to_sfixed(-1445.0/65536.0,1,-nbitq), 
to_sfixed(1743.0/65536.0,1,-nbitq), 
to_sfixed(-5205.0/65536.0,1,-nbitq), 
to_sfixed(-1674.0/65536.0,1,-nbitq), 
to_sfixed(-2688.0/65536.0,1,-nbitq), 
to_sfixed(-5057.0/65536.0,1,-nbitq), 
to_sfixed(-539.0/65536.0,1,-nbitq), 
to_sfixed(626.0/65536.0,1,-nbitq), 
to_sfixed(824.0/65536.0,1,-nbitq), 
to_sfixed(5912.0/65536.0,1,-nbitq), 
to_sfixed(1422.0/65536.0,1,-nbitq), 
to_sfixed(1715.0/65536.0,1,-nbitq), 
to_sfixed(2342.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1392.0/65536.0,1,-nbitq), 
to_sfixed(1047.0/65536.0,1,-nbitq), 
to_sfixed(933.0/65536.0,1,-nbitq), 
to_sfixed(-1629.0/65536.0,1,-nbitq), 
to_sfixed(5170.0/65536.0,1,-nbitq), 
to_sfixed(575.0/65536.0,1,-nbitq), 
to_sfixed(132.0/65536.0,1,-nbitq), 
to_sfixed(-805.0/65536.0,1,-nbitq), 
to_sfixed(-889.0/65536.0,1,-nbitq), 
to_sfixed(-1157.0/65536.0,1,-nbitq), 
to_sfixed(-3353.0/65536.0,1,-nbitq), 
to_sfixed(5447.0/65536.0,1,-nbitq), 
to_sfixed(-823.0/65536.0,1,-nbitq), 
to_sfixed(4128.0/65536.0,1,-nbitq), 
to_sfixed(1565.0/65536.0,1,-nbitq), 
to_sfixed(-1265.0/65536.0,1,-nbitq), 
to_sfixed(-2755.0/65536.0,1,-nbitq), 
to_sfixed(-3710.0/65536.0,1,-nbitq), 
to_sfixed(2766.0/65536.0,1,-nbitq), 
to_sfixed(2110.0/65536.0,1,-nbitq), 
to_sfixed(-5852.0/65536.0,1,-nbitq), 
to_sfixed(384.0/65536.0,1,-nbitq), 
to_sfixed(2668.0/65536.0,1,-nbitq), 
to_sfixed(4555.0/65536.0,1,-nbitq), 
to_sfixed(1051.0/65536.0,1,-nbitq), 
to_sfixed(569.0/65536.0,1,-nbitq), 
to_sfixed(-1815.0/65536.0,1,-nbitq), 
to_sfixed(-1809.0/65536.0,1,-nbitq), 
to_sfixed(-3736.0/65536.0,1,-nbitq), 
to_sfixed(-2460.0/65536.0,1,-nbitq), 
to_sfixed(-2409.0/65536.0,1,-nbitq), 
to_sfixed(-1287.0/65536.0,1,-nbitq), 
to_sfixed(-38.0/65536.0,1,-nbitq), 
to_sfixed(-170.0/65536.0,1,-nbitq), 
to_sfixed(-372.0/65536.0,1,-nbitq), 
to_sfixed(-3227.0/65536.0,1,-nbitq), 
to_sfixed(2425.0/65536.0,1,-nbitq), 
to_sfixed(4602.0/65536.0,1,-nbitq), 
to_sfixed(-52.0/65536.0,1,-nbitq), 
to_sfixed(-784.0/65536.0,1,-nbitq), 
to_sfixed(-1644.0/65536.0,1,-nbitq), 
to_sfixed(-1483.0/65536.0,1,-nbitq), 
to_sfixed(-1283.0/65536.0,1,-nbitq), 
to_sfixed(-2247.0/65536.0,1,-nbitq), 
to_sfixed(-1331.0/65536.0,1,-nbitq), 
to_sfixed(393.0/65536.0,1,-nbitq), 
to_sfixed(-750.0/65536.0,1,-nbitq), 
to_sfixed(381.0/65536.0,1,-nbitq), 
to_sfixed(-780.0/65536.0,1,-nbitq), 
to_sfixed(438.0/65536.0,1,-nbitq), 
to_sfixed(-817.0/65536.0,1,-nbitq), 
to_sfixed(-2170.0/65536.0,1,-nbitq), 
to_sfixed(629.0/65536.0,1,-nbitq), 
to_sfixed(741.0/65536.0,1,-nbitq), 
to_sfixed(4118.0/65536.0,1,-nbitq), 
to_sfixed(603.0/65536.0,1,-nbitq), 
to_sfixed(-2026.0/65536.0,1,-nbitq), 
to_sfixed(-1087.0/65536.0,1,-nbitq), 
to_sfixed(1816.0/65536.0,1,-nbitq), 
to_sfixed(-558.0/65536.0,1,-nbitq), 
to_sfixed(-5622.0/65536.0,1,-nbitq), 
to_sfixed(60.0/65536.0,1,-nbitq), 
to_sfixed(1670.0/65536.0,1,-nbitq), 
to_sfixed(1054.0/65536.0,1,-nbitq), 
to_sfixed(1621.0/65536.0,1,-nbitq), 
to_sfixed(3064.0/65536.0,1,-nbitq), 
to_sfixed(699.0/65536.0,1,-nbitq), 
to_sfixed(-2275.0/65536.0,1,-nbitq), 
to_sfixed(3249.0/65536.0,1,-nbitq), 
to_sfixed(915.0/65536.0,1,-nbitq), 
to_sfixed(1509.0/65536.0,1,-nbitq), 
to_sfixed(387.0/65536.0,1,-nbitq), 
to_sfixed(-930.0/65536.0,1,-nbitq), 
to_sfixed(-486.0/65536.0,1,-nbitq), 
to_sfixed(-24.0/65536.0,1,-nbitq), 
to_sfixed(1157.0/65536.0,1,-nbitq), 
to_sfixed(5347.0/65536.0,1,-nbitq), 
to_sfixed(4.0/65536.0,1,-nbitq), 
to_sfixed(-467.0/65536.0,1,-nbitq), 
to_sfixed(-1592.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-991.0/65536.0,1,-nbitq), 
to_sfixed(-950.0/65536.0,1,-nbitq), 
to_sfixed(1317.0/65536.0,1,-nbitq), 
to_sfixed(-300.0/65536.0,1,-nbitq), 
to_sfixed(4463.0/65536.0,1,-nbitq), 
to_sfixed(424.0/65536.0,1,-nbitq), 
to_sfixed(1828.0/65536.0,1,-nbitq), 
to_sfixed(32.0/65536.0,1,-nbitq), 
to_sfixed(452.0/65536.0,1,-nbitq), 
to_sfixed(951.0/65536.0,1,-nbitq), 
to_sfixed(197.0/65536.0,1,-nbitq), 
to_sfixed(4542.0/65536.0,1,-nbitq), 
to_sfixed(940.0/65536.0,1,-nbitq), 
to_sfixed(-217.0/65536.0,1,-nbitq), 
to_sfixed(-2554.0/65536.0,1,-nbitq), 
to_sfixed(3217.0/65536.0,1,-nbitq), 
to_sfixed(1233.0/65536.0,1,-nbitq), 
to_sfixed(-1895.0/65536.0,1,-nbitq), 
to_sfixed(-754.0/65536.0,1,-nbitq), 
to_sfixed(2905.0/65536.0,1,-nbitq), 
to_sfixed(-4338.0/65536.0,1,-nbitq), 
to_sfixed(50.0/65536.0,1,-nbitq), 
to_sfixed(-1990.0/65536.0,1,-nbitq), 
to_sfixed(-707.0/65536.0,1,-nbitq), 
to_sfixed(-1236.0/65536.0,1,-nbitq), 
to_sfixed(-875.0/65536.0,1,-nbitq), 
to_sfixed(-1331.0/65536.0,1,-nbitq), 
to_sfixed(-1609.0/65536.0,1,-nbitq), 
to_sfixed(-3151.0/65536.0,1,-nbitq), 
to_sfixed(2013.0/65536.0,1,-nbitq), 
to_sfixed(161.0/65536.0,1,-nbitq), 
to_sfixed(336.0/65536.0,1,-nbitq), 
to_sfixed(-3056.0/65536.0,1,-nbitq), 
to_sfixed(22.0/65536.0,1,-nbitq), 
to_sfixed(-53.0/65536.0,1,-nbitq), 
to_sfixed(2104.0/65536.0,1,-nbitq), 
to_sfixed(4145.0/65536.0,1,-nbitq), 
to_sfixed(-347.0/65536.0,1,-nbitq), 
to_sfixed(1233.0/65536.0,1,-nbitq), 
to_sfixed(2002.0/65536.0,1,-nbitq), 
to_sfixed(-3108.0/65536.0,1,-nbitq), 
to_sfixed(-983.0/65536.0,1,-nbitq), 
to_sfixed(-7523.0/65536.0,1,-nbitq), 
to_sfixed(-1824.0/65536.0,1,-nbitq), 
to_sfixed(-1205.0/65536.0,1,-nbitq), 
to_sfixed(955.0/65536.0,1,-nbitq), 
to_sfixed(1098.0/65536.0,1,-nbitq), 
to_sfixed(-13.0/65536.0,1,-nbitq), 
to_sfixed(-1998.0/65536.0,1,-nbitq), 
to_sfixed(7.0/65536.0,1,-nbitq), 
to_sfixed(1891.0/65536.0,1,-nbitq), 
to_sfixed(-317.0/65536.0,1,-nbitq), 
to_sfixed(-1087.0/65536.0,1,-nbitq), 
to_sfixed(1840.0/65536.0,1,-nbitq), 
to_sfixed(865.0/65536.0,1,-nbitq), 
to_sfixed(3300.0/65536.0,1,-nbitq), 
to_sfixed(-2591.0/65536.0,1,-nbitq), 
to_sfixed(-2212.0/65536.0,1,-nbitq), 
to_sfixed(843.0/65536.0,1,-nbitq), 
to_sfixed(3809.0/65536.0,1,-nbitq), 
to_sfixed(3114.0/65536.0,1,-nbitq), 
to_sfixed(2402.0/65536.0,1,-nbitq), 
to_sfixed(472.0/65536.0,1,-nbitq), 
to_sfixed(-2675.0/65536.0,1,-nbitq), 
to_sfixed(1893.0/65536.0,1,-nbitq), 
to_sfixed(3068.0/65536.0,1,-nbitq), 
to_sfixed(-150.0/65536.0,1,-nbitq), 
to_sfixed(290.0/65536.0,1,-nbitq), 
to_sfixed(1134.0/65536.0,1,-nbitq), 
to_sfixed(-2476.0/65536.0,1,-nbitq), 
to_sfixed(2083.0/65536.0,1,-nbitq), 
to_sfixed(-3453.0/65536.0,1,-nbitq), 
to_sfixed(1262.0/65536.0,1,-nbitq), 
to_sfixed(-2362.0/65536.0,1,-nbitq), 
to_sfixed(1181.0/65536.0,1,-nbitq), 
to_sfixed(-1674.0/65536.0,1,-nbitq), 
to_sfixed(-2317.0/65536.0,1,-nbitq), 
to_sfixed(-127.0/65536.0,1,-nbitq), 
to_sfixed(-884.0/65536.0,1,-nbitq), 
to_sfixed(-392.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1878.0/65536.0,1,-nbitq), 
to_sfixed(-347.0/65536.0,1,-nbitq), 
to_sfixed(2789.0/65536.0,1,-nbitq), 
to_sfixed(-1625.0/65536.0,1,-nbitq), 
to_sfixed(-1140.0/65536.0,1,-nbitq), 
to_sfixed(822.0/65536.0,1,-nbitq), 
to_sfixed(337.0/65536.0,1,-nbitq), 
to_sfixed(-238.0/65536.0,1,-nbitq), 
to_sfixed(345.0/65536.0,1,-nbitq), 
to_sfixed(2038.0/65536.0,1,-nbitq), 
to_sfixed(2921.0/65536.0,1,-nbitq), 
to_sfixed(3616.0/65536.0,1,-nbitq), 
to_sfixed(1055.0/65536.0,1,-nbitq), 
to_sfixed(-891.0/65536.0,1,-nbitq), 
to_sfixed(-1639.0/65536.0,1,-nbitq), 
to_sfixed(-1415.0/65536.0,1,-nbitq), 
to_sfixed(2013.0/65536.0,1,-nbitq), 
to_sfixed(-1669.0/65536.0,1,-nbitq), 
to_sfixed(1401.0/65536.0,1,-nbitq), 
to_sfixed(-90.0/65536.0,1,-nbitq), 
to_sfixed(-1444.0/65536.0,1,-nbitq), 
to_sfixed(2135.0/65536.0,1,-nbitq), 
to_sfixed(1210.0/65536.0,1,-nbitq), 
to_sfixed(640.0/65536.0,1,-nbitq), 
to_sfixed(-3111.0/65536.0,1,-nbitq), 
to_sfixed(-1806.0/65536.0,1,-nbitq), 
to_sfixed(-2284.0/65536.0,1,-nbitq), 
to_sfixed(1804.0/65536.0,1,-nbitq), 
to_sfixed(-4187.0/65536.0,1,-nbitq), 
to_sfixed(2011.0/65536.0,1,-nbitq), 
to_sfixed(-3044.0/65536.0,1,-nbitq), 
to_sfixed(-1482.0/65536.0,1,-nbitq), 
to_sfixed(-2800.0/65536.0,1,-nbitq), 
to_sfixed(1372.0/65536.0,1,-nbitq), 
to_sfixed(-3064.0/65536.0,1,-nbitq), 
to_sfixed(1428.0/65536.0,1,-nbitq), 
to_sfixed(-42.0/65536.0,1,-nbitq), 
to_sfixed(-5507.0/65536.0,1,-nbitq), 
to_sfixed(-454.0/65536.0,1,-nbitq), 
to_sfixed(1592.0/65536.0,1,-nbitq), 
to_sfixed(-3898.0/65536.0,1,-nbitq), 
to_sfixed(-2534.0/65536.0,1,-nbitq), 
to_sfixed(-7546.0/65536.0,1,-nbitq), 
to_sfixed(1135.0/65536.0,1,-nbitq), 
to_sfixed(2524.0/65536.0,1,-nbitq), 
to_sfixed(624.0/65536.0,1,-nbitq), 
to_sfixed(1925.0/65536.0,1,-nbitq), 
to_sfixed(534.0/65536.0,1,-nbitq), 
to_sfixed(-1273.0/65536.0,1,-nbitq), 
to_sfixed(-227.0/65536.0,1,-nbitq), 
to_sfixed(2180.0/65536.0,1,-nbitq), 
to_sfixed(-2060.0/65536.0,1,-nbitq), 
to_sfixed(1801.0/65536.0,1,-nbitq), 
to_sfixed(-760.0/65536.0,1,-nbitq), 
to_sfixed(766.0/65536.0,1,-nbitq), 
to_sfixed(-1311.0/65536.0,1,-nbitq), 
to_sfixed(2860.0/65536.0,1,-nbitq), 
to_sfixed(2162.0/65536.0,1,-nbitq), 
to_sfixed(324.0/65536.0,1,-nbitq), 
to_sfixed(-246.0/65536.0,1,-nbitq), 
to_sfixed(1287.0/65536.0,1,-nbitq), 
to_sfixed(2571.0/65536.0,1,-nbitq), 
to_sfixed(1238.0/65536.0,1,-nbitq), 
to_sfixed(1749.0/65536.0,1,-nbitq), 
to_sfixed(-1787.0/65536.0,1,-nbitq), 
to_sfixed(479.0/65536.0,1,-nbitq), 
to_sfixed(-5288.0/65536.0,1,-nbitq), 
to_sfixed(1369.0/65536.0,1,-nbitq), 
to_sfixed(2371.0/65536.0,1,-nbitq), 
to_sfixed(2217.0/65536.0,1,-nbitq), 
to_sfixed(744.0/65536.0,1,-nbitq), 
to_sfixed(295.0/65536.0,1,-nbitq), 
to_sfixed(-41.0/65536.0,1,-nbitq), 
to_sfixed(-1477.0/65536.0,1,-nbitq), 
to_sfixed(-1525.0/65536.0,1,-nbitq), 
to_sfixed(-807.0/65536.0,1,-nbitq), 
to_sfixed(1181.0/65536.0,1,-nbitq), 
to_sfixed(-1303.0/65536.0,1,-nbitq), 
to_sfixed(-1843.0/65536.0,1,-nbitq), 
to_sfixed(2184.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3.0/65536.0,1,-nbitq), 
to_sfixed(-3257.0/65536.0,1,-nbitq), 
to_sfixed(4644.0/65536.0,1,-nbitq), 
to_sfixed(-3061.0/65536.0,1,-nbitq), 
to_sfixed(2341.0/65536.0,1,-nbitq), 
to_sfixed(321.0/65536.0,1,-nbitq), 
to_sfixed(2319.0/65536.0,1,-nbitq), 
to_sfixed(-3016.0/65536.0,1,-nbitq), 
to_sfixed(2355.0/65536.0,1,-nbitq), 
to_sfixed(2779.0/65536.0,1,-nbitq), 
to_sfixed(1463.0/65536.0,1,-nbitq), 
to_sfixed(4437.0/65536.0,1,-nbitq), 
to_sfixed(1281.0/65536.0,1,-nbitq), 
to_sfixed(586.0/65536.0,1,-nbitq), 
to_sfixed(2693.0/65536.0,1,-nbitq), 
to_sfixed(-1945.0/65536.0,1,-nbitq), 
to_sfixed(-2170.0/65536.0,1,-nbitq), 
to_sfixed(1886.0/65536.0,1,-nbitq), 
to_sfixed(4.0/65536.0,1,-nbitq), 
to_sfixed(2611.0/65536.0,1,-nbitq), 
to_sfixed(-437.0/65536.0,1,-nbitq), 
to_sfixed(-1418.0/65536.0,1,-nbitq), 
to_sfixed(-283.0/65536.0,1,-nbitq), 
to_sfixed(-1192.0/65536.0,1,-nbitq), 
to_sfixed(-2163.0/65536.0,1,-nbitq), 
to_sfixed(274.0/65536.0,1,-nbitq), 
to_sfixed(2160.0/65536.0,1,-nbitq), 
to_sfixed(-1702.0/65536.0,1,-nbitq), 
to_sfixed(722.0/65536.0,1,-nbitq), 
to_sfixed(139.0/65536.0,1,-nbitq), 
to_sfixed(345.0/65536.0,1,-nbitq), 
to_sfixed(-2068.0/65536.0,1,-nbitq), 
to_sfixed(936.0/65536.0,1,-nbitq), 
to_sfixed(1068.0/65536.0,1,-nbitq), 
to_sfixed(2177.0/65536.0,1,-nbitq), 
to_sfixed(-1465.0/65536.0,1,-nbitq), 
to_sfixed(-321.0/65536.0,1,-nbitq), 
to_sfixed(-4233.0/65536.0,1,-nbitq), 
to_sfixed(-2161.0/65536.0,1,-nbitq), 
to_sfixed(-1727.0/65536.0,1,-nbitq), 
to_sfixed(-482.0/65536.0,1,-nbitq), 
to_sfixed(748.0/65536.0,1,-nbitq), 
to_sfixed(-2399.0/65536.0,1,-nbitq), 
to_sfixed(1841.0/65536.0,1,-nbitq), 
to_sfixed(129.0/65536.0,1,-nbitq), 
to_sfixed(1079.0/65536.0,1,-nbitq), 
to_sfixed(-1844.0/65536.0,1,-nbitq), 
to_sfixed(363.0/65536.0,1,-nbitq), 
to_sfixed(-709.0/65536.0,1,-nbitq), 
to_sfixed(-56.0/65536.0,1,-nbitq), 
to_sfixed(9.0/65536.0,1,-nbitq), 
to_sfixed(570.0/65536.0,1,-nbitq), 
to_sfixed(-552.0/65536.0,1,-nbitq), 
to_sfixed(-1985.0/65536.0,1,-nbitq), 
to_sfixed(2914.0/65536.0,1,-nbitq), 
to_sfixed(2499.0/65536.0,1,-nbitq), 
to_sfixed(3079.0/65536.0,1,-nbitq), 
to_sfixed(2033.0/65536.0,1,-nbitq), 
to_sfixed(172.0/65536.0,1,-nbitq), 
to_sfixed(-60.0/65536.0,1,-nbitq), 
to_sfixed(-1865.0/65536.0,1,-nbitq), 
to_sfixed(-2918.0/65536.0,1,-nbitq), 
to_sfixed(-2435.0/65536.0,1,-nbitq), 
to_sfixed(-2420.0/65536.0,1,-nbitq), 
to_sfixed(1516.0/65536.0,1,-nbitq), 
to_sfixed(3197.0/65536.0,1,-nbitq), 
to_sfixed(-343.0/65536.0,1,-nbitq), 
to_sfixed(-824.0/65536.0,1,-nbitq), 
to_sfixed(2773.0/65536.0,1,-nbitq), 
to_sfixed(1999.0/65536.0,1,-nbitq), 
to_sfixed(-625.0/65536.0,1,-nbitq), 
to_sfixed(-1071.0/65536.0,1,-nbitq), 
to_sfixed(-1717.0/65536.0,1,-nbitq), 
to_sfixed(-2479.0/65536.0,1,-nbitq), 
to_sfixed(2540.0/65536.0,1,-nbitq), 
to_sfixed(3270.0/65536.0,1,-nbitq), 
to_sfixed(-1983.0/65536.0,1,-nbitq), 
to_sfixed(951.0/65536.0,1,-nbitq), 
to_sfixed(1209.0/65536.0,1,-nbitq), 
to_sfixed(4820.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1165.0/65536.0,1,-nbitq), 
to_sfixed(-2149.0/65536.0,1,-nbitq), 
to_sfixed(3647.0/65536.0,1,-nbitq), 
to_sfixed(-2751.0/65536.0,1,-nbitq), 
to_sfixed(2446.0/65536.0,1,-nbitq), 
to_sfixed(752.0/65536.0,1,-nbitq), 
to_sfixed(-3264.0/65536.0,1,-nbitq), 
to_sfixed(1287.0/65536.0,1,-nbitq), 
to_sfixed(236.0/65536.0,1,-nbitq), 
to_sfixed(343.0/65536.0,1,-nbitq), 
to_sfixed(1867.0/65536.0,1,-nbitq), 
to_sfixed(2036.0/65536.0,1,-nbitq), 
to_sfixed(941.0/65536.0,1,-nbitq), 
to_sfixed(2308.0/65536.0,1,-nbitq), 
to_sfixed(1437.0/65536.0,1,-nbitq), 
to_sfixed(-806.0/65536.0,1,-nbitq), 
to_sfixed(-1236.0/65536.0,1,-nbitq), 
to_sfixed(-997.0/65536.0,1,-nbitq), 
to_sfixed(2111.0/65536.0,1,-nbitq), 
to_sfixed(2330.0/65536.0,1,-nbitq), 
to_sfixed(-1573.0/65536.0,1,-nbitq), 
to_sfixed(1117.0/65536.0,1,-nbitq), 
to_sfixed(-185.0/65536.0,1,-nbitq), 
to_sfixed(3982.0/65536.0,1,-nbitq), 
to_sfixed(-2234.0/65536.0,1,-nbitq), 
to_sfixed(-812.0/65536.0,1,-nbitq), 
to_sfixed(-3312.0/65536.0,1,-nbitq), 
to_sfixed(2233.0/65536.0,1,-nbitq), 
to_sfixed(-1053.0/65536.0,1,-nbitq), 
to_sfixed(2457.0/65536.0,1,-nbitq), 
to_sfixed(-3201.0/65536.0,1,-nbitq), 
to_sfixed(-2312.0/65536.0,1,-nbitq), 
to_sfixed(598.0/65536.0,1,-nbitq), 
to_sfixed(-3146.0/65536.0,1,-nbitq), 
to_sfixed(-253.0/65536.0,1,-nbitq), 
to_sfixed(-1294.0/65536.0,1,-nbitq), 
to_sfixed(1747.0/65536.0,1,-nbitq), 
to_sfixed(-3045.0/65536.0,1,-nbitq), 
to_sfixed(1756.0/65536.0,1,-nbitq), 
to_sfixed(-1188.0/65536.0,1,-nbitq), 
to_sfixed(-1316.0/65536.0,1,-nbitq), 
to_sfixed(47.0/65536.0,1,-nbitq), 
to_sfixed(-5411.0/65536.0,1,-nbitq), 
to_sfixed(1710.0/65536.0,1,-nbitq), 
to_sfixed(2935.0/65536.0,1,-nbitq), 
to_sfixed(2794.0/65536.0,1,-nbitq), 
to_sfixed(91.0/65536.0,1,-nbitq), 
to_sfixed(-1100.0/65536.0,1,-nbitq), 
to_sfixed(1836.0/65536.0,1,-nbitq), 
to_sfixed(1002.0/65536.0,1,-nbitq), 
to_sfixed(819.0/65536.0,1,-nbitq), 
to_sfixed(-2721.0/65536.0,1,-nbitq), 
to_sfixed(323.0/65536.0,1,-nbitq), 
to_sfixed(-2481.0/65536.0,1,-nbitq), 
to_sfixed(982.0/65536.0,1,-nbitq), 
to_sfixed(3284.0/65536.0,1,-nbitq), 
to_sfixed(-347.0/65536.0,1,-nbitq), 
to_sfixed(1360.0/65536.0,1,-nbitq), 
to_sfixed(-2453.0/65536.0,1,-nbitq), 
to_sfixed(2838.0/65536.0,1,-nbitq), 
to_sfixed(1310.0/65536.0,1,-nbitq), 
to_sfixed(-1536.0/65536.0,1,-nbitq), 
to_sfixed(-1723.0/65536.0,1,-nbitq), 
to_sfixed(2293.0/65536.0,1,-nbitq), 
to_sfixed(2781.0/65536.0,1,-nbitq), 
to_sfixed(149.0/65536.0,1,-nbitq), 
to_sfixed(1878.0/65536.0,1,-nbitq), 
to_sfixed(193.0/65536.0,1,-nbitq), 
to_sfixed(-1568.0/65536.0,1,-nbitq), 
to_sfixed(-1199.0/65536.0,1,-nbitq), 
to_sfixed(-968.0/65536.0,1,-nbitq), 
to_sfixed(2430.0/65536.0,1,-nbitq), 
to_sfixed(2433.0/65536.0,1,-nbitq), 
to_sfixed(-192.0/65536.0,1,-nbitq), 
to_sfixed(2084.0/65536.0,1,-nbitq), 
to_sfixed(-499.0/65536.0,1,-nbitq), 
to_sfixed(3530.0/65536.0,1,-nbitq), 
to_sfixed(4095.0/65536.0,1,-nbitq), 
to_sfixed(-2686.0/65536.0,1,-nbitq), 
to_sfixed(2906.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-600.0/65536.0,1,-nbitq), 
to_sfixed(2290.0/65536.0,1,-nbitq), 
to_sfixed(3492.0/65536.0,1,-nbitq), 
to_sfixed(-2790.0/65536.0,1,-nbitq), 
to_sfixed(-3225.0/65536.0,1,-nbitq), 
to_sfixed(-3651.0/65536.0,1,-nbitq), 
to_sfixed(680.0/65536.0,1,-nbitq), 
to_sfixed(1560.0/65536.0,1,-nbitq), 
to_sfixed(-1260.0/65536.0,1,-nbitq), 
to_sfixed(339.0/65536.0,1,-nbitq), 
to_sfixed(-1975.0/65536.0,1,-nbitq), 
to_sfixed(-594.0/65536.0,1,-nbitq), 
to_sfixed(2493.0/65536.0,1,-nbitq), 
to_sfixed(59.0/65536.0,1,-nbitq), 
to_sfixed(2230.0/65536.0,1,-nbitq), 
to_sfixed(553.0/65536.0,1,-nbitq), 
to_sfixed(-1440.0/65536.0,1,-nbitq), 
to_sfixed(2969.0/65536.0,1,-nbitq), 
to_sfixed(-725.0/65536.0,1,-nbitq), 
to_sfixed(2750.0/65536.0,1,-nbitq), 
to_sfixed(-3047.0/65536.0,1,-nbitq), 
to_sfixed(3243.0/65536.0,1,-nbitq), 
to_sfixed(911.0/65536.0,1,-nbitq), 
to_sfixed(-226.0/65536.0,1,-nbitq), 
to_sfixed(97.0/65536.0,1,-nbitq), 
to_sfixed(2492.0/65536.0,1,-nbitq), 
to_sfixed(-425.0/65536.0,1,-nbitq), 
to_sfixed(1690.0/65536.0,1,-nbitq), 
to_sfixed(-3513.0/65536.0,1,-nbitq), 
to_sfixed(-2213.0/65536.0,1,-nbitq), 
to_sfixed(-2955.0/65536.0,1,-nbitq), 
to_sfixed(-2571.0/65536.0,1,-nbitq), 
to_sfixed(-3083.0/65536.0,1,-nbitq), 
to_sfixed(-4930.0/65536.0,1,-nbitq), 
to_sfixed(-1266.0/65536.0,1,-nbitq), 
to_sfixed(2050.0/65536.0,1,-nbitq), 
to_sfixed(287.0/65536.0,1,-nbitq), 
to_sfixed(-3804.0/65536.0,1,-nbitq), 
to_sfixed(468.0/65536.0,1,-nbitq), 
to_sfixed(-1979.0/65536.0,1,-nbitq), 
to_sfixed(-388.0/65536.0,1,-nbitq), 
to_sfixed(928.0/65536.0,1,-nbitq), 
to_sfixed(-672.0/65536.0,1,-nbitq), 
to_sfixed(1934.0/65536.0,1,-nbitq), 
to_sfixed(3035.0/65536.0,1,-nbitq), 
to_sfixed(5039.0/65536.0,1,-nbitq), 
to_sfixed(1575.0/65536.0,1,-nbitq), 
to_sfixed(-3.0/65536.0,1,-nbitq), 
to_sfixed(-98.0/65536.0,1,-nbitq), 
to_sfixed(624.0/65536.0,1,-nbitq), 
to_sfixed(-1335.0/65536.0,1,-nbitq), 
to_sfixed(1425.0/65536.0,1,-nbitq), 
to_sfixed(2950.0/65536.0,1,-nbitq), 
to_sfixed(-1139.0/65536.0,1,-nbitq), 
to_sfixed(3773.0/65536.0,1,-nbitq), 
to_sfixed(-2018.0/65536.0,1,-nbitq), 
to_sfixed(1599.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(-935.0/65536.0,1,-nbitq), 
to_sfixed(5643.0/65536.0,1,-nbitq), 
to_sfixed(539.0/65536.0,1,-nbitq), 
to_sfixed(2643.0/65536.0,1,-nbitq), 
to_sfixed(858.0/65536.0,1,-nbitq), 
to_sfixed(-2044.0/65536.0,1,-nbitq), 
to_sfixed(-903.0/65536.0,1,-nbitq), 
to_sfixed(205.0/65536.0,1,-nbitq), 
to_sfixed(-2257.0/65536.0,1,-nbitq), 
to_sfixed(-3189.0/65536.0,1,-nbitq), 
to_sfixed(2273.0/65536.0,1,-nbitq), 
to_sfixed(12.0/65536.0,1,-nbitq), 
to_sfixed(-95.0/65536.0,1,-nbitq), 
to_sfixed(-2726.0/65536.0,1,-nbitq), 
to_sfixed(180.0/65536.0,1,-nbitq), 
to_sfixed(860.0/65536.0,1,-nbitq), 
to_sfixed(1521.0/65536.0,1,-nbitq), 
to_sfixed(2335.0/65536.0,1,-nbitq), 
to_sfixed(2595.0/65536.0,1,-nbitq), 
to_sfixed(1610.0/65536.0,1,-nbitq), 
to_sfixed(-287.0/65536.0,1,-nbitq), 
to_sfixed(4718.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3.0/65536.0,1,-nbitq), 
to_sfixed(1113.0/65536.0,1,-nbitq), 
to_sfixed(2357.0/65536.0,1,-nbitq), 
to_sfixed(-104.0/65536.0,1,-nbitq), 
to_sfixed(779.0/65536.0,1,-nbitq), 
to_sfixed(117.0/65536.0,1,-nbitq), 
to_sfixed(-2163.0/65536.0,1,-nbitq), 
to_sfixed(2797.0/65536.0,1,-nbitq), 
to_sfixed(-2193.0/65536.0,1,-nbitq), 
to_sfixed(550.0/65536.0,1,-nbitq), 
to_sfixed(-669.0/65536.0,1,-nbitq), 
to_sfixed(24.0/65536.0,1,-nbitq), 
to_sfixed(1245.0/65536.0,1,-nbitq), 
to_sfixed(-1588.0/65536.0,1,-nbitq), 
to_sfixed(223.0/65536.0,1,-nbitq), 
to_sfixed(3175.0/65536.0,1,-nbitq), 
to_sfixed(-593.0/65536.0,1,-nbitq), 
to_sfixed(2397.0/65536.0,1,-nbitq), 
to_sfixed(-334.0/65536.0,1,-nbitq), 
to_sfixed(-2065.0/65536.0,1,-nbitq), 
to_sfixed(-4166.0/65536.0,1,-nbitq), 
to_sfixed(2808.0/65536.0,1,-nbitq), 
to_sfixed(-330.0/65536.0,1,-nbitq), 
to_sfixed(2490.0/65536.0,1,-nbitq), 
to_sfixed(1611.0/65536.0,1,-nbitq), 
to_sfixed(865.0/65536.0,1,-nbitq), 
to_sfixed(877.0/65536.0,1,-nbitq), 
to_sfixed(-720.0/65536.0,1,-nbitq), 
to_sfixed(-810.0/65536.0,1,-nbitq), 
to_sfixed(-2321.0/65536.0,1,-nbitq), 
to_sfixed(-1088.0/65536.0,1,-nbitq), 
to_sfixed(-946.0/65536.0,1,-nbitq), 
to_sfixed(-2653.0/65536.0,1,-nbitq), 
to_sfixed(30.0/65536.0,1,-nbitq), 
to_sfixed(-1938.0/65536.0,1,-nbitq), 
to_sfixed(-2301.0/65536.0,1,-nbitq), 
to_sfixed(-369.0/65536.0,1,-nbitq), 
to_sfixed(1572.0/65536.0,1,-nbitq), 
to_sfixed(-3077.0/65536.0,1,-nbitq), 
to_sfixed(2052.0/65536.0,1,-nbitq), 
to_sfixed(-1230.0/65536.0,1,-nbitq), 
to_sfixed(1016.0/65536.0,1,-nbitq), 
to_sfixed(-2155.0/65536.0,1,-nbitq), 
to_sfixed(2145.0/65536.0,1,-nbitq), 
to_sfixed(2803.0/65536.0,1,-nbitq), 
to_sfixed(2620.0/65536.0,1,-nbitq), 
to_sfixed(1778.0/65536.0,1,-nbitq), 
to_sfixed(-1557.0/65536.0,1,-nbitq), 
to_sfixed(-616.0/65536.0,1,-nbitq), 
to_sfixed(330.0/65536.0,1,-nbitq), 
to_sfixed(265.0/65536.0,1,-nbitq), 
to_sfixed(3324.0/65536.0,1,-nbitq), 
to_sfixed(-2280.0/65536.0,1,-nbitq), 
to_sfixed(-3103.0/65536.0,1,-nbitq), 
to_sfixed(95.0/65536.0,1,-nbitq), 
to_sfixed(1783.0/65536.0,1,-nbitq), 
to_sfixed(1064.0/65536.0,1,-nbitq), 
to_sfixed(-194.0/65536.0,1,-nbitq), 
to_sfixed(-2422.0/65536.0,1,-nbitq), 
to_sfixed(4963.0/65536.0,1,-nbitq), 
to_sfixed(-3529.0/65536.0,1,-nbitq), 
to_sfixed(1116.0/65536.0,1,-nbitq), 
to_sfixed(-2387.0/65536.0,1,-nbitq), 
to_sfixed(-1768.0/65536.0,1,-nbitq), 
to_sfixed(3415.0/65536.0,1,-nbitq), 
to_sfixed(3174.0/65536.0,1,-nbitq), 
to_sfixed(2822.0/65536.0,1,-nbitq), 
to_sfixed(1699.0/65536.0,1,-nbitq), 
to_sfixed(1562.0/65536.0,1,-nbitq), 
to_sfixed(-1052.0/65536.0,1,-nbitq), 
to_sfixed(-13.0/65536.0,1,-nbitq), 
to_sfixed(-2169.0/65536.0,1,-nbitq), 
to_sfixed(1598.0/65536.0,1,-nbitq), 
to_sfixed(-2045.0/65536.0,1,-nbitq), 
to_sfixed(-8.0/65536.0,1,-nbitq), 
to_sfixed(3313.0/65536.0,1,-nbitq), 
to_sfixed(-356.0/65536.0,1,-nbitq), 
to_sfixed(566.0/65536.0,1,-nbitq), 
to_sfixed(-2648.0/65536.0,1,-nbitq), 
to_sfixed(1720.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2651.0/65536.0,1,-nbitq), 
to_sfixed(2269.0/65536.0,1,-nbitq), 
to_sfixed(-1143.0/65536.0,1,-nbitq), 
to_sfixed(-1200.0/65536.0,1,-nbitq), 
to_sfixed(743.0/65536.0,1,-nbitq), 
to_sfixed(-2413.0/65536.0,1,-nbitq), 
to_sfixed(-69.0/65536.0,1,-nbitq), 
to_sfixed(-1908.0/65536.0,1,-nbitq), 
to_sfixed(-1644.0/65536.0,1,-nbitq), 
to_sfixed(-2526.0/65536.0,1,-nbitq), 
to_sfixed(-1905.0/65536.0,1,-nbitq), 
to_sfixed(4620.0/65536.0,1,-nbitq), 
to_sfixed(-2286.0/65536.0,1,-nbitq), 
to_sfixed(147.0/65536.0,1,-nbitq), 
to_sfixed(-71.0/65536.0,1,-nbitq), 
to_sfixed(686.0/65536.0,1,-nbitq), 
to_sfixed(672.0/65536.0,1,-nbitq), 
to_sfixed(-133.0/65536.0,1,-nbitq), 
to_sfixed(-356.0/65536.0,1,-nbitq), 
to_sfixed(96.0/65536.0,1,-nbitq), 
to_sfixed(-2784.0/65536.0,1,-nbitq), 
to_sfixed(1866.0/65536.0,1,-nbitq), 
to_sfixed(2640.0/65536.0,1,-nbitq), 
to_sfixed(-238.0/65536.0,1,-nbitq), 
to_sfixed(-2107.0/65536.0,1,-nbitq), 
to_sfixed(-605.0/65536.0,1,-nbitq), 
to_sfixed(1203.0/65536.0,1,-nbitq), 
to_sfixed(2933.0/65536.0,1,-nbitq), 
to_sfixed(898.0/65536.0,1,-nbitq), 
to_sfixed(2289.0/65536.0,1,-nbitq), 
to_sfixed(-2117.0/65536.0,1,-nbitq), 
to_sfixed(262.0/65536.0,1,-nbitq), 
to_sfixed(-2863.0/65536.0,1,-nbitq), 
to_sfixed(23.0/65536.0,1,-nbitq), 
to_sfixed(1263.0/65536.0,1,-nbitq), 
to_sfixed(567.0/65536.0,1,-nbitq), 
to_sfixed(-136.0/65536.0,1,-nbitq), 
to_sfixed(-1938.0/65536.0,1,-nbitq), 
to_sfixed(1447.0/65536.0,1,-nbitq), 
to_sfixed(-1308.0/65536.0,1,-nbitq), 
to_sfixed(-1456.0/65536.0,1,-nbitq), 
to_sfixed(-725.0/65536.0,1,-nbitq), 
to_sfixed(-994.0/65536.0,1,-nbitq), 
to_sfixed(978.0/65536.0,1,-nbitq), 
to_sfixed(-482.0/65536.0,1,-nbitq), 
to_sfixed(2235.0/65536.0,1,-nbitq), 
to_sfixed(-869.0/65536.0,1,-nbitq), 
to_sfixed(63.0/65536.0,1,-nbitq), 
to_sfixed(1576.0/65536.0,1,-nbitq), 
to_sfixed(2105.0/65536.0,1,-nbitq), 
to_sfixed(2855.0/65536.0,1,-nbitq), 
to_sfixed(1170.0/65536.0,1,-nbitq), 
to_sfixed(-2752.0/65536.0,1,-nbitq), 
to_sfixed(2498.0/65536.0,1,-nbitq), 
to_sfixed(2001.0/65536.0,1,-nbitq), 
to_sfixed(2636.0/65536.0,1,-nbitq), 
to_sfixed(-1396.0/65536.0,1,-nbitq), 
to_sfixed(-32.0/65536.0,1,-nbitq), 
to_sfixed(2617.0/65536.0,1,-nbitq), 
to_sfixed(3456.0/65536.0,1,-nbitq), 
to_sfixed(1212.0/65536.0,1,-nbitq), 
to_sfixed(-1037.0/65536.0,1,-nbitq), 
to_sfixed(491.0/65536.0,1,-nbitq), 
to_sfixed(-99.0/65536.0,1,-nbitq), 
to_sfixed(2370.0/65536.0,1,-nbitq), 
to_sfixed(1747.0/65536.0,1,-nbitq), 
to_sfixed(158.0/65536.0,1,-nbitq), 
to_sfixed(-3614.0/65536.0,1,-nbitq), 
to_sfixed(605.0/65536.0,1,-nbitq), 
to_sfixed(919.0/65536.0,1,-nbitq), 
to_sfixed(2406.0/65536.0,1,-nbitq), 
to_sfixed(-4699.0/65536.0,1,-nbitq), 
to_sfixed(2017.0/65536.0,1,-nbitq), 
to_sfixed(852.0/65536.0,1,-nbitq), 
to_sfixed(1484.0/65536.0,1,-nbitq), 
to_sfixed(-695.0/65536.0,1,-nbitq), 
to_sfixed(300.0/65536.0,1,-nbitq), 
to_sfixed(4393.0/65536.0,1,-nbitq), 
to_sfixed(-544.0/65536.0,1,-nbitq), 
to_sfixed(-202.0/65536.0,1,-nbitq)  ), 
( to_sfixed(636.0/65536.0,1,-nbitq), 
to_sfixed(2478.0/65536.0,1,-nbitq), 
to_sfixed(-1270.0/65536.0,1,-nbitq), 
to_sfixed(-4010.0/65536.0,1,-nbitq), 
to_sfixed(-3262.0/65536.0,1,-nbitq), 
to_sfixed(-2455.0/65536.0,1,-nbitq), 
to_sfixed(-422.0/65536.0,1,-nbitq), 
to_sfixed(-2863.0/65536.0,1,-nbitq), 
to_sfixed(457.0/65536.0,1,-nbitq), 
to_sfixed(2704.0/65536.0,1,-nbitq), 
to_sfixed(-1820.0/65536.0,1,-nbitq), 
to_sfixed(1660.0/65536.0,1,-nbitq), 
to_sfixed(2570.0/65536.0,1,-nbitq), 
to_sfixed(2542.0/65536.0,1,-nbitq), 
to_sfixed(-1587.0/65536.0,1,-nbitq), 
to_sfixed(2507.0/65536.0,1,-nbitq), 
to_sfixed(-1685.0/65536.0,1,-nbitq), 
to_sfixed(1472.0/65536.0,1,-nbitq), 
to_sfixed(3961.0/65536.0,1,-nbitq), 
to_sfixed(2943.0/65536.0,1,-nbitq), 
to_sfixed(-1286.0/65536.0,1,-nbitq), 
to_sfixed(3046.0/65536.0,1,-nbitq), 
to_sfixed(3925.0/65536.0,1,-nbitq), 
to_sfixed(87.0/65536.0,1,-nbitq), 
to_sfixed(980.0/65536.0,1,-nbitq), 
to_sfixed(-1348.0/65536.0,1,-nbitq), 
to_sfixed(-3901.0/65536.0,1,-nbitq), 
to_sfixed(-595.0/65536.0,1,-nbitq), 
to_sfixed(-2027.0/65536.0,1,-nbitq), 
to_sfixed(-185.0/65536.0,1,-nbitq), 
to_sfixed(-2092.0/65536.0,1,-nbitq), 
to_sfixed(-3174.0/65536.0,1,-nbitq), 
to_sfixed(-5659.0/65536.0,1,-nbitq), 
to_sfixed(-3650.0/65536.0,1,-nbitq), 
to_sfixed(1399.0/65536.0,1,-nbitq), 
to_sfixed(1456.0/65536.0,1,-nbitq), 
to_sfixed(1901.0/65536.0,1,-nbitq), 
to_sfixed(-156.0/65536.0,1,-nbitq), 
to_sfixed(1858.0/65536.0,1,-nbitq), 
to_sfixed(1237.0/65536.0,1,-nbitq), 
to_sfixed(372.0/65536.0,1,-nbitq), 
to_sfixed(595.0/65536.0,1,-nbitq), 
to_sfixed(-783.0/65536.0,1,-nbitq), 
to_sfixed(1316.0/65536.0,1,-nbitq), 
to_sfixed(2086.0/65536.0,1,-nbitq), 
to_sfixed(2152.0/65536.0,1,-nbitq), 
to_sfixed(1468.0/65536.0,1,-nbitq), 
to_sfixed(-522.0/65536.0,1,-nbitq), 
to_sfixed(2652.0/65536.0,1,-nbitq), 
to_sfixed(-111.0/65536.0,1,-nbitq), 
to_sfixed(-1060.0/65536.0,1,-nbitq), 
to_sfixed(-2533.0/65536.0,1,-nbitq), 
to_sfixed(-1876.0/65536.0,1,-nbitq), 
to_sfixed(1785.0/65536.0,1,-nbitq), 
to_sfixed(3387.0/65536.0,1,-nbitq), 
to_sfixed(-2290.0/65536.0,1,-nbitq), 
to_sfixed(1664.0/65536.0,1,-nbitq), 
to_sfixed(764.0/65536.0,1,-nbitq), 
to_sfixed(-144.0/65536.0,1,-nbitq), 
to_sfixed(2101.0/65536.0,1,-nbitq), 
to_sfixed(-2660.0/65536.0,1,-nbitq), 
to_sfixed(773.0/65536.0,1,-nbitq), 
to_sfixed(849.0/65536.0,1,-nbitq), 
to_sfixed(2521.0/65536.0,1,-nbitq), 
to_sfixed(-1604.0/65536.0,1,-nbitq), 
to_sfixed(1783.0/65536.0,1,-nbitq), 
to_sfixed(1765.0/65536.0,1,-nbitq), 
to_sfixed(-2691.0/65536.0,1,-nbitq), 
to_sfixed(-2004.0/65536.0,1,-nbitq), 
to_sfixed(-1699.0/65536.0,1,-nbitq), 
to_sfixed(-2435.0/65536.0,1,-nbitq), 
to_sfixed(-110.0/65536.0,1,-nbitq), 
to_sfixed(2676.0/65536.0,1,-nbitq), 
to_sfixed(-3052.0/65536.0,1,-nbitq), 
to_sfixed(-2353.0/65536.0,1,-nbitq), 
to_sfixed(-1180.0/65536.0,1,-nbitq), 
to_sfixed(3186.0/65536.0,1,-nbitq), 
to_sfixed(1631.0/65536.0,1,-nbitq), 
to_sfixed(152.0/65536.0,1,-nbitq), 
to_sfixed(4506.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-421.0/65536.0,1,-nbitq), 
to_sfixed(-2894.0/65536.0,1,-nbitq), 
to_sfixed(3317.0/65536.0,1,-nbitq), 
to_sfixed(56.0/65536.0,1,-nbitq), 
to_sfixed(-91.0/65536.0,1,-nbitq), 
to_sfixed(-4660.0/65536.0,1,-nbitq), 
to_sfixed(-108.0/65536.0,1,-nbitq), 
to_sfixed(-1930.0/65536.0,1,-nbitq), 
to_sfixed(321.0/65536.0,1,-nbitq), 
to_sfixed(-1601.0/65536.0,1,-nbitq), 
to_sfixed(-182.0/65536.0,1,-nbitq), 
to_sfixed(-129.0/65536.0,1,-nbitq), 
to_sfixed(-2700.0/65536.0,1,-nbitq), 
to_sfixed(282.0/65536.0,1,-nbitq), 
to_sfixed(3023.0/65536.0,1,-nbitq), 
to_sfixed(3217.0/65536.0,1,-nbitq), 
to_sfixed(1064.0/65536.0,1,-nbitq), 
to_sfixed(4698.0/65536.0,1,-nbitq), 
to_sfixed(2207.0/65536.0,1,-nbitq), 
to_sfixed(1644.0/65536.0,1,-nbitq), 
to_sfixed(-1880.0/65536.0,1,-nbitq), 
to_sfixed(-1073.0/65536.0,1,-nbitq), 
to_sfixed(2199.0/65536.0,1,-nbitq), 
to_sfixed(3266.0/65536.0,1,-nbitq), 
to_sfixed(-3345.0/65536.0,1,-nbitq), 
to_sfixed(1905.0/65536.0,1,-nbitq), 
to_sfixed(-3435.0/65536.0,1,-nbitq), 
to_sfixed(-1196.0/65536.0,1,-nbitq), 
to_sfixed(-3070.0/65536.0,1,-nbitq), 
to_sfixed(43.0/65536.0,1,-nbitq), 
to_sfixed(1217.0/65536.0,1,-nbitq), 
to_sfixed(-1910.0/65536.0,1,-nbitq), 
to_sfixed(-5180.0/65536.0,1,-nbitq), 
to_sfixed(-5409.0/65536.0,1,-nbitq), 
to_sfixed(-708.0/65536.0,1,-nbitq), 
to_sfixed(1360.0/65536.0,1,-nbitq), 
to_sfixed(2269.0/65536.0,1,-nbitq), 
to_sfixed(697.0/65536.0,1,-nbitq), 
to_sfixed(-3430.0/65536.0,1,-nbitq), 
to_sfixed(1633.0/65536.0,1,-nbitq), 
to_sfixed(1265.0/65536.0,1,-nbitq), 
to_sfixed(-191.0/65536.0,1,-nbitq), 
to_sfixed(-4741.0/65536.0,1,-nbitq), 
to_sfixed(206.0/65536.0,1,-nbitq), 
to_sfixed(1506.0/65536.0,1,-nbitq), 
to_sfixed(6345.0/65536.0,1,-nbitq), 
to_sfixed(1910.0/65536.0,1,-nbitq), 
to_sfixed(-222.0/65536.0,1,-nbitq), 
to_sfixed(2842.0/65536.0,1,-nbitq), 
to_sfixed(1120.0/65536.0,1,-nbitq), 
to_sfixed(3095.0/65536.0,1,-nbitq), 
to_sfixed(-18.0/65536.0,1,-nbitq), 
to_sfixed(-2153.0/65536.0,1,-nbitq), 
to_sfixed(3501.0/65536.0,1,-nbitq), 
to_sfixed(3666.0/65536.0,1,-nbitq), 
to_sfixed(-425.0/65536.0,1,-nbitq), 
to_sfixed(3046.0/65536.0,1,-nbitq), 
to_sfixed(-2197.0/65536.0,1,-nbitq), 
to_sfixed(-541.0/65536.0,1,-nbitq), 
to_sfixed(-488.0/65536.0,1,-nbitq), 
to_sfixed(-1010.0/65536.0,1,-nbitq), 
to_sfixed(-2651.0/65536.0,1,-nbitq), 
to_sfixed(-2684.0/65536.0,1,-nbitq), 
to_sfixed(-23.0/65536.0,1,-nbitq), 
to_sfixed(387.0/65536.0,1,-nbitq), 
to_sfixed(-550.0/65536.0,1,-nbitq), 
to_sfixed(-2152.0/65536.0,1,-nbitq), 
to_sfixed(-4325.0/65536.0,1,-nbitq), 
to_sfixed(2690.0/65536.0,1,-nbitq), 
to_sfixed(1659.0/65536.0,1,-nbitq), 
to_sfixed(-1127.0/65536.0,1,-nbitq), 
to_sfixed(-1818.0/65536.0,1,-nbitq), 
to_sfixed(-1378.0/65536.0,1,-nbitq), 
to_sfixed(2069.0/65536.0,1,-nbitq), 
to_sfixed(-724.0/65536.0,1,-nbitq), 
to_sfixed(1754.0/65536.0,1,-nbitq), 
to_sfixed(2105.0/65536.0,1,-nbitq), 
to_sfixed(30.0/65536.0,1,-nbitq), 
to_sfixed(-1089.0/65536.0,1,-nbitq), 
to_sfixed(3636.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1266.0/65536.0,1,-nbitq), 
to_sfixed(533.0/65536.0,1,-nbitq), 
to_sfixed(-358.0/65536.0,1,-nbitq), 
to_sfixed(-1434.0/65536.0,1,-nbitq), 
to_sfixed(-1732.0/65536.0,1,-nbitq), 
to_sfixed(-3035.0/65536.0,1,-nbitq), 
to_sfixed(-148.0/65536.0,1,-nbitq), 
to_sfixed(-4656.0/65536.0,1,-nbitq), 
to_sfixed(-3145.0/65536.0,1,-nbitq), 
to_sfixed(-2839.0/65536.0,1,-nbitq), 
to_sfixed(-2238.0/65536.0,1,-nbitq), 
to_sfixed(2746.0/65536.0,1,-nbitq), 
to_sfixed(1175.0/65536.0,1,-nbitq), 
to_sfixed(-3707.0/65536.0,1,-nbitq), 
to_sfixed(2590.0/65536.0,1,-nbitq), 
to_sfixed(198.0/65536.0,1,-nbitq), 
to_sfixed(-161.0/65536.0,1,-nbitq), 
to_sfixed(-1031.0/65536.0,1,-nbitq), 
to_sfixed(-730.0/65536.0,1,-nbitq), 
to_sfixed(294.0/65536.0,1,-nbitq), 
to_sfixed(-3071.0/65536.0,1,-nbitq), 
to_sfixed(1406.0/65536.0,1,-nbitq), 
to_sfixed(6601.0/65536.0,1,-nbitq), 
to_sfixed(3920.0/65536.0,1,-nbitq), 
to_sfixed(237.0/65536.0,1,-nbitq), 
to_sfixed(2296.0/65536.0,1,-nbitq), 
to_sfixed(-2736.0/65536.0,1,-nbitq), 
to_sfixed(158.0/65536.0,1,-nbitq), 
to_sfixed(-815.0/65536.0,1,-nbitq), 
to_sfixed(1867.0/65536.0,1,-nbitq), 
to_sfixed(-3279.0/65536.0,1,-nbitq), 
to_sfixed(1036.0/65536.0,1,-nbitq), 
to_sfixed(-5375.0/65536.0,1,-nbitq), 
to_sfixed(-4461.0/65536.0,1,-nbitq), 
to_sfixed(71.0/65536.0,1,-nbitq), 
to_sfixed(-2107.0/65536.0,1,-nbitq), 
to_sfixed(1192.0/65536.0,1,-nbitq), 
to_sfixed(-2518.0/65536.0,1,-nbitq), 
to_sfixed(1591.0/65536.0,1,-nbitq), 
to_sfixed(857.0/65536.0,1,-nbitq), 
to_sfixed(334.0/65536.0,1,-nbitq), 
to_sfixed(-719.0/65536.0,1,-nbitq), 
to_sfixed(-4277.0/65536.0,1,-nbitq), 
to_sfixed(1747.0/65536.0,1,-nbitq), 
to_sfixed(1726.0/65536.0,1,-nbitq), 
to_sfixed(7322.0/65536.0,1,-nbitq), 
to_sfixed(843.0/65536.0,1,-nbitq), 
to_sfixed(-3348.0/65536.0,1,-nbitq), 
to_sfixed(887.0/65536.0,1,-nbitq), 
to_sfixed(-386.0/65536.0,1,-nbitq), 
to_sfixed(-1747.0/65536.0,1,-nbitq), 
to_sfixed(-2828.0/65536.0,1,-nbitq), 
to_sfixed(1695.0/65536.0,1,-nbitq), 
to_sfixed(-664.0/65536.0,1,-nbitq), 
to_sfixed(-263.0/65536.0,1,-nbitq), 
to_sfixed(-115.0/65536.0,1,-nbitq), 
to_sfixed(2089.0/65536.0,1,-nbitq), 
to_sfixed(-743.0/65536.0,1,-nbitq), 
to_sfixed(1784.0/65536.0,1,-nbitq), 
to_sfixed(1417.0/65536.0,1,-nbitq), 
to_sfixed(1232.0/65536.0,1,-nbitq), 
to_sfixed(2343.0/65536.0,1,-nbitq), 
to_sfixed(-746.0/65536.0,1,-nbitq), 
to_sfixed(-134.0/65536.0,1,-nbitq), 
to_sfixed(3351.0/65536.0,1,-nbitq), 
to_sfixed(-1404.0/65536.0,1,-nbitq), 
to_sfixed(-1343.0/65536.0,1,-nbitq), 
to_sfixed(1644.0/65536.0,1,-nbitq), 
to_sfixed(1898.0/65536.0,1,-nbitq), 
to_sfixed(2506.0/65536.0,1,-nbitq), 
to_sfixed(-747.0/65536.0,1,-nbitq), 
to_sfixed(-838.0/65536.0,1,-nbitq), 
to_sfixed(-994.0/65536.0,1,-nbitq), 
to_sfixed(1668.0/65536.0,1,-nbitq), 
to_sfixed(-879.0/65536.0,1,-nbitq), 
to_sfixed(3187.0/65536.0,1,-nbitq), 
to_sfixed(-12.0/65536.0,1,-nbitq), 
to_sfixed(3106.0/65536.0,1,-nbitq), 
to_sfixed(-1294.0/65536.0,1,-nbitq), 
to_sfixed(812.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1152.0/65536.0,1,-nbitq), 
to_sfixed(715.0/65536.0,1,-nbitq), 
to_sfixed(26.0/65536.0,1,-nbitq), 
to_sfixed(-1240.0/65536.0,1,-nbitq), 
to_sfixed(543.0/65536.0,1,-nbitq), 
to_sfixed(-1809.0/65536.0,1,-nbitq), 
to_sfixed(2060.0/65536.0,1,-nbitq), 
to_sfixed(1055.0/65536.0,1,-nbitq), 
to_sfixed(1315.0/65536.0,1,-nbitq), 
to_sfixed(2354.0/65536.0,1,-nbitq), 
to_sfixed(-525.0/65536.0,1,-nbitq), 
to_sfixed(5007.0/65536.0,1,-nbitq), 
to_sfixed(907.0/65536.0,1,-nbitq), 
to_sfixed(-2928.0/65536.0,1,-nbitq), 
to_sfixed(1554.0/65536.0,1,-nbitq), 
to_sfixed(1900.0/65536.0,1,-nbitq), 
to_sfixed(-931.0/65536.0,1,-nbitq), 
to_sfixed(-192.0/65536.0,1,-nbitq), 
to_sfixed(1624.0/65536.0,1,-nbitq), 
to_sfixed(-1204.0/65536.0,1,-nbitq), 
to_sfixed(-273.0/65536.0,1,-nbitq), 
to_sfixed(-1592.0/65536.0,1,-nbitq), 
to_sfixed(1648.0/65536.0,1,-nbitq), 
to_sfixed(-539.0/65536.0,1,-nbitq), 
to_sfixed(904.0/65536.0,1,-nbitq), 
to_sfixed(1216.0/65536.0,1,-nbitq), 
to_sfixed(-3096.0/65536.0,1,-nbitq), 
to_sfixed(-1589.0/65536.0,1,-nbitq), 
to_sfixed(-2791.0/65536.0,1,-nbitq), 
to_sfixed(498.0/65536.0,1,-nbitq), 
to_sfixed(-3431.0/65536.0,1,-nbitq), 
to_sfixed(-2289.0/65536.0,1,-nbitq), 
to_sfixed(-3693.0/65536.0,1,-nbitq), 
to_sfixed(-1015.0/65536.0,1,-nbitq), 
to_sfixed(687.0/65536.0,1,-nbitq), 
to_sfixed(181.0/65536.0,1,-nbitq), 
to_sfixed(500.0/65536.0,1,-nbitq), 
to_sfixed(-404.0/65536.0,1,-nbitq), 
to_sfixed(973.0/65536.0,1,-nbitq), 
to_sfixed(333.0/65536.0,1,-nbitq), 
to_sfixed(-2490.0/65536.0,1,-nbitq), 
to_sfixed(-882.0/65536.0,1,-nbitq), 
to_sfixed(-3013.0/65536.0,1,-nbitq), 
to_sfixed(-2152.0/65536.0,1,-nbitq), 
to_sfixed(-623.0/65536.0,1,-nbitq), 
to_sfixed(8607.0/65536.0,1,-nbitq), 
to_sfixed(86.0/65536.0,1,-nbitq), 
to_sfixed(1090.0/65536.0,1,-nbitq), 
to_sfixed(349.0/65536.0,1,-nbitq), 
to_sfixed(1525.0/65536.0,1,-nbitq), 
to_sfixed(1868.0/65536.0,1,-nbitq), 
to_sfixed(-1620.0/65536.0,1,-nbitq), 
to_sfixed(-667.0/65536.0,1,-nbitq), 
to_sfixed(-1744.0/65536.0,1,-nbitq), 
to_sfixed(1072.0/65536.0,1,-nbitq), 
to_sfixed(-1489.0/65536.0,1,-nbitq), 
to_sfixed(679.0/65536.0,1,-nbitq), 
to_sfixed(-1273.0/65536.0,1,-nbitq), 
to_sfixed(-1284.0/65536.0,1,-nbitq), 
to_sfixed(2726.0/65536.0,1,-nbitq), 
to_sfixed(530.0/65536.0,1,-nbitq), 
to_sfixed(-2735.0/65536.0,1,-nbitq), 
to_sfixed(3175.0/65536.0,1,-nbitq), 
to_sfixed(459.0/65536.0,1,-nbitq), 
to_sfixed(3533.0/65536.0,1,-nbitq), 
to_sfixed(3270.0/65536.0,1,-nbitq), 
to_sfixed(573.0/65536.0,1,-nbitq), 
to_sfixed(923.0/65536.0,1,-nbitq), 
to_sfixed(4400.0/65536.0,1,-nbitq), 
to_sfixed(527.0/65536.0,1,-nbitq), 
to_sfixed(-419.0/65536.0,1,-nbitq), 
to_sfixed(-1886.0/65536.0,1,-nbitq), 
to_sfixed(-114.0/65536.0,1,-nbitq), 
to_sfixed(-3017.0/65536.0,1,-nbitq), 
to_sfixed(-2747.0/65536.0,1,-nbitq), 
to_sfixed(2266.0/65536.0,1,-nbitq), 
to_sfixed(1294.0/65536.0,1,-nbitq), 
to_sfixed(3174.0/65536.0,1,-nbitq), 
to_sfixed(924.0/65536.0,1,-nbitq), 
to_sfixed(4603.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2707.0/65536.0,1,-nbitq), 
to_sfixed(525.0/65536.0,1,-nbitq), 
to_sfixed(-656.0/65536.0,1,-nbitq), 
to_sfixed(-5400.0/65536.0,1,-nbitq), 
to_sfixed(-2667.0/65536.0,1,-nbitq), 
to_sfixed(-2180.0/65536.0,1,-nbitq), 
to_sfixed(377.0/65536.0,1,-nbitq), 
to_sfixed(546.0/65536.0,1,-nbitq), 
to_sfixed(-2716.0/65536.0,1,-nbitq), 
to_sfixed(1667.0/65536.0,1,-nbitq), 
to_sfixed(-971.0/65536.0,1,-nbitq), 
to_sfixed(4580.0/65536.0,1,-nbitq), 
to_sfixed(-621.0/65536.0,1,-nbitq), 
to_sfixed(-4164.0/65536.0,1,-nbitq), 
to_sfixed(-3252.0/65536.0,1,-nbitq), 
to_sfixed(580.0/65536.0,1,-nbitq), 
to_sfixed(1566.0/65536.0,1,-nbitq), 
to_sfixed(1564.0/65536.0,1,-nbitq), 
to_sfixed(3379.0/65536.0,1,-nbitq), 
to_sfixed(-668.0/65536.0,1,-nbitq), 
to_sfixed(1738.0/65536.0,1,-nbitq), 
to_sfixed(1539.0/65536.0,1,-nbitq), 
to_sfixed(1619.0/65536.0,1,-nbitq), 
to_sfixed(-1838.0/65536.0,1,-nbitq), 
to_sfixed(-2115.0/65536.0,1,-nbitq), 
to_sfixed(-1913.0/65536.0,1,-nbitq), 
to_sfixed(620.0/65536.0,1,-nbitq), 
to_sfixed(-1869.0/65536.0,1,-nbitq), 
to_sfixed(-1396.0/65536.0,1,-nbitq), 
to_sfixed(2017.0/65536.0,1,-nbitq), 
to_sfixed(-2595.0/65536.0,1,-nbitq), 
to_sfixed(-1720.0/65536.0,1,-nbitq), 
to_sfixed(-3167.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(1078.0/65536.0,1,-nbitq), 
to_sfixed(50.0/65536.0,1,-nbitq), 
to_sfixed(1877.0/65536.0,1,-nbitq), 
to_sfixed(-2194.0/65536.0,1,-nbitq), 
to_sfixed(4861.0/65536.0,1,-nbitq), 
to_sfixed(-557.0/65536.0,1,-nbitq), 
to_sfixed(-643.0/65536.0,1,-nbitq), 
to_sfixed(2528.0/65536.0,1,-nbitq), 
to_sfixed(-1052.0/65536.0,1,-nbitq), 
to_sfixed(507.0/65536.0,1,-nbitq), 
to_sfixed(1346.0/65536.0,1,-nbitq), 
to_sfixed(810.0/65536.0,1,-nbitq), 
to_sfixed(-270.0/65536.0,1,-nbitq), 
to_sfixed(-3733.0/65536.0,1,-nbitq), 
to_sfixed(1028.0/65536.0,1,-nbitq), 
to_sfixed(-943.0/65536.0,1,-nbitq), 
to_sfixed(-1680.0/65536.0,1,-nbitq), 
to_sfixed(36.0/65536.0,1,-nbitq), 
to_sfixed(-1138.0/65536.0,1,-nbitq), 
to_sfixed(-853.0/65536.0,1,-nbitq), 
to_sfixed(645.0/65536.0,1,-nbitq), 
to_sfixed(-3541.0/65536.0,1,-nbitq), 
to_sfixed(2960.0/65536.0,1,-nbitq), 
to_sfixed(3453.0/65536.0,1,-nbitq), 
to_sfixed(-125.0/65536.0,1,-nbitq), 
to_sfixed(-1843.0/65536.0,1,-nbitq), 
to_sfixed(1761.0/65536.0,1,-nbitq), 
to_sfixed(-2130.0/65536.0,1,-nbitq), 
to_sfixed(-1632.0/65536.0,1,-nbitq), 
to_sfixed(-563.0/65536.0,1,-nbitq), 
to_sfixed(3564.0/65536.0,1,-nbitq), 
to_sfixed(2496.0/65536.0,1,-nbitq), 
to_sfixed(5529.0/65536.0,1,-nbitq), 
to_sfixed(-1223.0/65536.0,1,-nbitq), 
to_sfixed(4160.0/65536.0,1,-nbitq), 
to_sfixed(3757.0/65536.0,1,-nbitq), 
to_sfixed(33.0/65536.0,1,-nbitq), 
to_sfixed(-4021.0/65536.0,1,-nbitq), 
to_sfixed(-2601.0/65536.0,1,-nbitq), 
to_sfixed(2000.0/65536.0,1,-nbitq), 
to_sfixed(477.0/65536.0,1,-nbitq), 
to_sfixed(503.0/65536.0,1,-nbitq), 
to_sfixed(1676.0/65536.0,1,-nbitq), 
to_sfixed(2878.0/65536.0,1,-nbitq), 
to_sfixed(1862.0/65536.0,1,-nbitq), 
to_sfixed(854.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1549.0/65536.0,1,-nbitq), 
to_sfixed(635.0/65536.0,1,-nbitq), 
to_sfixed(-978.0/65536.0,1,-nbitq), 
to_sfixed(-4543.0/65536.0,1,-nbitq), 
to_sfixed(-3125.0/65536.0,1,-nbitq), 
to_sfixed(-3765.0/65536.0,1,-nbitq), 
to_sfixed(761.0/65536.0,1,-nbitq), 
to_sfixed(2270.0/65536.0,1,-nbitq), 
to_sfixed(-2459.0/65536.0,1,-nbitq), 
to_sfixed(1186.0/65536.0,1,-nbitq), 
to_sfixed(161.0/65536.0,1,-nbitq), 
to_sfixed(6236.0/65536.0,1,-nbitq), 
to_sfixed(2450.0/65536.0,1,-nbitq), 
to_sfixed(-4106.0/65536.0,1,-nbitq), 
to_sfixed(-44.0/65536.0,1,-nbitq), 
to_sfixed(881.0/65536.0,1,-nbitq), 
to_sfixed(-1128.0/65536.0,1,-nbitq), 
to_sfixed(3337.0/65536.0,1,-nbitq), 
to_sfixed(-1895.0/65536.0,1,-nbitq), 
to_sfixed(-580.0/65536.0,1,-nbitq), 
to_sfixed(-1255.0/65536.0,1,-nbitq), 
to_sfixed(3363.0/65536.0,1,-nbitq), 
to_sfixed(4182.0/65536.0,1,-nbitq), 
to_sfixed(-981.0/65536.0,1,-nbitq), 
to_sfixed(1900.0/65536.0,1,-nbitq), 
to_sfixed(-2855.0/65536.0,1,-nbitq), 
to_sfixed(-1488.0/65536.0,1,-nbitq), 
to_sfixed(874.0/65536.0,1,-nbitq), 
to_sfixed(-3229.0/65536.0,1,-nbitq), 
to_sfixed(-1389.0/65536.0,1,-nbitq), 
to_sfixed(-2659.0/65536.0,1,-nbitq), 
to_sfixed(-1852.0/65536.0,1,-nbitq), 
to_sfixed(-4560.0/65536.0,1,-nbitq), 
to_sfixed(-3035.0/65536.0,1,-nbitq), 
to_sfixed(1095.0/65536.0,1,-nbitq), 
to_sfixed(-2899.0/65536.0,1,-nbitq), 
to_sfixed(-1859.0/65536.0,1,-nbitq), 
to_sfixed(1582.0/65536.0,1,-nbitq), 
to_sfixed(5464.0/65536.0,1,-nbitq), 
to_sfixed(647.0/65536.0,1,-nbitq), 
to_sfixed(-4200.0/65536.0,1,-nbitq), 
to_sfixed(2003.0/65536.0,1,-nbitq), 
to_sfixed(-450.0/65536.0,1,-nbitq), 
to_sfixed(-90.0/65536.0,1,-nbitq), 
to_sfixed(1055.0/65536.0,1,-nbitq), 
to_sfixed(4360.0/65536.0,1,-nbitq), 
to_sfixed(-3579.0/65536.0,1,-nbitq), 
to_sfixed(116.0/65536.0,1,-nbitq), 
to_sfixed(1819.0/65536.0,1,-nbitq), 
to_sfixed(4003.0/65536.0,1,-nbitq), 
to_sfixed(1716.0/65536.0,1,-nbitq), 
to_sfixed(-5003.0/65536.0,1,-nbitq), 
to_sfixed(-2072.0/65536.0,1,-nbitq), 
to_sfixed(1466.0/65536.0,1,-nbitq), 
to_sfixed(827.0/65536.0,1,-nbitq), 
to_sfixed(-5051.0/65536.0,1,-nbitq), 
to_sfixed(364.0/65536.0,1,-nbitq), 
to_sfixed(1641.0/65536.0,1,-nbitq), 
to_sfixed(1857.0/65536.0,1,-nbitq), 
to_sfixed(-4170.0/65536.0,1,-nbitq), 
to_sfixed(-2781.0/65536.0,1,-nbitq), 
to_sfixed(2675.0/65536.0,1,-nbitq), 
to_sfixed(-2632.0/65536.0,1,-nbitq), 
to_sfixed(-1958.0/65536.0,1,-nbitq), 
to_sfixed(3105.0/65536.0,1,-nbitq), 
to_sfixed(572.0/65536.0,1,-nbitq), 
to_sfixed(1548.0/65536.0,1,-nbitq), 
to_sfixed(-798.0/65536.0,1,-nbitq), 
to_sfixed(3628.0/65536.0,1,-nbitq), 
to_sfixed(8761.0/65536.0,1,-nbitq), 
to_sfixed(2882.0/65536.0,1,-nbitq), 
to_sfixed(-3771.0/65536.0,1,-nbitq), 
to_sfixed(-1274.0/65536.0,1,-nbitq), 
to_sfixed(-2689.0/65536.0,1,-nbitq), 
to_sfixed(-1984.0/65536.0,1,-nbitq), 
to_sfixed(-1440.0/65536.0,1,-nbitq), 
to_sfixed(2181.0/65536.0,1,-nbitq), 
to_sfixed(862.0/65536.0,1,-nbitq), 
to_sfixed(799.0/65536.0,1,-nbitq), 
to_sfixed(-994.0/65536.0,1,-nbitq)  ), 
( to_sfixed(700.0/65536.0,1,-nbitq), 
to_sfixed(3341.0/65536.0,1,-nbitq), 
to_sfixed(-4091.0/65536.0,1,-nbitq), 
to_sfixed(-4785.0/65536.0,1,-nbitq), 
to_sfixed(1756.0/65536.0,1,-nbitq), 
to_sfixed(-1354.0/65536.0,1,-nbitq), 
to_sfixed(-1739.0/65536.0,1,-nbitq), 
to_sfixed(447.0/65536.0,1,-nbitq), 
to_sfixed(1171.0/65536.0,1,-nbitq), 
to_sfixed(-2746.0/65536.0,1,-nbitq), 
to_sfixed(182.0/65536.0,1,-nbitq), 
to_sfixed(4099.0/65536.0,1,-nbitq), 
to_sfixed(-2181.0/65536.0,1,-nbitq), 
to_sfixed(731.0/65536.0,1,-nbitq), 
to_sfixed(1257.0/65536.0,1,-nbitq), 
to_sfixed(2280.0/65536.0,1,-nbitq), 
to_sfixed(2107.0/65536.0,1,-nbitq), 
to_sfixed(2441.0/65536.0,1,-nbitq), 
to_sfixed(230.0/65536.0,1,-nbitq), 
to_sfixed(456.0/65536.0,1,-nbitq), 
to_sfixed(142.0/65536.0,1,-nbitq), 
to_sfixed(601.0/65536.0,1,-nbitq), 
to_sfixed(4264.0/65536.0,1,-nbitq), 
to_sfixed(259.0/65536.0,1,-nbitq), 
to_sfixed(3023.0/65536.0,1,-nbitq), 
to_sfixed(-4438.0/65536.0,1,-nbitq), 
to_sfixed(-1535.0/65536.0,1,-nbitq), 
to_sfixed(-1937.0/65536.0,1,-nbitq), 
to_sfixed(2308.0/65536.0,1,-nbitq), 
to_sfixed(-1484.0/65536.0,1,-nbitq), 
to_sfixed(1719.0/65536.0,1,-nbitq), 
to_sfixed(-1636.0/65536.0,1,-nbitq), 
to_sfixed(641.0/65536.0,1,-nbitq), 
to_sfixed(838.0/65536.0,1,-nbitq), 
to_sfixed(-3099.0/65536.0,1,-nbitq), 
to_sfixed(2431.0/65536.0,1,-nbitq), 
to_sfixed(-648.0/65536.0,1,-nbitq), 
to_sfixed(843.0/65536.0,1,-nbitq), 
to_sfixed(2381.0/65536.0,1,-nbitq), 
to_sfixed(-3168.0/65536.0,1,-nbitq), 
to_sfixed(-3520.0/65536.0,1,-nbitq), 
to_sfixed(133.0/65536.0,1,-nbitq), 
to_sfixed(616.0/65536.0,1,-nbitq), 
to_sfixed(-1032.0/65536.0,1,-nbitq), 
to_sfixed(-561.0/65536.0,1,-nbitq), 
to_sfixed(230.0/65536.0,1,-nbitq), 
to_sfixed(-595.0/65536.0,1,-nbitq), 
to_sfixed(-4610.0/65536.0,1,-nbitq), 
to_sfixed(1154.0/65536.0,1,-nbitq), 
to_sfixed(-627.0/65536.0,1,-nbitq), 
to_sfixed(-1454.0/65536.0,1,-nbitq), 
to_sfixed(-3721.0/65536.0,1,-nbitq), 
to_sfixed(-4881.0/65536.0,1,-nbitq), 
to_sfixed(-3559.0/65536.0,1,-nbitq), 
to_sfixed(4703.0/65536.0,1,-nbitq), 
to_sfixed(-2250.0/65536.0,1,-nbitq), 
to_sfixed(2162.0/65536.0,1,-nbitq), 
to_sfixed(-1135.0/65536.0,1,-nbitq), 
to_sfixed(1881.0/65536.0,1,-nbitq), 
to_sfixed(-2949.0/65536.0,1,-nbitq), 
to_sfixed(325.0/65536.0,1,-nbitq), 
to_sfixed(-1033.0/65536.0,1,-nbitq), 
to_sfixed(-2793.0/65536.0,1,-nbitq), 
to_sfixed(2345.0/65536.0,1,-nbitq), 
to_sfixed(3278.0/65536.0,1,-nbitq), 
to_sfixed(-1259.0/65536.0,1,-nbitq), 
to_sfixed(3994.0/65536.0,1,-nbitq), 
to_sfixed(2630.0/65536.0,1,-nbitq), 
to_sfixed(334.0/65536.0,1,-nbitq), 
to_sfixed(7578.0/65536.0,1,-nbitq), 
to_sfixed(-2435.0/65536.0,1,-nbitq), 
to_sfixed(-3015.0/65536.0,1,-nbitq), 
to_sfixed(-1676.0/65536.0,1,-nbitq), 
to_sfixed(-491.0/65536.0,1,-nbitq), 
to_sfixed(2358.0/65536.0,1,-nbitq), 
to_sfixed(882.0/65536.0,1,-nbitq), 
to_sfixed(-507.0/65536.0,1,-nbitq), 
to_sfixed(3637.0/65536.0,1,-nbitq), 
to_sfixed(-3144.0/65536.0,1,-nbitq), 
to_sfixed(1749.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1827.0/65536.0,1,-nbitq), 
to_sfixed(1164.0/65536.0,1,-nbitq), 
to_sfixed(-3086.0/65536.0,1,-nbitq), 
to_sfixed(-1787.0/65536.0,1,-nbitq), 
to_sfixed(3381.0/65536.0,1,-nbitq), 
to_sfixed(-3539.0/65536.0,1,-nbitq), 
to_sfixed(963.0/65536.0,1,-nbitq), 
to_sfixed(-2389.0/65536.0,1,-nbitq), 
to_sfixed(1997.0/65536.0,1,-nbitq), 
to_sfixed(2399.0/65536.0,1,-nbitq), 
to_sfixed(-1921.0/65536.0,1,-nbitq), 
to_sfixed(3065.0/65536.0,1,-nbitq), 
to_sfixed(1303.0/65536.0,1,-nbitq), 
to_sfixed(-3886.0/65536.0,1,-nbitq), 
to_sfixed(400.0/65536.0,1,-nbitq), 
to_sfixed(-2130.0/65536.0,1,-nbitq), 
to_sfixed(-956.0/65536.0,1,-nbitq), 
to_sfixed(-2280.0/65536.0,1,-nbitq), 
to_sfixed(-1430.0/65536.0,1,-nbitq), 
to_sfixed(-2110.0/65536.0,1,-nbitq), 
to_sfixed(262.0/65536.0,1,-nbitq), 
to_sfixed(2478.0/65536.0,1,-nbitq), 
to_sfixed(3230.0/65536.0,1,-nbitq), 
to_sfixed(-1336.0/65536.0,1,-nbitq), 
to_sfixed(3285.0/65536.0,1,-nbitq), 
to_sfixed(-3575.0/65536.0,1,-nbitq), 
to_sfixed(-3750.0/65536.0,1,-nbitq), 
to_sfixed(-210.0/65536.0,1,-nbitq), 
to_sfixed(-1034.0/65536.0,1,-nbitq), 
to_sfixed(544.0/65536.0,1,-nbitq), 
to_sfixed(-3157.0/65536.0,1,-nbitq), 
to_sfixed(-2106.0/65536.0,1,-nbitq), 
to_sfixed(-4030.0/65536.0,1,-nbitq), 
to_sfixed(-3214.0/65536.0,1,-nbitq), 
to_sfixed(-2009.0/65536.0,1,-nbitq), 
to_sfixed(1508.0/65536.0,1,-nbitq), 
to_sfixed(299.0/65536.0,1,-nbitq), 
to_sfixed(-319.0/65536.0,1,-nbitq), 
to_sfixed(3058.0/65536.0,1,-nbitq), 
to_sfixed(-758.0/65536.0,1,-nbitq), 
to_sfixed(203.0/65536.0,1,-nbitq), 
to_sfixed(-128.0/65536.0,1,-nbitq), 
to_sfixed(1711.0/65536.0,1,-nbitq), 
to_sfixed(-3833.0/65536.0,1,-nbitq), 
to_sfixed(2042.0/65536.0,1,-nbitq), 
to_sfixed(791.0/65536.0,1,-nbitq), 
to_sfixed(-920.0/65536.0,1,-nbitq), 
to_sfixed(-524.0/65536.0,1,-nbitq), 
to_sfixed(2442.0/65536.0,1,-nbitq), 
to_sfixed(3877.0/65536.0,1,-nbitq), 
to_sfixed(-2509.0/65536.0,1,-nbitq), 
to_sfixed(760.0/65536.0,1,-nbitq), 
to_sfixed(-1412.0/65536.0,1,-nbitq), 
to_sfixed(-2624.0/65536.0,1,-nbitq), 
to_sfixed(761.0/65536.0,1,-nbitq), 
to_sfixed(-645.0/65536.0,1,-nbitq), 
to_sfixed(-1843.0/65536.0,1,-nbitq), 
to_sfixed(387.0/65536.0,1,-nbitq), 
to_sfixed(2692.0/65536.0,1,-nbitq), 
to_sfixed(-2353.0/65536.0,1,-nbitq), 
to_sfixed(391.0/65536.0,1,-nbitq), 
to_sfixed(374.0/65536.0,1,-nbitq), 
to_sfixed(1002.0/65536.0,1,-nbitq), 
to_sfixed(-1434.0/65536.0,1,-nbitq), 
to_sfixed(-1974.0/65536.0,1,-nbitq), 
to_sfixed(-1138.0/65536.0,1,-nbitq), 
to_sfixed(5589.0/65536.0,1,-nbitq), 
to_sfixed(789.0/65536.0,1,-nbitq), 
to_sfixed(714.0/65536.0,1,-nbitq), 
to_sfixed(3124.0/65536.0,1,-nbitq), 
to_sfixed(-1822.0/65536.0,1,-nbitq), 
to_sfixed(-3291.0/65536.0,1,-nbitq), 
to_sfixed(-363.0/65536.0,1,-nbitq), 
to_sfixed(1904.0/65536.0,1,-nbitq), 
to_sfixed(-2085.0/65536.0,1,-nbitq), 
to_sfixed(3801.0/65536.0,1,-nbitq), 
to_sfixed(-514.0/65536.0,1,-nbitq), 
to_sfixed(875.0/65536.0,1,-nbitq), 
to_sfixed(-1581.0/65536.0,1,-nbitq), 
to_sfixed(-506.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2150.0/65536.0,1,-nbitq), 
to_sfixed(-1646.0/65536.0,1,-nbitq), 
to_sfixed(-292.0/65536.0,1,-nbitq), 
to_sfixed(1460.0/65536.0,1,-nbitq), 
to_sfixed(1555.0/65536.0,1,-nbitq), 
to_sfixed(-1853.0/65536.0,1,-nbitq), 
to_sfixed(-337.0/65536.0,1,-nbitq), 
to_sfixed(-299.0/65536.0,1,-nbitq), 
to_sfixed(484.0/65536.0,1,-nbitq), 
to_sfixed(-2768.0/65536.0,1,-nbitq), 
to_sfixed(-1974.0/65536.0,1,-nbitq), 
to_sfixed(7411.0/65536.0,1,-nbitq), 
to_sfixed(-2333.0/65536.0,1,-nbitq), 
to_sfixed(-1563.0/65536.0,1,-nbitq), 
to_sfixed(967.0/65536.0,1,-nbitq), 
to_sfixed(-2126.0/65536.0,1,-nbitq), 
to_sfixed(-3050.0/65536.0,1,-nbitq), 
to_sfixed(1712.0/65536.0,1,-nbitq), 
to_sfixed(1717.0/65536.0,1,-nbitq), 
to_sfixed(1406.0/65536.0,1,-nbitq), 
to_sfixed(1514.0/65536.0,1,-nbitq), 
to_sfixed(-217.0/65536.0,1,-nbitq), 
to_sfixed(1743.0/65536.0,1,-nbitq), 
to_sfixed(1401.0/65536.0,1,-nbitq), 
to_sfixed(3490.0/65536.0,1,-nbitq), 
to_sfixed(-2596.0/65536.0,1,-nbitq), 
to_sfixed(-2094.0/65536.0,1,-nbitq), 
to_sfixed(2679.0/65536.0,1,-nbitq), 
to_sfixed(2586.0/65536.0,1,-nbitq), 
to_sfixed(1286.0/65536.0,1,-nbitq), 
to_sfixed(-2612.0/65536.0,1,-nbitq), 
to_sfixed(1652.0/65536.0,1,-nbitq), 
to_sfixed(65.0/65536.0,1,-nbitq), 
to_sfixed(-3222.0/65536.0,1,-nbitq), 
to_sfixed(208.0/65536.0,1,-nbitq), 
to_sfixed(-1157.0/65536.0,1,-nbitq), 
to_sfixed(3307.0/65536.0,1,-nbitq), 
to_sfixed(3512.0/65536.0,1,-nbitq), 
to_sfixed(-66.0/65536.0,1,-nbitq), 
to_sfixed(-2319.0/65536.0,1,-nbitq), 
to_sfixed(-2194.0/65536.0,1,-nbitq), 
to_sfixed(-1119.0/65536.0,1,-nbitq), 
to_sfixed(-3890.0/65536.0,1,-nbitq), 
to_sfixed(946.0/65536.0,1,-nbitq), 
to_sfixed(-2147.0/65536.0,1,-nbitq), 
to_sfixed(1285.0/65536.0,1,-nbitq), 
to_sfixed(955.0/65536.0,1,-nbitq), 
to_sfixed(-3461.0/65536.0,1,-nbitq), 
to_sfixed(-1608.0/65536.0,1,-nbitq), 
to_sfixed(3068.0/65536.0,1,-nbitq), 
to_sfixed(-1503.0/65536.0,1,-nbitq), 
to_sfixed(2792.0/65536.0,1,-nbitq), 
to_sfixed(-2350.0/65536.0,1,-nbitq), 
to_sfixed(-2521.0/65536.0,1,-nbitq), 
to_sfixed(4096.0/65536.0,1,-nbitq), 
to_sfixed(-107.0/65536.0,1,-nbitq), 
to_sfixed(-1181.0/65536.0,1,-nbitq), 
to_sfixed(-2157.0/65536.0,1,-nbitq), 
to_sfixed(1393.0/65536.0,1,-nbitq), 
to_sfixed(-2890.0/65536.0,1,-nbitq), 
to_sfixed(1780.0/65536.0,1,-nbitq), 
to_sfixed(-419.0/65536.0,1,-nbitq), 
to_sfixed(1516.0/65536.0,1,-nbitq), 
to_sfixed(-2962.0/65536.0,1,-nbitq), 
to_sfixed(-2097.0/65536.0,1,-nbitq), 
to_sfixed(-1868.0/65536.0,1,-nbitq), 
to_sfixed(5897.0/65536.0,1,-nbitq), 
to_sfixed(3458.0/65536.0,1,-nbitq), 
to_sfixed(2527.0/65536.0,1,-nbitq), 
to_sfixed(5619.0/65536.0,1,-nbitq), 
to_sfixed(-1566.0/65536.0,1,-nbitq), 
to_sfixed(-1756.0/65536.0,1,-nbitq), 
to_sfixed(-3332.0/65536.0,1,-nbitq), 
to_sfixed(1326.0/65536.0,1,-nbitq), 
to_sfixed(-2772.0/65536.0,1,-nbitq), 
to_sfixed(934.0/65536.0,1,-nbitq), 
to_sfixed(-1944.0/65536.0,1,-nbitq), 
to_sfixed(3197.0/65536.0,1,-nbitq), 
to_sfixed(-1378.0/65536.0,1,-nbitq), 
to_sfixed(-1455.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3425.0/65536.0,1,-nbitq), 
to_sfixed(-2888.0/65536.0,1,-nbitq), 
to_sfixed(6814.0/65536.0,1,-nbitq), 
to_sfixed(1889.0/65536.0,1,-nbitq), 
to_sfixed(2828.0/65536.0,1,-nbitq), 
to_sfixed(2123.0/65536.0,1,-nbitq), 
to_sfixed(1740.0/65536.0,1,-nbitq), 
to_sfixed(-3131.0/65536.0,1,-nbitq), 
to_sfixed(75.0/65536.0,1,-nbitq), 
to_sfixed(-211.0/65536.0,1,-nbitq), 
to_sfixed(-2088.0/65536.0,1,-nbitq), 
to_sfixed(6476.0/65536.0,1,-nbitq), 
to_sfixed(-1467.0/65536.0,1,-nbitq), 
to_sfixed(3552.0/65536.0,1,-nbitq), 
to_sfixed(-1822.0/65536.0,1,-nbitq), 
to_sfixed(-1939.0/65536.0,1,-nbitq), 
to_sfixed(1241.0/65536.0,1,-nbitq), 
to_sfixed(-7295.0/65536.0,1,-nbitq), 
to_sfixed(-1038.0/65536.0,1,-nbitq), 
to_sfixed(-596.0/65536.0,1,-nbitq), 
to_sfixed(-1807.0/65536.0,1,-nbitq), 
to_sfixed(-1135.0/65536.0,1,-nbitq), 
to_sfixed(-4436.0/65536.0,1,-nbitq), 
to_sfixed(3254.0/65536.0,1,-nbitq), 
to_sfixed(746.0/65536.0,1,-nbitq), 
to_sfixed(3872.0/65536.0,1,-nbitq), 
to_sfixed(-1917.0/65536.0,1,-nbitq), 
to_sfixed(325.0/65536.0,1,-nbitq), 
to_sfixed(2440.0/65536.0,1,-nbitq), 
to_sfixed(3250.0/65536.0,1,-nbitq), 
to_sfixed(-3215.0/65536.0,1,-nbitq), 
to_sfixed(1124.0/65536.0,1,-nbitq), 
to_sfixed(972.0/65536.0,1,-nbitq), 
to_sfixed(-2294.0/65536.0,1,-nbitq), 
to_sfixed(700.0/65536.0,1,-nbitq), 
to_sfixed(-1393.0/65536.0,1,-nbitq), 
to_sfixed(1457.0/65536.0,1,-nbitq), 
to_sfixed(1114.0/65536.0,1,-nbitq), 
to_sfixed(4852.0/65536.0,1,-nbitq), 
to_sfixed(3099.0/65536.0,1,-nbitq), 
to_sfixed(1132.0/65536.0,1,-nbitq), 
to_sfixed(1986.0/65536.0,1,-nbitq), 
to_sfixed(-3451.0/65536.0,1,-nbitq), 
to_sfixed(-1718.0/65536.0,1,-nbitq), 
to_sfixed(-244.0/65536.0,1,-nbitq), 
to_sfixed(3596.0/65536.0,1,-nbitq), 
to_sfixed(-2091.0/65536.0,1,-nbitq), 
to_sfixed(-1614.0/65536.0,1,-nbitq), 
to_sfixed(2871.0/65536.0,1,-nbitq), 
to_sfixed(2313.0/65536.0,1,-nbitq), 
to_sfixed(2105.0/65536.0,1,-nbitq), 
to_sfixed(654.0/65536.0,1,-nbitq), 
to_sfixed(2751.0/65536.0,1,-nbitq), 
to_sfixed(-2607.0/65536.0,1,-nbitq), 
to_sfixed(-1872.0/65536.0,1,-nbitq), 
to_sfixed(3216.0/65536.0,1,-nbitq), 
to_sfixed(1834.0/65536.0,1,-nbitq), 
to_sfixed(1665.0/65536.0,1,-nbitq), 
to_sfixed(2705.0/65536.0,1,-nbitq), 
to_sfixed(-1200.0/65536.0,1,-nbitq), 
to_sfixed(-898.0/65536.0,1,-nbitq), 
to_sfixed(-2989.0/65536.0,1,-nbitq), 
to_sfixed(-2077.0/65536.0,1,-nbitq), 
to_sfixed(461.0/65536.0,1,-nbitq), 
to_sfixed(425.0/65536.0,1,-nbitq), 
to_sfixed(-1890.0/65536.0,1,-nbitq), 
to_sfixed(2705.0/65536.0,1,-nbitq), 
to_sfixed(551.0/65536.0,1,-nbitq), 
to_sfixed(1784.0/65536.0,1,-nbitq), 
to_sfixed(3142.0/65536.0,1,-nbitq), 
to_sfixed(-3132.0/65536.0,1,-nbitq), 
to_sfixed(-3071.0/65536.0,1,-nbitq), 
to_sfixed(1107.0/65536.0,1,-nbitq), 
to_sfixed(-1317.0/65536.0,1,-nbitq), 
to_sfixed(13.0/65536.0,1,-nbitq), 
to_sfixed(2258.0/65536.0,1,-nbitq), 
to_sfixed(2692.0/65536.0,1,-nbitq), 
to_sfixed(-496.0/65536.0,1,-nbitq), 
to_sfixed(485.0/65536.0,1,-nbitq), 
to_sfixed(3865.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3237.0/65536.0,1,-nbitq), 
to_sfixed(-3430.0/65536.0,1,-nbitq), 
to_sfixed(4879.0/65536.0,1,-nbitq), 
to_sfixed(1786.0/65536.0,1,-nbitq), 
to_sfixed(2899.0/65536.0,1,-nbitq), 
to_sfixed(-707.0/65536.0,1,-nbitq), 
to_sfixed(3072.0/65536.0,1,-nbitq), 
to_sfixed(-3766.0/65536.0,1,-nbitq), 
to_sfixed(-1825.0/65536.0,1,-nbitq), 
to_sfixed(1391.0/65536.0,1,-nbitq), 
to_sfixed(-1807.0/65536.0,1,-nbitq), 
to_sfixed(3318.0/65536.0,1,-nbitq), 
to_sfixed(2251.0/65536.0,1,-nbitq), 
to_sfixed(3080.0/65536.0,1,-nbitq), 
to_sfixed(511.0/65536.0,1,-nbitq), 
to_sfixed(-1425.0/65536.0,1,-nbitq), 
to_sfixed(-898.0/65536.0,1,-nbitq), 
to_sfixed(-2108.0/65536.0,1,-nbitq), 
to_sfixed(4347.0/65536.0,1,-nbitq), 
to_sfixed(-1965.0/65536.0,1,-nbitq), 
to_sfixed(-5604.0/65536.0,1,-nbitq), 
to_sfixed(-2839.0/65536.0,1,-nbitq), 
to_sfixed(-3925.0/65536.0,1,-nbitq), 
to_sfixed(3118.0/65536.0,1,-nbitq), 
to_sfixed(-2058.0/65536.0,1,-nbitq), 
to_sfixed(4846.0/65536.0,1,-nbitq), 
to_sfixed(808.0/65536.0,1,-nbitq), 
to_sfixed(1147.0/65536.0,1,-nbitq), 
to_sfixed(-1829.0/65536.0,1,-nbitq), 
to_sfixed(1374.0/65536.0,1,-nbitq), 
to_sfixed(-3981.0/65536.0,1,-nbitq), 
to_sfixed(-3525.0/65536.0,1,-nbitq), 
to_sfixed(-444.0/65536.0,1,-nbitq), 
to_sfixed(-4958.0/65536.0,1,-nbitq), 
to_sfixed(-3606.0/65536.0,1,-nbitq), 
to_sfixed(-1779.0/65536.0,1,-nbitq), 
to_sfixed(2696.0/65536.0,1,-nbitq), 
to_sfixed(2076.0/65536.0,1,-nbitq), 
to_sfixed(7575.0/65536.0,1,-nbitq), 
to_sfixed(1151.0/65536.0,1,-nbitq), 
to_sfixed(3768.0/65536.0,1,-nbitq), 
to_sfixed(751.0/65536.0,1,-nbitq), 
to_sfixed(-3898.0/65536.0,1,-nbitq), 
to_sfixed(1608.0/65536.0,1,-nbitq), 
to_sfixed(1670.0/65536.0,1,-nbitq), 
to_sfixed(4291.0/65536.0,1,-nbitq), 
to_sfixed(-2712.0/65536.0,1,-nbitq), 
to_sfixed(2891.0/65536.0,1,-nbitq), 
to_sfixed(-2457.0/65536.0,1,-nbitq), 
to_sfixed(4840.0/65536.0,1,-nbitq), 
to_sfixed(-274.0/65536.0,1,-nbitq), 
to_sfixed(6152.0/65536.0,1,-nbitq), 
to_sfixed(2084.0/65536.0,1,-nbitq), 
to_sfixed(1246.0/65536.0,1,-nbitq), 
to_sfixed(3712.0/65536.0,1,-nbitq), 
to_sfixed(3485.0/65536.0,1,-nbitq), 
to_sfixed(2316.0/65536.0,1,-nbitq), 
to_sfixed(1646.0/65536.0,1,-nbitq), 
to_sfixed(-2912.0/65536.0,1,-nbitq), 
to_sfixed(-1953.0/65536.0,1,-nbitq), 
to_sfixed(-411.0/65536.0,1,-nbitq), 
to_sfixed(2457.0/65536.0,1,-nbitq), 
to_sfixed(-512.0/65536.0,1,-nbitq), 
to_sfixed(2243.0/65536.0,1,-nbitq), 
to_sfixed(4998.0/65536.0,1,-nbitq), 
to_sfixed(-307.0/65536.0,1,-nbitq), 
to_sfixed(4213.0/65536.0,1,-nbitq), 
to_sfixed(827.0/65536.0,1,-nbitq), 
to_sfixed(-754.0/65536.0,1,-nbitq), 
to_sfixed(-1489.0/65536.0,1,-nbitq), 
to_sfixed(1935.0/65536.0,1,-nbitq), 
to_sfixed(-776.0/65536.0,1,-nbitq), 
to_sfixed(-497.0/65536.0,1,-nbitq), 
to_sfixed(306.0/65536.0,1,-nbitq), 
to_sfixed(850.0/65536.0,1,-nbitq), 
to_sfixed(-1637.0/65536.0,1,-nbitq), 
to_sfixed(301.0/65536.0,1,-nbitq), 
to_sfixed(678.0/65536.0,1,-nbitq), 
to_sfixed(-1117.0/65536.0,1,-nbitq), 
to_sfixed(1361.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3524.0/65536.0,1,-nbitq), 
to_sfixed(-1201.0/65536.0,1,-nbitq), 
to_sfixed(2938.0/65536.0,1,-nbitq), 
to_sfixed(-1660.0/65536.0,1,-nbitq), 
to_sfixed(1126.0/65536.0,1,-nbitq), 
to_sfixed(-2917.0/65536.0,1,-nbitq), 
to_sfixed(2048.0/65536.0,1,-nbitq), 
to_sfixed(43.0/65536.0,1,-nbitq), 
to_sfixed(-1524.0/65536.0,1,-nbitq), 
to_sfixed(1110.0/65536.0,1,-nbitq), 
to_sfixed(969.0/65536.0,1,-nbitq), 
to_sfixed(5953.0/65536.0,1,-nbitq), 
to_sfixed(2141.0/65536.0,1,-nbitq), 
to_sfixed(-4270.0/65536.0,1,-nbitq), 
to_sfixed(2945.0/65536.0,1,-nbitq), 
to_sfixed(2092.0/65536.0,1,-nbitq), 
to_sfixed(-1818.0/65536.0,1,-nbitq), 
to_sfixed(-1380.0/65536.0,1,-nbitq), 
to_sfixed(4401.0/65536.0,1,-nbitq), 
to_sfixed(2299.0/65536.0,1,-nbitq), 
to_sfixed(-3730.0/65536.0,1,-nbitq), 
to_sfixed(1064.0/65536.0,1,-nbitq), 
to_sfixed(-2830.0/65536.0,1,-nbitq), 
to_sfixed(-1543.0/65536.0,1,-nbitq), 
to_sfixed(-792.0/65536.0,1,-nbitq), 
to_sfixed(2903.0/65536.0,1,-nbitq), 
to_sfixed(-3031.0/65536.0,1,-nbitq), 
to_sfixed(1993.0/65536.0,1,-nbitq), 
to_sfixed(-2839.0/65536.0,1,-nbitq), 
to_sfixed(-3891.0/65536.0,1,-nbitq), 
to_sfixed(70.0/65536.0,1,-nbitq), 
to_sfixed(-3383.0/65536.0,1,-nbitq), 
to_sfixed(-602.0/65536.0,1,-nbitq), 
to_sfixed(671.0/65536.0,1,-nbitq), 
to_sfixed(325.0/65536.0,1,-nbitq), 
to_sfixed(-2162.0/65536.0,1,-nbitq), 
to_sfixed(2783.0/65536.0,1,-nbitq), 
to_sfixed(2236.0/65536.0,1,-nbitq), 
to_sfixed(6641.0/65536.0,1,-nbitq), 
to_sfixed(3555.0/65536.0,1,-nbitq), 
to_sfixed(-1088.0/65536.0,1,-nbitq), 
to_sfixed(-1183.0/65536.0,1,-nbitq), 
to_sfixed(-311.0/65536.0,1,-nbitq), 
to_sfixed(1797.0/65536.0,1,-nbitq), 
to_sfixed(1414.0/65536.0,1,-nbitq), 
to_sfixed(1558.0/65536.0,1,-nbitq), 
to_sfixed(-2867.0/65536.0,1,-nbitq), 
to_sfixed(-1330.0/65536.0,1,-nbitq), 
to_sfixed(2995.0/65536.0,1,-nbitq), 
to_sfixed(1422.0/65536.0,1,-nbitq), 
to_sfixed(2104.0/65536.0,1,-nbitq), 
to_sfixed(-7.0/65536.0,1,-nbitq), 
to_sfixed(188.0/65536.0,1,-nbitq), 
to_sfixed(-3390.0/65536.0,1,-nbitq), 
to_sfixed(3115.0/65536.0,1,-nbitq), 
to_sfixed(-1653.0/65536.0,1,-nbitq), 
to_sfixed(205.0/65536.0,1,-nbitq), 
to_sfixed(2707.0/65536.0,1,-nbitq), 
to_sfixed(-3157.0/65536.0,1,-nbitq), 
to_sfixed(-146.0/65536.0,1,-nbitq), 
to_sfixed(-5736.0/65536.0,1,-nbitq), 
to_sfixed(2292.0/65536.0,1,-nbitq), 
to_sfixed(2160.0/65536.0,1,-nbitq), 
to_sfixed(1648.0/65536.0,1,-nbitq), 
to_sfixed(2598.0/65536.0,1,-nbitq), 
to_sfixed(1988.0/65536.0,1,-nbitq), 
to_sfixed(3575.0/65536.0,1,-nbitq), 
to_sfixed(4075.0/65536.0,1,-nbitq), 
to_sfixed(2521.0/65536.0,1,-nbitq), 
to_sfixed(-1105.0/65536.0,1,-nbitq), 
to_sfixed(-3187.0/65536.0,1,-nbitq), 
to_sfixed(-194.0/65536.0,1,-nbitq), 
to_sfixed(-1193.0/65536.0,1,-nbitq), 
to_sfixed(-670.0/65536.0,1,-nbitq), 
to_sfixed(457.0/65536.0,1,-nbitq), 
to_sfixed(-636.0/65536.0,1,-nbitq), 
to_sfixed(592.0/65536.0,1,-nbitq), 
to_sfixed(4532.0/65536.0,1,-nbitq), 
to_sfixed(-1899.0/65536.0,1,-nbitq), 
to_sfixed(2358.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1694.0/65536.0,1,-nbitq), 
to_sfixed(-547.0/65536.0,1,-nbitq), 
to_sfixed(-1620.0/65536.0,1,-nbitq), 
to_sfixed(-3671.0/65536.0,1,-nbitq), 
to_sfixed(-12.0/65536.0,1,-nbitq), 
to_sfixed(-746.0/65536.0,1,-nbitq), 
to_sfixed(2613.0/65536.0,1,-nbitq), 
to_sfixed(-3175.0/65536.0,1,-nbitq), 
to_sfixed(-1040.0/65536.0,1,-nbitq), 
to_sfixed(-1339.0/65536.0,1,-nbitq), 
to_sfixed(643.0/65536.0,1,-nbitq), 
to_sfixed(797.0/65536.0,1,-nbitq), 
to_sfixed(1177.0/65536.0,1,-nbitq), 
to_sfixed(927.0/65536.0,1,-nbitq), 
to_sfixed(-1131.0/65536.0,1,-nbitq), 
to_sfixed(962.0/65536.0,1,-nbitq), 
to_sfixed(373.0/65536.0,1,-nbitq), 
to_sfixed(-1341.0/65536.0,1,-nbitq), 
to_sfixed(3164.0/65536.0,1,-nbitq), 
to_sfixed(1906.0/65536.0,1,-nbitq), 
to_sfixed(-334.0/65536.0,1,-nbitq), 
to_sfixed(1438.0/65536.0,1,-nbitq), 
to_sfixed(2971.0/65536.0,1,-nbitq), 
to_sfixed(1562.0/65536.0,1,-nbitq), 
to_sfixed(674.0/65536.0,1,-nbitq), 
to_sfixed(-617.0/65536.0,1,-nbitq), 
to_sfixed(-3178.0/65536.0,1,-nbitq), 
to_sfixed(3086.0/65536.0,1,-nbitq), 
to_sfixed(-3540.0/65536.0,1,-nbitq), 
to_sfixed(-3426.0/65536.0,1,-nbitq), 
to_sfixed(1862.0/65536.0,1,-nbitq), 
to_sfixed(-2071.0/65536.0,1,-nbitq), 
to_sfixed(466.0/65536.0,1,-nbitq), 
to_sfixed(-1007.0/65536.0,1,-nbitq), 
to_sfixed(-701.0/65536.0,1,-nbitq), 
to_sfixed(-1678.0/65536.0,1,-nbitq), 
to_sfixed(1664.0/65536.0,1,-nbitq), 
to_sfixed(1404.0/65536.0,1,-nbitq), 
to_sfixed(1049.0/65536.0,1,-nbitq), 
to_sfixed(1631.0/65536.0,1,-nbitq), 
to_sfixed(113.0/65536.0,1,-nbitq), 
to_sfixed(-885.0/65536.0,1,-nbitq), 
to_sfixed(-1834.0/65536.0,1,-nbitq), 
to_sfixed(-531.0/65536.0,1,-nbitq), 
to_sfixed(-2585.0/65536.0,1,-nbitq), 
to_sfixed(3480.0/65536.0,1,-nbitq), 
to_sfixed(1383.0/65536.0,1,-nbitq), 
to_sfixed(3185.0/65536.0,1,-nbitq), 
to_sfixed(-49.0/65536.0,1,-nbitq), 
to_sfixed(408.0/65536.0,1,-nbitq), 
to_sfixed(-1196.0/65536.0,1,-nbitq), 
to_sfixed(910.0/65536.0,1,-nbitq), 
to_sfixed(-282.0/65536.0,1,-nbitq), 
to_sfixed(-4981.0/65536.0,1,-nbitq), 
to_sfixed(2774.0/65536.0,1,-nbitq), 
to_sfixed(2528.0/65536.0,1,-nbitq), 
to_sfixed(-478.0/65536.0,1,-nbitq), 
to_sfixed(3149.0/65536.0,1,-nbitq), 
to_sfixed(1920.0/65536.0,1,-nbitq), 
to_sfixed(-1158.0/65536.0,1,-nbitq), 
to_sfixed(-4696.0/65536.0,1,-nbitq), 
to_sfixed(2256.0/65536.0,1,-nbitq), 
to_sfixed(2584.0/65536.0,1,-nbitq), 
to_sfixed(-808.0/65536.0,1,-nbitq), 
to_sfixed(1331.0/65536.0,1,-nbitq), 
to_sfixed(-1012.0/65536.0,1,-nbitq), 
to_sfixed(-1263.0/65536.0,1,-nbitq), 
to_sfixed(1968.0/65536.0,1,-nbitq), 
to_sfixed(4011.0/65536.0,1,-nbitq), 
to_sfixed(2677.0/65536.0,1,-nbitq), 
to_sfixed(-2386.0/65536.0,1,-nbitq), 
to_sfixed(156.0/65536.0,1,-nbitq), 
to_sfixed(119.0/65536.0,1,-nbitq), 
to_sfixed(-857.0/65536.0,1,-nbitq), 
to_sfixed(-2070.0/65536.0,1,-nbitq), 
to_sfixed(4443.0/65536.0,1,-nbitq), 
to_sfixed(1160.0/65536.0,1,-nbitq), 
to_sfixed(4084.0/65536.0,1,-nbitq), 
to_sfixed(-1588.0/65536.0,1,-nbitq), 
to_sfixed(2174.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-510.0/65536.0,1,-nbitq), 
to_sfixed(2002.0/65536.0,1,-nbitq), 
to_sfixed(1492.0/65536.0,1,-nbitq), 
to_sfixed(-4346.0/65536.0,1,-nbitq), 
to_sfixed(-1054.0/65536.0,1,-nbitq), 
to_sfixed(-187.0/65536.0,1,-nbitq), 
to_sfixed(616.0/65536.0,1,-nbitq), 
to_sfixed(-1147.0/65536.0,1,-nbitq), 
to_sfixed(-2936.0/65536.0,1,-nbitq), 
to_sfixed(1765.0/65536.0,1,-nbitq), 
to_sfixed(27.0/65536.0,1,-nbitq), 
to_sfixed(4945.0/65536.0,1,-nbitq), 
to_sfixed(1338.0/65536.0,1,-nbitq), 
to_sfixed(-3397.0/65536.0,1,-nbitq), 
to_sfixed(3328.0/65536.0,1,-nbitq), 
to_sfixed(484.0/65536.0,1,-nbitq), 
to_sfixed(-896.0/65536.0,1,-nbitq), 
to_sfixed(1458.0/65536.0,1,-nbitq), 
to_sfixed(315.0/65536.0,1,-nbitq), 
to_sfixed(-2061.0/65536.0,1,-nbitq), 
to_sfixed(-5181.0/65536.0,1,-nbitq), 
to_sfixed(2174.0/65536.0,1,-nbitq), 
to_sfixed(3221.0/65536.0,1,-nbitq), 
to_sfixed(4066.0/65536.0,1,-nbitq), 
to_sfixed(-757.0/65536.0,1,-nbitq), 
to_sfixed(1655.0/65536.0,1,-nbitq), 
to_sfixed(-964.0/65536.0,1,-nbitq), 
to_sfixed(2866.0/65536.0,1,-nbitq), 
to_sfixed(-544.0/65536.0,1,-nbitq), 
to_sfixed(888.0/65536.0,1,-nbitq), 
to_sfixed(1088.0/65536.0,1,-nbitq), 
to_sfixed(-198.0/65536.0,1,-nbitq), 
to_sfixed(-4011.0/65536.0,1,-nbitq), 
to_sfixed(629.0/65536.0,1,-nbitq), 
to_sfixed(-132.0/65536.0,1,-nbitq), 
to_sfixed(-3493.0/65536.0,1,-nbitq), 
to_sfixed(-649.0/65536.0,1,-nbitq), 
to_sfixed(1416.0/65536.0,1,-nbitq), 
to_sfixed(4255.0/65536.0,1,-nbitq), 
to_sfixed(-1585.0/65536.0,1,-nbitq), 
to_sfixed(276.0/65536.0,1,-nbitq), 
to_sfixed(-2874.0/65536.0,1,-nbitq), 
to_sfixed(-918.0/65536.0,1,-nbitq), 
to_sfixed(-672.0/65536.0,1,-nbitq), 
to_sfixed(-2443.0/65536.0,1,-nbitq), 
to_sfixed(3407.0/65536.0,1,-nbitq), 
to_sfixed(185.0/65536.0,1,-nbitq), 
to_sfixed(-1440.0/65536.0,1,-nbitq), 
to_sfixed(2420.0/65536.0,1,-nbitq), 
to_sfixed(994.0/65536.0,1,-nbitq), 
to_sfixed(-961.0/65536.0,1,-nbitq), 
to_sfixed(139.0/65536.0,1,-nbitq), 
to_sfixed(-605.0/65536.0,1,-nbitq), 
to_sfixed(-445.0/65536.0,1,-nbitq), 
to_sfixed(3435.0/65536.0,1,-nbitq), 
to_sfixed(-2584.0/65536.0,1,-nbitq), 
to_sfixed(480.0/65536.0,1,-nbitq), 
to_sfixed(-2058.0/65536.0,1,-nbitq), 
to_sfixed(-1048.0/65536.0,1,-nbitq), 
to_sfixed(-1643.0/65536.0,1,-nbitq), 
to_sfixed(-6041.0/65536.0,1,-nbitq), 
to_sfixed(-385.0/65536.0,1,-nbitq), 
to_sfixed(1123.0/65536.0,1,-nbitq), 
to_sfixed(-1945.0/65536.0,1,-nbitq), 
to_sfixed(-1455.0/65536.0,1,-nbitq), 
to_sfixed(2776.0/65536.0,1,-nbitq), 
to_sfixed(1481.0/65536.0,1,-nbitq), 
to_sfixed(2175.0/65536.0,1,-nbitq), 
to_sfixed(595.0/65536.0,1,-nbitq), 
to_sfixed(-2725.0/65536.0,1,-nbitq), 
to_sfixed(-2077.0/65536.0,1,-nbitq), 
to_sfixed(-2346.0/65536.0,1,-nbitq), 
to_sfixed(586.0/65536.0,1,-nbitq), 
to_sfixed(1440.0/65536.0,1,-nbitq), 
to_sfixed(-264.0/65536.0,1,-nbitq), 
to_sfixed(2689.0/65536.0,1,-nbitq), 
to_sfixed(2745.0/65536.0,1,-nbitq), 
to_sfixed(-567.0/65536.0,1,-nbitq), 
to_sfixed(-1100.0/65536.0,1,-nbitq), 
to_sfixed(3709.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2679.0/65536.0,1,-nbitq), 
to_sfixed(-1310.0/65536.0,1,-nbitq), 
to_sfixed(2472.0/65536.0,1,-nbitq), 
to_sfixed(-3623.0/65536.0,1,-nbitq), 
to_sfixed(-2725.0/65536.0,1,-nbitq), 
to_sfixed(-424.0/65536.0,1,-nbitq), 
to_sfixed(-2407.0/65536.0,1,-nbitq), 
to_sfixed(-394.0/65536.0,1,-nbitq), 
to_sfixed(956.0/65536.0,1,-nbitq), 
to_sfixed(-1583.0/65536.0,1,-nbitq), 
to_sfixed(-1831.0/65536.0,1,-nbitq), 
to_sfixed(1866.0/65536.0,1,-nbitq), 
to_sfixed(-731.0/65536.0,1,-nbitq), 
to_sfixed(-3176.0/65536.0,1,-nbitq), 
to_sfixed(-497.0/65536.0,1,-nbitq), 
to_sfixed(2163.0/65536.0,1,-nbitq), 
to_sfixed(-2285.0/65536.0,1,-nbitq), 
to_sfixed(-2204.0/65536.0,1,-nbitq), 
to_sfixed(3273.0/65536.0,1,-nbitq), 
to_sfixed(2398.0/65536.0,1,-nbitq), 
to_sfixed(-463.0/65536.0,1,-nbitq), 
to_sfixed(2046.0/65536.0,1,-nbitq), 
to_sfixed(2168.0/65536.0,1,-nbitq), 
to_sfixed(3202.0/65536.0,1,-nbitq), 
to_sfixed(-2115.0/65536.0,1,-nbitq), 
to_sfixed(279.0/65536.0,1,-nbitq), 
to_sfixed(-401.0/65536.0,1,-nbitq), 
to_sfixed(-809.0/65536.0,1,-nbitq), 
to_sfixed(-2059.0/65536.0,1,-nbitq), 
to_sfixed(-7.0/65536.0,1,-nbitq), 
to_sfixed(2026.0/65536.0,1,-nbitq), 
to_sfixed(-2522.0/65536.0,1,-nbitq), 
to_sfixed(-1043.0/65536.0,1,-nbitq), 
to_sfixed(1036.0/65536.0,1,-nbitq), 
to_sfixed(244.0/65536.0,1,-nbitq), 
to_sfixed(976.0/65536.0,1,-nbitq), 
to_sfixed(718.0/65536.0,1,-nbitq), 
to_sfixed(-1334.0/65536.0,1,-nbitq), 
to_sfixed(-614.0/65536.0,1,-nbitq), 
to_sfixed(-2083.0/65536.0,1,-nbitq), 
to_sfixed(466.0/65536.0,1,-nbitq), 
to_sfixed(1107.0/65536.0,1,-nbitq), 
to_sfixed(-1626.0/65536.0,1,-nbitq), 
to_sfixed(3369.0/65536.0,1,-nbitq), 
to_sfixed(3183.0/65536.0,1,-nbitq), 
to_sfixed(1354.0/65536.0,1,-nbitq), 
to_sfixed(-2685.0/65536.0,1,-nbitq), 
to_sfixed(-1313.0/65536.0,1,-nbitq), 
to_sfixed(-78.0/65536.0,1,-nbitq), 
to_sfixed(-1143.0/65536.0,1,-nbitq), 
to_sfixed(1888.0/65536.0,1,-nbitq), 
to_sfixed(-1721.0/65536.0,1,-nbitq), 
to_sfixed(-17.0/65536.0,1,-nbitq), 
to_sfixed(1485.0/65536.0,1,-nbitq), 
to_sfixed(1635.0/65536.0,1,-nbitq), 
to_sfixed(-874.0/65536.0,1,-nbitq), 
to_sfixed(-2366.0/65536.0,1,-nbitq), 
to_sfixed(2966.0/65536.0,1,-nbitq), 
to_sfixed(1596.0/65536.0,1,-nbitq), 
to_sfixed(621.0/65536.0,1,-nbitq), 
to_sfixed(598.0/65536.0,1,-nbitq), 
to_sfixed(-1889.0/65536.0,1,-nbitq), 
to_sfixed(1345.0/65536.0,1,-nbitq), 
to_sfixed(-3336.0/65536.0,1,-nbitq), 
to_sfixed(2555.0/65536.0,1,-nbitq), 
to_sfixed(3333.0/65536.0,1,-nbitq), 
to_sfixed(1301.0/65536.0,1,-nbitq), 
to_sfixed(672.0/65536.0,1,-nbitq), 
to_sfixed(2176.0/65536.0,1,-nbitq), 
to_sfixed(-168.0/65536.0,1,-nbitq), 
to_sfixed(2680.0/65536.0,1,-nbitq), 
to_sfixed(1461.0/65536.0,1,-nbitq), 
to_sfixed(210.0/65536.0,1,-nbitq), 
to_sfixed(-1458.0/65536.0,1,-nbitq), 
to_sfixed(204.0/65536.0,1,-nbitq), 
to_sfixed(3072.0/65536.0,1,-nbitq), 
to_sfixed(8.0/65536.0,1,-nbitq), 
to_sfixed(-28.0/65536.0,1,-nbitq), 
to_sfixed(29.0/65536.0,1,-nbitq), 
to_sfixed(4981.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-7.0/65536.0,1,-nbitq), 
to_sfixed(1638.0/65536.0,1,-nbitq), 
to_sfixed(1001.0/65536.0,1,-nbitq), 
to_sfixed(-1711.0/65536.0,1,-nbitq), 
to_sfixed(-2629.0/65536.0,1,-nbitq), 
to_sfixed(-4188.0/65536.0,1,-nbitq), 
to_sfixed(-2542.0/65536.0,1,-nbitq), 
to_sfixed(-306.0/65536.0,1,-nbitq), 
to_sfixed(-1547.0/65536.0,1,-nbitq), 
to_sfixed(-2487.0/65536.0,1,-nbitq), 
to_sfixed(2088.0/65536.0,1,-nbitq), 
to_sfixed(1124.0/65536.0,1,-nbitq), 
to_sfixed(2069.0/65536.0,1,-nbitq), 
to_sfixed(-1764.0/65536.0,1,-nbitq), 
to_sfixed(1936.0/65536.0,1,-nbitq), 
to_sfixed(-2455.0/65536.0,1,-nbitq), 
to_sfixed(-740.0/65536.0,1,-nbitq), 
to_sfixed(1478.0/65536.0,1,-nbitq), 
to_sfixed(897.0/65536.0,1,-nbitq), 
to_sfixed(72.0/65536.0,1,-nbitq), 
to_sfixed(-4445.0/65536.0,1,-nbitq), 
to_sfixed(3508.0/65536.0,1,-nbitq), 
to_sfixed(-649.0/65536.0,1,-nbitq), 
to_sfixed(85.0/65536.0,1,-nbitq), 
to_sfixed(1343.0/65536.0,1,-nbitq), 
to_sfixed(3552.0/65536.0,1,-nbitq), 
to_sfixed(-1222.0/65536.0,1,-nbitq), 
to_sfixed(40.0/65536.0,1,-nbitq), 
to_sfixed(1503.0/65536.0,1,-nbitq), 
to_sfixed(1541.0/65536.0,1,-nbitq), 
to_sfixed(81.0/65536.0,1,-nbitq), 
to_sfixed(1290.0/65536.0,1,-nbitq), 
to_sfixed(-209.0/65536.0,1,-nbitq), 
to_sfixed(-2724.0/65536.0,1,-nbitq), 
to_sfixed(2411.0/65536.0,1,-nbitq), 
to_sfixed(1987.0/65536.0,1,-nbitq), 
to_sfixed(478.0/65536.0,1,-nbitq), 
to_sfixed(-4084.0/65536.0,1,-nbitq), 
to_sfixed(153.0/65536.0,1,-nbitq), 
to_sfixed(-41.0/65536.0,1,-nbitq), 
to_sfixed(271.0/65536.0,1,-nbitq), 
to_sfixed(-390.0/65536.0,1,-nbitq), 
to_sfixed(-3881.0/65536.0,1,-nbitq), 
to_sfixed(-1353.0/65536.0,1,-nbitq), 
to_sfixed(-770.0/65536.0,1,-nbitq), 
to_sfixed(-73.0/65536.0,1,-nbitq), 
to_sfixed(-238.0/65536.0,1,-nbitq), 
to_sfixed(1909.0/65536.0,1,-nbitq), 
to_sfixed(-1059.0/65536.0,1,-nbitq), 
to_sfixed(-304.0/65536.0,1,-nbitq), 
to_sfixed(1559.0/65536.0,1,-nbitq), 
to_sfixed(2325.0/65536.0,1,-nbitq), 
to_sfixed(997.0/65536.0,1,-nbitq), 
to_sfixed(415.0/65536.0,1,-nbitq), 
to_sfixed(3331.0/65536.0,1,-nbitq), 
to_sfixed(1760.0/65536.0,1,-nbitq), 
to_sfixed(-811.0/65536.0,1,-nbitq), 
to_sfixed(2055.0/65536.0,1,-nbitq), 
to_sfixed(-784.0/65536.0,1,-nbitq), 
to_sfixed(5309.0/65536.0,1,-nbitq), 
to_sfixed(1978.0/65536.0,1,-nbitq), 
to_sfixed(-784.0/65536.0,1,-nbitq), 
to_sfixed(-395.0/65536.0,1,-nbitq), 
to_sfixed(-2554.0/65536.0,1,-nbitq), 
to_sfixed(-2040.0/65536.0,1,-nbitq), 
to_sfixed(1254.0/65536.0,1,-nbitq), 
to_sfixed(-3318.0/65536.0,1,-nbitq), 
to_sfixed(753.0/65536.0,1,-nbitq), 
to_sfixed(-1814.0/65536.0,1,-nbitq), 
to_sfixed(-396.0/65536.0,1,-nbitq), 
to_sfixed(-1018.0/65536.0,1,-nbitq), 
to_sfixed(-1602.0/65536.0,1,-nbitq), 
to_sfixed(911.0/65536.0,1,-nbitq), 
to_sfixed(-1267.0/65536.0,1,-nbitq), 
to_sfixed(-1972.0/65536.0,1,-nbitq), 
to_sfixed(1454.0/65536.0,1,-nbitq), 
to_sfixed(-348.0/65536.0,1,-nbitq), 
to_sfixed(4080.0/65536.0,1,-nbitq), 
to_sfixed(500.0/65536.0,1,-nbitq), 
to_sfixed(5540.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1515.0/65536.0,1,-nbitq), 
to_sfixed(1213.0/65536.0,1,-nbitq), 
to_sfixed(-192.0/65536.0,1,-nbitq), 
to_sfixed(-2706.0/65536.0,1,-nbitq), 
to_sfixed(975.0/65536.0,1,-nbitq), 
to_sfixed(-891.0/65536.0,1,-nbitq), 
to_sfixed(1212.0/65536.0,1,-nbitq), 
to_sfixed(1634.0/65536.0,1,-nbitq), 
to_sfixed(-2433.0/65536.0,1,-nbitq), 
to_sfixed(-1867.0/65536.0,1,-nbitq), 
to_sfixed(-2258.0/65536.0,1,-nbitq), 
to_sfixed(341.0/65536.0,1,-nbitq), 
to_sfixed(2083.0/65536.0,1,-nbitq), 
to_sfixed(789.0/65536.0,1,-nbitq), 
to_sfixed(-473.0/65536.0,1,-nbitq), 
to_sfixed(1542.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(-1479.0/65536.0,1,-nbitq), 
to_sfixed(333.0/65536.0,1,-nbitq), 
to_sfixed(-718.0/65536.0,1,-nbitq), 
to_sfixed(49.0/65536.0,1,-nbitq), 
to_sfixed(435.0/65536.0,1,-nbitq), 
to_sfixed(218.0/65536.0,1,-nbitq), 
to_sfixed(1655.0/65536.0,1,-nbitq), 
to_sfixed(-2324.0/65536.0,1,-nbitq), 
to_sfixed(1659.0/65536.0,1,-nbitq), 
to_sfixed(-834.0/65536.0,1,-nbitq), 
to_sfixed(-1766.0/65536.0,1,-nbitq), 
to_sfixed(-3424.0/65536.0,1,-nbitq), 
to_sfixed(-2613.0/65536.0,1,-nbitq), 
to_sfixed(2610.0/65536.0,1,-nbitq), 
to_sfixed(170.0/65536.0,1,-nbitq), 
to_sfixed(-1736.0/65536.0,1,-nbitq), 
to_sfixed(-2149.0/65536.0,1,-nbitq), 
to_sfixed(-974.0/65536.0,1,-nbitq), 
to_sfixed(2500.0/65536.0,1,-nbitq), 
to_sfixed(871.0/65536.0,1,-nbitq), 
to_sfixed(-4011.0/65536.0,1,-nbitq), 
to_sfixed(520.0/65536.0,1,-nbitq), 
to_sfixed(2817.0/65536.0,1,-nbitq), 
to_sfixed(1598.0/65536.0,1,-nbitq), 
to_sfixed(1753.0/65536.0,1,-nbitq), 
to_sfixed(-1332.0/65536.0,1,-nbitq), 
to_sfixed(-1038.0/65536.0,1,-nbitq), 
to_sfixed(-2320.0/65536.0,1,-nbitq), 
to_sfixed(3033.0/65536.0,1,-nbitq), 
to_sfixed(1679.0/65536.0,1,-nbitq), 
to_sfixed(-1536.0/65536.0,1,-nbitq), 
to_sfixed(-253.0/65536.0,1,-nbitq), 
to_sfixed(3140.0/65536.0,1,-nbitq), 
to_sfixed(796.0/65536.0,1,-nbitq), 
to_sfixed(-1922.0/65536.0,1,-nbitq), 
to_sfixed(590.0/65536.0,1,-nbitq), 
to_sfixed(-1224.0/65536.0,1,-nbitq), 
to_sfixed(3675.0/65536.0,1,-nbitq), 
to_sfixed(-2046.0/65536.0,1,-nbitq), 
to_sfixed(-2339.0/65536.0,1,-nbitq), 
to_sfixed(3067.0/65536.0,1,-nbitq), 
to_sfixed(435.0/65536.0,1,-nbitq), 
to_sfixed(2245.0/65536.0,1,-nbitq), 
to_sfixed(2417.0/65536.0,1,-nbitq), 
to_sfixed(1827.0/65536.0,1,-nbitq), 
to_sfixed(1139.0/65536.0,1,-nbitq), 
to_sfixed(1600.0/65536.0,1,-nbitq), 
to_sfixed(-677.0/65536.0,1,-nbitq), 
to_sfixed(-1252.0/65536.0,1,-nbitq), 
to_sfixed(-1388.0/65536.0,1,-nbitq), 
to_sfixed(-2078.0/65536.0,1,-nbitq), 
to_sfixed(-1409.0/65536.0,1,-nbitq), 
to_sfixed(3061.0/65536.0,1,-nbitq), 
to_sfixed(-45.0/65536.0,1,-nbitq), 
to_sfixed(2741.0/65536.0,1,-nbitq), 
to_sfixed(3266.0/65536.0,1,-nbitq), 
to_sfixed(2227.0/65536.0,1,-nbitq), 
to_sfixed(804.0/65536.0,1,-nbitq), 
to_sfixed(3498.0/65536.0,1,-nbitq), 
to_sfixed(1733.0/65536.0,1,-nbitq), 
to_sfixed(1474.0/65536.0,1,-nbitq), 
to_sfixed(-2322.0/65536.0,1,-nbitq), 
to_sfixed(2388.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1623.0/65536.0,1,-nbitq), 
to_sfixed(246.0/65536.0,1,-nbitq), 
to_sfixed(3031.0/65536.0,1,-nbitq), 
to_sfixed(-950.0/65536.0,1,-nbitq), 
to_sfixed(2144.0/65536.0,1,-nbitq), 
to_sfixed(82.0/65536.0,1,-nbitq), 
to_sfixed(-2234.0/65536.0,1,-nbitq), 
to_sfixed(-1267.0/65536.0,1,-nbitq), 
to_sfixed(-2281.0/65536.0,1,-nbitq), 
to_sfixed(2234.0/65536.0,1,-nbitq), 
to_sfixed(896.0/65536.0,1,-nbitq), 
to_sfixed(-2500.0/65536.0,1,-nbitq), 
to_sfixed(-1370.0/65536.0,1,-nbitq), 
to_sfixed(1513.0/65536.0,1,-nbitq), 
to_sfixed(-548.0/65536.0,1,-nbitq), 
to_sfixed(2851.0/65536.0,1,-nbitq), 
to_sfixed(1764.0/65536.0,1,-nbitq), 
to_sfixed(3264.0/65536.0,1,-nbitq), 
to_sfixed(1702.0/65536.0,1,-nbitq), 
to_sfixed(-617.0/65536.0,1,-nbitq), 
to_sfixed(610.0/65536.0,1,-nbitq), 
to_sfixed(-2640.0/65536.0,1,-nbitq), 
to_sfixed(1628.0/65536.0,1,-nbitq), 
to_sfixed(709.0/65536.0,1,-nbitq), 
to_sfixed(444.0/65536.0,1,-nbitq), 
to_sfixed(620.0/65536.0,1,-nbitq), 
to_sfixed(-3615.0/65536.0,1,-nbitq), 
to_sfixed(-2461.0/65536.0,1,-nbitq), 
to_sfixed(-884.0/65536.0,1,-nbitq), 
to_sfixed(1967.0/65536.0,1,-nbitq), 
to_sfixed(1643.0/65536.0,1,-nbitq), 
to_sfixed(466.0/65536.0,1,-nbitq), 
to_sfixed(-637.0/65536.0,1,-nbitq), 
to_sfixed(338.0/65536.0,1,-nbitq), 
to_sfixed(-2220.0/65536.0,1,-nbitq), 
to_sfixed(-1305.0/65536.0,1,-nbitq), 
to_sfixed(1231.0/65536.0,1,-nbitq), 
to_sfixed(-716.0/65536.0,1,-nbitq), 
to_sfixed(-929.0/65536.0,1,-nbitq), 
to_sfixed(1767.0/65536.0,1,-nbitq), 
to_sfixed(-2434.0/65536.0,1,-nbitq), 
to_sfixed(-1557.0/65536.0,1,-nbitq), 
to_sfixed(-4.0/65536.0,1,-nbitq), 
to_sfixed(3783.0/65536.0,1,-nbitq), 
to_sfixed(440.0/65536.0,1,-nbitq), 
to_sfixed(699.0/65536.0,1,-nbitq), 
to_sfixed(-2797.0/65536.0,1,-nbitq), 
to_sfixed(-1797.0/65536.0,1,-nbitq), 
to_sfixed(-240.0/65536.0,1,-nbitq), 
to_sfixed(-497.0/65536.0,1,-nbitq), 
to_sfixed(2802.0/65536.0,1,-nbitq), 
to_sfixed(3057.0/65536.0,1,-nbitq), 
to_sfixed(-1568.0/65536.0,1,-nbitq), 
to_sfixed(-2942.0/65536.0,1,-nbitq), 
to_sfixed(4094.0/65536.0,1,-nbitq), 
to_sfixed(-1498.0/65536.0,1,-nbitq), 
to_sfixed(-734.0/65536.0,1,-nbitq), 
to_sfixed(1045.0/65536.0,1,-nbitq), 
to_sfixed(136.0/65536.0,1,-nbitq), 
to_sfixed(617.0/65536.0,1,-nbitq), 
to_sfixed(-204.0/65536.0,1,-nbitq), 
to_sfixed(-2597.0/65536.0,1,-nbitq), 
to_sfixed(1007.0/65536.0,1,-nbitq), 
to_sfixed(-411.0/65536.0,1,-nbitq), 
to_sfixed(-74.0/65536.0,1,-nbitq), 
to_sfixed(1253.0/65536.0,1,-nbitq), 
to_sfixed(-831.0/65536.0,1,-nbitq), 
to_sfixed(-3330.0/65536.0,1,-nbitq), 
to_sfixed(1642.0/65536.0,1,-nbitq), 
to_sfixed(-2413.0/65536.0,1,-nbitq), 
to_sfixed(900.0/65536.0,1,-nbitq), 
to_sfixed(-1936.0/65536.0,1,-nbitq), 
to_sfixed(3957.0/65536.0,1,-nbitq), 
to_sfixed(-2684.0/65536.0,1,-nbitq), 
to_sfixed(1926.0/65536.0,1,-nbitq), 
to_sfixed(1959.0/65536.0,1,-nbitq), 
to_sfixed(-2063.0/65536.0,1,-nbitq), 
to_sfixed(4427.0/65536.0,1,-nbitq), 
to_sfixed(1299.0/65536.0,1,-nbitq), 
to_sfixed(1109.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2969.0/65536.0,1,-nbitq), 
to_sfixed(-1380.0/65536.0,1,-nbitq), 
to_sfixed(917.0/65536.0,1,-nbitq), 
to_sfixed(-2628.0/65536.0,1,-nbitq), 
to_sfixed(806.0/65536.0,1,-nbitq), 
to_sfixed(-3709.0/65536.0,1,-nbitq), 
to_sfixed(2220.0/65536.0,1,-nbitq), 
to_sfixed(476.0/65536.0,1,-nbitq), 
to_sfixed(1872.0/65536.0,1,-nbitq), 
to_sfixed(-2484.0/65536.0,1,-nbitq), 
to_sfixed(-3453.0/65536.0,1,-nbitq), 
to_sfixed(-1729.0/65536.0,1,-nbitq), 
to_sfixed(-857.0/65536.0,1,-nbitq), 
to_sfixed(230.0/65536.0,1,-nbitq), 
to_sfixed(977.0/65536.0,1,-nbitq), 
to_sfixed(714.0/65536.0,1,-nbitq), 
to_sfixed(-913.0/65536.0,1,-nbitq), 
to_sfixed(1415.0/65536.0,1,-nbitq), 
to_sfixed(1250.0/65536.0,1,-nbitq), 
to_sfixed(2567.0/65536.0,1,-nbitq), 
to_sfixed(-2389.0/65536.0,1,-nbitq), 
to_sfixed(382.0/65536.0,1,-nbitq), 
to_sfixed(2701.0/65536.0,1,-nbitq), 
to_sfixed(4145.0/65536.0,1,-nbitq), 
to_sfixed(787.0/65536.0,1,-nbitq), 
to_sfixed(-1921.0/65536.0,1,-nbitq), 
to_sfixed(-3335.0/65536.0,1,-nbitq), 
to_sfixed(3053.0/65536.0,1,-nbitq), 
to_sfixed(-1716.0/65536.0,1,-nbitq), 
to_sfixed(-1343.0/65536.0,1,-nbitq), 
to_sfixed(1053.0/65536.0,1,-nbitq), 
to_sfixed(-290.0/65536.0,1,-nbitq), 
to_sfixed(-2663.0/65536.0,1,-nbitq), 
to_sfixed(-5218.0/65536.0,1,-nbitq), 
to_sfixed(1663.0/65536.0,1,-nbitq), 
to_sfixed(-2095.0/65536.0,1,-nbitq), 
to_sfixed(-25.0/65536.0,1,-nbitq), 
to_sfixed(-2794.0/65536.0,1,-nbitq), 
to_sfixed(-1345.0/65536.0,1,-nbitq), 
to_sfixed(-2487.0/65536.0,1,-nbitq), 
to_sfixed(1317.0/65536.0,1,-nbitq), 
to_sfixed(552.0/65536.0,1,-nbitq), 
to_sfixed(-453.0/65536.0,1,-nbitq), 
to_sfixed(-1224.0/65536.0,1,-nbitq), 
to_sfixed(-2012.0/65536.0,1,-nbitq), 
to_sfixed(2359.0/65536.0,1,-nbitq), 
to_sfixed(1149.0/65536.0,1,-nbitq), 
to_sfixed(194.0/65536.0,1,-nbitq), 
to_sfixed(1609.0/65536.0,1,-nbitq), 
to_sfixed(784.0/65536.0,1,-nbitq), 
to_sfixed(2116.0/65536.0,1,-nbitq), 
to_sfixed(-1399.0/65536.0,1,-nbitq), 
to_sfixed(-766.0/65536.0,1,-nbitq), 
to_sfixed(-2663.0/65536.0,1,-nbitq), 
to_sfixed(2512.0/65536.0,1,-nbitq), 
to_sfixed(1816.0/65536.0,1,-nbitq), 
to_sfixed(263.0/65536.0,1,-nbitq), 
to_sfixed(1293.0/65536.0,1,-nbitq), 
to_sfixed(2364.0/65536.0,1,-nbitq), 
to_sfixed(4008.0/65536.0,1,-nbitq), 
to_sfixed(-2434.0/65536.0,1,-nbitq), 
to_sfixed(-2585.0/65536.0,1,-nbitq), 
to_sfixed(587.0/65536.0,1,-nbitq), 
to_sfixed(-41.0/65536.0,1,-nbitq), 
to_sfixed(1260.0/65536.0,1,-nbitq), 
to_sfixed(-1058.0/65536.0,1,-nbitq), 
to_sfixed(3270.0/65536.0,1,-nbitq), 
to_sfixed(-2119.0/65536.0,1,-nbitq), 
to_sfixed(348.0/65536.0,1,-nbitq), 
to_sfixed(1525.0/65536.0,1,-nbitq), 
to_sfixed(1269.0/65536.0,1,-nbitq), 
to_sfixed(-1004.0/65536.0,1,-nbitq), 
to_sfixed(-1023.0/65536.0,1,-nbitq), 
to_sfixed(-3052.0/65536.0,1,-nbitq), 
to_sfixed(2036.0/65536.0,1,-nbitq), 
to_sfixed(97.0/65536.0,1,-nbitq), 
to_sfixed(2597.0/65536.0,1,-nbitq), 
to_sfixed(2688.0/65536.0,1,-nbitq), 
to_sfixed(1300.0/65536.0,1,-nbitq), 
to_sfixed(2371.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2622.0/65536.0,1,-nbitq), 
to_sfixed(-2573.0/65536.0,1,-nbitq), 
to_sfixed(3749.0/65536.0,1,-nbitq), 
to_sfixed(914.0/65536.0,1,-nbitq), 
to_sfixed(-2119.0/65536.0,1,-nbitq), 
to_sfixed(-3034.0/65536.0,1,-nbitq), 
to_sfixed(1656.0/65536.0,1,-nbitq), 
to_sfixed(-2905.0/65536.0,1,-nbitq), 
to_sfixed(-1769.0/65536.0,1,-nbitq), 
to_sfixed(541.0/65536.0,1,-nbitq), 
to_sfixed(1666.0/65536.0,1,-nbitq), 
to_sfixed(-509.0/65536.0,1,-nbitq), 
to_sfixed(98.0/65536.0,1,-nbitq), 
to_sfixed(-1033.0/65536.0,1,-nbitq), 
to_sfixed(-830.0/65536.0,1,-nbitq), 
to_sfixed(463.0/65536.0,1,-nbitq), 
to_sfixed(-2420.0/65536.0,1,-nbitq), 
to_sfixed(3983.0/65536.0,1,-nbitq), 
to_sfixed(-1282.0/65536.0,1,-nbitq), 
to_sfixed(3027.0/65536.0,1,-nbitq), 
to_sfixed(-217.0/65536.0,1,-nbitq), 
to_sfixed(-922.0/65536.0,1,-nbitq), 
to_sfixed(-1380.0/65536.0,1,-nbitq), 
to_sfixed(4449.0/65536.0,1,-nbitq), 
to_sfixed(-461.0/65536.0,1,-nbitq), 
to_sfixed(-1101.0/65536.0,1,-nbitq), 
to_sfixed(1494.0/65536.0,1,-nbitq), 
to_sfixed(-1896.0/65536.0,1,-nbitq), 
to_sfixed(1733.0/65536.0,1,-nbitq), 
to_sfixed(1709.0/65536.0,1,-nbitq), 
to_sfixed(2174.0/65536.0,1,-nbitq), 
to_sfixed(-1330.0/65536.0,1,-nbitq), 
to_sfixed(79.0/65536.0,1,-nbitq), 
to_sfixed(-3833.0/65536.0,1,-nbitq), 
to_sfixed(-1463.0/65536.0,1,-nbitq), 
to_sfixed(-245.0/65536.0,1,-nbitq), 
to_sfixed(-1315.0/65536.0,1,-nbitq), 
to_sfixed(1036.0/65536.0,1,-nbitq), 
to_sfixed(-4041.0/65536.0,1,-nbitq), 
to_sfixed(1660.0/65536.0,1,-nbitq), 
to_sfixed(-3640.0/65536.0,1,-nbitq), 
to_sfixed(-1881.0/65536.0,1,-nbitq), 
to_sfixed(694.0/65536.0,1,-nbitq), 
to_sfixed(3683.0/65536.0,1,-nbitq), 
to_sfixed(1098.0/65536.0,1,-nbitq), 
to_sfixed(5683.0/65536.0,1,-nbitq), 
to_sfixed(2940.0/65536.0,1,-nbitq), 
to_sfixed(-2169.0/65536.0,1,-nbitq), 
to_sfixed(-2241.0/65536.0,1,-nbitq), 
to_sfixed(-992.0/65536.0,1,-nbitq), 
to_sfixed(1427.0/65536.0,1,-nbitq), 
to_sfixed(2369.0/65536.0,1,-nbitq), 
to_sfixed(-699.0/65536.0,1,-nbitq), 
to_sfixed(-965.0/65536.0,1,-nbitq), 
to_sfixed(-1250.0/65536.0,1,-nbitq), 
to_sfixed(-1758.0/65536.0,1,-nbitq), 
to_sfixed(1440.0/65536.0,1,-nbitq), 
to_sfixed(792.0/65536.0,1,-nbitq), 
to_sfixed(1389.0/65536.0,1,-nbitq), 
to_sfixed(5087.0/65536.0,1,-nbitq), 
to_sfixed(-835.0/65536.0,1,-nbitq), 
to_sfixed(2378.0/65536.0,1,-nbitq), 
to_sfixed(-87.0/65536.0,1,-nbitq), 
to_sfixed(1885.0/65536.0,1,-nbitq), 
to_sfixed(-326.0/65536.0,1,-nbitq), 
to_sfixed(-553.0/65536.0,1,-nbitq), 
to_sfixed(-2023.0/65536.0,1,-nbitq), 
to_sfixed(362.0/65536.0,1,-nbitq), 
to_sfixed(-224.0/65536.0,1,-nbitq), 
to_sfixed(-1253.0/65536.0,1,-nbitq), 
to_sfixed(2259.0/65536.0,1,-nbitq), 
to_sfixed(-769.0/65536.0,1,-nbitq), 
to_sfixed(-33.0/65536.0,1,-nbitq), 
to_sfixed(1230.0/65536.0,1,-nbitq), 
to_sfixed(2442.0/65536.0,1,-nbitq), 
to_sfixed(2465.0/65536.0,1,-nbitq), 
to_sfixed(-2242.0/65536.0,1,-nbitq), 
to_sfixed(3375.0/65536.0,1,-nbitq), 
to_sfixed(-1129.0/65536.0,1,-nbitq), 
to_sfixed(977.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(134.0/65536.0,1,-nbitq), 
to_sfixed(-690.0/65536.0,1,-nbitq), 
to_sfixed(3767.0/65536.0,1,-nbitq), 
to_sfixed(-1472.0/65536.0,1,-nbitq), 
to_sfixed(717.0/65536.0,1,-nbitq), 
to_sfixed(-4465.0/65536.0,1,-nbitq), 
to_sfixed(1996.0/65536.0,1,-nbitq), 
to_sfixed(-3517.0/65536.0,1,-nbitq), 
to_sfixed(1127.0/65536.0,1,-nbitq), 
to_sfixed(-1884.0/65536.0,1,-nbitq), 
to_sfixed(117.0/65536.0,1,-nbitq), 
to_sfixed(-837.0/65536.0,1,-nbitq), 
to_sfixed(-1681.0/65536.0,1,-nbitq), 
to_sfixed(-2673.0/65536.0,1,-nbitq), 
to_sfixed(249.0/65536.0,1,-nbitq), 
to_sfixed(-717.0/65536.0,1,-nbitq), 
to_sfixed(-2039.0/65536.0,1,-nbitq), 
to_sfixed(1819.0/65536.0,1,-nbitq), 
to_sfixed(1762.0/65536.0,1,-nbitq), 
to_sfixed(-1099.0/65536.0,1,-nbitq), 
to_sfixed(-104.0/65536.0,1,-nbitq), 
to_sfixed(-1763.0/65536.0,1,-nbitq), 
to_sfixed(1655.0/65536.0,1,-nbitq), 
to_sfixed(420.0/65536.0,1,-nbitq), 
to_sfixed(-951.0/65536.0,1,-nbitq), 
to_sfixed(972.0/65536.0,1,-nbitq), 
to_sfixed(-582.0/65536.0,1,-nbitq), 
to_sfixed(2931.0/65536.0,1,-nbitq), 
to_sfixed(-1435.0/65536.0,1,-nbitq), 
to_sfixed(-1941.0/65536.0,1,-nbitq), 
to_sfixed(1436.0/65536.0,1,-nbitq), 
to_sfixed(-1007.0/65536.0,1,-nbitq), 
to_sfixed(-4419.0/65536.0,1,-nbitq), 
to_sfixed(-247.0/65536.0,1,-nbitq), 
to_sfixed(-1071.0/65536.0,1,-nbitq), 
to_sfixed(-1804.0/65536.0,1,-nbitq), 
to_sfixed(-1739.0/65536.0,1,-nbitq), 
to_sfixed(1415.0/65536.0,1,-nbitq), 
to_sfixed(-47.0/65536.0,1,-nbitq), 
to_sfixed(276.0/65536.0,1,-nbitq), 
to_sfixed(617.0/65536.0,1,-nbitq), 
to_sfixed(-1660.0/65536.0,1,-nbitq), 
to_sfixed(-2858.0/65536.0,1,-nbitq), 
to_sfixed(1052.0/65536.0,1,-nbitq), 
to_sfixed(2346.0/65536.0,1,-nbitq), 
to_sfixed(4676.0/65536.0,1,-nbitq), 
to_sfixed(3.0/65536.0,1,-nbitq), 
to_sfixed(1801.0/65536.0,1,-nbitq), 
to_sfixed(2136.0/65536.0,1,-nbitq), 
to_sfixed(3704.0/65536.0,1,-nbitq), 
to_sfixed(823.0/65536.0,1,-nbitq), 
to_sfixed(-2501.0/65536.0,1,-nbitq), 
to_sfixed(569.0/65536.0,1,-nbitq), 
to_sfixed(-2205.0/65536.0,1,-nbitq), 
to_sfixed(4108.0/65536.0,1,-nbitq), 
to_sfixed(-2419.0/65536.0,1,-nbitq), 
to_sfixed(2501.0/65536.0,1,-nbitq), 
to_sfixed(-1456.0/65536.0,1,-nbitq), 
to_sfixed(3013.0/65536.0,1,-nbitq), 
to_sfixed(1942.0/65536.0,1,-nbitq), 
to_sfixed(1952.0/65536.0,1,-nbitq), 
to_sfixed(-2192.0/65536.0,1,-nbitq), 
to_sfixed(1269.0/65536.0,1,-nbitq), 
to_sfixed(1017.0/65536.0,1,-nbitq), 
to_sfixed(1318.0/65536.0,1,-nbitq), 
to_sfixed(-672.0/65536.0,1,-nbitq), 
to_sfixed(-1123.0/65536.0,1,-nbitq), 
to_sfixed(-1429.0/65536.0,1,-nbitq), 
to_sfixed(1365.0/65536.0,1,-nbitq), 
to_sfixed(-822.0/65536.0,1,-nbitq), 
to_sfixed(-2555.0/65536.0,1,-nbitq), 
to_sfixed(-1983.0/65536.0,1,-nbitq), 
to_sfixed(1605.0/65536.0,1,-nbitq), 
to_sfixed(-1376.0/65536.0,1,-nbitq), 
to_sfixed(-2515.0/65536.0,1,-nbitq), 
to_sfixed(661.0/65536.0,1,-nbitq), 
to_sfixed(-1430.0/65536.0,1,-nbitq), 
to_sfixed(3551.0/65536.0,1,-nbitq), 
to_sfixed(2559.0/65536.0,1,-nbitq), 
to_sfixed(4715.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3584.0/65536.0,1,-nbitq), 
to_sfixed(203.0/65536.0,1,-nbitq), 
to_sfixed(118.0/65536.0,1,-nbitq), 
to_sfixed(-1203.0/65536.0,1,-nbitq), 
to_sfixed(-1406.0/65536.0,1,-nbitq), 
to_sfixed(930.0/65536.0,1,-nbitq), 
to_sfixed(494.0/65536.0,1,-nbitq), 
to_sfixed(-1170.0/65536.0,1,-nbitq), 
to_sfixed(2123.0/65536.0,1,-nbitq), 
to_sfixed(1875.0/65536.0,1,-nbitq), 
to_sfixed(966.0/65536.0,1,-nbitq), 
to_sfixed(-1911.0/65536.0,1,-nbitq), 
to_sfixed(-72.0/65536.0,1,-nbitq), 
to_sfixed(-3534.0/65536.0,1,-nbitq), 
to_sfixed(-210.0/65536.0,1,-nbitq), 
to_sfixed(-523.0/65536.0,1,-nbitq), 
to_sfixed(792.0/65536.0,1,-nbitq), 
to_sfixed(943.0/65536.0,1,-nbitq), 
to_sfixed(-198.0/65536.0,1,-nbitq), 
to_sfixed(-770.0/65536.0,1,-nbitq), 
to_sfixed(140.0/65536.0,1,-nbitq), 
to_sfixed(-1529.0/65536.0,1,-nbitq), 
to_sfixed(2315.0/65536.0,1,-nbitq), 
to_sfixed(4003.0/65536.0,1,-nbitq), 
to_sfixed(414.0/65536.0,1,-nbitq), 
to_sfixed(3645.0/65536.0,1,-nbitq), 
to_sfixed(-3327.0/65536.0,1,-nbitq), 
to_sfixed(-438.0/65536.0,1,-nbitq), 
to_sfixed(2221.0/65536.0,1,-nbitq), 
to_sfixed(-1624.0/65536.0,1,-nbitq), 
to_sfixed(-922.0/65536.0,1,-nbitq), 
to_sfixed(-1627.0/65536.0,1,-nbitq), 
to_sfixed(-3982.0/65536.0,1,-nbitq), 
to_sfixed(-4281.0/65536.0,1,-nbitq), 
to_sfixed(-2462.0/65536.0,1,-nbitq), 
to_sfixed(-1868.0/65536.0,1,-nbitq), 
to_sfixed(-2880.0/65536.0,1,-nbitq), 
to_sfixed(1102.0/65536.0,1,-nbitq), 
to_sfixed(-1906.0/65536.0,1,-nbitq), 
to_sfixed(1591.0/65536.0,1,-nbitq), 
to_sfixed(-599.0/65536.0,1,-nbitq), 
to_sfixed(2234.0/65536.0,1,-nbitq), 
to_sfixed(-3310.0/65536.0,1,-nbitq), 
to_sfixed(-292.0/65536.0,1,-nbitq), 
to_sfixed(1862.0/65536.0,1,-nbitq), 
to_sfixed(2430.0/65536.0,1,-nbitq), 
to_sfixed(1274.0/65536.0,1,-nbitq), 
to_sfixed(-1135.0/65536.0,1,-nbitq), 
to_sfixed(-1302.0/65536.0,1,-nbitq), 
to_sfixed(432.0/65536.0,1,-nbitq), 
to_sfixed(3109.0/65536.0,1,-nbitq), 
to_sfixed(2375.0/65536.0,1,-nbitq), 
to_sfixed(-4005.0/65536.0,1,-nbitq), 
to_sfixed(-827.0/65536.0,1,-nbitq), 
to_sfixed(-810.0/65536.0,1,-nbitq), 
to_sfixed(-1290.0/65536.0,1,-nbitq), 
to_sfixed(2054.0/65536.0,1,-nbitq), 
to_sfixed(-501.0/65536.0,1,-nbitq), 
to_sfixed(2268.0/65536.0,1,-nbitq), 
to_sfixed(895.0/65536.0,1,-nbitq), 
to_sfixed(-494.0/65536.0,1,-nbitq), 
to_sfixed(-2753.0/65536.0,1,-nbitq), 
to_sfixed(1295.0/65536.0,1,-nbitq), 
to_sfixed(1296.0/65536.0,1,-nbitq), 
to_sfixed(3747.0/65536.0,1,-nbitq), 
to_sfixed(34.0/65536.0,1,-nbitq), 
to_sfixed(-1433.0/65536.0,1,-nbitq), 
to_sfixed(324.0/65536.0,1,-nbitq), 
to_sfixed(2713.0/65536.0,1,-nbitq), 
to_sfixed(1707.0/65536.0,1,-nbitq), 
to_sfixed(299.0/65536.0,1,-nbitq), 
to_sfixed(-1184.0/65536.0,1,-nbitq), 
to_sfixed(-859.0/65536.0,1,-nbitq), 
to_sfixed(-222.0/65536.0,1,-nbitq), 
to_sfixed(-2908.0/65536.0,1,-nbitq), 
to_sfixed(144.0/65536.0,1,-nbitq), 
to_sfixed(2610.0/65536.0,1,-nbitq), 
to_sfixed(4336.0/65536.0,1,-nbitq), 
to_sfixed(731.0/65536.0,1,-nbitq), 
to_sfixed(946.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2077.0/65536.0,1,-nbitq), 
to_sfixed(-265.0/65536.0,1,-nbitq), 
to_sfixed(2345.0/65536.0,1,-nbitq), 
to_sfixed(824.0/65536.0,1,-nbitq), 
to_sfixed(-2394.0/65536.0,1,-nbitq), 
to_sfixed(438.0/65536.0,1,-nbitq), 
to_sfixed(-2358.0/65536.0,1,-nbitq), 
to_sfixed(187.0/65536.0,1,-nbitq), 
to_sfixed(2198.0/65536.0,1,-nbitq), 
to_sfixed(-639.0/65536.0,1,-nbitq), 
to_sfixed(-3959.0/65536.0,1,-nbitq), 
to_sfixed(1809.0/65536.0,1,-nbitq), 
to_sfixed(782.0/65536.0,1,-nbitq), 
to_sfixed(-3982.0/65536.0,1,-nbitq), 
to_sfixed(772.0/65536.0,1,-nbitq), 
to_sfixed(-1862.0/65536.0,1,-nbitq), 
to_sfixed(-2381.0/65536.0,1,-nbitq), 
to_sfixed(-906.0/65536.0,1,-nbitq), 
to_sfixed(3231.0/65536.0,1,-nbitq), 
to_sfixed(2261.0/65536.0,1,-nbitq), 
to_sfixed(-4635.0/65536.0,1,-nbitq), 
to_sfixed(-2533.0/65536.0,1,-nbitq), 
to_sfixed(428.0/65536.0,1,-nbitq), 
to_sfixed(1412.0/65536.0,1,-nbitq), 
to_sfixed(-1755.0/65536.0,1,-nbitq), 
to_sfixed(2722.0/65536.0,1,-nbitq), 
to_sfixed(-1813.0/65536.0,1,-nbitq), 
to_sfixed(-685.0/65536.0,1,-nbitq), 
to_sfixed(488.0/65536.0,1,-nbitq), 
to_sfixed(-1704.0/65536.0,1,-nbitq), 
to_sfixed(-2481.0/65536.0,1,-nbitq), 
to_sfixed(-1596.0/65536.0,1,-nbitq), 
to_sfixed(-8.0/65536.0,1,-nbitq), 
to_sfixed(-4687.0/65536.0,1,-nbitq), 
to_sfixed(2183.0/65536.0,1,-nbitq), 
to_sfixed(-559.0/65536.0,1,-nbitq), 
to_sfixed(-1441.0/65536.0,1,-nbitq), 
to_sfixed(543.0/65536.0,1,-nbitq), 
to_sfixed(-2504.0/65536.0,1,-nbitq), 
to_sfixed(3705.0/65536.0,1,-nbitq), 
to_sfixed(-1244.0/65536.0,1,-nbitq), 
to_sfixed(-2032.0/65536.0,1,-nbitq), 
to_sfixed(-133.0/65536.0,1,-nbitq), 
to_sfixed(-2410.0/65536.0,1,-nbitq), 
to_sfixed(296.0/65536.0,1,-nbitq), 
to_sfixed(597.0/65536.0,1,-nbitq), 
to_sfixed(-730.0/65536.0,1,-nbitq), 
to_sfixed(-1489.0/65536.0,1,-nbitq), 
to_sfixed(2925.0/65536.0,1,-nbitq), 
to_sfixed(1094.0/65536.0,1,-nbitq), 
to_sfixed(-1569.0/65536.0,1,-nbitq), 
to_sfixed(1578.0/65536.0,1,-nbitq), 
to_sfixed(-3865.0/65536.0,1,-nbitq), 
to_sfixed(45.0/65536.0,1,-nbitq), 
to_sfixed(470.0/65536.0,1,-nbitq), 
to_sfixed(1789.0/65536.0,1,-nbitq), 
to_sfixed(-1157.0/65536.0,1,-nbitq), 
to_sfixed(-2099.0/65536.0,1,-nbitq), 
to_sfixed(-746.0/65536.0,1,-nbitq), 
to_sfixed(3608.0/65536.0,1,-nbitq), 
to_sfixed(-470.0/65536.0,1,-nbitq), 
to_sfixed(2165.0/65536.0,1,-nbitq), 
to_sfixed(-2327.0/65536.0,1,-nbitq), 
to_sfixed(-634.0/65536.0,1,-nbitq), 
to_sfixed(67.0/65536.0,1,-nbitq), 
to_sfixed(1032.0/65536.0,1,-nbitq), 
to_sfixed(2903.0/65536.0,1,-nbitq), 
to_sfixed(-1232.0/65536.0,1,-nbitq), 
to_sfixed(1791.0/65536.0,1,-nbitq), 
to_sfixed(2185.0/65536.0,1,-nbitq), 
to_sfixed(-910.0/65536.0,1,-nbitq), 
to_sfixed(-322.0/65536.0,1,-nbitq), 
to_sfixed(407.0/65536.0,1,-nbitq), 
to_sfixed(-416.0/65536.0,1,-nbitq), 
to_sfixed(987.0/65536.0,1,-nbitq), 
to_sfixed(827.0/65536.0,1,-nbitq), 
to_sfixed(1274.0/65536.0,1,-nbitq), 
to_sfixed(4519.0/65536.0,1,-nbitq), 
to_sfixed(726.0/65536.0,1,-nbitq), 
to_sfixed(2296.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2438.0/65536.0,1,-nbitq), 
to_sfixed(1549.0/65536.0,1,-nbitq), 
to_sfixed(-611.0/65536.0,1,-nbitq), 
to_sfixed(333.0/65536.0,1,-nbitq), 
to_sfixed(753.0/65536.0,1,-nbitq), 
to_sfixed(-4086.0/65536.0,1,-nbitq), 
to_sfixed(-1228.0/65536.0,1,-nbitq), 
to_sfixed(-2433.0/65536.0,1,-nbitq), 
to_sfixed(-558.0/65536.0,1,-nbitq), 
to_sfixed(2480.0/65536.0,1,-nbitq), 
to_sfixed(-1902.0/65536.0,1,-nbitq), 
to_sfixed(3223.0/65536.0,1,-nbitq), 
to_sfixed(-1512.0/65536.0,1,-nbitq), 
to_sfixed(1154.0/65536.0,1,-nbitq), 
to_sfixed(3068.0/65536.0,1,-nbitq), 
to_sfixed(2737.0/65536.0,1,-nbitq), 
to_sfixed(1509.0/65536.0,1,-nbitq), 
to_sfixed(3727.0/65536.0,1,-nbitq), 
to_sfixed(1362.0/65536.0,1,-nbitq), 
to_sfixed(1371.0/65536.0,1,-nbitq), 
to_sfixed(-2337.0/65536.0,1,-nbitq), 
to_sfixed(-2499.0/65536.0,1,-nbitq), 
to_sfixed(2362.0/65536.0,1,-nbitq), 
to_sfixed(1300.0/65536.0,1,-nbitq), 
to_sfixed(446.0/65536.0,1,-nbitq), 
to_sfixed(668.0/65536.0,1,-nbitq), 
to_sfixed(-2323.0/65536.0,1,-nbitq), 
to_sfixed(26.0/65536.0,1,-nbitq), 
to_sfixed(1313.0/65536.0,1,-nbitq), 
to_sfixed(947.0/65536.0,1,-nbitq), 
to_sfixed(1755.0/65536.0,1,-nbitq), 
to_sfixed(1302.0/65536.0,1,-nbitq), 
to_sfixed(-3450.0/65536.0,1,-nbitq), 
to_sfixed(-2150.0/65536.0,1,-nbitq), 
to_sfixed(-2618.0/65536.0,1,-nbitq), 
to_sfixed(1997.0/65536.0,1,-nbitq), 
to_sfixed(-2505.0/65536.0,1,-nbitq), 
to_sfixed(724.0/65536.0,1,-nbitq), 
to_sfixed(2300.0/65536.0,1,-nbitq), 
to_sfixed(1290.0/65536.0,1,-nbitq), 
to_sfixed(-2650.0/65536.0,1,-nbitq), 
to_sfixed(59.0/65536.0,1,-nbitq), 
to_sfixed(-3287.0/65536.0,1,-nbitq), 
to_sfixed(-2485.0/65536.0,1,-nbitq), 
to_sfixed(-1577.0/65536.0,1,-nbitq), 
to_sfixed(6787.0/65536.0,1,-nbitq), 
to_sfixed(1692.0/65536.0,1,-nbitq), 
to_sfixed(1488.0/65536.0,1,-nbitq), 
to_sfixed(1276.0/65536.0,1,-nbitq), 
to_sfixed(-162.0/65536.0,1,-nbitq), 
to_sfixed(1135.0/65536.0,1,-nbitq), 
to_sfixed(1761.0/65536.0,1,-nbitq), 
to_sfixed(331.0/65536.0,1,-nbitq), 
to_sfixed(3501.0/65536.0,1,-nbitq), 
to_sfixed(1573.0/65536.0,1,-nbitq), 
to_sfixed(76.0/65536.0,1,-nbitq), 
to_sfixed(-1871.0/65536.0,1,-nbitq), 
to_sfixed(-61.0/65536.0,1,-nbitq), 
to_sfixed(1867.0/65536.0,1,-nbitq), 
to_sfixed(3796.0/65536.0,1,-nbitq), 
to_sfixed(1382.0/65536.0,1,-nbitq), 
to_sfixed(2061.0/65536.0,1,-nbitq), 
to_sfixed(1202.0/65536.0,1,-nbitq), 
to_sfixed(894.0/65536.0,1,-nbitq), 
to_sfixed(2298.0/65536.0,1,-nbitq), 
to_sfixed(-501.0/65536.0,1,-nbitq), 
to_sfixed(502.0/65536.0,1,-nbitq), 
to_sfixed(1389.0/65536.0,1,-nbitq), 
to_sfixed(157.0/65536.0,1,-nbitq), 
to_sfixed(-713.0/65536.0,1,-nbitq), 
to_sfixed(1982.0/65536.0,1,-nbitq), 
to_sfixed(-2880.0/65536.0,1,-nbitq), 
to_sfixed(-1908.0/65536.0,1,-nbitq), 
to_sfixed(-2085.0/65536.0,1,-nbitq), 
to_sfixed(433.0/65536.0,1,-nbitq), 
to_sfixed(-1181.0/65536.0,1,-nbitq), 
to_sfixed(2478.0/65536.0,1,-nbitq), 
to_sfixed(2981.0/65536.0,1,-nbitq), 
to_sfixed(1294.0/65536.0,1,-nbitq), 
to_sfixed(3152.0/65536.0,1,-nbitq)  ), 
( to_sfixed(977.0/65536.0,1,-nbitq), 
to_sfixed(494.0/65536.0,1,-nbitq), 
to_sfixed(2740.0/65536.0,1,-nbitq), 
to_sfixed(1404.0/65536.0,1,-nbitq), 
to_sfixed(518.0/65536.0,1,-nbitq), 
to_sfixed(-2310.0/65536.0,1,-nbitq), 
to_sfixed(-1763.0/65536.0,1,-nbitq), 
to_sfixed(-180.0/65536.0,1,-nbitq), 
to_sfixed(-2829.0/65536.0,1,-nbitq), 
to_sfixed(576.0/65536.0,1,-nbitq), 
to_sfixed(-2165.0/65536.0,1,-nbitq), 
to_sfixed(865.0/65536.0,1,-nbitq), 
to_sfixed(-88.0/65536.0,1,-nbitq), 
to_sfixed(-2275.0/65536.0,1,-nbitq), 
to_sfixed(-674.0/65536.0,1,-nbitq), 
to_sfixed(-1373.0/65536.0,1,-nbitq), 
to_sfixed(-1349.0/65536.0,1,-nbitq), 
to_sfixed(3794.0/65536.0,1,-nbitq), 
to_sfixed(4178.0/65536.0,1,-nbitq), 
to_sfixed(2135.0/65536.0,1,-nbitq), 
to_sfixed(1305.0/65536.0,1,-nbitq), 
to_sfixed(-1591.0/65536.0,1,-nbitq), 
to_sfixed(5497.0/65536.0,1,-nbitq), 
to_sfixed(892.0/65536.0,1,-nbitq), 
to_sfixed(-2428.0/65536.0,1,-nbitq), 
to_sfixed(1315.0/65536.0,1,-nbitq), 
to_sfixed(-3642.0/65536.0,1,-nbitq), 
to_sfixed(-191.0/65536.0,1,-nbitq), 
to_sfixed(-1869.0/65536.0,1,-nbitq), 
to_sfixed(2555.0/65536.0,1,-nbitq), 
to_sfixed(-2002.0/65536.0,1,-nbitq), 
to_sfixed(-1018.0/65536.0,1,-nbitq), 
to_sfixed(-243.0/65536.0,1,-nbitq), 
to_sfixed(-5534.0/65536.0,1,-nbitq), 
to_sfixed(-2408.0/65536.0,1,-nbitq), 
to_sfixed(1137.0/65536.0,1,-nbitq), 
to_sfixed(1345.0/65536.0,1,-nbitq), 
to_sfixed(854.0/65536.0,1,-nbitq), 
to_sfixed(-2016.0/65536.0,1,-nbitq), 
to_sfixed(2170.0/65536.0,1,-nbitq), 
to_sfixed(-3091.0/65536.0,1,-nbitq), 
to_sfixed(2000.0/65536.0,1,-nbitq), 
to_sfixed(-1917.0/65536.0,1,-nbitq), 
to_sfixed(467.0/65536.0,1,-nbitq), 
to_sfixed(-26.0/65536.0,1,-nbitq), 
to_sfixed(4701.0/65536.0,1,-nbitq), 
to_sfixed(1129.0/65536.0,1,-nbitq), 
to_sfixed(-1084.0/65536.0,1,-nbitq), 
to_sfixed(2520.0/65536.0,1,-nbitq), 
to_sfixed(246.0/65536.0,1,-nbitq), 
to_sfixed(2820.0/65536.0,1,-nbitq), 
to_sfixed(1558.0/65536.0,1,-nbitq), 
to_sfixed(-3742.0/65536.0,1,-nbitq), 
to_sfixed(386.0/65536.0,1,-nbitq), 
to_sfixed(2276.0/65536.0,1,-nbitq), 
to_sfixed(218.0/65536.0,1,-nbitq), 
to_sfixed(486.0/65536.0,1,-nbitq), 
to_sfixed(-1010.0/65536.0,1,-nbitq), 
to_sfixed(873.0/65536.0,1,-nbitq), 
to_sfixed(2363.0/65536.0,1,-nbitq), 
to_sfixed(-340.0/65536.0,1,-nbitq), 
to_sfixed(-571.0/65536.0,1,-nbitq), 
to_sfixed(2111.0/65536.0,1,-nbitq), 
to_sfixed(85.0/65536.0,1,-nbitq), 
to_sfixed(-8.0/65536.0,1,-nbitq), 
to_sfixed(-1052.0/65536.0,1,-nbitq), 
to_sfixed(2752.0/65536.0,1,-nbitq), 
to_sfixed(1594.0/65536.0,1,-nbitq), 
to_sfixed(2066.0/65536.0,1,-nbitq), 
to_sfixed(822.0/65536.0,1,-nbitq), 
to_sfixed(3066.0/65536.0,1,-nbitq), 
to_sfixed(-3264.0/65536.0,1,-nbitq), 
to_sfixed(-1781.0/65536.0,1,-nbitq), 
to_sfixed(-2766.0/65536.0,1,-nbitq), 
to_sfixed(-2712.0/65536.0,1,-nbitq), 
to_sfixed(1208.0/65536.0,1,-nbitq), 
to_sfixed(-2054.0/65536.0,1,-nbitq), 
to_sfixed(1586.0/65536.0,1,-nbitq), 
to_sfixed(79.0/65536.0,1,-nbitq), 
to_sfixed(1305.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-449.0/65536.0,1,-nbitq), 
to_sfixed(-435.0/65536.0,1,-nbitq), 
to_sfixed(2659.0/65536.0,1,-nbitq), 
to_sfixed(-1316.0/65536.0,1,-nbitq), 
to_sfixed(-520.0/65536.0,1,-nbitq), 
to_sfixed(1073.0/65536.0,1,-nbitq), 
to_sfixed(-283.0/65536.0,1,-nbitq), 
to_sfixed(1683.0/65536.0,1,-nbitq), 
to_sfixed(774.0/65536.0,1,-nbitq), 
to_sfixed(2391.0/65536.0,1,-nbitq), 
to_sfixed(-3625.0/65536.0,1,-nbitq), 
to_sfixed(4039.0/65536.0,1,-nbitq), 
to_sfixed(1984.0/65536.0,1,-nbitq), 
to_sfixed(1309.0/65536.0,1,-nbitq), 
to_sfixed(-21.0/65536.0,1,-nbitq), 
to_sfixed(-2520.0/65536.0,1,-nbitq), 
to_sfixed(1850.0/65536.0,1,-nbitq), 
to_sfixed(4646.0/65536.0,1,-nbitq), 
to_sfixed(2020.0/65536.0,1,-nbitq), 
to_sfixed(2533.0/65536.0,1,-nbitq), 
to_sfixed(-3622.0/65536.0,1,-nbitq), 
to_sfixed(4425.0/65536.0,1,-nbitq), 
to_sfixed(2150.0/65536.0,1,-nbitq), 
to_sfixed(-590.0/65536.0,1,-nbitq), 
to_sfixed(-3323.0/65536.0,1,-nbitq), 
to_sfixed(-2026.0/65536.0,1,-nbitq), 
to_sfixed(1178.0/65536.0,1,-nbitq), 
to_sfixed(-1791.0/65536.0,1,-nbitq), 
to_sfixed(-1959.0/65536.0,1,-nbitq), 
to_sfixed(1863.0/65536.0,1,-nbitq), 
to_sfixed(-1882.0/65536.0,1,-nbitq), 
to_sfixed(-628.0/65536.0,1,-nbitq), 
to_sfixed(-5476.0/65536.0,1,-nbitq), 
to_sfixed(-4101.0/65536.0,1,-nbitq), 
to_sfixed(1037.0/65536.0,1,-nbitq), 
to_sfixed(-752.0/65536.0,1,-nbitq), 
to_sfixed(2777.0/65536.0,1,-nbitq), 
to_sfixed(269.0/65536.0,1,-nbitq), 
to_sfixed(5919.0/65536.0,1,-nbitq), 
to_sfixed(1491.0/65536.0,1,-nbitq), 
to_sfixed(-1078.0/65536.0,1,-nbitq), 
to_sfixed(-945.0/65536.0,1,-nbitq), 
to_sfixed(-4675.0/65536.0,1,-nbitq), 
to_sfixed(-1153.0/65536.0,1,-nbitq), 
to_sfixed(-910.0/65536.0,1,-nbitq), 
to_sfixed(5379.0/65536.0,1,-nbitq), 
to_sfixed(-544.0/65536.0,1,-nbitq), 
to_sfixed(3056.0/65536.0,1,-nbitq), 
to_sfixed(1172.0/65536.0,1,-nbitq), 
to_sfixed(1752.0/65536.0,1,-nbitq), 
to_sfixed(-1293.0/65536.0,1,-nbitq), 
to_sfixed(-749.0/65536.0,1,-nbitq), 
to_sfixed(-1204.0/65536.0,1,-nbitq), 
to_sfixed(1789.0/65536.0,1,-nbitq), 
to_sfixed(2056.0/65536.0,1,-nbitq), 
to_sfixed(673.0/65536.0,1,-nbitq), 
to_sfixed(3063.0/65536.0,1,-nbitq), 
to_sfixed(2110.0/65536.0,1,-nbitq), 
to_sfixed(-2575.0/65536.0,1,-nbitq), 
to_sfixed(2252.0/65536.0,1,-nbitq), 
to_sfixed(-3448.0/65536.0,1,-nbitq), 
to_sfixed(-1760.0/65536.0,1,-nbitq), 
to_sfixed(1522.0/65536.0,1,-nbitq), 
to_sfixed(1883.0/65536.0,1,-nbitq), 
to_sfixed(-393.0/65536.0,1,-nbitq), 
to_sfixed(-796.0/65536.0,1,-nbitq), 
to_sfixed(2829.0/65536.0,1,-nbitq), 
to_sfixed(401.0/65536.0,1,-nbitq), 
to_sfixed(2426.0/65536.0,1,-nbitq), 
to_sfixed(-699.0/65536.0,1,-nbitq), 
to_sfixed(400.0/65536.0,1,-nbitq), 
to_sfixed(130.0/65536.0,1,-nbitq), 
to_sfixed(972.0/65536.0,1,-nbitq), 
to_sfixed(1817.0/65536.0,1,-nbitq), 
to_sfixed(1058.0/65536.0,1,-nbitq), 
to_sfixed(-3018.0/65536.0,1,-nbitq), 
to_sfixed(-274.0/65536.0,1,-nbitq), 
to_sfixed(1413.0/65536.0,1,-nbitq), 
to_sfixed(-1864.0/65536.0,1,-nbitq), 
to_sfixed(3688.0/65536.0,1,-nbitq)  ), 
( to_sfixed(169.0/65536.0,1,-nbitq), 
to_sfixed(-519.0/65536.0,1,-nbitq), 
to_sfixed(-1160.0/65536.0,1,-nbitq), 
to_sfixed(-854.0/65536.0,1,-nbitq), 
to_sfixed(1101.0/65536.0,1,-nbitq), 
to_sfixed(-2636.0/65536.0,1,-nbitq), 
to_sfixed(2348.0/65536.0,1,-nbitq), 
to_sfixed(-2964.0/65536.0,1,-nbitq), 
to_sfixed(348.0/65536.0,1,-nbitq), 
to_sfixed(2376.0/65536.0,1,-nbitq), 
to_sfixed(-4966.0/65536.0,1,-nbitq), 
to_sfixed(2705.0/65536.0,1,-nbitq), 
to_sfixed(1838.0/65536.0,1,-nbitq), 
to_sfixed(-897.0/65536.0,1,-nbitq), 
to_sfixed(3247.0/65536.0,1,-nbitq), 
to_sfixed(1356.0/65536.0,1,-nbitq), 
to_sfixed(-1860.0/65536.0,1,-nbitq), 
to_sfixed(2944.0/65536.0,1,-nbitq), 
to_sfixed(22.0/65536.0,1,-nbitq), 
to_sfixed(-942.0/65536.0,1,-nbitq), 
to_sfixed(353.0/65536.0,1,-nbitq), 
to_sfixed(164.0/65536.0,1,-nbitq), 
to_sfixed(338.0/65536.0,1,-nbitq), 
to_sfixed(549.0/65536.0,1,-nbitq), 
to_sfixed(-185.0/65536.0,1,-nbitq), 
to_sfixed(-2566.0/65536.0,1,-nbitq), 
to_sfixed(-982.0/65536.0,1,-nbitq), 
to_sfixed(648.0/65536.0,1,-nbitq), 
to_sfixed(-3295.0/65536.0,1,-nbitq), 
to_sfixed(2962.0/65536.0,1,-nbitq), 
to_sfixed(582.0/65536.0,1,-nbitq), 
to_sfixed(-770.0/65536.0,1,-nbitq), 
to_sfixed(-1951.0/65536.0,1,-nbitq), 
to_sfixed(-2675.0/65536.0,1,-nbitq), 
to_sfixed(-2043.0/65536.0,1,-nbitq), 
to_sfixed(521.0/65536.0,1,-nbitq), 
to_sfixed(2718.0/65536.0,1,-nbitq), 
to_sfixed(-1716.0/65536.0,1,-nbitq), 
to_sfixed(5541.0/65536.0,1,-nbitq), 
to_sfixed(-601.0/65536.0,1,-nbitq), 
to_sfixed(1934.0/65536.0,1,-nbitq), 
to_sfixed(-399.0/65536.0,1,-nbitq), 
to_sfixed(-1979.0/65536.0,1,-nbitq), 
to_sfixed(-2357.0/65536.0,1,-nbitq), 
to_sfixed(1596.0/65536.0,1,-nbitq), 
to_sfixed(3549.0/65536.0,1,-nbitq), 
to_sfixed(2714.0/65536.0,1,-nbitq), 
to_sfixed(-1733.0/65536.0,1,-nbitq), 
to_sfixed(2061.0/65536.0,1,-nbitq), 
to_sfixed(2281.0/65536.0,1,-nbitq), 
to_sfixed(863.0/65536.0,1,-nbitq), 
to_sfixed(-4041.0/65536.0,1,-nbitq), 
to_sfixed(-2674.0/65536.0,1,-nbitq), 
to_sfixed(1141.0/65536.0,1,-nbitq), 
to_sfixed(2056.0/65536.0,1,-nbitq), 
to_sfixed(101.0/65536.0,1,-nbitq), 
to_sfixed(1801.0/65536.0,1,-nbitq), 
to_sfixed(-1422.0/65536.0,1,-nbitq), 
to_sfixed(683.0/65536.0,1,-nbitq), 
to_sfixed(1230.0/65536.0,1,-nbitq), 
to_sfixed(228.0/65536.0,1,-nbitq), 
to_sfixed(-570.0/65536.0,1,-nbitq), 
to_sfixed(1875.0/65536.0,1,-nbitq), 
to_sfixed(-2692.0/65536.0,1,-nbitq), 
to_sfixed(-17.0/65536.0,1,-nbitq), 
to_sfixed(4653.0/65536.0,1,-nbitq), 
to_sfixed(3275.0/65536.0,1,-nbitq), 
to_sfixed(2014.0/65536.0,1,-nbitq), 
to_sfixed(-656.0/65536.0,1,-nbitq), 
to_sfixed(466.0/65536.0,1,-nbitq), 
to_sfixed(354.0/65536.0,1,-nbitq), 
to_sfixed(-1465.0/65536.0,1,-nbitq), 
to_sfixed(-1672.0/65536.0,1,-nbitq), 
to_sfixed(591.0/65536.0,1,-nbitq), 
to_sfixed(-1501.0/65536.0,1,-nbitq), 
to_sfixed(903.0/65536.0,1,-nbitq), 
to_sfixed(-981.0/65536.0,1,-nbitq), 
to_sfixed(2844.0/65536.0,1,-nbitq), 
to_sfixed(2567.0/65536.0,1,-nbitq), 
to_sfixed(-835.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-821.0/65536.0,1,-nbitq), 
to_sfixed(2052.0/65536.0,1,-nbitq), 
to_sfixed(-528.0/65536.0,1,-nbitq), 
to_sfixed(-3407.0/65536.0,1,-nbitq), 
to_sfixed(-724.0/65536.0,1,-nbitq), 
to_sfixed(-3570.0/65536.0,1,-nbitq), 
to_sfixed(-398.0/65536.0,1,-nbitq), 
to_sfixed(-1951.0/65536.0,1,-nbitq), 
to_sfixed(1085.0/65536.0,1,-nbitq), 
to_sfixed(-419.0/65536.0,1,-nbitq), 
to_sfixed(-3294.0/65536.0,1,-nbitq), 
to_sfixed(3969.0/65536.0,1,-nbitq), 
to_sfixed(1066.0/65536.0,1,-nbitq), 
to_sfixed(1683.0/65536.0,1,-nbitq), 
to_sfixed(-537.0/65536.0,1,-nbitq), 
to_sfixed(-576.0/65536.0,1,-nbitq), 
to_sfixed(2472.0/65536.0,1,-nbitq), 
to_sfixed(3923.0/65536.0,1,-nbitq), 
to_sfixed(4528.0/65536.0,1,-nbitq), 
to_sfixed(-392.0/65536.0,1,-nbitq), 
to_sfixed(-1693.0/65536.0,1,-nbitq), 
to_sfixed(1219.0/65536.0,1,-nbitq), 
to_sfixed(-107.0/65536.0,1,-nbitq), 
to_sfixed(-214.0/65536.0,1,-nbitq), 
to_sfixed(-2688.0/65536.0,1,-nbitq), 
to_sfixed(-1584.0/65536.0,1,-nbitq), 
to_sfixed(-899.0/65536.0,1,-nbitq), 
to_sfixed(-49.0/65536.0,1,-nbitq), 
to_sfixed(-2001.0/65536.0,1,-nbitq), 
to_sfixed(-1493.0/65536.0,1,-nbitq), 
to_sfixed(-1327.0/65536.0,1,-nbitq), 
to_sfixed(-3168.0/65536.0,1,-nbitq), 
to_sfixed(-5788.0/65536.0,1,-nbitq), 
to_sfixed(-3788.0/65536.0,1,-nbitq), 
to_sfixed(1004.0/65536.0,1,-nbitq), 
to_sfixed(-215.0/65536.0,1,-nbitq), 
to_sfixed(3301.0/65536.0,1,-nbitq), 
to_sfixed(1985.0/65536.0,1,-nbitq), 
to_sfixed(1583.0/65536.0,1,-nbitq), 
to_sfixed(1005.0/65536.0,1,-nbitq), 
to_sfixed(2928.0/65536.0,1,-nbitq), 
to_sfixed(174.0/65536.0,1,-nbitq), 
to_sfixed(-3583.0/65536.0,1,-nbitq), 
to_sfixed(-1643.0/65536.0,1,-nbitq), 
to_sfixed(-34.0/65536.0,1,-nbitq), 
to_sfixed(2210.0/65536.0,1,-nbitq), 
to_sfixed(1574.0/65536.0,1,-nbitq), 
to_sfixed(-1123.0/65536.0,1,-nbitq), 
to_sfixed(3013.0/65536.0,1,-nbitq), 
to_sfixed(3555.0/65536.0,1,-nbitq), 
to_sfixed(773.0/65536.0,1,-nbitq), 
to_sfixed(846.0/65536.0,1,-nbitq), 
to_sfixed(-3515.0/65536.0,1,-nbitq), 
to_sfixed(2449.0/65536.0,1,-nbitq), 
to_sfixed(5168.0/65536.0,1,-nbitq), 
to_sfixed(-1801.0/65536.0,1,-nbitq), 
to_sfixed(2927.0/65536.0,1,-nbitq), 
to_sfixed(-2354.0/65536.0,1,-nbitq), 
to_sfixed(422.0/65536.0,1,-nbitq), 
to_sfixed(468.0/65536.0,1,-nbitq), 
to_sfixed(102.0/65536.0,1,-nbitq), 
to_sfixed(1544.0/65536.0,1,-nbitq), 
to_sfixed(2179.0/65536.0,1,-nbitq), 
to_sfixed(1487.0/65536.0,1,-nbitq), 
to_sfixed(-1731.0/65536.0,1,-nbitq), 
to_sfixed(106.0/65536.0,1,-nbitq), 
to_sfixed(-570.0/65536.0,1,-nbitq), 
to_sfixed(-1057.0/65536.0,1,-nbitq), 
to_sfixed(1848.0/65536.0,1,-nbitq), 
to_sfixed(-197.0/65536.0,1,-nbitq), 
to_sfixed(831.0/65536.0,1,-nbitq), 
to_sfixed(3139.0/65536.0,1,-nbitq), 
to_sfixed(-1003.0/65536.0,1,-nbitq), 
to_sfixed(-1747.0/65536.0,1,-nbitq), 
to_sfixed(-718.0/65536.0,1,-nbitq), 
to_sfixed(1307.0/65536.0,1,-nbitq), 
to_sfixed(1200.0/65536.0,1,-nbitq), 
to_sfixed(5008.0/65536.0,1,-nbitq), 
to_sfixed(876.0/65536.0,1,-nbitq), 
to_sfixed(-305.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1441.0/65536.0,1,-nbitq), 
to_sfixed(-2419.0/65536.0,1,-nbitq), 
to_sfixed(-1574.0/65536.0,1,-nbitq), 
to_sfixed(-2320.0/65536.0,1,-nbitq), 
to_sfixed(-4217.0/65536.0,1,-nbitq), 
to_sfixed(-853.0/65536.0,1,-nbitq), 
to_sfixed(-2285.0/65536.0,1,-nbitq), 
to_sfixed(-1618.0/65536.0,1,-nbitq), 
to_sfixed(-3327.0/65536.0,1,-nbitq), 
to_sfixed(-883.0/65536.0,1,-nbitq), 
to_sfixed(-4348.0/65536.0,1,-nbitq), 
to_sfixed(1718.0/65536.0,1,-nbitq), 
to_sfixed(-2299.0/65536.0,1,-nbitq), 
to_sfixed(-2206.0/65536.0,1,-nbitq), 
to_sfixed(-172.0/65536.0,1,-nbitq), 
to_sfixed(303.0/65536.0,1,-nbitq), 
to_sfixed(-695.0/65536.0,1,-nbitq), 
to_sfixed(2181.0/65536.0,1,-nbitq), 
to_sfixed(967.0/65536.0,1,-nbitq), 
to_sfixed(-47.0/65536.0,1,-nbitq), 
to_sfixed(-359.0/65536.0,1,-nbitq), 
to_sfixed(-1008.0/65536.0,1,-nbitq), 
to_sfixed(3816.0/65536.0,1,-nbitq), 
to_sfixed(3119.0/65536.0,1,-nbitq), 
to_sfixed(1137.0/65536.0,1,-nbitq), 
to_sfixed(2653.0/65536.0,1,-nbitq), 
to_sfixed(-345.0/65536.0,1,-nbitq), 
to_sfixed(1240.0/65536.0,1,-nbitq), 
to_sfixed(-2713.0/65536.0,1,-nbitq), 
to_sfixed(-265.0/65536.0,1,-nbitq), 
to_sfixed(-2975.0/65536.0,1,-nbitq), 
to_sfixed(1172.0/65536.0,1,-nbitq), 
to_sfixed(-2935.0/65536.0,1,-nbitq), 
to_sfixed(-2549.0/65536.0,1,-nbitq), 
to_sfixed(324.0/65536.0,1,-nbitq), 
to_sfixed(731.0/65536.0,1,-nbitq), 
to_sfixed(-2155.0/65536.0,1,-nbitq), 
to_sfixed(2107.0/65536.0,1,-nbitq), 
to_sfixed(4846.0/65536.0,1,-nbitq), 
to_sfixed(219.0/65536.0,1,-nbitq), 
to_sfixed(1580.0/65536.0,1,-nbitq), 
to_sfixed(-3205.0/65536.0,1,-nbitq), 
to_sfixed(-5375.0/65536.0,1,-nbitq), 
to_sfixed(-2377.0/65536.0,1,-nbitq), 
to_sfixed(3307.0/65536.0,1,-nbitq), 
to_sfixed(4172.0/65536.0,1,-nbitq), 
to_sfixed(-2934.0/65536.0,1,-nbitq), 
to_sfixed(-73.0/65536.0,1,-nbitq), 
to_sfixed(199.0/65536.0,1,-nbitq), 
to_sfixed(2101.0/65536.0,1,-nbitq), 
to_sfixed(-2325.0/65536.0,1,-nbitq), 
to_sfixed(1571.0/65536.0,1,-nbitq), 
to_sfixed(-628.0/65536.0,1,-nbitq), 
to_sfixed(-209.0/65536.0,1,-nbitq), 
to_sfixed(2477.0/65536.0,1,-nbitq), 
to_sfixed(219.0/65536.0,1,-nbitq), 
to_sfixed(1520.0/65536.0,1,-nbitq), 
to_sfixed(1643.0/65536.0,1,-nbitq), 
to_sfixed(1823.0/65536.0,1,-nbitq), 
to_sfixed(-392.0/65536.0,1,-nbitq), 
to_sfixed(883.0/65536.0,1,-nbitq), 
to_sfixed(-1380.0/65536.0,1,-nbitq), 
to_sfixed(2839.0/65536.0,1,-nbitq), 
to_sfixed(-2641.0/65536.0,1,-nbitq), 
to_sfixed(3071.0/65536.0,1,-nbitq), 
to_sfixed(2834.0/65536.0,1,-nbitq), 
to_sfixed(3076.0/65536.0,1,-nbitq), 
to_sfixed(-2597.0/65536.0,1,-nbitq), 
to_sfixed(1.0/65536.0,1,-nbitq), 
to_sfixed(188.0/65536.0,1,-nbitq), 
to_sfixed(-1686.0/65536.0,1,-nbitq), 
to_sfixed(-425.0/65536.0,1,-nbitq), 
to_sfixed(-394.0/65536.0,1,-nbitq), 
to_sfixed(-820.0/65536.0,1,-nbitq), 
to_sfixed(1872.0/65536.0,1,-nbitq), 
to_sfixed(-2210.0/65536.0,1,-nbitq), 
to_sfixed(1428.0/65536.0,1,-nbitq), 
to_sfixed(2818.0/65536.0,1,-nbitq), 
to_sfixed(2697.0/65536.0,1,-nbitq), 
to_sfixed(-166.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2914.0/65536.0,1,-nbitq), 
to_sfixed(1938.0/65536.0,1,-nbitq), 
to_sfixed(10.0/65536.0,1,-nbitq), 
to_sfixed(-3893.0/65536.0,1,-nbitq), 
to_sfixed(1111.0/65536.0,1,-nbitq), 
to_sfixed(1095.0/65536.0,1,-nbitq), 
to_sfixed(841.0/65536.0,1,-nbitq), 
to_sfixed(-727.0/65536.0,1,-nbitq), 
to_sfixed(1782.0/65536.0,1,-nbitq), 
to_sfixed(-278.0/65536.0,1,-nbitq), 
to_sfixed(-3171.0/65536.0,1,-nbitq), 
to_sfixed(3788.0/65536.0,1,-nbitq), 
to_sfixed(-1857.0/65536.0,1,-nbitq), 
to_sfixed(-3675.0/65536.0,1,-nbitq), 
to_sfixed(-105.0/65536.0,1,-nbitq), 
to_sfixed(-2514.0/65536.0,1,-nbitq), 
to_sfixed(1817.0/65536.0,1,-nbitq), 
to_sfixed(4052.0/65536.0,1,-nbitq), 
to_sfixed(1995.0/65536.0,1,-nbitq), 
to_sfixed(410.0/65536.0,1,-nbitq), 
to_sfixed(-1063.0/65536.0,1,-nbitq), 
to_sfixed(3742.0/65536.0,1,-nbitq), 
to_sfixed(3552.0/65536.0,1,-nbitq), 
to_sfixed(2283.0/65536.0,1,-nbitq), 
to_sfixed(-1951.0/65536.0,1,-nbitq), 
to_sfixed(914.0/65536.0,1,-nbitq), 
to_sfixed(1171.0/65536.0,1,-nbitq), 
to_sfixed(604.0/65536.0,1,-nbitq), 
to_sfixed(-3099.0/65536.0,1,-nbitq), 
to_sfixed(-1324.0/65536.0,1,-nbitq), 
to_sfixed(54.0/65536.0,1,-nbitq), 
to_sfixed(-2942.0/65536.0,1,-nbitq), 
to_sfixed(-1440.0/65536.0,1,-nbitq), 
to_sfixed(-2156.0/65536.0,1,-nbitq), 
to_sfixed(-1019.0/65536.0,1,-nbitq), 
to_sfixed(-2440.0/65536.0,1,-nbitq), 
to_sfixed(3387.0/65536.0,1,-nbitq), 
to_sfixed(-3482.0/65536.0,1,-nbitq), 
to_sfixed(6734.0/65536.0,1,-nbitq), 
to_sfixed(-946.0/65536.0,1,-nbitq), 
to_sfixed(3100.0/65536.0,1,-nbitq), 
to_sfixed(-2666.0/65536.0,1,-nbitq), 
to_sfixed(-633.0/65536.0,1,-nbitq), 
to_sfixed(206.0/65536.0,1,-nbitq), 
to_sfixed(3111.0/65536.0,1,-nbitq), 
to_sfixed(2749.0/65536.0,1,-nbitq), 
to_sfixed(1778.0/65536.0,1,-nbitq), 
to_sfixed(1722.0/65536.0,1,-nbitq), 
to_sfixed(2326.0/65536.0,1,-nbitq), 
to_sfixed(421.0/65536.0,1,-nbitq), 
to_sfixed(1489.0/65536.0,1,-nbitq), 
to_sfixed(1489.0/65536.0,1,-nbitq), 
to_sfixed(-4016.0/65536.0,1,-nbitq), 
to_sfixed(683.0/65536.0,1,-nbitq), 
to_sfixed(2969.0/65536.0,1,-nbitq), 
to_sfixed(1681.0/65536.0,1,-nbitq), 
to_sfixed(-782.0/65536.0,1,-nbitq), 
to_sfixed(-2546.0/65536.0,1,-nbitq), 
to_sfixed(1053.0/65536.0,1,-nbitq), 
to_sfixed(-787.0/65536.0,1,-nbitq), 
to_sfixed(1431.0/65536.0,1,-nbitq), 
to_sfixed(1862.0/65536.0,1,-nbitq), 
to_sfixed(3079.0/65536.0,1,-nbitq), 
to_sfixed(1639.0/65536.0,1,-nbitq), 
to_sfixed(-1761.0/65536.0,1,-nbitq), 
to_sfixed(3688.0/65536.0,1,-nbitq), 
to_sfixed(728.0/65536.0,1,-nbitq), 
to_sfixed(-2579.0/65536.0,1,-nbitq), 
to_sfixed(3269.0/65536.0,1,-nbitq), 
to_sfixed(2434.0/65536.0,1,-nbitq), 
to_sfixed(2151.0/65536.0,1,-nbitq), 
to_sfixed(-1221.0/65536.0,1,-nbitq), 
to_sfixed(1311.0/65536.0,1,-nbitq), 
to_sfixed(-2211.0/65536.0,1,-nbitq), 
to_sfixed(66.0/65536.0,1,-nbitq), 
to_sfixed(1707.0/65536.0,1,-nbitq), 
to_sfixed(-741.0/65536.0,1,-nbitq), 
to_sfixed(5414.0/65536.0,1,-nbitq), 
to_sfixed(1950.0/65536.0,1,-nbitq), 
to_sfixed(2047.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1432.0/65536.0,1,-nbitq), 
to_sfixed(-1327.0/65536.0,1,-nbitq), 
to_sfixed(1141.0/65536.0,1,-nbitq), 
to_sfixed(-798.0/65536.0,1,-nbitq), 
to_sfixed(-3179.0/65536.0,1,-nbitq), 
to_sfixed(-760.0/65536.0,1,-nbitq), 
to_sfixed(1044.0/65536.0,1,-nbitq), 
to_sfixed(-810.0/65536.0,1,-nbitq), 
to_sfixed(2214.0/65536.0,1,-nbitq), 
to_sfixed(-1629.0/65536.0,1,-nbitq), 
to_sfixed(-4309.0/65536.0,1,-nbitq), 
to_sfixed(1741.0/65536.0,1,-nbitq), 
to_sfixed(-1004.0/65536.0,1,-nbitq), 
to_sfixed(1015.0/65536.0,1,-nbitq), 
to_sfixed(1157.0/65536.0,1,-nbitq), 
to_sfixed(2642.0/65536.0,1,-nbitq), 
to_sfixed(-2550.0/65536.0,1,-nbitq), 
to_sfixed(1816.0/65536.0,1,-nbitq), 
to_sfixed(1884.0/65536.0,1,-nbitq), 
to_sfixed(-1969.0/65536.0,1,-nbitq), 
to_sfixed(-5581.0/65536.0,1,-nbitq), 
to_sfixed(-3453.0/65536.0,1,-nbitq), 
to_sfixed(-884.0/65536.0,1,-nbitq), 
to_sfixed(-80.0/65536.0,1,-nbitq), 
to_sfixed(-1552.0/65536.0,1,-nbitq), 
to_sfixed(-1764.0/65536.0,1,-nbitq), 
to_sfixed(620.0/65536.0,1,-nbitq), 
to_sfixed(2281.0/65536.0,1,-nbitq), 
to_sfixed(-2996.0/65536.0,1,-nbitq), 
to_sfixed(4553.0/65536.0,1,-nbitq), 
to_sfixed(-1572.0/65536.0,1,-nbitq), 
to_sfixed(-3588.0/65536.0,1,-nbitq), 
to_sfixed(-2689.0/65536.0,1,-nbitq), 
to_sfixed(-3257.0/65536.0,1,-nbitq), 
to_sfixed(-1757.0/65536.0,1,-nbitq), 
to_sfixed(-2144.0/65536.0,1,-nbitq), 
to_sfixed(-1944.0/65536.0,1,-nbitq), 
to_sfixed(-730.0/65536.0,1,-nbitq), 
to_sfixed(4790.0/65536.0,1,-nbitq), 
to_sfixed(2720.0/65536.0,1,-nbitq), 
to_sfixed(464.0/65536.0,1,-nbitq), 
to_sfixed(113.0/65536.0,1,-nbitq), 
to_sfixed(-4030.0/65536.0,1,-nbitq), 
to_sfixed(860.0/65536.0,1,-nbitq), 
to_sfixed(19.0/65536.0,1,-nbitq), 
to_sfixed(5026.0/65536.0,1,-nbitq), 
to_sfixed(1167.0/65536.0,1,-nbitq), 
to_sfixed(375.0/65536.0,1,-nbitq), 
to_sfixed(-1815.0/65536.0,1,-nbitq), 
to_sfixed(3089.0/65536.0,1,-nbitq), 
to_sfixed(3043.0/65536.0,1,-nbitq), 
to_sfixed(-578.0/65536.0,1,-nbitq), 
to_sfixed(-3741.0/65536.0,1,-nbitq), 
to_sfixed(-2590.0/65536.0,1,-nbitq), 
to_sfixed(299.0/65536.0,1,-nbitq), 
to_sfixed(2406.0/65536.0,1,-nbitq), 
to_sfixed(321.0/65536.0,1,-nbitq), 
to_sfixed(510.0/65536.0,1,-nbitq), 
to_sfixed(1519.0/65536.0,1,-nbitq), 
to_sfixed(962.0/65536.0,1,-nbitq), 
to_sfixed(2450.0/65536.0,1,-nbitq), 
to_sfixed(-890.0/65536.0,1,-nbitq), 
to_sfixed(582.0/65536.0,1,-nbitq), 
to_sfixed(-2730.0/65536.0,1,-nbitq), 
to_sfixed(2901.0/65536.0,1,-nbitq), 
to_sfixed(484.0/65536.0,1,-nbitq), 
to_sfixed(2886.0/65536.0,1,-nbitq), 
to_sfixed(1132.0/65536.0,1,-nbitq), 
to_sfixed(-2050.0/65536.0,1,-nbitq), 
to_sfixed(1890.0/65536.0,1,-nbitq), 
to_sfixed(2820.0/65536.0,1,-nbitq), 
to_sfixed(2458.0/65536.0,1,-nbitq), 
to_sfixed(-2161.0/65536.0,1,-nbitq), 
to_sfixed(-1417.0/65536.0,1,-nbitq), 
to_sfixed(-635.0/65536.0,1,-nbitq), 
to_sfixed(-1341.0/65536.0,1,-nbitq), 
to_sfixed(-1269.0/65536.0,1,-nbitq), 
to_sfixed(355.0/65536.0,1,-nbitq), 
to_sfixed(-776.0/65536.0,1,-nbitq), 
to_sfixed(4844.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-759.0/65536.0,1,-nbitq), 
to_sfixed(-2203.0/65536.0,1,-nbitq), 
to_sfixed(-1087.0/65536.0,1,-nbitq), 
to_sfixed(-4936.0/65536.0,1,-nbitq), 
to_sfixed(-3858.0/65536.0,1,-nbitq), 
to_sfixed(-3143.0/65536.0,1,-nbitq), 
to_sfixed(1456.0/65536.0,1,-nbitq), 
to_sfixed(-3821.0/65536.0,1,-nbitq), 
to_sfixed(1852.0/65536.0,1,-nbitq), 
to_sfixed(-605.0/65536.0,1,-nbitq), 
to_sfixed(-3799.0/65536.0,1,-nbitq), 
to_sfixed(3823.0/65536.0,1,-nbitq), 
to_sfixed(-562.0/65536.0,1,-nbitq), 
to_sfixed(-779.0/65536.0,1,-nbitq), 
to_sfixed(2932.0/65536.0,1,-nbitq), 
to_sfixed(3185.0/65536.0,1,-nbitq), 
to_sfixed(-2221.0/65536.0,1,-nbitq), 
to_sfixed(308.0/65536.0,1,-nbitq), 
to_sfixed(3409.0/65536.0,1,-nbitq), 
to_sfixed(3087.0/65536.0,1,-nbitq), 
to_sfixed(-5083.0/65536.0,1,-nbitq), 
to_sfixed(-2916.0/65536.0,1,-nbitq), 
to_sfixed(2172.0/65536.0,1,-nbitq), 
to_sfixed(-311.0/65536.0,1,-nbitq), 
to_sfixed(-961.0/65536.0,1,-nbitq), 
to_sfixed(1059.0/65536.0,1,-nbitq), 
to_sfixed(-678.0/65536.0,1,-nbitq), 
to_sfixed(-1708.0/65536.0,1,-nbitq), 
to_sfixed(87.0/65536.0,1,-nbitq), 
to_sfixed(3547.0/65536.0,1,-nbitq), 
to_sfixed(1759.0/65536.0,1,-nbitq), 
to_sfixed(-2628.0/65536.0,1,-nbitq), 
to_sfixed(-4271.0/65536.0,1,-nbitq), 
to_sfixed(-2780.0/65536.0,1,-nbitq), 
to_sfixed(2548.0/65536.0,1,-nbitq), 
to_sfixed(1690.0/65536.0,1,-nbitq), 
to_sfixed(-1583.0/65536.0,1,-nbitq), 
to_sfixed(1526.0/65536.0,1,-nbitq), 
to_sfixed(2038.0/65536.0,1,-nbitq), 
to_sfixed(-147.0/65536.0,1,-nbitq), 
to_sfixed(1177.0/65536.0,1,-nbitq), 
to_sfixed(-2868.0/65536.0,1,-nbitq), 
to_sfixed(-637.0/65536.0,1,-nbitq), 
to_sfixed(1793.0/65536.0,1,-nbitq), 
to_sfixed(3038.0/65536.0,1,-nbitq), 
to_sfixed(2034.0/65536.0,1,-nbitq), 
to_sfixed(-290.0/65536.0,1,-nbitq), 
to_sfixed(1951.0/65536.0,1,-nbitq), 
to_sfixed(2453.0/65536.0,1,-nbitq), 
to_sfixed(3437.0/65536.0,1,-nbitq), 
to_sfixed(678.0/65536.0,1,-nbitq), 
to_sfixed(3496.0/65536.0,1,-nbitq), 
to_sfixed(820.0/65536.0,1,-nbitq), 
to_sfixed(200.0/65536.0,1,-nbitq), 
to_sfixed(2384.0/65536.0,1,-nbitq), 
to_sfixed(-705.0/65536.0,1,-nbitq), 
to_sfixed(1502.0/65536.0,1,-nbitq), 
to_sfixed(1274.0/65536.0,1,-nbitq), 
to_sfixed(1984.0/65536.0,1,-nbitq), 
to_sfixed(3417.0/65536.0,1,-nbitq), 
to_sfixed(-338.0/65536.0,1,-nbitq), 
to_sfixed(2591.0/65536.0,1,-nbitq), 
to_sfixed(619.0/65536.0,1,-nbitq), 
to_sfixed(-1237.0/65536.0,1,-nbitq), 
to_sfixed(286.0/65536.0,1,-nbitq), 
to_sfixed(1614.0/65536.0,1,-nbitq), 
to_sfixed(-905.0/65536.0,1,-nbitq), 
to_sfixed(268.0/65536.0,1,-nbitq), 
to_sfixed(3337.0/65536.0,1,-nbitq), 
to_sfixed(1960.0/65536.0,1,-nbitq), 
to_sfixed(-2127.0/65536.0,1,-nbitq), 
to_sfixed(-98.0/65536.0,1,-nbitq), 
to_sfixed(659.0/65536.0,1,-nbitq), 
to_sfixed(1534.0/65536.0,1,-nbitq), 
to_sfixed(1986.0/65536.0,1,-nbitq), 
to_sfixed(936.0/65536.0,1,-nbitq), 
to_sfixed(3219.0/65536.0,1,-nbitq), 
to_sfixed(2937.0/65536.0,1,-nbitq), 
to_sfixed(376.0/65536.0,1,-nbitq), 
to_sfixed(2387.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2897.0/65536.0,1,-nbitq), 
to_sfixed(-1278.0/65536.0,1,-nbitq), 
to_sfixed(3995.0/65536.0,1,-nbitq), 
to_sfixed(-1903.0/65536.0,1,-nbitq), 
to_sfixed(-2120.0/65536.0,1,-nbitq), 
to_sfixed(-1073.0/65536.0,1,-nbitq), 
to_sfixed(-843.0/65536.0,1,-nbitq), 
to_sfixed(-354.0/65536.0,1,-nbitq), 
to_sfixed(83.0/65536.0,1,-nbitq), 
to_sfixed(-530.0/65536.0,1,-nbitq), 
to_sfixed(-3774.0/65536.0,1,-nbitq), 
to_sfixed(895.0/65536.0,1,-nbitq), 
to_sfixed(1092.0/65536.0,1,-nbitq), 
to_sfixed(-499.0/65536.0,1,-nbitq), 
to_sfixed(3024.0/65536.0,1,-nbitq), 
to_sfixed(-2609.0/65536.0,1,-nbitq), 
to_sfixed(-1221.0/65536.0,1,-nbitq), 
to_sfixed(-1344.0/65536.0,1,-nbitq), 
to_sfixed(-100.0/65536.0,1,-nbitq), 
to_sfixed(-1844.0/65536.0,1,-nbitq), 
to_sfixed(-4349.0/65536.0,1,-nbitq), 
to_sfixed(2862.0/65536.0,1,-nbitq), 
to_sfixed(533.0/65536.0,1,-nbitq), 
to_sfixed(-513.0/65536.0,1,-nbitq), 
to_sfixed(-632.0/65536.0,1,-nbitq), 
to_sfixed(166.0/65536.0,1,-nbitq), 
to_sfixed(-240.0/65536.0,1,-nbitq), 
to_sfixed(-1956.0/65536.0,1,-nbitq), 
to_sfixed(462.0/65536.0,1,-nbitq), 
to_sfixed(1976.0/65536.0,1,-nbitq), 
to_sfixed(-2513.0/65536.0,1,-nbitq), 
to_sfixed(-1927.0/65536.0,1,-nbitq), 
to_sfixed(-1129.0/65536.0,1,-nbitq), 
to_sfixed(1173.0/65536.0,1,-nbitq), 
to_sfixed(-625.0/65536.0,1,-nbitq), 
to_sfixed(-9.0/65536.0,1,-nbitq), 
to_sfixed(-517.0/65536.0,1,-nbitq), 
to_sfixed(1028.0/65536.0,1,-nbitq), 
to_sfixed(3057.0/65536.0,1,-nbitq), 
to_sfixed(2308.0/65536.0,1,-nbitq), 
to_sfixed(-679.0/65536.0,1,-nbitq), 
to_sfixed(-941.0/65536.0,1,-nbitq), 
to_sfixed(-364.0/65536.0,1,-nbitq), 
to_sfixed(753.0/65536.0,1,-nbitq), 
to_sfixed(330.0/65536.0,1,-nbitq), 
to_sfixed(4835.0/65536.0,1,-nbitq), 
to_sfixed(1646.0/65536.0,1,-nbitq), 
to_sfixed(3333.0/65536.0,1,-nbitq), 
to_sfixed(1638.0/65536.0,1,-nbitq), 
to_sfixed(-349.0/65536.0,1,-nbitq), 
to_sfixed(1303.0/65536.0,1,-nbitq), 
to_sfixed(944.0/65536.0,1,-nbitq), 
to_sfixed(-1640.0/65536.0,1,-nbitq), 
to_sfixed(-2180.0/65536.0,1,-nbitq), 
to_sfixed(5077.0/65536.0,1,-nbitq), 
to_sfixed(1030.0/65536.0,1,-nbitq), 
to_sfixed(-1035.0/65536.0,1,-nbitq), 
to_sfixed(1627.0/65536.0,1,-nbitq), 
to_sfixed(435.0/65536.0,1,-nbitq), 
to_sfixed(3074.0/65536.0,1,-nbitq), 
to_sfixed(-5008.0/65536.0,1,-nbitq), 
to_sfixed(-2236.0/65536.0,1,-nbitq), 
to_sfixed(1688.0/65536.0,1,-nbitq), 
to_sfixed(509.0/65536.0,1,-nbitq), 
to_sfixed(4019.0/65536.0,1,-nbitq), 
to_sfixed(3055.0/65536.0,1,-nbitq), 
to_sfixed(-999.0/65536.0,1,-nbitq), 
to_sfixed(1119.0/65536.0,1,-nbitq), 
to_sfixed(3112.0/65536.0,1,-nbitq), 
to_sfixed(-468.0/65536.0,1,-nbitq), 
to_sfixed(2850.0/65536.0,1,-nbitq), 
to_sfixed(640.0/65536.0,1,-nbitq), 
to_sfixed(163.0/65536.0,1,-nbitq), 
to_sfixed(1696.0/65536.0,1,-nbitq), 
to_sfixed(-2711.0/65536.0,1,-nbitq), 
to_sfixed(-597.0/65536.0,1,-nbitq), 
to_sfixed(-467.0/65536.0,1,-nbitq), 
to_sfixed(2214.0/65536.0,1,-nbitq), 
to_sfixed(-1257.0/65536.0,1,-nbitq), 
to_sfixed(1273.0/65536.0,1,-nbitq)  ), 
( to_sfixed(28.0/65536.0,1,-nbitq), 
to_sfixed(-2383.0/65536.0,1,-nbitq), 
to_sfixed(-237.0/65536.0,1,-nbitq), 
to_sfixed(-3015.0/65536.0,1,-nbitq), 
to_sfixed(-1266.0/65536.0,1,-nbitq), 
to_sfixed(862.0/65536.0,1,-nbitq), 
to_sfixed(43.0/65536.0,1,-nbitq), 
to_sfixed(-623.0/65536.0,1,-nbitq), 
to_sfixed(263.0/65536.0,1,-nbitq), 
to_sfixed(-2852.0/65536.0,1,-nbitq), 
to_sfixed(-3458.0/65536.0,1,-nbitq), 
to_sfixed(-677.0/65536.0,1,-nbitq), 
to_sfixed(-2541.0/65536.0,1,-nbitq), 
to_sfixed(294.0/65536.0,1,-nbitq), 
to_sfixed(1475.0/65536.0,1,-nbitq), 
to_sfixed(613.0/65536.0,1,-nbitq), 
to_sfixed(-3044.0/65536.0,1,-nbitq), 
to_sfixed(2138.0/65536.0,1,-nbitq), 
to_sfixed(2171.0/65536.0,1,-nbitq), 
to_sfixed(967.0/65536.0,1,-nbitq), 
to_sfixed(-559.0/65536.0,1,-nbitq), 
to_sfixed(-1207.0/65536.0,1,-nbitq), 
to_sfixed(2167.0/65536.0,1,-nbitq), 
to_sfixed(-1027.0/65536.0,1,-nbitq), 
to_sfixed(-187.0/65536.0,1,-nbitq), 
to_sfixed(2161.0/65536.0,1,-nbitq), 
to_sfixed(-2472.0/65536.0,1,-nbitq), 
to_sfixed(649.0/65536.0,1,-nbitq), 
to_sfixed(-416.0/65536.0,1,-nbitq), 
to_sfixed(-2664.0/65536.0,1,-nbitq), 
to_sfixed(1274.0/65536.0,1,-nbitq), 
to_sfixed(-3180.0/65536.0,1,-nbitq), 
to_sfixed(-1229.0/65536.0,1,-nbitq), 
to_sfixed(434.0/65536.0,1,-nbitq), 
to_sfixed(2970.0/65536.0,1,-nbitq), 
to_sfixed(-2858.0/65536.0,1,-nbitq), 
to_sfixed(103.0/65536.0,1,-nbitq), 
to_sfixed(-143.0/65536.0,1,-nbitq), 
to_sfixed(591.0/65536.0,1,-nbitq), 
to_sfixed(277.0/65536.0,1,-nbitq), 
to_sfixed(-2614.0/65536.0,1,-nbitq), 
to_sfixed(-543.0/65536.0,1,-nbitq), 
to_sfixed(-3225.0/65536.0,1,-nbitq), 
to_sfixed(863.0/65536.0,1,-nbitq), 
to_sfixed(171.0/65536.0,1,-nbitq), 
to_sfixed(35.0/65536.0,1,-nbitq), 
to_sfixed(-1993.0/65536.0,1,-nbitq), 
to_sfixed(230.0/65536.0,1,-nbitq), 
to_sfixed(2524.0/65536.0,1,-nbitq), 
to_sfixed(-1147.0/65536.0,1,-nbitq), 
to_sfixed(2156.0/65536.0,1,-nbitq), 
to_sfixed(-2243.0/65536.0,1,-nbitq), 
to_sfixed(-1692.0/65536.0,1,-nbitq), 
to_sfixed(-3206.0/65536.0,1,-nbitq), 
to_sfixed(488.0/65536.0,1,-nbitq), 
to_sfixed(315.0/65536.0,1,-nbitq), 
to_sfixed(2251.0/65536.0,1,-nbitq), 
to_sfixed(2827.0/65536.0,1,-nbitq), 
to_sfixed(-2759.0/65536.0,1,-nbitq), 
to_sfixed(541.0/65536.0,1,-nbitq), 
to_sfixed(-1794.0/65536.0,1,-nbitq), 
to_sfixed(-1498.0/65536.0,1,-nbitq), 
to_sfixed(1948.0/65536.0,1,-nbitq), 
to_sfixed(-2871.0/65536.0,1,-nbitq), 
to_sfixed(-255.0/65536.0,1,-nbitq), 
to_sfixed(9.0/65536.0,1,-nbitq), 
to_sfixed(164.0/65536.0,1,-nbitq), 
to_sfixed(938.0/65536.0,1,-nbitq), 
to_sfixed(556.0/65536.0,1,-nbitq), 
to_sfixed(-2005.0/65536.0,1,-nbitq), 
to_sfixed(2780.0/65536.0,1,-nbitq), 
to_sfixed(-1622.0/65536.0,1,-nbitq), 
to_sfixed(2630.0/65536.0,1,-nbitq), 
to_sfixed(-1073.0/65536.0,1,-nbitq), 
to_sfixed(-1094.0/65536.0,1,-nbitq), 
to_sfixed(4062.0/65536.0,1,-nbitq), 
to_sfixed(28.0/65536.0,1,-nbitq), 
to_sfixed(2034.0/65536.0,1,-nbitq), 
to_sfixed(-1075.0/65536.0,1,-nbitq), 
to_sfixed(2242.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-395.0/65536.0,1,-nbitq), 
to_sfixed(-1397.0/65536.0,1,-nbitq), 
to_sfixed(4414.0/65536.0,1,-nbitq), 
to_sfixed(-1092.0/65536.0,1,-nbitq), 
to_sfixed(266.0/65536.0,1,-nbitq), 
to_sfixed(-4437.0/65536.0,1,-nbitq), 
to_sfixed(1965.0/65536.0,1,-nbitq), 
to_sfixed(-840.0/65536.0,1,-nbitq), 
to_sfixed(-745.0/65536.0,1,-nbitq), 
to_sfixed(-2403.0/65536.0,1,-nbitq), 
to_sfixed(-2475.0/65536.0,1,-nbitq), 
to_sfixed(333.0/65536.0,1,-nbitq), 
to_sfixed(-1910.0/65536.0,1,-nbitq), 
to_sfixed(-2970.0/65536.0,1,-nbitq), 
to_sfixed(2014.0/65536.0,1,-nbitq), 
to_sfixed(-1736.0/65536.0,1,-nbitq), 
to_sfixed(-2183.0/65536.0,1,-nbitq), 
to_sfixed(1121.0/65536.0,1,-nbitq), 
to_sfixed(-1260.0/65536.0,1,-nbitq), 
to_sfixed(2035.0/65536.0,1,-nbitq), 
to_sfixed(-2027.0/65536.0,1,-nbitq), 
to_sfixed(1953.0/65536.0,1,-nbitq), 
to_sfixed(1106.0/65536.0,1,-nbitq), 
to_sfixed(-648.0/65536.0,1,-nbitq), 
to_sfixed(-515.0/65536.0,1,-nbitq), 
to_sfixed(2251.0/65536.0,1,-nbitq), 
to_sfixed(-2152.0/65536.0,1,-nbitq), 
to_sfixed(2312.0/65536.0,1,-nbitq), 
to_sfixed(-1296.0/65536.0,1,-nbitq), 
to_sfixed(1671.0/65536.0,1,-nbitq), 
to_sfixed(1237.0/65536.0,1,-nbitq), 
to_sfixed(507.0/65536.0,1,-nbitq), 
to_sfixed(-3702.0/65536.0,1,-nbitq), 
to_sfixed(614.0/65536.0,1,-nbitq), 
to_sfixed(2967.0/65536.0,1,-nbitq), 
to_sfixed(-1647.0/65536.0,1,-nbitq), 
to_sfixed(2669.0/65536.0,1,-nbitq), 
to_sfixed(-2373.0/65536.0,1,-nbitq), 
to_sfixed(396.0/65536.0,1,-nbitq), 
to_sfixed(-373.0/65536.0,1,-nbitq), 
to_sfixed(-1657.0/65536.0,1,-nbitq), 
to_sfixed(1238.0/65536.0,1,-nbitq), 
to_sfixed(-1254.0/65536.0,1,-nbitq), 
to_sfixed(-837.0/65536.0,1,-nbitq), 
to_sfixed(1690.0/65536.0,1,-nbitq), 
to_sfixed(2238.0/65536.0,1,-nbitq), 
to_sfixed(295.0/65536.0,1,-nbitq), 
to_sfixed(-1550.0/65536.0,1,-nbitq), 
to_sfixed(2237.0/65536.0,1,-nbitq), 
to_sfixed(718.0/65536.0,1,-nbitq), 
to_sfixed(2270.0/65536.0,1,-nbitq), 
to_sfixed(-1412.0/65536.0,1,-nbitq), 
to_sfixed(-2285.0/65536.0,1,-nbitq), 
to_sfixed(-1562.0/65536.0,1,-nbitq), 
to_sfixed(4969.0/65536.0,1,-nbitq), 
to_sfixed(-1403.0/65536.0,1,-nbitq), 
to_sfixed(-2173.0/65536.0,1,-nbitq), 
to_sfixed(1910.0/65536.0,1,-nbitq), 
to_sfixed(-2833.0/65536.0,1,-nbitq), 
to_sfixed(1401.0/65536.0,1,-nbitq), 
to_sfixed(-6118.0/65536.0,1,-nbitq), 
to_sfixed(-50.0/65536.0,1,-nbitq), 
to_sfixed(1651.0/65536.0,1,-nbitq), 
to_sfixed(-1050.0/65536.0,1,-nbitq), 
to_sfixed(2062.0/65536.0,1,-nbitq), 
to_sfixed(-101.0/65536.0,1,-nbitq), 
to_sfixed(-1020.0/65536.0,1,-nbitq), 
to_sfixed(-1357.0/65536.0,1,-nbitq), 
to_sfixed(-70.0/65536.0,1,-nbitq), 
to_sfixed(-1874.0/65536.0,1,-nbitq), 
to_sfixed(-2331.0/65536.0,1,-nbitq), 
to_sfixed(-492.0/65536.0,1,-nbitq), 
to_sfixed(3114.0/65536.0,1,-nbitq), 
to_sfixed(-1662.0/65536.0,1,-nbitq), 
to_sfixed(2314.0/65536.0,1,-nbitq), 
to_sfixed(1220.0/65536.0,1,-nbitq), 
to_sfixed(3055.0/65536.0,1,-nbitq), 
to_sfixed(4138.0/65536.0,1,-nbitq), 
to_sfixed(567.0/65536.0,1,-nbitq), 
to_sfixed(3507.0/65536.0,1,-nbitq)  ), 
( to_sfixed(542.0/65536.0,1,-nbitq), 
to_sfixed(-1934.0/65536.0,1,-nbitq), 
to_sfixed(-400.0/65536.0,1,-nbitq), 
to_sfixed(-1599.0/65536.0,1,-nbitq), 
to_sfixed(-3038.0/65536.0,1,-nbitq), 
to_sfixed(-9.0/65536.0,1,-nbitq), 
to_sfixed(-821.0/65536.0,1,-nbitq), 
to_sfixed(-3265.0/65536.0,1,-nbitq), 
to_sfixed(-1796.0/65536.0,1,-nbitq), 
to_sfixed(449.0/65536.0,1,-nbitq), 
to_sfixed(1778.0/65536.0,1,-nbitq), 
to_sfixed(2661.0/65536.0,1,-nbitq), 
to_sfixed(-88.0/65536.0,1,-nbitq), 
to_sfixed(618.0/65536.0,1,-nbitq), 
to_sfixed(761.0/65536.0,1,-nbitq), 
to_sfixed(-2763.0/65536.0,1,-nbitq), 
to_sfixed(-597.0/65536.0,1,-nbitq), 
to_sfixed(1209.0/65536.0,1,-nbitq), 
to_sfixed(-1366.0/65536.0,1,-nbitq), 
to_sfixed(405.0/65536.0,1,-nbitq), 
to_sfixed(400.0/65536.0,1,-nbitq), 
to_sfixed(-1120.0/65536.0,1,-nbitq), 
to_sfixed(3832.0/65536.0,1,-nbitq), 
to_sfixed(2010.0/65536.0,1,-nbitq), 
to_sfixed(-4143.0/65536.0,1,-nbitq), 
to_sfixed(1833.0/65536.0,1,-nbitq), 
to_sfixed(-136.0/65536.0,1,-nbitq), 
to_sfixed(-1384.0/65536.0,1,-nbitq), 
to_sfixed(-279.0/65536.0,1,-nbitq), 
to_sfixed(2854.0/65536.0,1,-nbitq), 
to_sfixed(-2214.0/65536.0,1,-nbitq), 
to_sfixed(1295.0/65536.0,1,-nbitq), 
to_sfixed(-376.0/65536.0,1,-nbitq), 
to_sfixed(-4114.0/65536.0,1,-nbitq), 
to_sfixed(-645.0/65536.0,1,-nbitq), 
to_sfixed(1242.0/65536.0,1,-nbitq), 
to_sfixed(2784.0/65536.0,1,-nbitq), 
to_sfixed(-2957.0/65536.0,1,-nbitq), 
to_sfixed(-1735.0/65536.0,1,-nbitq), 
to_sfixed(1228.0/65536.0,1,-nbitq), 
to_sfixed(-2297.0/65536.0,1,-nbitq), 
to_sfixed(1978.0/65536.0,1,-nbitq), 
to_sfixed(-2504.0/65536.0,1,-nbitq), 
to_sfixed(3022.0/65536.0,1,-nbitq), 
to_sfixed(-1250.0/65536.0,1,-nbitq), 
to_sfixed(4923.0/65536.0,1,-nbitq), 
to_sfixed(-382.0/65536.0,1,-nbitq), 
to_sfixed(-493.0/65536.0,1,-nbitq), 
to_sfixed(1611.0/65536.0,1,-nbitq), 
to_sfixed(885.0/65536.0,1,-nbitq), 
to_sfixed(1358.0/65536.0,1,-nbitq), 
to_sfixed(-1103.0/65536.0,1,-nbitq), 
to_sfixed(-3500.0/65536.0,1,-nbitq), 
to_sfixed(1738.0/65536.0,1,-nbitq), 
to_sfixed(-805.0/65536.0,1,-nbitq), 
to_sfixed(2046.0/65536.0,1,-nbitq), 
to_sfixed(755.0/65536.0,1,-nbitq), 
to_sfixed(3069.0/65536.0,1,-nbitq), 
to_sfixed(2002.0/65536.0,1,-nbitq), 
to_sfixed(-546.0/65536.0,1,-nbitq), 
to_sfixed(-706.0/65536.0,1,-nbitq), 
to_sfixed(-1933.0/65536.0,1,-nbitq), 
to_sfixed(2463.0/65536.0,1,-nbitq), 
to_sfixed(-1592.0/65536.0,1,-nbitq), 
to_sfixed(-1583.0/65536.0,1,-nbitq), 
to_sfixed(-1418.0/65536.0,1,-nbitq), 
to_sfixed(-520.0/65536.0,1,-nbitq), 
to_sfixed(-3193.0/65536.0,1,-nbitq), 
to_sfixed(796.0/65536.0,1,-nbitq), 
to_sfixed(887.0/65536.0,1,-nbitq), 
to_sfixed(804.0/65536.0,1,-nbitq), 
to_sfixed(-3429.0/65536.0,1,-nbitq), 
to_sfixed(999.0/65536.0,1,-nbitq), 
to_sfixed(-3206.0/65536.0,1,-nbitq), 
to_sfixed(2159.0/65536.0,1,-nbitq), 
to_sfixed(1823.0/65536.0,1,-nbitq), 
to_sfixed(88.0/65536.0,1,-nbitq), 
to_sfixed(3641.0/65536.0,1,-nbitq), 
to_sfixed(-407.0/65536.0,1,-nbitq), 
to_sfixed(2237.0/65536.0,1,-nbitq)  ), 
( to_sfixed(1553.0/65536.0,1,-nbitq), 
to_sfixed(2673.0/65536.0,1,-nbitq), 
to_sfixed(2061.0/65536.0,1,-nbitq), 
to_sfixed(-262.0/65536.0,1,-nbitq), 
to_sfixed(463.0/65536.0,1,-nbitq), 
to_sfixed(-4557.0/65536.0,1,-nbitq), 
to_sfixed(-3213.0/65536.0,1,-nbitq), 
to_sfixed(1145.0/65536.0,1,-nbitq), 
to_sfixed(1973.0/65536.0,1,-nbitq), 
to_sfixed(904.0/65536.0,1,-nbitq), 
to_sfixed(-167.0/65536.0,1,-nbitq), 
to_sfixed(833.0/65536.0,1,-nbitq), 
to_sfixed(542.0/65536.0,1,-nbitq), 
to_sfixed(-3197.0/65536.0,1,-nbitq), 
to_sfixed(-1815.0/65536.0,1,-nbitq), 
to_sfixed(-694.0/65536.0,1,-nbitq), 
to_sfixed(-2404.0/65536.0,1,-nbitq), 
to_sfixed(3313.0/65536.0,1,-nbitq), 
to_sfixed(923.0/65536.0,1,-nbitq), 
to_sfixed(2466.0/65536.0,1,-nbitq), 
to_sfixed(-2740.0/65536.0,1,-nbitq), 
to_sfixed(2521.0/65536.0,1,-nbitq), 
to_sfixed(73.0/65536.0,1,-nbitq), 
to_sfixed(884.0/65536.0,1,-nbitq), 
to_sfixed(1244.0/65536.0,1,-nbitq), 
to_sfixed(389.0/65536.0,1,-nbitq), 
to_sfixed(-3818.0/65536.0,1,-nbitq), 
to_sfixed(2784.0/65536.0,1,-nbitq), 
to_sfixed(-2669.0/65536.0,1,-nbitq), 
to_sfixed(2600.0/65536.0,1,-nbitq), 
to_sfixed(-2410.0/65536.0,1,-nbitq), 
to_sfixed(2056.0/65536.0,1,-nbitq), 
to_sfixed(-2096.0/65536.0,1,-nbitq), 
to_sfixed(-2996.0/65536.0,1,-nbitq), 
to_sfixed(-2829.0/65536.0,1,-nbitq), 
to_sfixed(2536.0/65536.0,1,-nbitq), 
to_sfixed(224.0/65536.0,1,-nbitq), 
to_sfixed(-2639.0/65536.0,1,-nbitq), 
to_sfixed(-3025.0/65536.0,1,-nbitq), 
to_sfixed(55.0/65536.0,1,-nbitq), 
to_sfixed(-2915.0/65536.0,1,-nbitq), 
to_sfixed(-2879.0/65536.0,1,-nbitq), 
to_sfixed(-3339.0/65536.0,1,-nbitq), 
to_sfixed(140.0/65536.0,1,-nbitq), 
to_sfixed(-611.0/65536.0,1,-nbitq), 
to_sfixed(2329.0/65536.0,1,-nbitq), 
to_sfixed(-1887.0/65536.0,1,-nbitq), 
to_sfixed(-1758.0/65536.0,1,-nbitq), 
to_sfixed(3388.0/65536.0,1,-nbitq), 
to_sfixed(12.0/65536.0,1,-nbitq), 
to_sfixed(2785.0/65536.0,1,-nbitq), 
to_sfixed(2528.0/65536.0,1,-nbitq), 
to_sfixed(-911.0/65536.0,1,-nbitq), 
to_sfixed(-1044.0/65536.0,1,-nbitq), 
to_sfixed(4271.0/65536.0,1,-nbitq), 
to_sfixed(1581.0/65536.0,1,-nbitq), 
to_sfixed(-1369.0/65536.0,1,-nbitq), 
to_sfixed(-1456.0/65536.0,1,-nbitq), 
to_sfixed(1122.0/65536.0,1,-nbitq), 
to_sfixed(369.0/65536.0,1,-nbitq), 
to_sfixed(1274.0/65536.0,1,-nbitq), 
to_sfixed(-938.0/65536.0,1,-nbitq), 
to_sfixed(1099.0/65536.0,1,-nbitq), 
to_sfixed(-670.0/65536.0,1,-nbitq), 
to_sfixed(24.0/65536.0,1,-nbitq), 
to_sfixed(1303.0/65536.0,1,-nbitq), 
to_sfixed(847.0/65536.0,1,-nbitq), 
to_sfixed(-3269.0/65536.0,1,-nbitq), 
to_sfixed(2442.0/65536.0,1,-nbitq), 
to_sfixed(-1081.0/65536.0,1,-nbitq), 
to_sfixed(-1324.0/65536.0,1,-nbitq), 
to_sfixed(510.0/65536.0,1,-nbitq), 
to_sfixed(335.0/65536.0,1,-nbitq), 
to_sfixed(-2930.0/65536.0,1,-nbitq), 
to_sfixed(-2168.0/65536.0,1,-nbitq), 
to_sfixed(3871.0/65536.0,1,-nbitq), 
to_sfixed(1989.0/65536.0,1,-nbitq), 
to_sfixed(2375.0/65536.0,1,-nbitq), 
to_sfixed(1257.0/65536.0,1,-nbitq), 
to_sfixed(203.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ), 
( to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq), 
to_sfixed(0.0/65536.0,1,-nbitq)  ) 
 ) ;

constant coef2 : typtabcnf2 := ( ( to_sfixed(-18377.0/65536.0,1,-nbitq), 
to_sfixed(-12879.0/65536.0,1,-nbitq), 
to_sfixed(14730.0/65536.0,1,-nbitq), 
to_sfixed(-8614.0/65536.0,1,-nbitq), 
to_sfixed(-9980.0/65536.0,1,-nbitq), 
to_sfixed(-10912.0/65536.0,1,-nbitq), 
to_sfixed(-15730.0/65536.0,1,-nbitq), 
to_sfixed(-10538.0/65536.0,1,-nbitq), 
to_sfixed(3632.0/65536.0,1,-nbitq), 
to_sfixed(-10428.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-17136.0/65536.0,1,-nbitq), 
to_sfixed(10990.0/65536.0,1,-nbitq), 
to_sfixed(15967.0/65536.0,1,-nbitq), 
to_sfixed(-16399.0/65536.0,1,-nbitq), 
to_sfixed(9058.0/65536.0,1,-nbitq), 
to_sfixed(2128.0/65536.0,1,-nbitq), 
to_sfixed(8046.0/65536.0,1,-nbitq), 
to_sfixed(8975.0/65536.0,1,-nbitq), 
to_sfixed(10135.0/65536.0,1,-nbitq), 
to_sfixed(4377.0/65536.0,1,-nbitq)  ), 
( to_sfixed(28448.0/65536.0,1,-nbitq), 
to_sfixed(7879.0/65536.0,1,-nbitq), 
to_sfixed(-15105.0/65536.0,1,-nbitq), 
to_sfixed(14547.0/65536.0,1,-nbitq), 
to_sfixed(-21157.0/65536.0,1,-nbitq), 
to_sfixed(11050.0/65536.0,1,-nbitq), 
to_sfixed(28557.0/65536.0,1,-nbitq), 
to_sfixed(-15363.0/65536.0,1,-nbitq), 
to_sfixed(-24922.0/65536.0,1,-nbitq), 
to_sfixed(12071.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-5765.0/65536.0,1,-nbitq), 
to_sfixed(-24259.0/65536.0,1,-nbitq), 
to_sfixed(-16543.0/65536.0,1,-nbitq), 
to_sfixed(16043.0/65536.0,1,-nbitq), 
to_sfixed(-3605.0/65536.0,1,-nbitq), 
to_sfixed(10212.0/65536.0,1,-nbitq), 
to_sfixed(-5895.0/65536.0,1,-nbitq), 
to_sfixed(16936.0/65536.0,1,-nbitq), 
to_sfixed(14894.0/65536.0,1,-nbitq), 
to_sfixed(9711.0/65536.0,1,-nbitq)  ), 
( to_sfixed(19256.0/65536.0,1,-nbitq), 
to_sfixed(1734.0/65536.0,1,-nbitq), 
to_sfixed(31573.0/65536.0,1,-nbitq), 
to_sfixed(22628.0/65536.0,1,-nbitq), 
to_sfixed(-7473.0/65536.0,1,-nbitq), 
to_sfixed(-363.0/65536.0,1,-nbitq), 
to_sfixed(-25922.0/65536.0,1,-nbitq), 
to_sfixed(-16356.0/65536.0,1,-nbitq), 
to_sfixed(4881.0/65536.0,1,-nbitq), 
to_sfixed(-14448.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-37658.0/65536.0,1,-nbitq), 
to_sfixed(-25372.0/65536.0,1,-nbitq), 
to_sfixed(-2992.0/65536.0,1,-nbitq), 
to_sfixed(-8023.0/65536.0,1,-nbitq), 
to_sfixed(10861.0/65536.0,1,-nbitq), 
to_sfixed(43024.0/65536.0,1,-nbitq), 
to_sfixed(-25327.0/65536.0,1,-nbitq), 
to_sfixed(11443.0/65536.0,1,-nbitq), 
to_sfixed(-9133.0/65536.0,1,-nbitq), 
to_sfixed(23836.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-11275.0/65536.0,1,-nbitq), 
to_sfixed(11898.0/65536.0,1,-nbitq), 
to_sfixed(17063.0/65536.0,1,-nbitq), 
to_sfixed(-10587.0/65536.0,1,-nbitq), 
to_sfixed(-5864.0/65536.0,1,-nbitq), 
to_sfixed(-20709.0/65536.0,1,-nbitq), 
to_sfixed(12368.0/65536.0,1,-nbitq), 
to_sfixed(-1925.0/65536.0,1,-nbitq), 
to_sfixed(18329.0/65536.0,1,-nbitq), 
to_sfixed(7252.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-24886.0/65536.0,1,-nbitq), 
to_sfixed(-5806.0/65536.0,1,-nbitq), 
to_sfixed(-19426.0/65536.0,1,-nbitq), 
to_sfixed(-14014.0/65536.0,1,-nbitq), 
to_sfixed(16223.0/65536.0,1,-nbitq), 
to_sfixed(-481.0/65536.0,1,-nbitq), 
to_sfixed(-14410.0/65536.0,1,-nbitq), 
to_sfixed(18772.0/65536.0,1,-nbitq), 
to_sfixed(7207.0/65536.0,1,-nbitq), 
to_sfixed(-3502.0/65536.0,1,-nbitq)  ), 
( to_sfixed(15905.0/65536.0,1,-nbitq), 
to_sfixed(15791.0/65536.0,1,-nbitq), 
to_sfixed(-9605.0/65536.0,1,-nbitq), 
to_sfixed(-7174.0/65536.0,1,-nbitq), 
to_sfixed(1793.0/65536.0,1,-nbitq), 
to_sfixed(14975.0/65536.0,1,-nbitq), 
to_sfixed(-18979.0/65536.0,1,-nbitq), 
to_sfixed(13577.0/65536.0,1,-nbitq), 
to_sfixed(-11097.0/65536.0,1,-nbitq), 
to_sfixed(-6125.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-837.0/65536.0,1,-nbitq), 
to_sfixed(-5401.0/65536.0,1,-nbitq), 
to_sfixed(826.0/65536.0,1,-nbitq), 
to_sfixed(-6662.0/65536.0,1,-nbitq), 
to_sfixed(-10303.0/65536.0,1,-nbitq), 
to_sfixed(101.0/65536.0,1,-nbitq), 
to_sfixed(-9594.0/65536.0,1,-nbitq), 
to_sfixed(11943.0/65536.0,1,-nbitq), 
to_sfixed(15898.0/65536.0,1,-nbitq), 
to_sfixed(-688.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-16589.0/65536.0,1,-nbitq), 
to_sfixed(4055.0/65536.0,1,-nbitq), 
to_sfixed(-5922.0/65536.0,1,-nbitq), 
to_sfixed(-2101.0/65536.0,1,-nbitq), 
to_sfixed(-12444.0/65536.0,1,-nbitq), 
to_sfixed(16305.0/65536.0,1,-nbitq), 
to_sfixed(-11732.0/65536.0,1,-nbitq), 
to_sfixed(11419.0/65536.0,1,-nbitq), 
to_sfixed(20672.0/65536.0,1,-nbitq), 
to_sfixed(-16592.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-29611.0/65536.0,1,-nbitq), 
to_sfixed(20768.0/65536.0,1,-nbitq), 
to_sfixed(16502.0/65536.0,1,-nbitq), 
to_sfixed(23524.0/65536.0,1,-nbitq), 
to_sfixed(-4592.0/65536.0,1,-nbitq), 
to_sfixed(16995.0/65536.0,1,-nbitq), 
to_sfixed(-14616.0/65536.0,1,-nbitq), 
to_sfixed(26590.0/65536.0,1,-nbitq), 
to_sfixed(-26683.0/65536.0,1,-nbitq), 
to_sfixed(-31516.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4320.0/65536.0,1,-nbitq), 
to_sfixed(-14944.0/65536.0,1,-nbitq), 
to_sfixed(-10346.0/65536.0,1,-nbitq), 
to_sfixed(-12931.0/65536.0,1,-nbitq), 
to_sfixed(-9263.0/65536.0,1,-nbitq), 
to_sfixed(11608.0/65536.0,1,-nbitq), 
to_sfixed(6832.0/65536.0,1,-nbitq), 
to_sfixed(16975.0/65536.0,1,-nbitq), 
to_sfixed(7526.0/65536.0,1,-nbitq), 
to_sfixed(-13757.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-28674.0/65536.0,1,-nbitq), 
to_sfixed(13476.0/65536.0,1,-nbitq), 
to_sfixed(-15207.0/65536.0,1,-nbitq), 
to_sfixed(15975.0/65536.0,1,-nbitq), 
to_sfixed(-5126.0/65536.0,1,-nbitq), 
to_sfixed(13066.0/65536.0,1,-nbitq), 
to_sfixed(-25882.0/65536.0,1,-nbitq), 
to_sfixed(114.0/65536.0,1,-nbitq), 
to_sfixed(18779.0/65536.0,1,-nbitq), 
to_sfixed(-13857.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5478.0/65536.0,1,-nbitq), 
to_sfixed(-14679.0/65536.0,1,-nbitq), 
to_sfixed(10419.0/65536.0,1,-nbitq), 
to_sfixed(-3700.0/65536.0,1,-nbitq), 
to_sfixed(-6607.0/65536.0,1,-nbitq), 
to_sfixed(10662.0/65536.0,1,-nbitq), 
to_sfixed(-846.0/65536.0,1,-nbitq), 
to_sfixed(-13726.0/65536.0,1,-nbitq), 
to_sfixed(-12474.0/65536.0,1,-nbitq), 
to_sfixed(19530.0/65536.0,1,-nbitq)  ), 
( to_sfixed(493.0/65536.0,1,-nbitq), 
to_sfixed(-7637.0/65536.0,1,-nbitq), 
to_sfixed(-14378.0/65536.0,1,-nbitq), 
to_sfixed(-4812.0/65536.0,1,-nbitq), 
to_sfixed(-9956.0/65536.0,1,-nbitq), 
to_sfixed(-1574.0/65536.0,1,-nbitq), 
to_sfixed(-4933.0/65536.0,1,-nbitq), 
to_sfixed(-8323.0/65536.0,1,-nbitq), 
to_sfixed(-3256.0/65536.0,1,-nbitq), 
to_sfixed(-6326.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-10207.0/65536.0,1,-nbitq), 
to_sfixed(2273.0/65536.0,1,-nbitq), 
to_sfixed(-10694.0/65536.0,1,-nbitq), 
to_sfixed(-10628.0/65536.0,1,-nbitq), 
to_sfixed(-10349.0/65536.0,1,-nbitq), 
to_sfixed(-17745.0/65536.0,1,-nbitq), 
to_sfixed(12888.0/65536.0,1,-nbitq), 
to_sfixed(1331.0/65536.0,1,-nbitq), 
to_sfixed(-16236.0/65536.0,1,-nbitq), 
to_sfixed(-13853.0/65536.0,1,-nbitq)  ), 
( to_sfixed(15021.0/65536.0,1,-nbitq), 
to_sfixed(-7093.0/65536.0,1,-nbitq), 
to_sfixed(-17406.0/65536.0,1,-nbitq), 
to_sfixed(-16554.0/65536.0,1,-nbitq), 
to_sfixed(13309.0/65536.0,1,-nbitq), 
to_sfixed(8307.0/65536.0,1,-nbitq), 
to_sfixed(-15216.0/65536.0,1,-nbitq), 
to_sfixed(12643.0/65536.0,1,-nbitq), 
to_sfixed(21167.0/65536.0,1,-nbitq), 
to_sfixed(20918.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-10444.0/65536.0,1,-nbitq), 
to_sfixed(3549.0/65536.0,1,-nbitq), 
to_sfixed(-20059.0/65536.0,1,-nbitq), 
to_sfixed(2785.0/65536.0,1,-nbitq), 
to_sfixed(-1427.0/65536.0,1,-nbitq), 
to_sfixed(1611.0/65536.0,1,-nbitq), 
to_sfixed(-18365.0/65536.0,1,-nbitq), 
to_sfixed(-18741.0/65536.0,1,-nbitq), 
to_sfixed(3552.0/65536.0,1,-nbitq), 
to_sfixed(24301.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5722.0/65536.0,1,-nbitq), 
to_sfixed(15018.0/65536.0,1,-nbitq), 
to_sfixed(-8483.0/65536.0,1,-nbitq), 
to_sfixed(-6296.0/65536.0,1,-nbitq), 
to_sfixed(12222.0/65536.0,1,-nbitq), 
to_sfixed(-12276.0/65536.0,1,-nbitq), 
to_sfixed(581.0/65536.0,1,-nbitq), 
to_sfixed(7896.0/65536.0,1,-nbitq), 
to_sfixed(950.0/65536.0,1,-nbitq), 
to_sfixed(5200.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-10871.0/65536.0,1,-nbitq), 
to_sfixed(-16391.0/65536.0,1,-nbitq), 
to_sfixed(15912.0/65536.0,1,-nbitq), 
to_sfixed(-24344.0/65536.0,1,-nbitq), 
to_sfixed(-7696.0/65536.0,1,-nbitq), 
to_sfixed(11970.0/65536.0,1,-nbitq), 
to_sfixed(68.0/65536.0,1,-nbitq), 
to_sfixed(755.0/65536.0,1,-nbitq), 
to_sfixed(15009.0/65536.0,1,-nbitq), 
to_sfixed(4288.0/65536.0,1,-nbitq)  ), 
( to_sfixed(21953.0/65536.0,1,-nbitq), 
to_sfixed(23870.0/65536.0,1,-nbitq), 
to_sfixed(-7924.0/65536.0,1,-nbitq), 
to_sfixed(-21939.0/65536.0,1,-nbitq), 
to_sfixed(-15149.0/65536.0,1,-nbitq), 
to_sfixed(-18915.0/65536.0,1,-nbitq), 
to_sfixed(15255.0/65536.0,1,-nbitq), 
to_sfixed(3947.0/65536.0,1,-nbitq), 
to_sfixed(-30063.0/65536.0,1,-nbitq), 
to_sfixed(19026.0/65536.0,1,-nbitq)  ), 
( to_sfixed(15354.0/65536.0,1,-nbitq), 
to_sfixed(37347.0/65536.0,1,-nbitq), 
to_sfixed(-17103.0/65536.0,1,-nbitq), 
to_sfixed(-8439.0/65536.0,1,-nbitq), 
to_sfixed(7660.0/65536.0,1,-nbitq), 
to_sfixed(-14329.0/65536.0,1,-nbitq), 
to_sfixed(16107.0/65536.0,1,-nbitq), 
to_sfixed(-18558.0/65536.0,1,-nbitq), 
to_sfixed(-25375.0/65536.0,1,-nbitq), 
to_sfixed(5597.0/65536.0,1,-nbitq)  ), 
( to_sfixed(17970.0/65536.0,1,-nbitq), 
to_sfixed(-11539.0/65536.0,1,-nbitq), 
to_sfixed(-30269.0/65536.0,1,-nbitq), 
to_sfixed(13847.0/65536.0,1,-nbitq), 
to_sfixed(7231.0/65536.0,1,-nbitq), 
to_sfixed(6075.0/65536.0,1,-nbitq), 
to_sfixed(-27106.0/65536.0,1,-nbitq), 
to_sfixed(-6568.0/65536.0,1,-nbitq), 
to_sfixed(-27771.0/65536.0,1,-nbitq), 
to_sfixed(6863.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-19738.0/65536.0,1,-nbitq), 
to_sfixed(-12997.0/65536.0,1,-nbitq), 
to_sfixed(-5110.0/65536.0,1,-nbitq), 
to_sfixed(-19690.0/65536.0,1,-nbitq), 
to_sfixed(20993.0/65536.0,1,-nbitq), 
to_sfixed(10697.0/65536.0,1,-nbitq), 
to_sfixed(4765.0/65536.0,1,-nbitq), 
to_sfixed(1097.0/65536.0,1,-nbitq), 
to_sfixed(625.0/65536.0,1,-nbitq), 
to_sfixed(2694.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-25938.0/65536.0,1,-nbitq), 
to_sfixed(-24424.0/65536.0,1,-nbitq), 
to_sfixed(-46949.0/65536.0,1,-nbitq), 
to_sfixed(25871.0/65536.0,1,-nbitq), 
to_sfixed(11051.0/65536.0,1,-nbitq), 
to_sfixed(37530.0/65536.0,1,-nbitq), 
to_sfixed(-7859.0/65536.0,1,-nbitq), 
to_sfixed(-12463.0/65536.0,1,-nbitq), 
to_sfixed(-8077.0/65536.0,1,-nbitq), 
to_sfixed(4426.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-4006.0/65536.0,1,-nbitq), 
to_sfixed(-30392.0/65536.0,1,-nbitq), 
to_sfixed(-5650.0/65536.0,1,-nbitq), 
to_sfixed(-1188.0/65536.0,1,-nbitq), 
to_sfixed(-27374.0/65536.0,1,-nbitq), 
to_sfixed(21693.0/65536.0,1,-nbitq), 
to_sfixed(-22461.0/65536.0,1,-nbitq), 
to_sfixed(26455.0/65536.0,1,-nbitq), 
to_sfixed(-12394.0/65536.0,1,-nbitq), 
to_sfixed(22797.0/65536.0,1,-nbitq)  ), 
( to_sfixed(15378.0/65536.0,1,-nbitq), 
to_sfixed(1255.0/65536.0,1,-nbitq), 
to_sfixed(-3075.0/65536.0,1,-nbitq), 
to_sfixed(9578.0/65536.0,1,-nbitq), 
to_sfixed(-3626.0/65536.0,1,-nbitq), 
to_sfixed(13050.0/65536.0,1,-nbitq), 
to_sfixed(-9650.0/65536.0,1,-nbitq), 
to_sfixed(13617.0/65536.0,1,-nbitq), 
to_sfixed(-4110.0/65536.0,1,-nbitq), 
to_sfixed(103.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-5148.0/65536.0,1,-nbitq), 
to_sfixed(-18883.0/65536.0,1,-nbitq), 
to_sfixed(25256.0/65536.0,1,-nbitq), 
to_sfixed(-8256.0/65536.0,1,-nbitq), 
to_sfixed(-13619.0/65536.0,1,-nbitq), 
to_sfixed(6419.0/65536.0,1,-nbitq), 
to_sfixed(-22709.0/65536.0,1,-nbitq), 
to_sfixed(6595.0/65536.0,1,-nbitq), 
to_sfixed(13887.0/65536.0,1,-nbitq), 
to_sfixed(30896.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-13114.0/65536.0,1,-nbitq), 
to_sfixed(8884.0/65536.0,1,-nbitq), 
to_sfixed(-4552.0/65536.0,1,-nbitq), 
to_sfixed(18202.0/65536.0,1,-nbitq), 
to_sfixed(-17431.0/65536.0,1,-nbitq), 
to_sfixed(10876.0/65536.0,1,-nbitq), 
to_sfixed(-7478.0/65536.0,1,-nbitq), 
to_sfixed(-11120.0/65536.0,1,-nbitq), 
to_sfixed(-13305.0/65536.0,1,-nbitq), 
to_sfixed(-2604.0/65536.0,1,-nbitq)  ), 
( to_sfixed(12735.0/65536.0,1,-nbitq), 
to_sfixed(-18883.0/65536.0,1,-nbitq), 
to_sfixed(12064.0/65536.0,1,-nbitq), 
to_sfixed(-2525.0/65536.0,1,-nbitq), 
to_sfixed(18996.0/65536.0,1,-nbitq), 
to_sfixed(17417.0/65536.0,1,-nbitq), 
to_sfixed(15290.0/65536.0,1,-nbitq), 
to_sfixed(-12512.0/65536.0,1,-nbitq), 
to_sfixed(3948.0/65536.0,1,-nbitq), 
to_sfixed(-10586.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4639.0/65536.0,1,-nbitq), 
to_sfixed(-15706.0/65536.0,1,-nbitq), 
to_sfixed(-17586.0/65536.0,1,-nbitq), 
to_sfixed(10039.0/65536.0,1,-nbitq), 
to_sfixed(8434.0/65536.0,1,-nbitq), 
to_sfixed(30629.0/65536.0,1,-nbitq), 
to_sfixed(-2583.0/65536.0,1,-nbitq), 
to_sfixed(-199.0/65536.0,1,-nbitq), 
to_sfixed(-25314.0/65536.0,1,-nbitq), 
to_sfixed(-3560.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-27236.0/65536.0,1,-nbitq), 
to_sfixed(-8128.0/65536.0,1,-nbitq), 
to_sfixed(-16375.0/65536.0,1,-nbitq), 
to_sfixed(-19063.0/65536.0,1,-nbitq), 
to_sfixed(-5590.0/65536.0,1,-nbitq), 
to_sfixed(6529.0/65536.0,1,-nbitq), 
to_sfixed(-14957.0/65536.0,1,-nbitq), 
to_sfixed(26197.0/65536.0,1,-nbitq), 
to_sfixed(-5392.0/65536.0,1,-nbitq), 
to_sfixed(3759.0/65536.0,1,-nbitq)  ), 
( to_sfixed(10926.0/65536.0,1,-nbitq), 
to_sfixed(2037.0/65536.0,1,-nbitq), 
to_sfixed(6077.0/65536.0,1,-nbitq), 
to_sfixed(-156.0/65536.0,1,-nbitq), 
to_sfixed(23622.0/65536.0,1,-nbitq), 
to_sfixed(-16194.0/65536.0,1,-nbitq), 
to_sfixed(-25524.0/65536.0,1,-nbitq), 
to_sfixed(36031.0/65536.0,1,-nbitq), 
to_sfixed(-19708.0/65536.0,1,-nbitq), 
to_sfixed(-28471.0/65536.0,1,-nbitq)  ), 
( to_sfixed(12204.0/65536.0,1,-nbitq), 
to_sfixed(12681.0/65536.0,1,-nbitq), 
to_sfixed(1409.0/65536.0,1,-nbitq), 
to_sfixed(2533.0/65536.0,1,-nbitq), 
to_sfixed(5997.0/65536.0,1,-nbitq), 
to_sfixed(10228.0/65536.0,1,-nbitq), 
to_sfixed(13473.0/65536.0,1,-nbitq), 
to_sfixed(-10404.0/65536.0,1,-nbitq), 
to_sfixed(-10271.0/65536.0,1,-nbitq), 
to_sfixed(-12466.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-8790.0/65536.0,1,-nbitq), 
to_sfixed(13409.0/65536.0,1,-nbitq), 
to_sfixed(-9593.0/65536.0,1,-nbitq), 
to_sfixed(7233.0/65536.0,1,-nbitq), 
to_sfixed(10244.0/65536.0,1,-nbitq), 
to_sfixed(-8814.0/65536.0,1,-nbitq), 
to_sfixed(13755.0/65536.0,1,-nbitq), 
to_sfixed(1797.0/65536.0,1,-nbitq), 
to_sfixed(-1714.0/65536.0,1,-nbitq), 
to_sfixed(4390.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4768.0/65536.0,1,-nbitq), 
to_sfixed(23579.0/65536.0,1,-nbitq), 
to_sfixed(33748.0/65536.0,1,-nbitq), 
to_sfixed(2338.0/65536.0,1,-nbitq), 
to_sfixed(-1956.0/65536.0,1,-nbitq), 
to_sfixed(-19470.0/65536.0,1,-nbitq), 
to_sfixed(21618.0/65536.0,1,-nbitq), 
to_sfixed(-21186.0/65536.0,1,-nbitq), 
to_sfixed(-22706.0/65536.0,1,-nbitq), 
to_sfixed(-14885.0/65536.0,1,-nbitq)  ), 
( to_sfixed(2574.0/65536.0,1,-nbitq), 
to_sfixed(18611.0/65536.0,1,-nbitq), 
to_sfixed(2775.0/65536.0,1,-nbitq), 
to_sfixed(-14717.0/65536.0,1,-nbitq), 
to_sfixed(23646.0/65536.0,1,-nbitq), 
to_sfixed(-2661.0/65536.0,1,-nbitq), 
to_sfixed(1369.0/65536.0,1,-nbitq), 
to_sfixed(22929.0/65536.0,1,-nbitq), 
to_sfixed(7335.0/65536.0,1,-nbitq), 
to_sfixed(-13501.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-30277.0/65536.0,1,-nbitq), 
to_sfixed(26576.0/65536.0,1,-nbitq), 
to_sfixed(5566.0/65536.0,1,-nbitq), 
to_sfixed(-1827.0/65536.0,1,-nbitq), 
to_sfixed(29707.0/65536.0,1,-nbitq), 
to_sfixed(-25113.0/65536.0,1,-nbitq), 
to_sfixed(23598.0/65536.0,1,-nbitq), 
to_sfixed(-11629.0/65536.0,1,-nbitq), 
to_sfixed(-16109.0/65536.0,1,-nbitq), 
to_sfixed(-18642.0/65536.0,1,-nbitq)  ), 
( to_sfixed(14814.0/65536.0,1,-nbitq), 
to_sfixed(14415.0/65536.0,1,-nbitq), 
to_sfixed(17151.0/65536.0,1,-nbitq), 
to_sfixed(6376.0/65536.0,1,-nbitq), 
to_sfixed(-16692.0/65536.0,1,-nbitq), 
to_sfixed(-14698.0/65536.0,1,-nbitq), 
to_sfixed(15949.0/65536.0,1,-nbitq), 
to_sfixed(-16817.0/65536.0,1,-nbitq), 
to_sfixed(-9545.0/65536.0,1,-nbitq), 
to_sfixed(-7160.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-24914.0/65536.0,1,-nbitq), 
to_sfixed(-7380.0/65536.0,1,-nbitq), 
to_sfixed(-26337.0/65536.0,1,-nbitq), 
to_sfixed(1218.0/65536.0,1,-nbitq), 
to_sfixed(685.0/65536.0,1,-nbitq), 
to_sfixed(2241.0/65536.0,1,-nbitq), 
to_sfixed(30080.0/65536.0,1,-nbitq), 
to_sfixed(-19704.0/65536.0,1,-nbitq), 
to_sfixed(15857.0/65536.0,1,-nbitq), 
to_sfixed(19058.0/65536.0,1,-nbitq)  ), 
( to_sfixed(958.0/65536.0,1,-nbitq), 
to_sfixed(-5454.0/65536.0,1,-nbitq), 
to_sfixed(5884.0/65536.0,1,-nbitq), 
to_sfixed(-6730.0/65536.0,1,-nbitq), 
to_sfixed(-12790.0/65536.0,1,-nbitq), 
to_sfixed(-12675.0/65536.0,1,-nbitq), 
to_sfixed(-14475.0/65536.0,1,-nbitq), 
to_sfixed(-14458.0/65536.0,1,-nbitq), 
to_sfixed(-10315.0/65536.0,1,-nbitq), 
to_sfixed(4521.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-15984.0/65536.0,1,-nbitq), 
to_sfixed(-10510.0/65536.0,1,-nbitq), 
to_sfixed(24522.0/65536.0,1,-nbitq), 
to_sfixed(-28355.0/65536.0,1,-nbitq), 
to_sfixed(772.0/65536.0,1,-nbitq), 
to_sfixed(19699.0/65536.0,1,-nbitq), 
to_sfixed(3321.0/65536.0,1,-nbitq), 
to_sfixed(16457.0/65536.0,1,-nbitq), 
to_sfixed(-1912.0/65536.0,1,-nbitq), 
to_sfixed(14239.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-8512.0/65536.0,1,-nbitq), 
to_sfixed(-14551.0/65536.0,1,-nbitq), 
to_sfixed(11489.0/65536.0,1,-nbitq), 
to_sfixed(-4071.0/65536.0,1,-nbitq), 
to_sfixed(15093.0/65536.0,1,-nbitq), 
to_sfixed(25964.0/65536.0,1,-nbitq), 
to_sfixed(-3969.0/65536.0,1,-nbitq), 
to_sfixed(-12464.0/65536.0,1,-nbitq), 
to_sfixed(-7249.0/65536.0,1,-nbitq), 
to_sfixed(-20983.0/65536.0,1,-nbitq)  ), 
( to_sfixed(3607.0/65536.0,1,-nbitq), 
to_sfixed(7157.0/65536.0,1,-nbitq), 
to_sfixed(-13336.0/65536.0,1,-nbitq), 
to_sfixed(-17266.0/65536.0,1,-nbitq), 
to_sfixed(7285.0/65536.0,1,-nbitq), 
to_sfixed(1810.0/65536.0,1,-nbitq), 
to_sfixed(-9749.0/65536.0,1,-nbitq), 
to_sfixed(3014.0/65536.0,1,-nbitq), 
to_sfixed(-1637.0/65536.0,1,-nbitq), 
to_sfixed(-6956.0/65536.0,1,-nbitq)  ), 
( to_sfixed(22300.0/65536.0,1,-nbitq), 
to_sfixed(-27094.0/65536.0,1,-nbitq), 
to_sfixed(-14739.0/65536.0,1,-nbitq), 
to_sfixed(9437.0/65536.0,1,-nbitq), 
to_sfixed(-35354.0/65536.0,1,-nbitq), 
to_sfixed(7044.0/65536.0,1,-nbitq), 
to_sfixed(25398.0/65536.0,1,-nbitq), 
to_sfixed(-13698.0/65536.0,1,-nbitq), 
to_sfixed(-18163.0/65536.0,1,-nbitq), 
to_sfixed(41388.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-1705.0/65536.0,1,-nbitq), 
to_sfixed(-2538.0/65536.0,1,-nbitq), 
to_sfixed(3229.0/65536.0,1,-nbitq), 
to_sfixed(1795.0/65536.0,1,-nbitq), 
to_sfixed(-4671.0/65536.0,1,-nbitq), 
to_sfixed(13624.0/65536.0,1,-nbitq), 
to_sfixed(-6176.0/65536.0,1,-nbitq), 
to_sfixed(-12631.0/65536.0,1,-nbitq), 
to_sfixed(-14305.0/65536.0,1,-nbitq), 
to_sfixed(5314.0/65536.0,1,-nbitq)  ), 
( to_sfixed(20576.0/65536.0,1,-nbitq), 
to_sfixed(-1093.0/65536.0,1,-nbitq), 
to_sfixed(-3185.0/65536.0,1,-nbitq), 
to_sfixed(18622.0/65536.0,1,-nbitq), 
to_sfixed(-9797.0/65536.0,1,-nbitq), 
to_sfixed(-607.0/65536.0,1,-nbitq), 
to_sfixed(-14576.0/65536.0,1,-nbitq), 
to_sfixed(22668.0/65536.0,1,-nbitq), 
to_sfixed(-5510.0/65536.0,1,-nbitq), 
to_sfixed(-1658.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-11055.0/65536.0,1,-nbitq), 
to_sfixed(1580.0/65536.0,1,-nbitq), 
to_sfixed(-4535.0/65536.0,1,-nbitq), 
to_sfixed(13379.0/65536.0,1,-nbitq), 
to_sfixed(-12258.0/65536.0,1,-nbitq), 
to_sfixed(-11026.0/65536.0,1,-nbitq), 
to_sfixed(-1563.0/65536.0,1,-nbitq), 
to_sfixed(-2084.0/65536.0,1,-nbitq), 
to_sfixed(-11976.0/65536.0,1,-nbitq), 
to_sfixed(-8589.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-975.0/65536.0,1,-nbitq), 
to_sfixed(-569.0/65536.0,1,-nbitq), 
to_sfixed(-6711.0/65536.0,1,-nbitq), 
to_sfixed(-444.0/65536.0,1,-nbitq), 
to_sfixed(12189.0/65536.0,1,-nbitq), 
to_sfixed(-2517.0/65536.0,1,-nbitq), 
to_sfixed(3294.0/65536.0,1,-nbitq), 
to_sfixed(11233.0/65536.0,1,-nbitq), 
to_sfixed(-3383.0/65536.0,1,-nbitq), 
to_sfixed(15165.0/65536.0,1,-nbitq)  ), 
( to_sfixed(400.0/65536.0,1,-nbitq), 
to_sfixed(-16650.0/65536.0,1,-nbitq), 
to_sfixed(16218.0/65536.0,1,-nbitq), 
to_sfixed(4500.0/65536.0,1,-nbitq), 
to_sfixed(6362.0/65536.0,1,-nbitq), 
to_sfixed(-13868.0/65536.0,1,-nbitq), 
to_sfixed(9190.0/65536.0,1,-nbitq), 
to_sfixed(-4197.0/65536.0,1,-nbitq), 
to_sfixed(-10341.0/65536.0,1,-nbitq), 
to_sfixed(-7065.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-18577.0/65536.0,1,-nbitq), 
to_sfixed(-16013.0/65536.0,1,-nbitq), 
to_sfixed(-4285.0/65536.0,1,-nbitq), 
to_sfixed(10890.0/65536.0,1,-nbitq), 
to_sfixed(-5053.0/65536.0,1,-nbitq), 
to_sfixed(13078.0/65536.0,1,-nbitq), 
to_sfixed(9916.0/65536.0,1,-nbitq), 
to_sfixed(-14848.0/65536.0,1,-nbitq), 
to_sfixed(32710.0/65536.0,1,-nbitq), 
to_sfixed(-12991.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-11025.0/65536.0,1,-nbitq), 
to_sfixed(-8608.0/65536.0,1,-nbitq), 
to_sfixed(17912.0/65536.0,1,-nbitq), 
to_sfixed(14491.0/65536.0,1,-nbitq), 
to_sfixed(14704.0/65536.0,1,-nbitq), 
to_sfixed(19223.0/65536.0,1,-nbitq), 
to_sfixed(9827.0/65536.0,1,-nbitq), 
to_sfixed(3500.0/65536.0,1,-nbitq), 
to_sfixed(-13639.0/65536.0,1,-nbitq), 
to_sfixed(-18300.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-7613.0/65536.0,1,-nbitq), 
to_sfixed(13600.0/65536.0,1,-nbitq), 
to_sfixed(-26529.0/65536.0,1,-nbitq), 
to_sfixed(5324.0/65536.0,1,-nbitq), 
to_sfixed(-12288.0/65536.0,1,-nbitq), 
to_sfixed(-7785.0/65536.0,1,-nbitq), 
to_sfixed(-18718.0/65536.0,1,-nbitq), 
to_sfixed(12669.0/65536.0,1,-nbitq), 
to_sfixed(15825.0/65536.0,1,-nbitq), 
to_sfixed(26762.0/65536.0,1,-nbitq)  ), 
( to_sfixed(21531.0/65536.0,1,-nbitq), 
to_sfixed(-147.0/65536.0,1,-nbitq), 
to_sfixed(7393.0/65536.0,1,-nbitq), 
to_sfixed(5233.0/65536.0,1,-nbitq), 
to_sfixed(12879.0/65536.0,1,-nbitq), 
to_sfixed(-15322.0/65536.0,1,-nbitq), 
to_sfixed(-9598.0/65536.0,1,-nbitq), 
to_sfixed(4236.0/65536.0,1,-nbitq), 
to_sfixed(-16367.0/65536.0,1,-nbitq), 
to_sfixed(-22343.0/65536.0,1,-nbitq)  ), 
( to_sfixed(11595.0/65536.0,1,-nbitq), 
to_sfixed(-5510.0/65536.0,1,-nbitq), 
to_sfixed(-4808.0/65536.0,1,-nbitq), 
to_sfixed(-5415.0/65536.0,1,-nbitq), 
to_sfixed(-11077.0/65536.0,1,-nbitq), 
to_sfixed(24936.0/65536.0,1,-nbitq), 
to_sfixed(2446.0/65536.0,1,-nbitq), 
to_sfixed(-32296.0/65536.0,1,-nbitq), 
to_sfixed(-22498.0/65536.0,1,-nbitq), 
to_sfixed(10211.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-6797.0/65536.0,1,-nbitq), 
to_sfixed(10444.0/65536.0,1,-nbitq), 
to_sfixed(-6372.0/65536.0,1,-nbitq), 
to_sfixed(9895.0/65536.0,1,-nbitq), 
to_sfixed(15284.0/65536.0,1,-nbitq), 
to_sfixed(-14585.0/65536.0,1,-nbitq), 
to_sfixed(3137.0/65536.0,1,-nbitq), 
to_sfixed(15924.0/65536.0,1,-nbitq), 
to_sfixed(-15104.0/65536.0,1,-nbitq), 
to_sfixed(-12091.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4408.0/65536.0,1,-nbitq), 
to_sfixed(11442.0/65536.0,1,-nbitq), 
to_sfixed(11324.0/65536.0,1,-nbitq), 
to_sfixed(-5079.0/65536.0,1,-nbitq), 
to_sfixed(-7738.0/65536.0,1,-nbitq), 
to_sfixed(-12241.0/65536.0,1,-nbitq), 
to_sfixed(-9367.0/65536.0,1,-nbitq), 
to_sfixed(-1870.0/65536.0,1,-nbitq), 
to_sfixed(14528.0/65536.0,1,-nbitq), 
to_sfixed(5564.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-8582.0/65536.0,1,-nbitq), 
to_sfixed(14825.0/65536.0,1,-nbitq), 
to_sfixed(10660.0/65536.0,1,-nbitq), 
to_sfixed(13517.0/65536.0,1,-nbitq), 
to_sfixed(-2270.0/65536.0,1,-nbitq), 
to_sfixed(-10318.0/65536.0,1,-nbitq), 
to_sfixed(-1418.0/65536.0,1,-nbitq), 
to_sfixed(-2800.0/65536.0,1,-nbitq), 
to_sfixed(-13495.0/65536.0,1,-nbitq), 
to_sfixed(8633.0/65536.0,1,-nbitq)  ), 
( to_sfixed(4799.0/65536.0,1,-nbitq), 
to_sfixed(-19046.0/65536.0,1,-nbitq), 
to_sfixed(-13966.0/65536.0,1,-nbitq), 
to_sfixed(25989.0/65536.0,1,-nbitq), 
to_sfixed(-18200.0/65536.0,1,-nbitq), 
to_sfixed(21400.0/65536.0,1,-nbitq), 
to_sfixed(-27992.0/65536.0,1,-nbitq), 
to_sfixed(1631.0/65536.0,1,-nbitq), 
to_sfixed(-9390.0/65536.0,1,-nbitq), 
to_sfixed(-17113.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-38175.0/65536.0,1,-nbitq), 
to_sfixed(8059.0/65536.0,1,-nbitq), 
to_sfixed(-5478.0/65536.0,1,-nbitq), 
to_sfixed(16095.0/65536.0,1,-nbitq), 
to_sfixed(-11462.0/65536.0,1,-nbitq), 
to_sfixed(-10057.0/65536.0,1,-nbitq), 
to_sfixed(22414.0/65536.0,1,-nbitq), 
to_sfixed(822.0/65536.0,1,-nbitq), 
to_sfixed(-3604.0/65536.0,1,-nbitq), 
to_sfixed(-13818.0/65536.0,1,-nbitq)  ), 
( to_sfixed(15132.0/65536.0,1,-nbitq), 
to_sfixed(-11526.0/65536.0,1,-nbitq), 
to_sfixed(-16056.0/65536.0,1,-nbitq), 
to_sfixed(7703.0/65536.0,1,-nbitq), 
to_sfixed(591.0/65536.0,1,-nbitq), 
to_sfixed(-11412.0/65536.0,1,-nbitq), 
to_sfixed(-14132.0/65536.0,1,-nbitq), 
to_sfixed(10931.0/65536.0,1,-nbitq), 
to_sfixed(13420.0/65536.0,1,-nbitq), 
to_sfixed(15841.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-15852.0/65536.0,1,-nbitq), 
to_sfixed(1684.0/65536.0,1,-nbitq), 
to_sfixed(-1772.0/65536.0,1,-nbitq), 
to_sfixed(-59.0/65536.0,1,-nbitq), 
to_sfixed(8958.0/65536.0,1,-nbitq), 
to_sfixed(-1613.0/65536.0,1,-nbitq), 
to_sfixed(-7570.0/65536.0,1,-nbitq), 
to_sfixed(3804.0/65536.0,1,-nbitq), 
to_sfixed(-1746.0/65536.0,1,-nbitq), 
to_sfixed(1086.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-3818.0/65536.0,1,-nbitq), 
to_sfixed(-2.0/65536.0,1,-nbitq), 
to_sfixed(12176.0/65536.0,1,-nbitq), 
to_sfixed(-7286.0/65536.0,1,-nbitq), 
to_sfixed(6484.0/65536.0,1,-nbitq), 
to_sfixed(-7897.0/65536.0,1,-nbitq), 
to_sfixed(8060.0/65536.0,1,-nbitq), 
to_sfixed(-16608.0/65536.0,1,-nbitq), 
to_sfixed(13902.0/65536.0,1,-nbitq), 
to_sfixed(-917.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-12201.0/65536.0,1,-nbitq), 
to_sfixed(5042.0/65536.0,1,-nbitq), 
to_sfixed(3253.0/65536.0,1,-nbitq), 
to_sfixed(9175.0/65536.0,1,-nbitq), 
to_sfixed(-1080.0/65536.0,1,-nbitq), 
to_sfixed(4282.0/65536.0,1,-nbitq), 
to_sfixed(25856.0/65536.0,1,-nbitq), 
to_sfixed(-31649.0/65536.0,1,-nbitq), 
to_sfixed(-16628.0/65536.0,1,-nbitq), 
to_sfixed(-732.0/65536.0,1,-nbitq)  ), 
( to_sfixed(23234.0/65536.0,1,-nbitq), 
to_sfixed(-14036.0/65536.0,1,-nbitq), 
to_sfixed(-14253.0/65536.0,1,-nbitq), 
to_sfixed(6249.0/65536.0,1,-nbitq), 
to_sfixed(24085.0/65536.0,1,-nbitq), 
to_sfixed(24257.0/65536.0,1,-nbitq), 
to_sfixed(-19557.0/65536.0,1,-nbitq), 
to_sfixed(-15298.0/65536.0,1,-nbitq), 
to_sfixed(-38103.0/65536.0,1,-nbitq), 
to_sfixed(31728.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-7446.0/65536.0,1,-nbitq), 
to_sfixed(-11284.0/65536.0,1,-nbitq), 
to_sfixed(7397.0/65536.0,1,-nbitq), 
to_sfixed(-18981.0/65536.0,1,-nbitq), 
to_sfixed(7207.0/65536.0,1,-nbitq), 
to_sfixed(-11519.0/65536.0,1,-nbitq), 
to_sfixed(18154.0/65536.0,1,-nbitq), 
to_sfixed(-18185.0/65536.0,1,-nbitq), 
to_sfixed(6933.0/65536.0,1,-nbitq), 
to_sfixed(16643.0/65536.0,1,-nbitq)  ), 
( to_sfixed(19088.0/65536.0,1,-nbitq), 
to_sfixed(-20106.0/65536.0,1,-nbitq), 
to_sfixed(4825.0/65536.0,1,-nbitq), 
to_sfixed(-26691.0/65536.0,1,-nbitq), 
to_sfixed(16428.0/65536.0,1,-nbitq), 
to_sfixed(28695.0/65536.0,1,-nbitq), 
to_sfixed(-8775.0/65536.0,1,-nbitq), 
to_sfixed(15270.0/65536.0,1,-nbitq), 
to_sfixed(2001.0/65536.0,1,-nbitq), 
to_sfixed(7449.0/65536.0,1,-nbitq)  ), 
( to_sfixed(24333.0/65536.0,1,-nbitq), 
to_sfixed(15260.0/65536.0,1,-nbitq), 
to_sfixed(3117.0/65536.0,1,-nbitq), 
to_sfixed(-12833.0/65536.0,1,-nbitq), 
to_sfixed(-19782.0/65536.0,1,-nbitq), 
to_sfixed(-7916.0/65536.0,1,-nbitq), 
to_sfixed(34835.0/65536.0,1,-nbitq), 
to_sfixed(-15492.0/65536.0,1,-nbitq), 
to_sfixed(7188.0/65536.0,1,-nbitq), 
to_sfixed(-7826.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-16774.0/65536.0,1,-nbitq), 
to_sfixed(15407.0/65536.0,1,-nbitq), 
to_sfixed(7268.0/65536.0,1,-nbitq), 
to_sfixed(-18645.0/65536.0,1,-nbitq), 
to_sfixed(-19329.0/65536.0,1,-nbitq), 
to_sfixed(-20152.0/65536.0,1,-nbitq), 
to_sfixed(867.0/65536.0,1,-nbitq), 
to_sfixed(14351.0/65536.0,1,-nbitq), 
to_sfixed(27129.0/65536.0,1,-nbitq), 
to_sfixed(-2924.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-2124.0/65536.0,1,-nbitq), 
to_sfixed(-9180.0/65536.0,1,-nbitq), 
to_sfixed(12226.0/65536.0,1,-nbitq), 
to_sfixed(3428.0/65536.0,1,-nbitq), 
to_sfixed(-5064.0/65536.0,1,-nbitq), 
to_sfixed(7222.0/65536.0,1,-nbitq), 
to_sfixed(-15293.0/65536.0,1,-nbitq), 
to_sfixed(-7553.0/65536.0,1,-nbitq), 
to_sfixed(-14817.0/65536.0,1,-nbitq), 
to_sfixed(-13525.0/65536.0,1,-nbitq)  ), 
( to_sfixed(15723.0/65536.0,1,-nbitq), 
to_sfixed(-20731.0/65536.0,1,-nbitq), 
to_sfixed(-9639.0/65536.0,1,-nbitq), 
to_sfixed(11984.0/65536.0,1,-nbitq), 
to_sfixed(16952.0/65536.0,1,-nbitq), 
to_sfixed(-11359.0/65536.0,1,-nbitq), 
to_sfixed(7736.0/65536.0,1,-nbitq), 
to_sfixed(-20681.0/65536.0,1,-nbitq), 
to_sfixed(-7961.0/65536.0,1,-nbitq), 
to_sfixed(20146.0/65536.0,1,-nbitq)  ), 
( to_sfixed(5590.0/65536.0,1,-nbitq), 
to_sfixed(-15494.0/65536.0,1,-nbitq), 
to_sfixed(-77.0/65536.0,1,-nbitq), 
to_sfixed(28457.0/65536.0,1,-nbitq), 
to_sfixed(-34842.0/65536.0,1,-nbitq), 
to_sfixed(-31896.0/65536.0,1,-nbitq), 
to_sfixed(12009.0/65536.0,1,-nbitq), 
to_sfixed(-26938.0/65536.0,1,-nbitq), 
to_sfixed(7029.0/65536.0,1,-nbitq), 
to_sfixed(-20382.0/65536.0,1,-nbitq)  ), 
( to_sfixed(16126.0/65536.0,1,-nbitq), 
to_sfixed(-4499.0/65536.0,1,-nbitq), 
to_sfixed(-6830.0/65536.0,1,-nbitq), 
to_sfixed(-227.0/65536.0,1,-nbitq), 
to_sfixed(5524.0/65536.0,1,-nbitq), 
to_sfixed(-16826.0/65536.0,1,-nbitq), 
to_sfixed(6964.0/65536.0,1,-nbitq), 
to_sfixed(5327.0/65536.0,1,-nbitq), 
to_sfixed(-13688.0/65536.0,1,-nbitq), 
to_sfixed(-2800.0/65536.0,1,-nbitq)  ), 
( to_sfixed(8865.0/65536.0,1,-nbitq), 
to_sfixed(-1245.0/65536.0,1,-nbitq), 
to_sfixed(-4864.0/65536.0,1,-nbitq), 
to_sfixed(4184.0/65536.0,1,-nbitq), 
to_sfixed(-2236.0/65536.0,1,-nbitq), 
to_sfixed(4847.0/65536.0,1,-nbitq), 
to_sfixed(-15009.0/65536.0,1,-nbitq), 
to_sfixed(-1304.0/65536.0,1,-nbitq), 
to_sfixed(308.0/65536.0,1,-nbitq), 
to_sfixed(7911.0/65536.0,1,-nbitq)  ), 
( to_sfixed(30335.0/65536.0,1,-nbitq), 
to_sfixed(-16181.0/65536.0,1,-nbitq), 
to_sfixed(13631.0/65536.0,1,-nbitq), 
to_sfixed(-10651.0/65536.0,1,-nbitq), 
to_sfixed(-20302.0/65536.0,1,-nbitq), 
to_sfixed(-7781.0/65536.0,1,-nbitq), 
to_sfixed(-8577.0/65536.0,1,-nbitq), 
to_sfixed(10058.0/65536.0,1,-nbitq), 
to_sfixed(-11436.0/65536.0,1,-nbitq), 
to_sfixed(-29.0/65536.0,1,-nbitq)  ), 
( to_sfixed(24521.0/65536.0,1,-nbitq), 
to_sfixed(17571.0/65536.0,1,-nbitq), 
to_sfixed(14201.0/65536.0,1,-nbitq), 
to_sfixed(13272.0/65536.0,1,-nbitq), 
to_sfixed(12121.0/65536.0,1,-nbitq), 
to_sfixed(-11170.0/65536.0,1,-nbitq), 
to_sfixed(-16617.0/65536.0,1,-nbitq), 
to_sfixed(-21267.0/65536.0,1,-nbitq), 
to_sfixed(-16775.0/65536.0,1,-nbitq), 
to_sfixed(-7275.0/65536.0,1,-nbitq)  ), 
( to_sfixed(25381.0/65536.0,1,-nbitq), 
to_sfixed(-23029.0/65536.0,1,-nbitq), 
to_sfixed(14282.0/65536.0,1,-nbitq), 
to_sfixed(-6033.0/65536.0,1,-nbitq), 
to_sfixed(-2664.0/65536.0,1,-nbitq), 
to_sfixed(-23610.0/65536.0,1,-nbitq), 
to_sfixed(10784.0/65536.0,1,-nbitq), 
to_sfixed(-28647.0/65536.0,1,-nbitq), 
to_sfixed(-14558.0/65536.0,1,-nbitq), 
to_sfixed(11760.0/65536.0,1,-nbitq)  ), 
( to_sfixed(-11471.0/65536.0,1,-nbitq), 
to_sfixed(-693.0/65536.0,1,-nbitq), 
to_sfixed(-15258.0/65536.0,1,-nbitq), 
to_sfixed(13695.0/65536.0,1,-nbitq), 
to_sfixed(14054.0/65536.0,1,-nbitq), 
to_sfixed(-16886.0/65536.0,1,-nbitq), 
to_sfixed(13335.0/65536.0,1,-nbitq), 
to_sfixed(1842.0/65536.0,1,-nbitq), 
to_sfixed(8129.0/65536.0,1,-nbitq), 
to_sfixed(-1049.0/65536.0,1,-nbitq)  ), 
( to_sfixed(27312.0/65536.0,1,-nbitq), 
to_sfixed(11124.0/65536.0,1,-nbitq), 
to_sfixed(15612.0/65536.0,1,-nbitq), 
to_sfixed(17992.0/65536.0,1,-nbitq), 
to_sfixed(-10407.0/65536.0,1,-nbitq), 
to_sfixed(-8401.0/65536.0,1,-nbitq), 
to_sfixed(24327.0/65536.0,1,-nbitq), 
to_sfixed(-17107.0/65536.0,1,-nbitq), 
to_sfixed(7533.0/65536.0,1,-nbitq), 
to_sfixed(5548.0/65536.0,1,-nbitq)  ) 
 ) ;
end package coeff;
