LIBRARY ieee, work;
USE ieee.std_logic_1164.all;
use IEEE.numeric_std.ALL;
use std.textio.all;
use ieee.fixed_pkg.all;
use ieee.fixed_float_types.all;

package coeff is
 
constant lngimag : integer := 784 ; 
constant lngfilt : integer := 784 ; 
constant nbneuron : integer := 80 ; 
constant nbsymbol : integer := 10 ; 
constant nbitq : integer := 32 ; 

constant ccf : integer := 2 ; 
constant ccf2 : integer := 4 ; 
constant cct : integer := 32 ; 
constant cct2 : integer := 1 ;

type typtabup is array(0 to lngimag-1) of std_logic ;								-- tableau indiquant les pixels effectivement utilisés lors des calculs
type typtabmul is array(natural range <>) of sfixed(3 downto -nbitq);
type typtabcst is array(natural range <>) of sfixed(1 downto -nbitq);
type typtabcnf1 is array(0 to lngimag-1, 0 to nbneuron-1) of sfixed(1 downto -nbitq);
type typtabcnf2 is array(0 to nbneuron-1, 0 to nbsymbol-1) of sfixed(1 downto -nbitq);
type typtabaccu is array(0 to nbneuron-1) of sfixed(8 downto -2*nbitq) ;
type typtabaccu2 is array(0 to nbsymbol-1) of sfixed(8 downto -2*nbitq) ;
subtype usng4 is unsigned(3 downto 0) ;
type typlabel is array(0 to 4) of usng4 ;

constant usedpix : typtabup := ( '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1'  ) ; 

constant cst1 : typtabcst := ( to_sfixed(-251483974.0/4294967296.0,1,-nbitq), to_sfixed(-58348487.0/4294967296.0,1,-nbitq), to_sfixed(132303994.0/4294967296.0,1,-nbitq), to_sfixed(177716109.0/4294967296.0,1,-nbitq), to_sfixed(-31935958.0/4294967296.0,1,-nbitq), to_sfixed(10177649.0/4294967296.0,1,-nbitq), to_sfixed(-295188506.0/4294967296.0,1,-nbitq), to_sfixed(-116662224.0/4294967296.0,1,-nbitq), to_sfixed(342447877.0/4294967296.0,1,-nbitq), to_sfixed(-608854209.0/4294967296.0,1,-nbitq), to_sfixed(-116118655.0/4294967296.0,1,-nbitq), to_sfixed(44666523.0/4294967296.0,1,-nbitq), to_sfixed(-324990993.0/4294967296.0,1,-nbitq), to_sfixed(396977518.0/4294967296.0,1,-nbitq), to_sfixed(93061357.0/4294967296.0,1,-nbitq), to_sfixed(151748345.0/4294967296.0,1,-nbitq), to_sfixed(653678427.0/4294967296.0,1,-nbitq), to_sfixed(-472526708.0/4294967296.0,1,-nbitq), to_sfixed(-31703772.0/4294967296.0,1,-nbitq), to_sfixed(-835001184.0/4294967296.0,1,-nbitq), to_sfixed(723344418.0/4294967296.0,1,-nbitq), to_sfixed(69816678.0/4294967296.0,1,-nbitq), to_sfixed(-281338060.0/4294967296.0,1,-nbitq), to_sfixed(255600017.0/4294967296.0,1,-nbitq), to_sfixed(-960376859.0/4294967296.0,1,-nbitq), to_sfixed(-289633948.0/4294967296.0,1,-nbitq), to_sfixed(1114847633.0/4294967296.0,1,-nbitq), to_sfixed(459781674.0/4294967296.0,1,-nbitq), to_sfixed(39710522.0/4294967296.0,1,-nbitq), to_sfixed(-373422413.0/4294967296.0,1,-nbitq), to_sfixed(281202646.0/4294967296.0,1,-nbitq), to_sfixed(-61980685.0/4294967296.0,1,-nbitq), to_sfixed(-436260966.0/4294967296.0,1,-nbitq), to_sfixed(-1096426691.0/4294967296.0,1,-nbitq), to_sfixed(-517352549.0/4294967296.0,1,-nbitq), to_sfixed(150641188.0/4294967296.0,1,-nbitq), to_sfixed(-168455825.0/4294967296.0,1,-nbitq), to_sfixed(150321410.0/4294967296.0,1,-nbitq), to_sfixed(485476355.0/4294967296.0,1,-nbitq), to_sfixed(-2166157525.0/4294967296.0,1,-nbitq), to_sfixed(82628214.0/4294967296.0,1,-nbitq), to_sfixed(-465636296.0/4294967296.0,1,-nbitq), to_sfixed(36129021.0/4294967296.0,1,-nbitq), to_sfixed(110049548.0/4294967296.0,1,-nbitq), to_sfixed(1471431780.0/4294967296.0,1,-nbitq), to_sfixed(435888314.0/4294967296.0,1,-nbitq), to_sfixed(887559283.0/4294967296.0,1,-nbitq), to_sfixed(39455771.0/4294967296.0,1,-nbitq), to_sfixed(1209347034.0/4294967296.0,1,-nbitq), to_sfixed(-273059483.0/4294967296.0,1,-nbitq), to_sfixed(720669509.0/4294967296.0,1,-nbitq), to_sfixed(423434590.0/4294967296.0,1,-nbitq), to_sfixed(294524908.0/4294967296.0,1,-nbitq), to_sfixed(235415051.0/4294967296.0,1,-nbitq), to_sfixed(-236912431.0/4294967296.0,1,-nbitq), to_sfixed(406132104.0/4294967296.0,1,-nbitq), to_sfixed(36869849.0/4294967296.0,1,-nbitq), to_sfixed(-59001443.0/4294967296.0,1,-nbitq), to_sfixed(-702221616.0/4294967296.0,1,-nbitq), to_sfixed(-736199128.0/4294967296.0,1,-nbitq), to_sfixed(199553092.0/4294967296.0,1,-nbitq), to_sfixed(181652087.0/4294967296.0,1,-nbitq), to_sfixed(296743504.0/4294967296.0,1,-nbitq), to_sfixed(-413916802.0/4294967296.0,1,-nbitq), to_sfixed(789121946.0/4294967296.0,1,-nbitq), to_sfixed(1329396571.0/4294967296.0,1,-nbitq), to_sfixed(-74711997.0/4294967296.0,1,-nbitq), to_sfixed(-139403285.0/4294967296.0,1,-nbitq), to_sfixed(-1019811361.0/4294967296.0,1,-nbitq), to_sfixed(96366034.0/4294967296.0,1,-nbitq), to_sfixed(-415243319.0/4294967296.0,1,-nbitq), to_sfixed(267951787.0/4294967296.0,1,-nbitq), to_sfixed(631032986.0/4294967296.0,1,-nbitq), to_sfixed(-1051453246.0/4294967296.0,1,-nbitq), to_sfixed(-1927534284.0/4294967296.0,1,-nbitq), to_sfixed(65082278.0/4294967296.0,1,-nbitq), to_sfixed(308326540.0/4294967296.0,1,-nbitq), to_sfixed(190930982.0/4294967296.0,1,-nbitq), to_sfixed(276441797.0/4294967296.0,1,-nbitq), to_sfixed(-398889616.0/4294967296.0,1,-nbitq)  ) ;
constant cst2 : typtabcst := ( to_sfixed(943154976.0/4294967296.0,1,-nbitq), to_sfixed(1258370405.0/4294967296.0,1,-nbitq), to_sfixed(3738704969.0/4294967296.0,1,-nbitq), to_sfixed(-1476405394.0/4294967296.0,1,-nbitq), to_sfixed(635989430.0/4294967296.0,1,-nbitq), to_sfixed(-3996997765.0/4294967296.0,1,-nbitq), to_sfixed(136989074.0/4294967296.0,1,-nbitq), to_sfixed(3358502798.0/4294967296.0,1,-nbitq), to_sfixed(-4176634186.0/4294967296.0,1,-nbitq), to_sfixed(-3460585768.0/4294967296.0,1,-nbitq)  ) ;

constant coef1 : typtabcnf1 := ( ( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(260848925.0/4294967296.0,1,-nbitq), 
to_sfixed(-250512075.0/4294967296.0,1,-nbitq), 
to_sfixed(336198333.0/4294967296.0,1,-nbitq), 
to_sfixed(-94661758.0/4294967296.0,1,-nbitq), 
to_sfixed(345404611.0/4294967296.0,1,-nbitq), 
to_sfixed(-250028936.0/4294967296.0,1,-nbitq), 
to_sfixed(255555929.0/4294967296.0,1,-nbitq), 
to_sfixed(175410730.0/4294967296.0,1,-nbitq), 
to_sfixed(-256147356.0/4294967296.0,1,-nbitq), 
to_sfixed(280025850.0/4294967296.0,1,-nbitq), 
to_sfixed(-83534354.0/4294967296.0,1,-nbitq), 
to_sfixed(-166704516.0/4294967296.0,1,-nbitq), 
to_sfixed(52533460.0/4294967296.0,1,-nbitq), 
to_sfixed(-16679065.0/4294967296.0,1,-nbitq), 
to_sfixed(-308237530.0/4294967296.0,1,-nbitq), 
to_sfixed(320466917.0/4294967296.0,1,-nbitq), 
to_sfixed(-175990608.0/4294967296.0,1,-nbitq), 
to_sfixed(208422812.0/4294967296.0,1,-nbitq), 
to_sfixed(313138581.0/4294967296.0,1,-nbitq), 
to_sfixed(-13026275.0/4294967296.0,1,-nbitq), 
to_sfixed(-207386683.0/4294967296.0,1,-nbitq), 
to_sfixed(229716215.0/4294967296.0,1,-nbitq), 
to_sfixed(199971870.0/4294967296.0,1,-nbitq), 
to_sfixed(155241360.0/4294967296.0,1,-nbitq), 
to_sfixed(103126870.0/4294967296.0,1,-nbitq), 
to_sfixed(-85924021.0/4294967296.0,1,-nbitq), 
to_sfixed(412029102.0/4294967296.0,1,-nbitq), 
to_sfixed(-135613410.0/4294967296.0,1,-nbitq), 
to_sfixed(-190534367.0/4294967296.0,1,-nbitq), 
to_sfixed(326598366.0/4294967296.0,1,-nbitq), 
to_sfixed(-359121683.0/4294967296.0,1,-nbitq), 
to_sfixed(-519111836.0/4294967296.0,1,-nbitq), 
to_sfixed(140188288.0/4294967296.0,1,-nbitq), 
to_sfixed(-368618329.0/4294967296.0,1,-nbitq), 
to_sfixed(339074466.0/4294967296.0,1,-nbitq), 
to_sfixed(-97906525.0/4294967296.0,1,-nbitq), 
to_sfixed(-243139923.0/4294967296.0,1,-nbitq), 
to_sfixed(374814893.0/4294967296.0,1,-nbitq), 
to_sfixed(-3228573.0/4294967296.0,1,-nbitq), 
to_sfixed(228091493.0/4294967296.0,1,-nbitq), 
to_sfixed(-226091253.0/4294967296.0,1,-nbitq), 
to_sfixed(177682387.0/4294967296.0,1,-nbitq), 
to_sfixed(52964445.0/4294967296.0,1,-nbitq), 
to_sfixed(52853398.0/4294967296.0,1,-nbitq), 
to_sfixed(98360231.0/4294967296.0,1,-nbitq), 
to_sfixed(59645195.0/4294967296.0,1,-nbitq), 
to_sfixed(-19588143.0/4294967296.0,1,-nbitq), 
to_sfixed(-218036453.0/4294967296.0,1,-nbitq), 
to_sfixed(-395953990.0/4294967296.0,1,-nbitq), 
to_sfixed(-85767429.0/4294967296.0,1,-nbitq), 
to_sfixed(92385464.0/4294967296.0,1,-nbitq), 
to_sfixed(31890279.0/4294967296.0,1,-nbitq), 
to_sfixed(63750476.0/4294967296.0,1,-nbitq), 
to_sfixed(204949674.0/4294967296.0,1,-nbitq), 
to_sfixed(284214914.0/4294967296.0,1,-nbitq), 
to_sfixed(377469286.0/4294967296.0,1,-nbitq), 
to_sfixed(263007549.0/4294967296.0,1,-nbitq), 
to_sfixed(61176393.0/4294967296.0,1,-nbitq), 
to_sfixed(-247671837.0/4294967296.0,1,-nbitq), 
to_sfixed(192378437.0/4294967296.0,1,-nbitq), 
to_sfixed(23957303.0/4294967296.0,1,-nbitq), 
to_sfixed(376463586.0/4294967296.0,1,-nbitq), 
to_sfixed(-159585521.0/4294967296.0,1,-nbitq), 
to_sfixed(76477573.0/4294967296.0,1,-nbitq), 
to_sfixed(68906188.0/4294967296.0,1,-nbitq), 
to_sfixed(60806674.0/4294967296.0,1,-nbitq), 
to_sfixed(209044260.0/4294967296.0,1,-nbitq), 
to_sfixed(-19392475.0/4294967296.0,1,-nbitq), 
to_sfixed(-38236542.0/4294967296.0,1,-nbitq), 
to_sfixed(120095327.0/4294967296.0,1,-nbitq), 
to_sfixed(-245651409.0/4294967296.0,1,-nbitq), 
to_sfixed(21705471.0/4294967296.0,1,-nbitq), 
to_sfixed(17196966.0/4294967296.0,1,-nbitq), 
to_sfixed(225792957.0/4294967296.0,1,-nbitq), 
to_sfixed(428910202.0/4294967296.0,1,-nbitq), 
to_sfixed(19892955.0/4294967296.0,1,-nbitq), 
to_sfixed(249171197.0/4294967296.0,1,-nbitq), 
to_sfixed(-434349569.0/4294967296.0,1,-nbitq), 
to_sfixed(-510256105.0/4294967296.0,1,-nbitq), 
to_sfixed(-285953118.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-402374978.0/4294967296.0,1,-nbitq), 
to_sfixed(-571232199.0/4294967296.0,1,-nbitq), 
to_sfixed(392349789.0/4294967296.0,1,-nbitq), 
to_sfixed(128898493.0/4294967296.0,1,-nbitq), 
to_sfixed(269736794.0/4294967296.0,1,-nbitq), 
to_sfixed(-133278331.0/4294967296.0,1,-nbitq), 
to_sfixed(347726238.0/4294967296.0,1,-nbitq), 
to_sfixed(-148377990.0/4294967296.0,1,-nbitq), 
to_sfixed(-125994708.0/4294967296.0,1,-nbitq), 
to_sfixed(73491543.0/4294967296.0,1,-nbitq), 
to_sfixed(256095362.0/4294967296.0,1,-nbitq), 
to_sfixed(573507318.0/4294967296.0,1,-nbitq), 
to_sfixed(-370376949.0/4294967296.0,1,-nbitq), 
to_sfixed(111013878.0/4294967296.0,1,-nbitq), 
to_sfixed(-8383519.0/4294967296.0,1,-nbitq), 
to_sfixed(140060221.0/4294967296.0,1,-nbitq), 
to_sfixed(-204533907.0/4294967296.0,1,-nbitq), 
to_sfixed(212331720.0/4294967296.0,1,-nbitq), 
to_sfixed(142704758.0/4294967296.0,1,-nbitq), 
to_sfixed(241909629.0/4294967296.0,1,-nbitq), 
to_sfixed(143701291.0/4294967296.0,1,-nbitq), 
to_sfixed(-158032523.0/4294967296.0,1,-nbitq), 
to_sfixed(567835832.0/4294967296.0,1,-nbitq), 
to_sfixed(-134022054.0/4294967296.0,1,-nbitq), 
to_sfixed(233182776.0/4294967296.0,1,-nbitq), 
to_sfixed(-72877655.0/4294967296.0,1,-nbitq), 
to_sfixed(418867071.0/4294967296.0,1,-nbitq), 
to_sfixed(-309935363.0/4294967296.0,1,-nbitq), 
to_sfixed(380186309.0/4294967296.0,1,-nbitq), 
to_sfixed(317926134.0/4294967296.0,1,-nbitq), 
to_sfixed(-596745821.0/4294967296.0,1,-nbitq), 
to_sfixed(-361540926.0/4294967296.0,1,-nbitq), 
to_sfixed(233731393.0/4294967296.0,1,-nbitq), 
to_sfixed(-365613522.0/4294967296.0,1,-nbitq), 
to_sfixed(458569504.0/4294967296.0,1,-nbitq), 
to_sfixed(150383694.0/4294967296.0,1,-nbitq), 
to_sfixed(357586132.0/4294967296.0,1,-nbitq), 
to_sfixed(406851917.0/4294967296.0,1,-nbitq), 
to_sfixed(-276438093.0/4294967296.0,1,-nbitq), 
to_sfixed(129572848.0/4294967296.0,1,-nbitq), 
to_sfixed(-409574631.0/4294967296.0,1,-nbitq), 
to_sfixed(120223475.0/4294967296.0,1,-nbitq), 
to_sfixed(-245670441.0/4294967296.0,1,-nbitq), 
to_sfixed(42234279.0/4294967296.0,1,-nbitq), 
to_sfixed(255730540.0/4294967296.0,1,-nbitq), 
to_sfixed(104767973.0/4294967296.0,1,-nbitq), 
to_sfixed(-204410980.0/4294967296.0,1,-nbitq), 
to_sfixed(48751701.0/4294967296.0,1,-nbitq), 
to_sfixed(74188721.0/4294967296.0,1,-nbitq), 
to_sfixed(176270664.0/4294967296.0,1,-nbitq), 
to_sfixed(260890101.0/4294967296.0,1,-nbitq), 
to_sfixed(66616811.0/4294967296.0,1,-nbitq), 
to_sfixed(29453455.0/4294967296.0,1,-nbitq), 
to_sfixed(-18051629.0/4294967296.0,1,-nbitq), 
to_sfixed(151206713.0/4294967296.0,1,-nbitq), 
to_sfixed(80293001.0/4294967296.0,1,-nbitq), 
to_sfixed(335461647.0/4294967296.0,1,-nbitq), 
to_sfixed(66755244.0/4294967296.0,1,-nbitq), 
to_sfixed(158161893.0/4294967296.0,1,-nbitq), 
to_sfixed(-248343592.0/4294967296.0,1,-nbitq), 
to_sfixed(-176948386.0/4294967296.0,1,-nbitq), 
to_sfixed(8275010.0/4294967296.0,1,-nbitq), 
to_sfixed(-529172188.0/4294967296.0,1,-nbitq), 
to_sfixed(393504978.0/4294967296.0,1,-nbitq), 
to_sfixed(-147160965.0/4294967296.0,1,-nbitq), 
to_sfixed(-419434203.0/4294967296.0,1,-nbitq), 
to_sfixed(657884485.0/4294967296.0,1,-nbitq), 
to_sfixed(191297137.0/4294967296.0,1,-nbitq), 
to_sfixed(216490318.0/4294967296.0,1,-nbitq), 
to_sfixed(315254580.0/4294967296.0,1,-nbitq), 
to_sfixed(69032030.0/4294967296.0,1,-nbitq), 
to_sfixed(-173901688.0/4294967296.0,1,-nbitq), 
to_sfixed(38301738.0/4294967296.0,1,-nbitq), 
to_sfixed(3119837.0/4294967296.0,1,-nbitq), 
to_sfixed(224177463.0/4294967296.0,1,-nbitq), 
to_sfixed(-111661049.0/4294967296.0,1,-nbitq), 
to_sfixed(429864604.0/4294967296.0,1,-nbitq), 
to_sfixed(-172369824.0/4294967296.0,1,-nbitq), 
to_sfixed(-395566617.0/4294967296.0,1,-nbitq), 
to_sfixed(-324634697.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-25510979.0/4294967296.0,1,-nbitq), 
to_sfixed(34376355.0/4294967296.0,1,-nbitq), 
to_sfixed(21698315.0/4294967296.0,1,-nbitq), 
to_sfixed(41837925.0/4294967296.0,1,-nbitq), 
to_sfixed(-197256590.0/4294967296.0,1,-nbitq), 
to_sfixed(301789700.0/4294967296.0,1,-nbitq), 
to_sfixed(375866833.0/4294967296.0,1,-nbitq), 
to_sfixed(-47510182.0/4294967296.0,1,-nbitq), 
to_sfixed(-11974987.0/4294967296.0,1,-nbitq), 
to_sfixed(296805530.0/4294967296.0,1,-nbitq), 
to_sfixed(-20927461.0/4294967296.0,1,-nbitq), 
to_sfixed(462973093.0/4294967296.0,1,-nbitq), 
to_sfixed(233775459.0/4294967296.0,1,-nbitq), 
to_sfixed(-223635162.0/4294967296.0,1,-nbitq), 
to_sfixed(-65317311.0/4294967296.0,1,-nbitq), 
to_sfixed(47397316.0/4294967296.0,1,-nbitq), 
to_sfixed(42184980.0/4294967296.0,1,-nbitq), 
to_sfixed(-394518129.0/4294967296.0,1,-nbitq), 
to_sfixed(-328111843.0/4294967296.0,1,-nbitq), 
to_sfixed(-411954858.0/4294967296.0,1,-nbitq), 
to_sfixed(230995298.0/4294967296.0,1,-nbitq), 
to_sfixed(411775088.0/4294967296.0,1,-nbitq), 
to_sfixed(408000622.0/4294967296.0,1,-nbitq), 
to_sfixed(-153390023.0/4294967296.0,1,-nbitq), 
to_sfixed(-57377792.0/4294967296.0,1,-nbitq), 
to_sfixed(62173879.0/4294967296.0,1,-nbitq), 
to_sfixed(-189232303.0/4294967296.0,1,-nbitq), 
to_sfixed(-534520802.0/4294967296.0,1,-nbitq), 
to_sfixed(312804670.0/4294967296.0,1,-nbitq), 
to_sfixed(-198904223.0/4294967296.0,1,-nbitq), 
to_sfixed(-314187940.0/4294967296.0,1,-nbitq), 
to_sfixed(57918682.0/4294967296.0,1,-nbitq), 
to_sfixed(-102039677.0/4294967296.0,1,-nbitq), 
to_sfixed(-172094382.0/4294967296.0,1,-nbitq), 
to_sfixed(68501327.0/4294967296.0,1,-nbitq), 
to_sfixed(-243695799.0/4294967296.0,1,-nbitq), 
to_sfixed(400838096.0/4294967296.0,1,-nbitq), 
to_sfixed(331254035.0/4294967296.0,1,-nbitq), 
to_sfixed(-59708637.0/4294967296.0,1,-nbitq), 
to_sfixed(416184702.0/4294967296.0,1,-nbitq), 
to_sfixed(-94707050.0/4294967296.0,1,-nbitq), 
to_sfixed(-1002780.0/4294967296.0,1,-nbitq), 
to_sfixed(-216093432.0/4294967296.0,1,-nbitq), 
to_sfixed(310911808.0/4294967296.0,1,-nbitq), 
to_sfixed(-121917193.0/4294967296.0,1,-nbitq), 
to_sfixed(79813241.0/4294967296.0,1,-nbitq), 
to_sfixed(66966335.0/4294967296.0,1,-nbitq), 
to_sfixed(-212738259.0/4294967296.0,1,-nbitq), 
to_sfixed(148975666.0/4294967296.0,1,-nbitq), 
to_sfixed(-131669791.0/4294967296.0,1,-nbitq), 
to_sfixed(71588180.0/4294967296.0,1,-nbitq), 
to_sfixed(-92015688.0/4294967296.0,1,-nbitq), 
to_sfixed(-263785419.0/4294967296.0,1,-nbitq), 
to_sfixed(34733652.0/4294967296.0,1,-nbitq), 
to_sfixed(-140768930.0/4294967296.0,1,-nbitq), 
to_sfixed(-112507795.0/4294967296.0,1,-nbitq), 
to_sfixed(-248790457.0/4294967296.0,1,-nbitq), 
to_sfixed(-523570410.0/4294967296.0,1,-nbitq), 
to_sfixed(347655114.0/4294967296.0,1,-nbitq), 
to_sfixed(-35680772.0/4294967296.0,1,-nbitq), 
to_sfixed(214498900.0/4294967296.0,1,-nbitq), 
to_sfixed(186866434.0/4294967296.0,1,-nbitq), 
to_sfixed(-228826450.0/4294967296.0,1,-nbitq), 
to_sfixed(186900557.0/4294967296.0,1,-nbitq), 
to_sfixed(-208134022.0/4294967296.0,1,-nbitq), 
to_sfixed(322045941.0/4294967296.0,1,-nbitq), 
to_sfixed(751264919.0/4294967296.0,1,-nbitq), 
to_sfixed(-147458604.0/4294967296.0,1,-nbitq), 
to_sfixed(24548029.0/4294967296.0,1,-nbitq), 
to_sfixed(-74619896.0/4294967296.0,1,-nbitq), 
to_sfixed(383230242.0/4294967296.0,1,-nbitq), 
to_sfixed(-169093700.0/4294967296.0,1,-nbitq), 
to_sfixed(-550180907.0/4294967296.0,1,-nbitq), 
to_sfixed(119057571.0/4294967296.0,1,-nbitq), 
to_sfixed(128313469.0/4294967296.0,1,-nbitq), 
to_sfixed(-195393515.0/4294967296.0,1,-nbitq), 
to_sfixed(-23711021.0/4294967296.0,1,-nbitq), 
to_sfixed(-158657484.0/4294967296.0,1,-nbitq), 
to_sfixed(-121337871.0/4294967296.0,1,-nbitq), 
to_sfixed(366666424.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(363772230.0/4294967296.0,1,-nbitq), 
to_sfixed(142309078.0/4294967296.0,1,-nbitq), 
to_sfixed(147930640.0/4294967296.0,1,-nbitq), 
to_sfixed(-173080545.0/4294967296.0,1,-nbitq), 
to_sfixed(340323424.0/4294967296.0,1,-nbitq), 
to_sfixed(257753679.0/4294967296.0,1,-nbitq), 
to_sfixed(89529008.0/4294967296.0,1,-nbitq), 
to_sfixed(213031097.0/4294967296.0,1,-nbitq), 
to_sfixed(-58258732.0/4294967296.0,1,-nbitq), 
to_sfixed(122984138.0/4294967296.0,1,-nbitq), 
to_sfixed(-398103012.0/4294967296.0,1,-nbitq), 
to_sfixed(178623706.0/4294967296.0,1,-nbitq), 
to_sfixed(101540398.0/4294967296.0,1,-nbitq), 
to_sfixed(424594022.0/4294967296.0,1,-nbitq), 
to_sfixed(358769568.0/4294967296.0,1,-nbitq), 
to_sfixed(-293057753.0/4294967296.0,1,-nbitq), 
to_sfixed(-249466800.0/4294967296.0,1,-nbitq), 
to_sfixed(-215435262.0/4294967296.0,1,-nbitq), 
to_sfixed(134640813.0/4294967296.0,1,-nbitq), 
to_sfixed(115275876.0/4294967296.0,1,-nbitq), 
to_sfixed(148066879.0/4294967296.0,1,-nbitq), 
to_sfixed(424405566.0/4294967296.0,1,-nbitq), 
to_sfixed(-2632965.0/4294967296.0,1,-nbitq), 
to_sfixed(-150212404.0/4294967296.0,1,-nbitq), 
to_sfixed(281771042.0/4294967296.0,1,-nbitq), 
to_sfixed(295271950.0/4294967296.0,1,-nbitq), 
to_sfixed(248465058.0/4294967296.0,1,-nbitq), 
to_sfixed(-268185023.0/4294967296.0,1,-nbitq), 
to_sfixed(468227658.0/4294967296.0,1,-nbitq), 
to_sfixed(-194317707.0/4294967296.0,1,-nbitq), 
to_sfixed(-585837797.0/4294967296.0,1,-nbitq), 
to_sfixed(-457121717.0/4294967296.0,1,-nbitq), 
to_sfixed(143973440.0/4294967296.0,1,-nbitq), 
to_sfixed(32877961.0/4294967296.0,1,-nbitq), 
to_sfixed(414843873.0/4294967296.0,1,-nbitq), 
to_sfixed(309852880.0/4294967296.0,1,-nbitq), 
to_sfixed(521599374.0/4294967296.0,1,-nbitq), 
to_sfixed(339383864.0/4294967296.0,1,-nbitq), 
to_sfixed(-195452131.0/4294967296.0,1,-nbitq), 
to_sfixed(93717022.0/4294967296.0,1,-nbitq), 
to_sfixed(-296835130.0/4294967296.0,1,-nbitq), 
to_sfixed(-137380432.0/4294967296.0,1,-nbitq), 
to_sfixed(112169290.0/4294967296.0,1,-nbitq), 
to_sfixed(-123222097.0/4294967296.0,1,-nbitq), 
to_sfixed(-60431422.0/4294967296.0,1,-nbitq), 
to_sfixed(360363034.0/4294967296.0,1,-nbitq), 
to_sfixed(-415041476.0/4294967296.0,1,-nbitq), 
to_sfixed(-379496981.0/4294967296.0,1,-nbitq), 
to_sfixed(-213958578.0/4294967296.0,1,-nbitq), 
to_sfixed(449859423.0/4294967296.0,1,-nbitq), 
to_sfixed(-276308212.0/4294967296.0,1,-nbitq), 
to_sfixed(-253202897.0/4294967296.0,1,-nbitq), 
to_sfixed(-172355243.0/4294967296.0,1,-nbitq), 
to_sfixed(230541102.0/4294967296.0,1,-nbitq), 
to_sfixed(-180409123.0/4294967296.0,1,-nbitq), 
to_sfixed(-332984234.0/4294967296.0,1,-nbitq), 
to_sfixed(348190620.0/4294967296.0,1,-nbitq), 
to_sfixed(-14861134.0/4294967296.0,1,-nbitq), 
to_sfixed(-323909606.0/4294967296.0,1,-nbitq), 
to_sfixed(-305530336.0/4294967296.0,1,-nbitq), 
to_sfixed(162104443.0/4294967296.0,1,-nbitq), 
to_sfixed(-155611534.0/4294967296.0,1,-nbitq), 
to_sfixed(94795659.0/4294967296.0,1,-nbitq), 
to_sfixed(437789587.0/4294967296.0,1,-nbitq), 
to_sfixed(99346290.0/4294967296.0,1,-nbitq), 
to_sfixed(-274921813.0/4294967296.0,1,-nbitq), 
to_sfixed(63136805.0/4294967296.0,1,-nbitq), 
to_sfixed(-7816079.0/4294967296.0,1,-nbitq), 
to_sfixed(361603137.0/4294967296.0,1,-nbitq), 
to_sfixed(479532835.0/4294967296.0,1,-nbitq), 
to_sfixed(-35021405.0/4294967296.0,1,-nbitq), 
to_sfixed(-224074259.0/4294967296.0,1,-nbitq), 
to_sfixed(105025020.0/4294967296.0,1,-nbitq), 
to_sfixed(167871865.0/4294967296.0,1,-nbitq), 
to_sfixed(378053996.0/4294967296.0,1,-nbitq), 
to_sfixed(36745903.0/4294967296.0,1,-nbitq), 
to_sfixed(153186766.0/4294967296.0,1,-nbitq), 
to_sfixed(-195100622.0/4294967296.0,1,-nbitq), 
to_sfixed(-436378062.0/4294967296.0,1,-nbitq), 
to_sfixed(-97815047.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(26988181.0/4294967296.0,1,-nbitq), 
to_sfixed(-378061365.0/4294967296.0,1,-nbitq), 
to_sfixed(455141739.0/4294967296.0,1,-nbitq), 
to_sfixed(310325604.0/4294967296.0,1,-nbitq), 
to_sfixed(311069190.0/4294967296.0,1,-nbitq), 
to_sfixed(94439702.0/4294967296.0,1,-nbitq), 
to_sfixed(401143581.0/4294967296.0,1,-nbitq), 
to_sfixed(115071041.0/4294967296.0,1,-nbitq), 
to_sfixed(-19141580.0/4294967296.0,1,-nbitq), 
to_sfixed(74633271.0/4294967296.0,1,-nbitq), 
to_sfixed(415032261.0/4294967296.0,1,-nbitq), 
to_sfixed(421884398.0/4294967296.0,1,-nbitq), 
to_sfixed(148646202.0/4294967296.0,1,-nbitq), 
to_sfixed(577956412.0/4294967296.0,1,-nbitq), 
to_sfixed(-92735209.0/4294967296.0,1,-nbitq), 
to_sfixed(283819557.0/4294967296.0,1,-nbitq), 
to_sfixed(-193803829.0/4294967296.0,1,-nbitq), 
to_sfixed(364300726.0/4294967296.0,1,-nbitq), 
to_sfixed(-158814309.0/4294967296.0,1,-nbitq), 
to_sfixed(-385524108.0/4294967296.0,1,-nbitq), 
to_sfixed(20580488.0/4294967296.0,1,-nbitq), 
to_sfixed(-102321045.0/4294967296.0,1,-nbitq), 
to_sfixed(558886372.0/4294967296.0,1,-nbitq), 
to_sfixed(-109449320.0/4294967296.0,1,-nbitq), 
to_sfixed(408954007.0/4294967296.0,1,-nbitq), 
to_sfixed(-121148869.0/4294967296.0,1,-nbitq), 
to_sfixed(-135675373.0/4294967296.0,1,-nbitq), 
to_sfixed(-51210641.0/4294967296.0,1,-nbitq), 
to_sfixed(-32500638.0/4294967296.0,1,-nbitq), 
to_sfixed(126474529.0/4294967296.0,1,-nbitq), 
to_sfixed(-512020306.0/4294967296.0,1,-nbitq), 
to_sfixed(-445321895.0/4294967296.0,1,-nbitq), 
to_sfixed(186751306.0/4294967296.0,1,-nbitq), 
to_sfixed(59797934.0/4294967296.0,1,-nbitq), 
to_sfixed(-79695518.0/4294967296.0,1,-nbitq), 
to_sfixed(204588178.0/4294967296.0,1,-nbitq), 
to_sfixed(-191448363.0/4294967296.0,1,-nbitq), 
to_sfixed(450005570.0/4294967296.0,1,-nbitq), 
to_sfixed(315068184.0/4294967296.0,1,-nbitq), 
to_sfixed(371290977.0/4294967296.0,1,-nbitq), 
to_sfixed(-421391337.0/4294967296.0,1,-nbitq), 
to_sfixed(89578209.0/4294967296.0,1,-nbitq), 
to_sfixed(-158631339.0/4294967296.0,1,-nbitq), 
to_sfixed(-257116817.0/4294967296.0,1,-nbitq), 
to_sfixed(179894612.0/4294967296.0,1,-nbitq), 
to_sfixed(268972213.0/4294967296.0,1,-nbitq), 
to_sfixed(-276586371.0/4294967296.0,1,-nbitq), 
to_sfixed(66362677.0/4294967296.0,1,-nbitq), 
to_sfixed(293116092.0/4294967296.0,1,-nbitq), 
to_sfixed(335259136.0/4294967296.0,1,-nbitq), 
to_sfixed(-327878423.0/4294967296.0,1,-nbitq), 
to_sfixed(-10684045.0/4294967296.0,1,-nbitq), 
to_sfixed(-663221132.0/4294967296.0,1,-nbitq), 
to_sfixed(-87583833.0/4294967296.0,1,-nbitq), 
to_sfixed(78624437.0/4294967296.0,1,-nbitq), 
to_sfixed(-275093647.0/4294967296.0,1,-nbitq), 
to_sfixed(-323488039.0/4294967296.0,1,-nbitq), 
to_sfixed(111005380.0/4294967296.0,1,-nbitq), 
to_sfixed(-7492145.0/4294967296.0,1,-nbitq), 
to_sfixed(232580817.0/4294967296.0,1,-nbitq), 
to_sfixed(24231074.0/4294967296.0,1,-nbitq), 
to_sfixed(-95767554.0/4294967296.0,1,-nbitq), 
to_sfixed(102815335.0/4294967296.0,1,-nbitq), 
to_sfixed(74367455.0/4294967296.0,1,-nbitq), 
to_sfixed(321556551.0/4294967296.0,1,-nbitq), 
to_sfixed(-100442076.0/4294967296.0,1,-nbitq), 
to_sfixed(749025401.0/4294967296.0,1,-nbitq), 
to_sfixed(-235795663.0/4294967296.0,1,-nbitq), 
to_sfixed(54320555.0/4294967296.0,1,-nbitq), 
to_sfixed(481293187.0/4294967296.0,1,-nbitq), 
to_sfixed(-318996382.0/4294967296.0,1,-nbitq), 
to_sfixed(119123605.0/4294967296.0,1,-nbitq), 
to_sfixed(166695021.0/4294967296.0,1,-nbitq), 
to_sfixed(-94582710.0/4294967296.0,1,-nbitq), 
to_sfixed(438469197.0/4294967296.0,1,-nbitq), 
to_sfixed(-382046868.0/4294967296.0,1,-nbitq), 
to_sfixed(-324865161.0/4294967296.0,1,-nbitq), 
to_sfixed(-440795410.0/4294967296.0,1,-nbitq), 
to_sfixed(-81748943.0/4294967296.0,1,-nbitq), 
to_sfixed(-39793455.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(248875802.0/4294967296.0,1,-nbitq), 
to_sfixed(147556723.0/4294967296.0,1,-nbitq), 
to_sfixed(-312172639.0/4294967296.0,1,-nbitq), 
to_sfixed(198165970.0/4294967296.0,1,-nbitq), 
to_sfixed(-214072651.0/4294967296.0,1,-nbitq), 
to_sfixed(228011614.0/4294967296.0,1,-nbitq), 
to_sfixed(-125990091.0/4294967296.0,1,-nbitq), 
to_sfixed(226355551.0/4294967296.0,1,-nbitq), 
to_sfixed(244769669.0/4294967296.0,1,-nbitq), 
to_sfixed(-153656900.0/4294967296.0,1,-nbitq), 
to_sfixed(-137867132.0/4294967296.0,1,-nbitq), 
to_sfixed(451646888.0/4294967296.0,1,-nbitq), 
to_sfixed(-372843920.0/4294967296.0,1,-nbitq), 
to_sfixed(392317406.0/4294967296.0,1,-nbitq), 
to_sfixed(254486312.0/4294967296.0,1,-nbitq), 
to_sfixed(-839082.0/4294967296.0,1,-nbitq), 
to_sfixed(-334074953.0/4294967296.0,1,-nbitq), 
to_sfixed(364110947.0/4294967296.0,1,-nbitq), 
to_sfixed(-34489144.0/4294967296.0,1,-nbitq), 
to_sfixed(-249792437.0/4294967296.0,1,-nbitq), 
to_sfixed(143187097.0/4294967296.0,1,-nbitq), 
to_sfixed(-144487582.0/4294967296.0,1,-nbitq), 
to_sfixed(-54480743.0/4294967296.0,1,-nbitq), 
to_sfixed(-133215275.0/4294967296.0,1,-nbitq), 
to_sfixed(364930322.0/4294967296.0,1,-nbitq), 
to_sfixed(-174952796.0/4294967296.0,1,-nbitq), 
to_sfixed(161422666.0/4294967296.0,1,-nbitq), 
to_sfixed(66808898.0/4294967296.0,1,-nbitq), 
to_sfixed(352527446.0/4294967296.0,1,-nbitq), 
to_sfixed(418062069.0/4294967296.0,1,-nbitq), 
to_sfixed(-176796775.0/4294967296.0,1,-nbitq), 
to_sfixed(130747928.0/4294967296.0,1,-nbitq), 
to_sfixed(-145928488.0/4294967296.0,1,-nbitq), 
to_sfixed(-437412649.0/4294967296.0,1,-nbitq), 
to_sfixed(330369872.0/4294967296.0,1,-nbitq), 
to_sfixed(110361846.0/4294967296.0,1,-nbitq), 
to_sfixed(-236302026.0/4294967296.0,1,-nbitq), 
to_sfixed(-141543050.0/4294967296.0,1,-nbitq), 
to_sfixed(-347142241.0/4294967296.0,1,-nbitq), 
to_sfixed(318182997.0/4294967296.0,1,-nbitq), 
to_sfixed(-456521414.0/4294967296.0,1,-nbitq), 
to_sfixed(395074648.0/4294967296.0,1,-nbitq), 
to_sfixed(220331652.0/4294967296.0,1,-nbitq), 
to_sfixed(376065360.0/4294967296.0,1,-nbitq), 
to_sfixed(424506222.0/4294967296.0,1,-nbitq), 
to_sfixed(275560625.0/4294967296.0,1,-nbitq), 
to_sfixed(-212495056.0/4294967296.0,1,-nbitq), 
to_sfixed(-314013778.0/4294967296.0,1,-nbitq), 
to_sfixed(156832076.0/4294967296.0,1,-nbitq), 
to_sfixed(450716119.0/4294967296.0,1,-nbitq), 
to_sfixed(55722043.0/4294967296.0,1,-nbitq), 
to_sfixed(419617348.0/4294967296.0,1,-nbitq), 
to_sfixed(-475034602.0/4294967296.0,1,-nbitq), 
to_sfixed(274822360.0/4294967296.0,1,-nbitq), 
to_sfixed(315366835.0/4294967296.0,1,-nbitq), 
to_sfixed(-40754538.0/4294967296.0,1,-nbitq), 
to_sfixed(43690732.0/4294967296.0,1,-nbitq), 
to_sfixed(-279180937.0/4294967296.0,1,-nbitq), 
to_sfixed(425969649.0/4294967296.0,1,-nbitq), 
to_sfixed(-42847427.0/4294967296.0,1,-nbitq), 
to_sfixed(-12604144.0/4294967296.0,1,-nbitq), 
to_sfixed(408215396.0/4294967296.0,1,-nbitq), 
to_sfixed(-262332180.0/4294967296.0,1,-nbitq), 
to_sfixed(261750797.0/4294967296.0,1,-nbitq), 
to_sfixed(-50572060.0/4294967296.0,1,-nbitq), 
to_sfixed(-131502034.0/4294967296.0,1,-nbitq), 
to_sfixed(552186882.0/4294967296.0,1,-nbitq), 
to_sfixed(-354278945.0/4294967296.0,1,-nbitq), 
to_sfixed(191994870.0/4294967296.0,1,-nbitq), 
to_sfixed(-205619104.0/4294967296.0,1,-nbitq), 
to_sfixed(-202491597.0/4294967296.0,1,-nbitq), 
to_sfixed(-84131478.0/4294967296.0,1,-nbitq), 
to_sfixed(-547744679.0/4294967296.0,1,-nbitq), 
to_sfixed(-208684466.0/4294967296.0,1,-nbitq), 
to_sfixed(28949731.0/4294967296.0,1,-nbitq), 
to_sfixed(-444918197.0/4294967296.0,1,-nbitq), 
to_sfixed(121755952.0/4294967296.0,1,-nbitq), 
to_sfixed(36107263.0/4294967296.0,1,-nbitq), 
to_sfixed(200210529.0/4294967296.0,1,-nbitq), 
to_sfixed(354474903.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-290658408.0/4294967296.0,1,-nbitq), 
to_sfixed(68121589.0/4294967296.0,1,-nbitq), 
to_sfixed(-210596141.0/4294967296.0,1,-nbitq), 
to_sfixed(-211425620.0/4294967296.0,1,-nbitq), 
to_sfixed(369794427.0/4294967296.0,1,-nbitq), 
to_sfixed(-386710695.0/4294967296.0,1,-nbitq), 
to_sfixed(373466330.0/4294967296.0,1,-nbitq), 
to_sfixed(-328658701.0/4294967296.0,1,-nbitq), 
to_sfixed(366091721.0/4294967296.0,1,-nbitq), 
to_sfixed(-248949859.0/4294967296.0,1,-nbitq), 
to_sfixed(-9623226.0/4294967296.0,1,-nbitq), 
to_sfixed(117936536.0/4294967296.0,1,-nbitq), 
to_sfixed(-318129493.0/4294967296.0,1,-nbitq), 
to_sfixed(531229524.0/4294967296.0,1,-nbitq), 
to_sfixed(-321857974.0/4294967296.0,1,-nbitq), 
to_sfixed(265085384.0/4294967296.0,1,-nbitq), 
to_sfixed(-57164069.0/4294967296.0,1,-nbitq), 
to_sfixed(132700035.0/4294967296.0,1,-nbitq), 
to_sfixed(-405363706.0/4294967296.0,1,-nbitq), 
to_sfixed(114396136.0/4294967296.0,1,-nbitq), 
to_sfixed(-187543475.0/4294967296.0,1,-nbitq), 
to_sfixed(-172357194.0/4294967296.0,1,-nbitq), 
to_sfixed(288304501.0/4294967296.0,1,-nbitq), 
to_sfixed(-414186519.0/4294967296.0,1,-nbitq), 
to_sfixed(-316310651.0/4294967296.0,1,-nbitq), 
to_sfixed(366603225.0/4294967296.0,1,-nbitq), 
to_sfixed(266525382.0/4294967296.0,1,-nbitq), 
to_sfixed(63065521.0/4294967296.0,1,-nbitq), 
to_sfixed(129552416.0/4294967296.0,1,-nbitq), 
to_sfixed(-222171850.0/4294967296.0,1,-nbitq), 
to_sfixed(117763565.0/4294967296.0,1,-nbitq), 
to_sfixed(-417243371.0/4294967296.0,1,-nbitq), 
to_sfixed(67789265.0/4294967296.0,1,-nbitq), 
to_sfixed(-516402501.0/4294967296.0,1,-nbitq), 
to_sfixed(-198693666.0/4294967296.0,1,-nbitq), 
to_sfixed(-200385510.0/4294967296.0,1,-nbitq), 
to_sfixed(70600603.0/4294967296.0,1,-nbitq), 
to_sfixed(48296367.0/4294967296.0,1,-nbitq), 
to_sfixed(-437679202.0/4294967296.0,1,-nbitq), 
to_sfixed(-63320637.0/4294967296.0,1,-nbitq), 
to_sfixed(8760996.0/4294967296.0,1,-nbitq), 
to_sfixed(-193581729.0/4294967296.0,1,-nbitq), 
to_sfixed(-78163681.0/4294967296.0,1,-nbitq), 
to_sfixed(-318201011.0/4294967296.0,1,-nbitq), 
to_sfixed(183980706.0/4294967296.0,1,-nbitq), 
to_sfixed(291288153.0/4294967296.0,1,-nbitq), 
to_sfixed(161378334.0/4294967296.0,1,-nbitq), 
to_sfixed(152236282.0/4294967296.0,1,-nbitq), 
to_sfixed(12270284.0/4294967296.0,1,-nbitq), 
to_sfixed(106848005.0/4294967296.0,1,-nbitq), 
to_sfixed(238858480.0/4294967296.0,1,-nbitq), 
to_sfixed(48902231.0/4294967296.0,1,-nbitq), 
to_sfixed(-124280482.0/4294967296.0,1,-nbitq), 
to_sfixed(153934792.0/4294967296.0,1,-nbitq), 
to_sfixed(-90300636.0/4294967296.0,1,-nbitq), 
to_sfixed(-290671430.0/4294967296.0,1,-nbitq), 
to_sfixed(389721980.0/4294967296.0,1,-nbitq), 
to_sfixed(224051027.0/4294967296.0,1,-nbitq), 
to_sfixed(371312911.0/4294967296.0,1,-nbitq), 
to_sfixed(361299146.0/4294967296.0,1,-nbitq), 
to_sfixed(177430387.0/4294967296.0,1,-nbitq), 
to_sfixed(165919576.0/4294967296.0,1,-nbitq), 
to_sfixed(-129868924.0/4294967296.0,1,-nbitq), 
to_sfixed(-76862499.0/4294967296.0,1,-nbitq), 
to_sfixed(-37712980.0/4294967296.0,1,-nbitq), 
to_sfixed(-316335224.0/4294967296.0,1,-nbitq), 
to_sfixed(777902411.0/4294967296.0,1,-nbitq), 
to_sfixed(39356131.0/4294967296.0,1,-nbitq), 
to_sfixed(-177321180.0/4294967296.0,1,-nbitq), 
to_sfixed(-1605205.0/4294967296.0,1,-nbitq), 
to_sfixed(-61285996.0/4294967296.0,1,-nbitq), 
to_sfixed(463381667.0/4294967296.0,1,-nbitq), 
to_sfixed(-2083262.0/4294967296.0,1,-nbitq), 
to_sfixed(-316398673.0/4294967296.0,1,-nbitq), 
to_sfixed(289922624.0/4294967296.0,1,-nbitq), 
to_sfixed(61461391.0/4294967296.0,1,-nbitq), 
to_sfixed(-245251367.0/4294967296.0,1,-nbitq), 
to_sfixed(-120237291.0/4294967296.0,1,-nbitq), 
to_sfixed(-578602323.0/4294967296.0,1,-nbitq), 
to_sfixed(91959700.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(215489130.0/4294967296.0,1,-nbitq), 
to_sfixed(-152644966.0/4294967296.0,1,-nbitq), 
to_sfixed(395262050.0/4294967296.0,1,-nbitq), 
to_sfixed(302855733.0/4294967296.0,1,-nbitq), 
to_sfixed(429804709.0/4294967296.0,1,-nbitq), 
to_sfixed(-144932734.0/4294967296.0,1,-nbitq), 
to_sfixed(354781973.0/4294967296.0,1,-nbitq), 
to_sfixed(-466826571.0/4294967296.0,1,-nbitq), 
to_sfixed(-263583770.0/4294967296.0,1,-nbitq), 
to_sfixed(387646930.0/4294967296.0,1,-nbitq), 
to_sfixed(-245876225.0/4294967296.0,1,-nbitq), 
to_sfixed(579598059.0/4294967296.0,1,-nbitq), 
to_sfixed(-615490219.0/4294967296.0,1,-nbitq), 
to_sfixed(395215537.0/4294967296.0,1,-nbitq), 
to_sfixed(-309735194.0/4294967296.0,1,-nbitq), 
to_sfixed(-439034717.0/4294967296.0,1,-nbitq), 
to_sfixed(-378294287.0/4294967296.0,1,-nbitq), 
to_sfixed(-345252907.0/4294967296.0,1,-nbitq), 
to_sfixed(-269398547.0/4294967296.0,1,-nbitq), 
to_sfixed(-202212668.0/4294967296.0,1,-nbitq), 
to_sfixed(329122283.0/4294967296.0,1,-nbitq), 
to_sfixed(-129653893.0/4294967296.0,1,-nbitq), 
to_sfixed(422379158.0/4294967296.0,1,-nbitq), 
to_sfixed(-424972183.0/4294967296.0,1,-nbitq), 
to_sfixed(-38293140.0/4294967296.0,1,-nbitq), 
to_sfixed(97705923.0/4294967296.0,1,-nbitq), 
to_sfixed(29573837.0/4294967296.0,1,-nbitq), 
to_sfixed(118537073.0/4294967296.0,1,-nbitq), 
to_sfixed(271601100.0/4294967296.0,1,-nbitq), 
to_sfixed(13053676.0/4294967296.0,1,-nbitq), 
to_sfixed(-277929155.0/4294967296.0,1,-nbitq), 
to_sfixed(-196658216.0/4294967296.0,1,-nbitq), 
to_sfixed(80595559.0/4294967296.0,1,-nbitq), 
to_sfixed(108964771.0/4294967296.0,1,-nbitq), 
to_sfixed(425474149.0/4294967296.0,1,-nbitq), 
to_sfixed(286392165.0/4294967296.0,1,-nbitq), 
to_sfixed(520986378.0/4294967296.0,1,-nbitq), 
to_sfixed(172870636.0/4294967296.0,1,-nbitq), 
to_sfixed(107591465.0/4294967296.0,1,-nbitq), 
to_sfixed(219455494.0/4294967296.0,1,-nbitq), 
to_sfixed(-341208082.0/4294967296.0,1,-nbitq), 
to_sfixed(140504992.0/4294967296.0,1,-nbitq), 
to_sfixed(-102348391.0/4294967296.0,1,-nbitq), 
to_sfixed(-72180948.0/4294967296.0,1,-nbitq), 
to_sfixed(208813970.0/4294967296.0,1,-nbitq), 
to_sfixed(24233198.0/4294967296.0,1,-nbitq), 
to_sfixed(96782188.0/4294967296.0,1,-nbitq), 
to_sfixed(-219858327.0/4294967296.0,1,-nbitq), 
to_sfixed(265392670.0/4294967296.0,1,-nbitq), 
to_sfixed(285780727.0/4294967296.0,1,-nbitq), 
to_sfixed(161812006.0/4294967296.0,1,-nbitq), 
to_sfixed(-224605001.0/4294967296.0,1,-nbitq), 
to_sfixed(-648970220.0/4294967296.0,1,-nbitq), 
to_sfixed(448053904.0/4294967296.0,1,-nbitq), 
to_sfixed(495375687.0/4294967296.0,1,-nbitq), 
to_sfixed(98352009.0/4294967296.0,1,-nbitq), 
to_sfixed(363993148.0/4294967296.0,1,-nbitq), 
to_sfixed(76792468.0/4294967296.0,1,-nbitq), 
to_sfixed(234745543.0/4294967296.0,1,-nbitq), 
to_sfixed(154060766.0/4294967296.0,1,-nbitq), 
to_sfixed(-67749612.0/4294967296.0,1,-nbitq), 
to_sfixed(-318689806.0/4294967296.0,1,-nbitq), 
to_sfixed(268413396.0/4294967296.0,1,-nbitq), 
to_sfixed(158372563.0/4294967296.0,1,-nbitq), 
to_sfixed(-41909315.0/4294967296.0,1,-nbitq), 
to_sfixed(18008571.0/4294967296.0,1,-nbitq), 
to_sfixed(511362636.0/4294967296.0,1,-nbitq), 
to_sfixed(3554585.0/4294967296.0,1,-nbitq), 
to_sfixed(342615444.0/4294967296.0,1,-nbitq), 
to_sfixed(-340033359.0/4294967296.0,1,-nbitq), 
to_sfixed(-485114554.0/4294967296.0,1,-nbitq), 
to_sfixed(399105450.0/4294967296.0,1,-nbitq), 
to_sfixed(-332683536.0/4294967296.0,1,-nbitq), 
to_sfixed(-282121134.0/4294967296.0,1,-nbitq), 
to_sfixed(-196596663.0/4294967296.0,1,-nbitq), 
to_sfixed(-436915166.0/4294967296.0,1,-nbitq), 
to_sfixed(-548183973.0/4294967296.0,1,-nbitq), 
to_sfixed(-414734958.0/4294967296.0,1,-nbitq), 
to_sfixed(-480799748.0/4294967296.0,1,-nbitq), 
to_sfixed(-307007061.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(515370414.0/4294967296.0,1,-nbitq), 
to_sfixed(280535766.0/4294967296.0,1,-nbitq), 
to_sfixed(-261220835.0/4294967296.0,1,-nbitq), 
to_sfixed(-157360204.0/4294967296.0,1,-nbitq), 
to_sfixed(-191933001.0/4294967296.0,1,-nbitq), 
to_sfixed(-430666865.0/4294967296.0,1,-nbitq), 
to_sfixed(-233343592.0/4294967296.0,1,-nbitq), 
to_sfixed(-26767741.0/4294967296.0,1,-nbitq), 
to_sfixed(464737235.0/4294967296.0,1,-nbitq), 
to_sfixed(-71059709.0/4294967296.0,1,-nbitq), 
to_sfixed(86322979.0/4294967296.0,1,-nbitq), 
to_sfixed(390374451.0/4294967296.0,1,-nbitq), 
to_sfixed(21080020.0/4294967296.0,1,-nbitq), 
to_sfixed(68775338.0/4294967296.0,1,-nbitq), 
to_sfixed(-294418485.0/4294967296.0,1,-nbitq), 
to_sfixed(106809842.0/4294967296.0,1,-nbitq), 
to_sfixed(-241065545.0/4294967296.0,1,-nbitq), 
to_sfixed(-249034268.0/4294967296.0,1,-nbitq), 
to_sfixed(-18830222.0/4294967296.0,1,-nbitq), 
to_sfixed(308141743.0/4294967296.0,1,-nbitq), 
to_sfixed(136886092.0/4294967296.0,1,-nbitq), 
to_sfixed(416953201.0/4294967296.0,1,-nbitq), 
to_sfixed(-110696710.0/4294967296.0,1,-nbitq), 
to_sfixed(-458116179.0/4294967296.0,1,-nbitq), 
to_sfixed(352742380.0/4294967296.0,1,-nbitq), 
to_sfixed(-235642242.0/4294967296.0,1,-nbitq), 
to_sfixed(114564057.0/4294967296.0,1,-nbitq), 
to_sfixed(75490884.0/4294967296.0,1,-nbitq), 
to_sfixed(-25630669.0/4294967296.0,1,-nbitq), 
to_sfixed(-245870644.0/4294967296.0,1,-nbitq), 
to_sfixed(207908300.0/4294967296.0,1,-nbitq), 
to_sfixed(-396307251.0/4294967296.0,1,-nbitq), 
to_sfixed(-131866340.0/4294967296.0,1,-nbitq), 
to_sfixed(-35805567.0/4294967296.0,1,-nbitq), 
to_sfixed(-34570706.0/4294967296.0,1,-nbitq), 
to_sfixed(31448546.0/4294967296.0,1,-nbitq), 
to_sfixed(464435228.0/4294967296.0,1,-nbitq), 
to_sfixed(84379087.0/4294967296.0,1,-nbitq), 
to_sfixed(-28701417.0/4294967296.0,1,-nbitq), 
to_sfixed(-289724881.0/4294967296.0,1,-nbitq), 
to_sfixed(-67658402.0/4294967296.0,1,-nbitq), 
to_sfixed(309642909.0/4294967296.0,1,-nbitq), 
to_sfixed(-3525964.0/4294967296.0,1,-nbitq), 
to_sfixed(215117156.0/4294967296.0,1,-nbitq), 
to_sfixed(281065742.0/4294967296.0,1,-nbitq), 
to_sfixed(-107805148.0/4294967296.0,1,-nbitq), 
to_sfixed(132042426.0/4294967296.0,1,-nbitq), 
to_sfixed(-44551221.0/4294967296.0,1,-nbitq), 
to_sfixed(94173826.0/4294967296.0,1,-nbitq), 
to_sfixed(341601293.0/4294967296.0,1,-nbitq), 
to_sfixed(162822661.0/4294967296.0,1,-nbitq), 
to_sfixed(-143436358.0/4294967296.0,1,-nbitq), 
to_sfixed(-549886601.0/4294967296.0,1,-nbitq), 
to_sfixed(169097299.0/4294967296.0,1,-nbitq), 
to_sfixed(432552195.0/4294967296.0,1,-nbitq), 
to_sfixed(-9439636.0/4294967296.0,1,-nbitq), 
to_sfixed(181409604.0/4294967296.0,1,-nbitq), 
to_sfixed(-317638806.0/4294967296.0,1,-nbitq), 
to_sfixed(-10938379.0/4294967296.0,1,-nbitq), 
to_sfixed(154469938.0/4294967296.0,1,-nbitq), 
to_sfixed(-285428402.0/4294967296.0,1,-nbitq), 
to_sfixed(76737368.0/4294967296.0,1,-nbitq), 
to_sfixed(-156103287.0/4294967296.0,1,-nbitq), 
to_sfixed(199982373.0/4294967296.0,1,-nbitq), 
to_sfixed(337092683.0/4294967296.0,1,-nbitq), 
to_sfixed(77580127.0/4294967296.0,1,-nbitq), 
to_sfixed(554273322.0/4294967296.0,1,-nbitq), 
to_sfixed(-7914221.0/4294967296.0,1,-nbitq), 
to_sfixed(301087591.0/4294967296.0,1,-nbitq), 
to_sfixed(-128730802.0/4294967296.0,1,-nbitq), 
to_sfixed(182799194.0/4294967296.0,1,-nbitq), 
to_sfixed(-246359512.0/4294967296.0,1,-nbitq), 
to_sfixed(-193461447.0/4294967296.0,1,-nbitq), 
to_sfixed(-220029101.0/4294967296.0,1,-nbitq), 
to_sfixed(20369055.0/4294967296.0,1,-nbitq), 
to_sfixed(4539441.0/4294967296.0,1,-nbitq), 
to_sfixed(-476952449.0/4294967296.0,1,-nbitq), 
to_sfixed(-493021270.0/4294967296.0,1,-nbitq), 
to_sfixed(-126944382.0/4294967296.0,1,-nbitq), 
to_sfixed(-365434691.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(74272072.0/4294967296.0,1,-nbitq), 
to_sfixed(417735439.0/4294967296.0,1,-nbitq), 
to_sfixed(303590583.0/4294967296.0,1,-nbitq), 
to_sfixed(-282058865.0/4294967296.0,1,-nbitq), 
to_sfixed(468594619.0/4294967296.0,1,-nbitq), 
to_sfixed(-164350203.0/4294967296.0,1,-nbitq), 
to_sfixed(-223024891.0/4294967296.0,1,-nbitq), 
to_sfixed(204636729.0/4294967296.0,1,-nbitq), 
to_sfixed(421567682.0/4294967296.0,1,-nbitq), 
to_sfixed(-65366712.0/4294967296.0,1,-nbitq), 
to_sfixed(-80764410.0/4294967296.0,1,-nbitq), 
to_sfixed(376765876.0/4294967296.0,1,-nbitq), 
to_sfixed(-389148119.0/4294967296.0,1,-nbitq), 
to_sfixed(482470367.0/4294967296.0,1,-nbitq), 
to_sfixed(382241732.0/4294967296.0,1,-nbitq), 
to_sfixed(-384228819.0/4294967296.0,1,-nbitq), 
to_sfixed(-30833193.0/4294967296.0,1,-nbitq), 
to_sfixed(352118701.0/4294967296.0,1,-nbitq), 
to_sfixed(187788401.0/4294967296.0,1,-nbitq), 
to_sfixed(-166793480.0/4294967296.0,1,-nbitq), 
to_sfixed(165349818.0/4294967296.0,1,-nbitq), 
to_sfixed(-285091468.0/4294967296.0,1,-nbitq), 
to_sfixed(-170388673.0/4294967296.0,1,-nbitq), 
to_sfixed(-163086310.0/4294967296.0,1,-nbitq), 
to_sfixed(-64071022.0/4294967296.0,1,-nbitq), 
to_sfixed(-351100192.0/4294967296.0,1,-nbitq), 
to_sfixed(-50263395.0/4294967296.0,1,-nbitq), 
to_sfixed(-381409505.0/4294967296.0,1,-nbitq), 
to_sfixed(334326323.0/4294967296.0,1,-nbitq), 
to_sfixed(477165157.0/4294967296.0,1,-nbitq), 
to_sfixed(-508248428.0/4294967296.0,1,-nbitq), 
to_sfixed(49100593.0/4294967296.0,1,-nbitq), 
to_sfixed(-186444544.0/4294967296.0,1,-nbitq), 
to_sfixed(217232618.0/4294967296.0,1,-nbitq), 
to_sfixed(454997626.0/4294967296.0,1,-nbitq), 
to_sfixed(-142569656.0/4294967296.0,1,-nbitq), 
to_sfixed(176312524.0/4294967296.0,1,-nbitq), 
to_sfixed(294608631.0/4294967296.0,1,-nbitq), 
to_sfixed(-380311904.0/4294967296.0,1,-nbitq), 
to_sfixed(-220393514.0/4294967296.0,1,-nbitq), 
to_sfixed(218942284.0/4294967296.0,1,-nbitq), 
to_sfixed(286938537.0/4294967296.0,1,-nbitq), 
to_sfixed(74885614.0/4294967296.0,1,-nbitq), 
to_sfixed(-166508421.0/4294967296.0,1,-nbitq), 
to_sfixed(-351387006.0/4294967296.0,1,-nbitq), 
to_sfixed(536003270.0/4294967296.0,1,-nbitq), 
to_sfixed(-32551959.0/4294967296.0,1,-nbitq), 
to_sfixed(152009690.0/4294967296.0,1,-nbitq), 
to_sfixed(307374042.0/4294967296.0,1,-nbitq), 
to_sfixed(75648774.0/4294967296.0,1,-nbitq), 
to_sfixed(-511194841.0/4294967296.0,1,-nbitq), 
to_sfixed(220460115.0/4294967296.0,1,-nbitq), 
to_sfixed(-322033497.0/4294967296.0,1,-nbitq), 
to_sfixed(104865487.0/4294967296.0,1,-nbitq), 
to_sfixed(-290906757.0/4294967296.0,1,-nbitq), 
to_sfixed(-17907005.0/4294967296.0,1,-nbitq), 
to_sfixed(22406606.0/4294967296.0,1,-nbitq), 
to_sfixed(-228462119.0/4294967296.0,1,-nbitq), 
to_sfixed(327057995.0/4294967296.0,1,-nbitq), 
to_sfixed(-32768954.0/4294967296.0,1,-nbitq), 
to_sfixed(-109109390.0/4294967296.0,1,-nbitq), 
to_sfixed(-61716876.0/4294967296.0,1,-nbitq), 
to_sfixed(180297087.0/4294967296.0,1,-nbitq), 
to_sfixed(143620910.0/4294967296.0,1,-nbitq), 
to_sfixed(111263216.0/4294967296.0,1,-nbitq), 
to_sfixed(66516756.0/4294967296.0,1,-nbitq), 
to_sfixed(201833565.0/4294967296.0,1,-nbitq), 
to_sfixed(-229467325.0/4294967296.0,1,-nbitq), 
to_sfixed(-287874469.0/4294967296.0,1,-nbitq), 
to_sfixed(-150090136.0/4294967296.0,1,-nbitq), 
to_sfixed(-188365590.0/4294967296.0,1,-nbitq), 
to_sfixed(37885312.0/4294967296.0,1,-nbitq), 
to_sfixed(-359112531.0/4294967296.0,1,-nbitq), 
to_sfixed(-70082805.0/4294967296.0,1,-nbitq), 
to_sfixed(50898782.0/4294967296.0,1,-nbitq), 
to_sfixed(-112902457.0/4294967296.0,1,-nbitq), 
to_sfixed(-614012742.0/4294967296.0,1,-nbitq), 
to_sfixed(-162730679.0/4294967296.0,1,-nbitq), 
to_sfixed(-427441973.0/4294967296.0,1,-nbitq), 
to_sfixed(-166157412.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(186561047.0/4294967296.0,1,-nbitq), 
to_sfixed(57655837.0/4294967296.0,1,-nbitq), 
to_sfixed(-111698453.0/4294967296.0,1,-nbitq), 
to_sfixed(162956095.0/4294967296.0,1,-nbitq), 
to_sfixed(-273431035.0/4294967296.0,1,-nbitq), 
to_sfixed(272221338.0/4294967296.0,1,-nbitq), 
to_sfixed(108985945.0/4294967296.0,1,-nbitq), 
to_sfixed(189849172.0/4294967296.0,1,-nbitq), 
to_sfixed(231678740.0/4294967296.0,1,-nbitq), 
to_sfixed(-233001482.0/4294967296.0,1,-nbitq), 
to_sfixed(75111915.0/4294967296.0,1,-nbitq), 
to_sfixed(522411586.0/4294967296.0,1,-nbitq), 
to_sfixed(-308328767.0/4294967296.0,1,-nbitq), 
to_sfixed(48266964.0/4294967296.0,1,-nbitq), 
to_sfixed(-415143464.0/4294967296.0,1,-nbitq), 
to_sfixed(-332957495.0/4294967296.0,1,-nbitq), 
to_sfixed(234125826.0/4294967296.0,1,-nbitq), 
to_sfixed(-216004978.0/4294967296.0,1,-nbitq), 
to_sfixed(-27188014.0/4294967296.0,1,-nbitq), 
to_sfixed(-331046747.0/4294967296.0,1,-nbitq), 
to_sfixed(-392318825.0/4294967296.0,1,-nbitq), 
to_sfixed(-34816831.0/4294967296.0,1,-nbitq), 
to_sfixed(283660256.0/4294967296.0,1,-nbitq), 
to_sfixed(-76678850.0/4294967296.0,1,-nbitq), 
to_sfixed(158911765.0/4294967296.0,1,-nbitq), 
to_sfixed(-446837080.0/4294967296.0,1,-nbitq), 
to_sfixed(183151006.0/4294967296.0,1,-nbitq), 
to_sfixed(-489441854.0/4294967296.0,1,-nbitq), 
to_sfixed(-54891294.0/4294967296.0,1,-nbitq), 
to_sfixed(368534468.0/4294967296.0,1,-nbitq), 
to_sfixed(-435016253.0/4294967296.0,1,-nbitq), 
to_sfixed(320288681.0/4294967296.0,1,-nbitq), 
to_sfixed(287407035.0/4294967296.0,1,-nbitq), 
to_sfixed(-244159507.0/4294967296.0,1,-nbitq), 
to_sfixed(230604029.0/4294967296.0,1,-nbitq), 
to_sfixed(-498197675.0/4294967296.0,1,-nbitq), 
to_sfixed(366013223.0/4294967296.0,1,-nbitq), 
to_sfixed(-211864342.0/4294967296.0,1,-nbitq), 
to_sfixed(-394420642.0/4294967296.0,1,-nbitq), 
to_sfixed(360800991.0/4294967296.0,1,-nbitq), 
to_sfixed(127416848.0/4294967296.0,1,-nbitq), 
to_sfixed(-133030343.0/4294967296.0,1,-nbitq), 
to_sfixed(381886389.0/4294967296.0,1,-nbitq), 
to_sfixed(-138171257.0/4294967296.0,1,-nbitq), 
to_sfixed(269905655.0/4294967296.0,1,-nbitq), 
to_sfixed(277483497.0/4294967296.0,1,-nbitq), 
to_sfixed(240994999.0/4294967296.0,1,-nbitq), 
to_sfixed(261206798.0/4294967296.0,1,-nbitq), 
to_sfixed(303015497.0/4294967296.0,1,-nbitq), 
to_sfixed(411830174.0/4294967296.0,1,-nbitq), 
to_sfixed(71554010.0/4294967296.0,1,-nbitq), 
to_sfixed(178766064.0/4294967296.0,1,-nbitq), 
to_sfixed(-86760518.0/4294967296.0,1,-nbitq), 
to_sfixed(94333445.0/4294967296.0,1,-nbitq), 
to_sfixed(-263323279.0/4294967296.0,1,-nbitq), 
to_sfixed(164076676.0/4294967296.0,1,-nbitq), 
to_sfixed(-90453170.0/4294967296.0,1,-nbitq), 
to_sfixed(185413942.0/4294967296.0,1,-nbitq), 
to_sfixed(224028719.0/4294967296.0,1,-nbitq), 
to_sfixed(422834609.0/4294967296.0,1,-nbitq), 
to_sfixed(-343838272.0/4294967296.0,1,-nbitq), 
to_sfixed(92644851.0/4294967296.0,1,-nbitq), 
to_sfixed(-39970214.0/4294967296.0,1,-nbitq), 
to_sfixed(-227667015.0/4294967296.0,1,-nbitq), 
to_sfixed(433545010.0/4294967296.0,1,-nbitq), 
to_sfixed(240357836.0/4294967296.0,1,-nbitq), 
to_sfixed(805756335.0/4294967296.0,1,-nbitq), 
to_sfixed(-124882072.0/4294967296.0,1,-nbitq), 
to_sfixed(430877458.0/4294967296.0,1,-nbitq), 
to_sfixed(-266649525.0/4294967296.0,1,-nbitq), 
to_sfixed(142541247.0/4294967296.0,1,-nbitq), 
to_sfixed(394037875.0/4294967296.0,1,-nbitq), 
to_sfixed(-247940246.0/4294967296.0,1,-nbitq), 
to_sfixed(379300569.0/4294967296.0,1,-nbitq), 
to_sfixed(-162034401.0/4294967296.0,1,-nbitq), 
to_sfixed(-369317579.0/4294967296.0,1,-nbitq), 
to_sfixed(-614546085.0/4294967296.0,1,-nbitq), 
to_sfixed(152207410.0/4294967296.0,1,-nbitq), 
to_sfixed(-353816195.0/4294967296.0,1,-nbitq), 
to_sfixed(351597119.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(171945588.0/4294967296.0,1,-nbitq), 
to_sfixed(188384907.0/4294967296.0,1,-nbitq), 
to_sfixed(251918797.0/4294967296.0,1,-nbitq), 
to_sfixed(-412626990.0/4294967296.0,1,-nbitq), 
to_sfixed(-133549667.0/4294967296.0,1,-nbitq), 
to_sfixed(-71073874.0/4294967296.0,1,-nbitq), 
to_sfixed(-192623761.0/4294967296.0,1,-nbitq), 
to_sfixed(151548773.0/4294967296.0,1,-nbitq), 
to_sfixed(237845026.0/4294967296.0,1,-nbitq), 
to_sfixed(-201563345.0/4294967296.0,1,-nbitq), 
to_sfixed(360641668.0/4294967296.0,1,-nbitq), 
to_sfixed(-8405850.0/4294967296.0,1,-nbitq), 
to_sfixed(-323484524.0/4294967296.0,1,-nbitq), 
to_sfixed(380271273.0/4294967296.0,1,-nbitq), 
to_sfixed(122895200.0/4294967296.0,1,-nbitq), 
to_sfixed(-514621735.0/4294967296.0,1,-nbitq), 
to_sfixed(286048032.0/4294967296.0,1,-nbitq), 
to_sfixed(-80408641.0/4294967296.0,1,-nbitq), 
to_sfixed(65566349.0/4294967296.0,1,-nbitq), 
to_sfixed(-131162048.0/4294967296.0,1,-nbitq), 
to_sfixed(130484752.0/4294967296.0,1,-nbitq), 
to_sfixed(142653363.0/4294967296.0,1,-nbitq), 
to_sfixed(307653931.0/4294967296.0,1,-nbitq), 
to_sfixed(150319319.0/4294967296.0,1,-nbitq), 
to_sfixed(31159885.0/4294967296.0,1,-nbitq), 
to_sfixed(-31902444.0/4294967296.0,1,-nbitq), 
to_sfixed(-311647947.0/4294967296.0,1,-nbitq), 
to_sfixed(-176832553.0/4294967296.0,1,-nbitq), 
to_sfixed(-75855229.0/4294967296.0,1,-nbitq), 
to_sfixed(289355947.0/4294967296.0,1,-nbitq), 
to_sfixed(-494191126.0/4294967296.0,1,-nbitq), 
to_sfixed(259608256.0/4294967296.0,1,-nbitq), 
to_sfixed(143122502.0/4294967296.0,1,-nbitq), 
to_sfixed(71201756.0/4294967296.0,1,-nbitq), 
to_sfixed(-237616723.0/4294967296.0,1,-nbitq), 
to_sfixed(-234163369.0/4294967296.0,1,-nbitq), 
to_sfixed(284152177.0/4294967296.0,1,-nbitq), 
to_sfixed(187568900.0/4294967296.0,1,-nbitq), 
to_sfixed(-200726730.0/4294967296.0,1,-nbitq), 
to_sfixed(408757943.0/4294967296.0,1,-nbitq), 
to_sfixed(366330110.0/4294967296.0,1,-nbitq), 
to_sfixed(-260496717.0/4294967296.0,1,-nbitq), 
to_sfixed(-331619993.0/4294967296.0,1,-nbitq), 
to_sfixed(-95839380.0/4294967296.0,1,-nbitq), 
to_sfixed(-457622378.0/4294967296.0,1,-nbitq), 
to_sfixed(-108452697.0/4294967296.0,1,-nbitq), 
to_sfixed(45452572.0/4294967296.0,1,-nbitq), 
to_sfixed(304243879.0/4294967296.0,1,-nbitq), 
to_sfixed(408211760.0/4294967296.0,1,-nbitq), 
to_sfixed(167061327.0/4294967296.0,1,-nbitq), 
to_sfixed(-459895194.0/4294967296.0,1,-nbitq), 
to_sfixed(-77434381.0/4294967296.0,1,-nbitq), 
to_sfixed(-142638291.0/4294967296.0,1,-nbitq), 
to_sfixed(-120831399.0/4294967296.0,1,-nbitq), 
to_sfixed(74745597.0/4294967296.0,1,-nbitq), 
to_sfixed(-257919069.0/4294967296.0,1,-nbitq), 
to_sfixed(-234510245.0/4294967296.0,1,-nbitq), 
to_sfixed(-8159691.0/4294967296.0,1,-nbitq), 
to_sfixed(-185591518.0/4294967296.0,1,-nbitq), 
to_sfixed(139206278.0/4294967296.0,1,-nbitq), 
to_sfixed(-356923490.0/4294967296.0,1,-nbitq), 
to_sfixed(29987302.0/4294967296.0,1,-nbitq), 
to_sfixed(205553820.0/4294967296.0,1,-nbitq), 
to_sfixed(341044189.0/4294967296.0,1,-nbitq), 
to_sfixed(349107822.0/4294967296.0,1,-nbitq), 
to_sfixed(-409795228.0/4294967296.0,1,-nbitq), 
to_sfixed(666369544.0/4294967296.0,1,-nbitq), 
to_sfixed(-389147727.0/4294967296.0,1,-nbitq), 
to_sfixed(-49864004.0/4294967296.0,1,-nbitq), 
to_sfixed(-186043700.0/4294967296.0,1,-nbitq), 
to_sfixed(-308460890.0/4294967296.0,1,-nbitq), 
to_sfixed(169880851.0/4294967296.0,1,-nbitq), 
to_sfixed(170587898.0/4294967296.0,1,-nbitq), 
to_sfixed(338591497.0/4294967296.0,1,-nbitq), 
to_sfixed(-195758805.0/4294967296.0,1,-nbitq), 
to_sfixed(-219137735.0/4294967296.0,1,-nbitq), 
to_sfixed(-622353821.0/4294967296.0,1,-nbitq), 
to_sfixed(-500024773.0/4294967296.0,1,-nbitq), 
to_sfixed(-558500024.0/4294967296.0,1,-nbitq), 
to_sfixed(-95938374.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(22970473.0/4294967296.0,1,-nbitq), 
to_sfixed(-57734670.0/4294967296.0,1,-nbitq), 
to_sfixed(316553012.0/4294967296.0,1,-nbitq), 
to_sfixed(-387012613.0/4294967296.0,1,-nbitq), 
to_sfixed(286934665.0/4294967296.0,1,-nbitq), 
to_sfixed(174225876.0/4294967296.0,1,-nbitq), 
to_sfixed(-204859307.0/4294967296.0,1,-nbitq), 
to_sfixed(285302677.0/4294967296.0,1,-nbitq), 
to_sfixed(-152872322.0/4294967296.0,1,-nbitq), 
to_sfixed(138365437.0/4294967296.0,1,-nbitq), 
to_sfixed(310726298.0/4294967296.0,1,-nbitq), 
to_sfixed(270336482.0/4294967296.0,1,-nbitq), 
to_sfixed(-313056328.0/4294967296.0,1,-nbitq), 
to_sfixed(38474946.0/4294967296.0,1,-nbitq), 
to_sfixed(-44299321.0/4294967296.0,1,-nbitq), 
to_sfixed(-309090780.0/4294967296.0,1,-nbitq), 
to_sfixed(258797693.0/4294967296.0,1,-nbitq), 
to_sfixed(-63690741.0/4294967296.0,1,-nbitq), 
to_sfixed(205993441.0/4294967296.0,1,-nbitq), 
to_sfixed(-142621392.0/4294967296.0,1,-nbitq), 
to_sfixed(143519218.0/4294967296.0,1,-nbitq), 
to_sfixed(205971767.0/4294967296.0,1,-nbitq), 
to_sfixed(274962763.0/4294967296.0,1,-nbitq), 
to_sfixed(-145221420.0/4294967296.0,1,-nbitq), 
to_sfixed(115313137.0/4294967296.0,1,-nbitq), 
to_sfixed(214610836.0/4294967296.0,1,-nbitq), 
to_sfixed(-7620647.0/4294967296.0,1,-nbitq), 
to_sfixed(-221679726.0/4294967296.0,1,-nbitq), 
to_sfixed(393848100.0/4294967296.0,1,-nbitq), 
to_sfixed(493907187.0/4294967296.0,1,-nbitq), 
to_sfixed(-120300598.0/4294967296.0,1,-nbitq), 
to_sfixed(293856316.0/4294967296.0,1,-nbitq), 
to_sfixed(445712236.0/4294967296.0,1,-nbitq), 
to_sfixed(-319815731.0/4294967296.0,1,-nbitq), 
to_sfixed(323760260.0/4294967296.0,1,-nbitq), 
to_sfixed(257437071.0/4294967296.0,1,-nbitq), 
to_sfixed(46676954.0/4294967296.0,1,-nbitq), 
to_sfixed(91158596.0/4294967296.0,1,-nbitq), 
to_sfixed(-77773011.0/4294967296.0,1,-nbitq), 
to_sfixed(352827365.0/4294967296.0,1,-nbitq), 
to_sfixed(-13767797.0/4294967296.0,1,-nbitq), 
to_sfixed(-303956021.0/4294967296.0,1,-nbitq), 
to_sfixed(-113563481.0/4294967296.0,1,-nbitq), 
to_sfixed(-93698327.0/4294967296.0,1,-nbitq), 
to_sfixed(77245531.0/4294967296.0,1,-nbitq), 
to_sfixed(67723244.0/4294967296.0,1,-nbitq), 
to_sfixed(151696080.0/4294967296.0,1,-nbitq), 
to_sfixed(87697270.0/4294967296.0,1,-nbitq), 
to_sfixed(37459711.0/4294967296.0,1,-nbitq), 
to_sfixed(-21239321.0/4294967296.0,1,-nbitq), 
to_sfixed(-389487638.0/4294967296.0,1,-nbitq), 
to_sfixed(-68930157.0/4294967296.0,1,-nbitq), 
to_sfixed(-137105369.0/4294967296.0,1,-nbitq), 
to_sfixed(352689448.0/4294967296.0,1,-nbitq), 
to_sfixed(515481964.0/4294967296.0,1,-nbitq), 
to_sfixed(93644805.0/4294967296.0,1,-nbitq), 
to_sfixed(-332050065.0/4294967296.0,1,-nbitq), 
to_sfixed(221125060.0/4294967296.0,1,-nbitq), 
to_sfixed(323048576.0/4294967296.0,1,-nbitq), 
to_sfixed(346804769.0/4294967296.0,1,-nbitq), 
to_sfixed(326424351.0/4294967296.0,1,-nbitq), 
to_sfixed(163932827.0/4294967296.0,1,-nbitq), 
to_sfixed(171540371.0/4294967296.0,1,-nbitq), 
to_sfixed(113627211.0/4294967296.0,1,-nbitq), 
to_sfixed(186075809.0/4294967296.0,1,-nbitq), 
to_sfixed(-144220205.0/4294967296.0,1,-nbitq), 
to_sfixed(216684192.0/4294967296.0,1,-nbitq), 
to_sfixed(-103748980.0/4294967296.0,1,-nbitq), 
to_sfixed(-143126891.0/4294967296.0,1,-nbitq), 
to_sfixed(-477320426.0/4294967296.0,1,-nbitq), 
to_sfixed(-160795427.0/4294967296.0,1,-nbitq), 
to_sfixed(170687836.0/4294967296.0,1,-nbitq), 
to_sfixed(-235237395.0/4294967296.0,1,-nbitq), 
to_sfixed(-288561389.0/4294967296.0,1,-nbitq), 
to_sfixed(381228957.0/4294967296.0,1,-nbitq), 
to_sfixed(16927469.0/4294967296.0,1,-nbitq), 
to_sfixed(-537233725.0/4294967296.0,1,-nbitq), 
to_sfixed(-346026206.0/4294967296.0,1,-nbitq), 
to_sfixed(131598822.0/4294967296.0,1,-nbitq), 
to_sfixed(20066639.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-148777823.0/4294967296.0,1,-nbitq), 
to_sfixed(69318341.0/4294967296.0,1,-nbitq), 
to_sfixed(-386833226.0/4294967296.0,1,-nbitq), 
to_sfixed(90114555.0/4294967296.0,1,-nbitq), 
to_sfixed(-46010001.0/4294967296.0,1,-nbitq), 
to_sfixed(-141603.0/4294967296.0,1,-nbitq), 
to_sfixed(347496476.0/4294967296.0,1,-nbitq), 
to_sfixed(204315828.0/4294967296.0,1,-nbitq), 
to_sfixed(331093343.0/4294967296.0,1,-nbitq), 
to_sfixed(158290267.0/4294967296.0,1,-nbitq), 
to_sfixed(168465346.0/4294967296.0,1,-nbitq), 
to_sfixed(43411297.0/4294967296.0,1,-nbitq), 
to_sfixed(-724848954.0/4294967296.0,1,-nbitq), 
to_sfixed(647050385.0/4294967296.0,1,-nbitq), 
to_sfixed(225210243.0/4294967296.0,1,-nbitq), 
to_sfixed(149459760.0/4294967296.0,1,-nbitq), 
to_sfixed(46906285.0/4294967296.0,1,-nbitq), 
to_sfixed(412379402.0/4294967296.0,1,-nbitq), 
to_sfixed(8525522.0/4294967296.0,1,-nbitq), 
to_sfixed(-172255413.0/4294967296.0,1,-nbitq), 
to_sfixed(149894866.0/4294967296.0,1,-nbitq), 
to_sfixed(351126026.0/4294967296.0,1,-nbitq), 
to_sfixed(56192947.0/4294967296.0,1,-nbitq), 
to_sfixed(304133608.0/4294967296.0,1,-nbitq), 
to_sfixed(-46777910.0/4294967296.0,1,-nbitq), 
to_sfixed(232296627.0/4294967296.0,1,-nbitq), 
to_sfixed(149287559.0/4294967296.0,1,-nbitq), 
to_sfixed(21290854.0/4294967296.0,1,-nbitq), 
to_sfixed(546412059.0/4294967296.0,1,-nbitq), 
to_sfixed(24328810.0/4294967296.0,1,-nbitq), 
to_sfixed(-27206311.0/4294967296.0,1,-nbitq), 
to_sfixed(-13724982.0/4294967296.0,1,-nbitq), 
to_sfixed(373991721.0/4294967296.0,1,-nbitq), 
to_sfixed(-269416828.0/4294967296.0,1,-nbitq), 
to_sfixed(399774063.0/4294967296.0,1,-nbitq), 
to_sfixed(51180587.0/4294967296.0,1,-nbitq), 
to_sfixed(204609944.0/4294967296.0,1,-nbitq), 
to_sfixed(160986867.0/4294967296.0,1,-nbitq), 
to_sfixed(274685547.0/4294967296.0,1,-nbitq), 
to_sfixed(316016749.0/4294967296.0,1,-nbitq), 
to_sfixed(165447508.0/4294967296.0,1,-nbitq), 
to_sfixed(-189743941.0/4294967296.0,1,-nbitq), 
to_sfixed(193705638.0/4294967296.0,1,-nbitq), 
to_sfixed(95060323.0/4294967296.0,1,-nbitq), 
to_sfixed(259771452.0/4294967296.0,1,-nbitq), 
to_sfixed(28563098.0/4294967296.0,1,-nbitq), 
to_sfixed(-135514789.0/4294967296.0,1,-nbitq), 
to_sfixed(-38569324.0/4294967296.0,1,-nbitq), 
to_sfixed(363247158.0/4294967296.0,1,-nbitq), 
to_sfixed(-162742207.0/4294967296.0,1,-nbitq), 
to_sfixed(-31993968.0/4294967296.0,1,-nbitq), 
to_sfixed(21515236.0/4294967296.0,1,-nbitq), 
to_sfixed(-312521710.0/4294967296.0,1,-nbitq), 
to_sfixed(-44276624.0/4294967296.0,1,-nbitq), 
to_sfixed(-133192816.0/4294967296.0,1,-nbitq), 
to_sfixed(-105785400.0/4294967296.0,1,-nbitq), 
to_sfixed(344283444.0/4294967296.0,1,-nbitq), 
to_sfixed(-255396814.0/4294967296.0,1,-nbitq), 
to_sfixed(-250189366.0/4294967296.0,1,-nbitq), 
to_sfixed(255672610.0/4294967296.0,1,-nbitq), 
to_sfixed(-312914882.0/4294967296.0,1,-nbitq), 
to_sfixed(-159150753.0/4294967296.0,1,-nbitq), 
to_sfixed(-92638991.0/4294967296.0,1,-nbitq), 
to_sfixed(-320522973.0/4294967296.0,1,-nbitq), 
to_sfixed(109654628.0/4294967296.0,1,-nbitq), 
to_sfixed(52499464.0/4294967296.0,1,-nbitq), 
to_sfixed(569220984.0/4294967296.0,1,-nbitq), 
to_sfixed(-316283027.0/4294967296.0,1,-nbitq), 
to_sfixed(-200894714.0/4294967296.0,1,-nbitq), 
to_sfixed(251714775.0/4294967296.0,1,-nbitq), 
to_sfixed(19584489.0/4294967296.0,1,-nbitq), 
to_sfixed(128553955.0/4294967296.0,1,-nbitq), 
to_sfixed(115132.0/4294967296.0,1,-nbitq), 
to_sfixed(415936909.0/4294967296.0,1,-nbitq), 
to_sfixed(-125896600.0/4294967296.0,1,-nbitq), 
to_sfixed(-491683434.0/4294967296.0,1,-nbitq), 
to_sfixed(-189842291.0/4294967296.0,1,-nbitq), 
to_sfixed(-536582575.0/4294967296.0,1,-nbitq), 
to_sfixed(-513579502.0/4294967296.0,1,-nbitq), 
to_sfixed(-38442819.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(542130235.0/4294967296.0,1,-nbitq), 
to_sfixed(-105238909.0/4294967296.0,1,-nbitq), 
to_sfixed(373425198.0/4294967296.0,1,-nbitq), 
to_sfixed(-20250883.0/4294967296.0,1,-nbitq), 
to_sfixed(-44354825.0/4294967296.0,1,-nbitq), 
to_sfixed(250002062.0/4294967296.0,1,-nbitq), 
to_sfixed(39519274.0/4294967296.0,1,-nbitq), 
to_sfixed(-227725648.0/4294967296.0,1,-nbitq), 
to_sfixed(-26803315.0/4294967296.0,1,-nbitq), 
to_sfixed(-66132883.0/4294967296.0,1,-nbitq), 
to_sfixed(140259051.0/4294967296.0,1,-nbitq), 
to_sfixed(83464006.0/4294967296.0,1,-nbitq), 
to_sfixed(-561678556.0/4294967296.0,1,-nbitq), 
to_sfixed(76064397.0/4294967296.0,1,-nbitq), 
to_sfixed(-247994528.0/4294967296.0,1,-nbitq), 
to_sfixed(265626405.0/4294967296.0,1,-nbitq), 
to_sfixed(368996311.0/4294967296.0,1,-nbitq), 
to_sfixed(126805106.0/4294967296.0,1,-nbitq), 
to_sfixed(-348907599.0/4294967296.0,1,-nbitq), 
to_sfixed(-243700073.0/4294967296.0,1,-nbitq), 
to_sfixed(782158.0/4294967296.0,1,-nbitq), 
to_sfixed(47609013.0/4294967296.0,1,-nbitq), 
to_sfixed(-94397698.0/4294967296.0,1,-nbitq), 
to_sfixed(154581086.0/4294967296.0,1,-nbitq), 
to_sfixed(-33297247.0/4294967296.0,1,-nbitq), 
to_sfixed(158189586.0/4294967296.0,1,-nbitq), 
to_sfixed(-204271914.0/4294967296.0,1,-nbitq), 
to_sfixed(-397272846.0/4294967296.0,1,-nbitq), 
to_sfixed(166214066.0/4294967296.0,1,-nbitq), 
to_sfixed(408662950.0/4294967296.0,1,-nbitq), 
to_sfixed(-482465535.0/4294967296.0,1,-nbitq), 
to_sfixed(262683664.0/4294967296.0,1,-nbitq), 
to_sfixed(288944356.0/4294967296.0,1,-nbitq), 
to_sfixed(-515618612.0/4294967296.0,1,-nbitq), 
to_sfixed(-20805384.0/4294967296.0,1,-nbitq), 
to_sfixed(185280878.0/4294967296.0,1,-nbitq), 
to_sfixed(-40246967.0/4294967296.0,1,-nbitq), 
to_sfixed(-290615870.0/4294967296.0,1,-nbitq), 
to_sfixed(-332054512.0/4294967296.0,1,-nbitq), 
to_sfixed(83428179.0/4294967296.0,1,-nbitq), 
to_sfixed(186471680.0/4294967296.0,1,-nbitq), 
to_sfixed(400262022.0/4294967296.0,1,-nbitq), 
to_sfixed(-354032221.0/4294967296.0,1,-nbitq), 
to_sfixed(443620704.0/4294967296.0,1,-nbitq), 
to_sfixed(-10330260.0/4294967296.0,1,-nbitq), 
to_sfixed(111725937.0/4294967296.0,1,-nbitq), 
to_sfixed(-310104362.0/4294967296.0,1,-nbitq), 
to_sfixed(-294704929.0/4294967296.0,1,-nbitq), 
to_sfixed(-375296406.0/4294967296.0,1,-nbitq), 
to_sfixed(-263919964.0/4294967296.0,1,-nbitq), 
to_sfixed(-671491203.0/4294967296.0,1,-nbitq), 
to_sfixed(-207416889.0/4294967296.0,1,-nbitq), 
to_sfixed(-653189016.0/4294967296.0,1,-nbitq), 
to_sfixed(270936067.0/4294967296.0,1,-nbitq), 
to_sfixed(420029708.0/4294967296.0,1,-nbitq), 
to_sfixed(324754088.0/4294967296.0,1,-nbitq), 
to_sfixed(166179162.0/4294967296.0,1,-nbitq), 
to_sfixed(120673945.0/4294967296.0,1,-nbitq), 
to_sfixed(220884142.0/4294967296.0,1,-nbitq), 
to_sfixed(-267304081.0/4294967296.0,1,-nbitq), 
to_sfixed(-313305793.0/4294967296.0,1,-nbitq), 
to_sfixed(347249138.0/4294967296.0,1,-nbitq), 
to_sfixed(-281509076.0/4294967296.0,1,-nbitq), 
to_sfixed(-281211069.0/4294967296.0,1,-nbitq), 
to_sfixed(-176486720.0/4294967296.0,1,-nbitq), 
to_sfixed(-426437867.0/4294967296.0,1,-nbitq), 
to_sfixed(797350303.0/4294967296.0,1,-nbitq), 
to_sfixed(-447765188.0/4294967296.0,1,-nbitq), 
to_sfixed(176137144.0/4294967296.0,1,-nbitq), 
to_sfixed(-24788414.0/4294967296.0,1,-nbitq), 
to_sfixed(-80192781.0/4294967296.0,1,-nbitq), 
to_sfixed(-170033462.0/4294967296.0,1,-nbitq), 
to_sfixed(-551109292.0/4294967296.0,1,-nbitq), 
to_sfixed(-253454720.0/4294967296.0,1,-nbitq), 
to_sfixed(-90918782.0/4294967296.0,1,-nbitq), 
to_sfixed(-471758103.0/4294967296.0,1,-nbitq), 
to_sfixed(-397120693.0/4294967296.0,1,-nbitq), 
to_sfixed(94282604.0/4294967296.0,1,-nbitq), 
to_sfixed(-29150455.0/4294967296.0,1,-nbitq), 
to_sfixed(73765319.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(17540848.0/4294967296.0,1,-nbitq), 
to_sfixed(-82647659.0/4294967296.0,1,-nbitq), 
to_sfixed(-43459499.0/4294967296.0,1,-nbitq), 
to_sfixed(402708434.0/4294967296.0,1,-nbitq), 
to_sfixed(85368102.0/4294967296.0,1,-nbitq), 
to_sfixed(-187269485.0/4294967296.0,1,-nbitq), 
to_sfixed(-164977036.0/4294967296.0,1,-nbitq), 
to_sfixed(106846051.0/4294967296.0,1,-nbitq), 
to_sfixed(54445008.0/4294967296.0,1,-nbitq), 
to_sfixed(-313419610.0/4294967296.0,1,-nbitq), 
to_sfixed(-166926612.0/4294967296.0,1,-nbitq), 
to_sfixed(395504499.0/4294967296.0,1,-nbitq), 
to_sfixed(-310228186.0/4294967296.0,1,-nbitq), 
to_sfixed(194428318.0/4294967296.0,1,-nbitq), 
to_sfixed(25189759.0/4294967296.0,1,-nbitq), 
to_sfixed(-378194614.0/4294967296.0,1,-nbitq), 
to_sfixed(121545783.0/4294967296.0,1,-nbitq), 
to_sfixed(-244542217.0/4294967296.0,1,-nbitq), 
to_sfixed(-401946149.0/4294967296.0,1,-nbitq), 
to_sfixed(317824559.0/4294967296.0,1,-nbitq), 
to_sfixed(-291282383.0/4294967296.0,1,-nbitq), 
to_sfixed(-100345914.0/4294967296.0,1,-nbitq), 
to_sfixed(-76608197.0/4294967296.0,1,-nbitq), 
to_sfixed(217104339.0/4294967296.0,1,-nbitq), 
to_sfixed(353821154.0/4294967296.0,1,-nbitq), 
to_sfixed(-346524787.0/4294967296.0,1,-nbitq), 
to_sfixed(-374674385.0/4294967296.0,1,-nbitq), 
to_sfixed(-545731026.0/4294967296.0,1,-nbitq), 
to_sfixed(481189254.0/4294967296.0,1,-nbitq), 
to_sfixed(226940519.0/4294967296.0,1,-nbitq), 
to_sfixed(-311911268.0/4294967296.0,1,-nbitq), 
to_sfixed(-26533237.0/4294967296.0,1,-nbitq), 
to_sfixed(-282619983.0/4294967296.0,1,-nbitq), 
to_sfixed(-174482688.0/4294967296.0,1,-nbitq), 
to_sfixed(195636839.0/4294967296.0,1,-nbitq), 
to_sfixed(351615681.0/4294967296.0,1,-nbitq), 
to_sfixed(289199408.0/4294967296.0,1,-nbitq), 
to_sfixed(-316926904.0/4294967296.0,1,-nbitq), 
to_sfixed(99838139.0/4294967296.0,1,-nbitq), 
to_sfixed(262257980.0/4294967296.0,1,-nbitq), 
to_sfixed(-166240704.0/4294967296.0,1,-nbitq), 
to_sfixed(180723186.0/4294967296.0,1,-nbitq), 
to_sfixed(-232099269.0/4294967296.0,1,-nbitq), 
to_sfixed(-1893802.0/4294967296.0,1,-nbitq), 
to_sfixed(85896900.0/4294967296.0,1,-nbitq), 
to_sfixed(219499802.0/4294967296.0,1,-nbitq), 
to_sfixed(-260520155.0/4294967296.0,1,-nbitq), 
to_sfixed(189597554.0/4294967296.0,1,-nbitq), 
to_sfixed(290946584.0/4294967296.0,1,-nbitq), 
to_sfixed(-201061362.0/4294967296.0,1,-nbitq), 
to_sfixed(-73930816.0/4294967296.0,1,-nbitq), 
to_sfixed(40939136.0/4294967296.0,1,-nbitq), 
to_sfixed(-119160962.0/4294967296.0,1,-nbitq), 
to_sfixed(351037547.0/4294967296.0,1,-nbitq), 
to_sfixed(382045509.0/4294967296.0,1,-nbitq), 
to_sfixed(88226787.0/4294967296.0,1,-nbitq), 
to_sfixed(205306242.0/4294967296.0,1,-nbitq), 
to_sfixed(21843100.0/4294967296.0,1,-nbitq), 
to_sfixed(-335253707.0/4294967296.0,1,-nbitq), 
to_sfixed(-226528257.0/4294967296.0,1,-nbitq), 
to_sfixed(50442284.0/4294967296.0,1,-nbitq), 
to_sfixed(131178180.0/4294967296.0,1,-nbitq), 
to_sfixed(162570077.0/4294967296.0,1,-nbitq), 
to_sfixed(-209726345.0/4294967296.0,1,-nbitq), 
to_sfixed(317185014.0/4294967296.0,1,-nbitq), 
to_sfixed(-184166149.0/4294967296.0,1,-nbitq), 
to_sfixed(140836138.0/4294967296.0,1,-nbitq), 
to_sfixed(299514683.0/4294967296.0,1,-nbitq), 
to_sfixed(-317171904.0/4294967296.0,1,-nbitq), 
to_sfixed(-183577536.0/4294967296.0,1,-nbitq), 
to_sfixed(-264558708.0/4294967296.0,1,-nbitq), 
to_sfixed(374546972.0/4294967296.0,1,-nbitq), 
to_sfixed(213221559.0/4294967296.0,1,-nbitq), 
to_sfixed(-110892134.0/4294967296.0,1,-nbitq), 
to_sfixed(501861347.0/4294967296.0,1,-nbitq), 
to_sfixed(79710551.0/4294967296.0,1,-nbitq), 
to_sfixed(8593855.0/4294967296.0,1,-nbitq), 
to_sfixed(-263798529.0/4294967296.0,1,-nbitq), 
to_sfixed(-150378817.0/4294967296.0,1,-nbitq), 
to_sfixed(-108579418.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(15890818.0/4294967296.0,1,-nbitq), 
to_sfixed(-187300442.0/4294967296.0,1,-nbitq), 
to_sfixed(-267403718.0/4294967296.0,1,-nbitq), 
to_sfixed(-327486273.0/4294967296.0,1,-nbitq), 
to_sfixed(283852052.0/4294967296.0,1,-nbitq), 
to_sfixed(-177853545.0/4294967296.0,1,-nbitq), 
to_sfixed(-271044138.0/4294967296.0,1,-nbitq), 
to_sfixed(85981899.0/4294967296.0,1,-nbitq), 
to_sfixed(-253494439.0/4294967296.0,1,-nbitq), 
to_sfixed(-223716758.0/4294967296.0,1,-nbitq), 
to_sfixed(-62476361.0/4294967296.0,1,-nbitq), 
to_sfixed(538244525.0/4294967296.0,1,-nbitq), 
to_sfixed(31750280.0/4294967296.0,1,-nbitq), 
to_sfixed(-84494239.0/4294967296.0,1,-nbitq), 
to_sfixed(12155345.0/4294967296.0,1,-nbitq), 
to_sfixed(169054889.0/4294967296.0,1,-nbitq), 
to_sfixed(-100810013.0/4294967296.0,1,-nbitq), 
to_sfixed(-314304153.0/4294967296.0,1,-nbitq), 
to_sfixed(245172029.0/4294967296.0,1,-nbitq), 
to_sfixed(-429937915.0/4294967296.0,1,-nbitq), 
to_sfixed(192121289.0/4294967296.0,1,-nbitq), 
to_sfixed(202695818.0/4294967296.0,1,-nbitq), 
to_sfixed(304151256.0/4294967296.0,1,-nbitq), 
to_sfixed(-333369899.0/4294967296.0,1,-nbitq), 
to_sfixed(356194463.0/4294967296.0,1,-nbitq), 
to_sfixed(404286866.0/4294967296.0,1,-nbitq), 
to_sfixed(212289018.0/4294967296.0,1,-nbitq), 
to_sfixed(94989643.0/4294967296.0,1,-nbitq), 
to_sfixed(299647610.0/4294967296.0,1,-nbitq), 
to_sfixed(-26519925.0/4294967296.0,1,-nbitq), 
to_sfixed(-403434965.0/4294967296.0,1,-nbitq), 
to_sfixed(-205714782.0/4294967296.0,1,-nbitq), 
to_sfixed(295529201.0/4294967296.0,1,-nbitq), 
to_sfixed(191336518.0/4294967296.0,1,-nbitq), 
to_sfixed(177135717.0/4294967296.0,1,-nbitq), 
to_sfixed(-37151970.0/4294967296.0,1,-nbitq), 
to_sfixed(-147302785.0/4294967296.0,1,-nbitq), 
to_sfixed(156538408.0/4294967296.0,1,-nbitq), 
to_sfixed(-383686963.0/4294967296.0,1,-nbitq), 
to_sfixed(-278408420.0/4294967296.0,1,-nbitq), 
to_sfixed(148355292.0/4294967296.0,1,-nbitq), 
to_sfixed(526842084.0/4294967296.0,1,-nbitq), 
to_sfixed(-230291947.0/4294967296.0,1,-nbitq), 
to_sfixed(-287406528.0/4294967296.0,1,-nbitq), 
to_sfixed(-359476129.0/4294967296.0,1,-nbitq), 
to_sfixed(-96304175.0/4294967296.0,1,-nbitq), 
to_sfixed(49848025.0/4294967296.0,1,-nbitq), 
to_sfixed(-123489889.0/4294967296.0,1,-nbitq), 
to_sfixed(-129850308.0/4294967296.0,1,-nbitq), 
to_sfixed(-223774147.0/4294967296.0,1,-nbitq), 
to_sfixed(-204169907.0/4294967296.0,1,-nbitq), 
to_sfixed(444236154.0/4294967296.0,1,-nbitq), 
to_sfixed(66998576.0/4294967296.0,1,-nbitq), 
to_sfixed(-234214890.0/4294967296.0,1,-nbitq), 
to_sfixed(-212694432.0/4294967296.0,1,-nbitq), 
to_sfixed(-232559049.0/4294967296.0,1,-nbitq), 
to_sfixed(-81050713.0/4294967296.0,1,-nbitq), 
to_sfixed(-18850527.0/4294967296.0,1,-nbitq), 
to_sfixed(152246053.0/4294967296.0,1,-nbitq), 
to_sfixed(-96992248.0/4294967296.0,1,-nbitq), 
to_sfixed(110724150.0/4294967296.0,1,-nbitq), 
to_sfixed(-179606449.0/4294967296.0,1,-nbitq), 
to_sfixed(-205662697.0/4294967296.0,1,-nbitq), 
to_sfixed(-193929189.0/4294967296.0,1,-nbitq), 
to_sfixed(235370080.0/4294967296.0,1,-nbitq), 
to_sfixed(-275018185.0/4294967296.0,1,-nbitq), 
to_sfixed(443512103.0/4294967296.0,1,-nbitq), 
to_sfixed(-258741161.0/4294967296.0,1,-nbitq), 
to_sfixed(385653917.0/4294967296.0,1,-nbitq), 
to_sfixed(645438313.0/4294967296.0,1,-nbitq), 
to_sfixed(-247755507.0/4294967296.0,1,-nbitq), 
to_sfixed(251562459.0/4294967296.0,1,-nbitq), 
to_sfixed(-536028184.0/4294967296.0,1,-nbitq), 
to_sfixed(-99516036.0/4294967296.0,1,-nbitq), 
to_sfixed(98609021.0/4294967296.0,1,-nbitq), 
to_sfixed(-172479910.0/4294967296.0,1,-nbitq), 
to_sfixed(-24115463.0/4294967296.0,1,-nbitq), 
to_sfixed(136459828.0/4294967296.0,1,-nbitq), 
to_sfixed(7865030.0/4294967296.0,1,-nbitq), 
to_sfixed(-24833518.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(360200712.0/4294967296.0,1,-nbitq), 
to_sfixed(52340407.0/4294967296.0,1,-nbitq), 
to_sfixed(-44003275.0/4294967296.0,1,-nbitq), 
to_sfixed(265740972.0/4294967296.0,1,-nbitq), 
to_sfixed(365025027.0/4294967296.0,1,-nbitq), 
to_sfixed(-230517821.0/4294967296.0,1,-nbitq), 
to_sfixed(129025319.0/4294967296.0,1,-nbitq), 
to_sfixed(-163665916.0/4294967296.0,1,-nbitq), 
to_sfixed(112936833.0/4294967296.0,1,-nbitq), 
to_sfixed(93524780.0/4294967296.0,1,-nbitq), 
to_sfixed(-279945566.0/4294967296.0,1,-nbitq), 
to_sfixed(-44128299.0/4294967296.0,1,-nbitq), 
to_sfixed(106728821.0/4294967296.0,1,-nbitq), 
to_sfixed(-223048438.0/4294967296.0,1,-nbitq), 
to_sfixed(-155579305.0/4294967296.0,1,-nbitq), 
to_sfixed(-344967990.0/4294967296.0,1,-nbitq), 
to_sfixed(22956589.0/4294967296.0,1,-nbitq), 
to_sfixed(-293673163.0/4294967296.0,1,-nbitq), 
to_sfixed(-482638276.0/4294967296.0,1,-nbitq), 
to_sfixed(-387837549.0/4294967296.0,1,-nbitq), 
to_sfixed(144227850.0/4294967296.0,1,-nbitq), 
to_sfixed(185770927.0/4294967296.0,1,-nbitq), 
to_sfixed(-148669880.0/4294967296.0,1,-nbitq), 
to_sfixed(288732575.0/4294967296.0,1,-nbitq), 
to_sfixed(305214782.0/4294967296.0,1,-nbitq), 
to_sfixed(-121091728.0/4294967296.0,1,-nbitq), 
to_sfixed(75673225.0/4294967296.0,1,-nbitq), 
to_sfixed(-574567659.0/4294967296.0,1,-nbitq), 
to_sfixed(-38333504.0/4294967296.0,1,-nbitq), 
to_sfixed(-207321919.0/4294967296.0,1,-nbitq), 
to_sfixed(-232310118.0/4294967296.0,1,-nbitq), 
to_sfixed(-186729390.0/4294967296.0,1,-nbitq), 
to_sfixed(255509248.0/4294967296.0,1,-nbitq), 
to_sfixed(-107001169.0/4294967296.0,1,-nbitq), 
to_sfixed(15125521.0/4294967296.0,1,-nbitq), 
to_sfixed(-142123942.0/4294967296.0,1,-nbitq), 
to_sfixed(117408576.0/4294967296.0,1,-nbitq), 
to_sfixed(240010278.0/4294967296.0,1,-nbitq), 
to_sfixed(-92683911.0/4294967296.0,1,-nbitq), 
to_sfixed(479720635.0/4294967296.0,1,-nbitq), 
to_sfixed(-383494242.0/4294967296.0,1,-nbitq), 
to_sfixed(-12222820.0/4294967296.0,1,-nbitq), 
to_sfixed(119207615.0/4294967296.0,1,-nbitq), 
to_sfixed(-369549318.0/4294967296.0,1,-nbitq), 
to_sfixed(393565766.0/4294967296.0,1,-nbitq), 
to_sfixed(-254104555.0/4294967296.0,1,-nbitq), 
to_sfixed(-313870770.0/4294967296.0,1,-nbitq), 
to_sfixed(-460557897.0/4294967296.0,1,-nbitq), 
to_sfixed(227471452.0/4294967296.0,1,-nbitq), 
to_sfixed(103965327.0/4294967296.0,1,-nbitq), 
to_sfixed(-10560044.0/4294967296.0,1,-nbitq), 
to_sfixed(-157229577.0/4294967296.0,1,-nbitq), 
to_sfixed(-530119823.0/4294967296.0,1,-nbitq), 
to_sfixed(134056062.0/4294967296.0,1,-nbitq), 
to_sfixed(460892322.0/4294967296.0,1,-nbitq), 
to_sfixed(-140692536.0/4294967296.0,1,-nbitq), 
to_sfixed(257679190.0/4294967296.0,1,-nbitq), 
to_sfixed(-212482518.0/4294967296.0,1,-nbitq), 
to_sfixed(270144036.0/4294967296.0,1,-nbitq), 
to_sfixed(208262765.0/4294967296.0,1,-nbitq), 
to_sfixed(211622494.0/4294967296.0,1,-nbitq), 
to_sfixed(92609161.0/4294967296.0,1,-nbitq), 
to_sfixed(246965700.0/4294967296.0,1,-nbitq), 
to_sfixed(-239055446.0/4294967296.0,1,-nbitq), 
to_sfixed(421917870.0/4294967296.0,1,-nbitq), 
to_sfixed(-8378342.0/4294967296.0,1,-nbitq), 
to_sfixed(419155138.0/4294967296.0,1,-nbitq), 
to_sfixed(-108868735.0/4294967296.0,1,-nbitq), 
to_sfixed(59902205.0/4294967296.0,1,-nbitq), 
to_sfixed(405668355.0/4294967296.0,1,-nbitq), 
to_sfixed(60604088.0/4294967296.0,1,-nbitq), 
to_sfixed(-169520980.0/4294967296.0,1,-nbitq), 
to_sfixed(-284785468.0/4294967296.0,1,-nbitq), 
to_sfixed(-284742132.0/4294967296.0,1,-nbitq), 
to_sfixed(-3073668.0/4294967296.0,1,-nbitq), 
to_sfixed(280721585.0/4294967296.0,1,-nbitq), 
to_sfixed(-98605844.0/4294967296.0,1,-nbitq), 
to_sfixed(-130970193.0/4294967296.0,1,-nbitq), 
to_sfixed(-167187046.0/4294967296.0,1,-nbitq), 
to_sfixed(161403769.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-355692349.0/4294967296.0,1,-nbitq), 
to_sfixed(-102091277.0/4294967296.0,1,-nbitq), 
to_sfixed(389744455.0/4294967296.0,1,-nbitq), 
to_sfixed(-340318922.0/4294967296.0,1,-nbitq), 
to_sfixed(184817304.0/4294967296.0,1,-nbitq), 
to_sfixed(-286666171.0/4294967296.0,1,-nbitq), 
to_sfixed(152661219.0/4294967296.0,1,-nbitq), 
to_sfixed(324942872.0/4294967296.0,1,-nbitq), 
to_sfixed(257503065.0/4294967296.0,1,-nbitq), 
to_sfixed(-12009282.0/4294967296.0,1,-nbitq), 
to_sfixed(345204747.0/4294967296.0,1,-nbitq), 
to_sfixed(412059339.0/4294967296.0,1,-nbitq), 
to_sfixed(94660788.0/4294967296.0,1,-nbitq), 
to_sfixed(-151848832.0/4294967296.0,1,-nbitq), 
to_sfixed(5581111.0/4294967296.0,1,-nbitq), 
to_sfixed(191900074.0/4294967296.0,1,-nbitq), 
to_sfixed(-145326475.0/4294967296.0,1,-nbitq), 
to_sfixed(-166716898.0/4294967296.0,1,-nbitq), 
to_sfixed(-120710563.0/4294967296.0,1,-nbitq), 
to_sfixed(17222797.0/4294967296.0,1,-nbitq), 
to_sfixed(-405287014.0/4294967296.0,1,-nbitq), 
to_sfixed(100848300.0/4294967296.0,1,-nbitq), 
to_sfixed(595043025.0/4294967296.0,1,-nbitq), 
to_sfixed(-285336054.0/4294967296.0,1,-nbitq), 
to_sfixed(57044309.0/4294967296.0,1,-nbitq), 
to_sfixed(53847023.0/4294967296.0,1,-nbitq), 
to_sfixed(25913868.0/4294967296.0,1,-nbitq), 
to_sfixed(96684119.0/4294967296.0,1,-nbitq), 
to_sfixed(419547375.0/4294967296.0,1,-nbitq), 
to_sfixed(443631183.0/4294967296.0,1,-nbitq), 
to_sfixed(-116810202.0/4294967296.0,1,-nbitq), 
to_sfixed(-138465112.0/4294967296.0,1,-nbitq), 
to_sfixed(443626328.0/4294967296.0,1,-nbitq), 
to_sfixed(-351559184.0/4294967296.0,1,-nbitq), 
to_sfixed(261725886.0/4294967296.0,1,-nbitq), 
to_sfixed(-63681483.0/4294967296.0,1,-nbitq), 
to_sfixed(-43280670.0/4294967296.0,1,-nbitq), 
to_sfixed(-66888101.0/4294967296.0,1,-nbitq), 
to_sfixed(-398943818.0/4294967296.0,1,-nbitq), 
to_sfixed(423408986.0/4294967296.0,1,-nbitq), 
to_sfixed(-306757608.0/4294967296.0,1,-nbitq), 
to_sfixed(494922851.0/4294967296.0,1,-nbitq), 
to_sfixed(248134572.0/4294967296.0,1,-nbitq), 
to_sfixed(242694614.0/4294967296.0,1,-nbitq), 
to_sfixed(-349229718.0/4294967296.0,1,-nbitq), 
to_sfixed(431399284.0/4294967296.0,1,-nbitq), 
to_sfixed(-75028997.0/4294967296.0,1,-nbitq), 
to_sfixed(-438544824.0/4294967296.0,1,-nbitq), 
to_sfixed(322260743.0/4294967296.0,1,-nbitq), 
to_sfixed(347852699.0/4294967296.0,1,-nbitq), 
to_sfixed(19310807.0/4294967296.0,1,-nbitq), 
to_sfixed(-118560092.0/4294967296.0,1,-nbitq), 
to_sfixed(153914833.0/4294967296.0,1,-nbitq), 
to_sfixed(-73477096.0/4294967296.0,1,-nbitq), 
to_sfixed(-105971240.0/4294967296.0,1,-nbitq), 
to_sfixed(137941290.0/4294967296.0,1,-nbitq), 
to_sfixed(-323061606.0/4294967296.0,1,-nbitq), 
to_sfixed(-141557607.0/4294967296.0,1,-nbitq), 
to_sfixed(422022749.0/4294967296.0,1,-nbitq), 
to_sfixed(132288346.0/4294967296.0,1,-nbitq), 
to_sfixed(-305911770.0/4294967296.0,1,-nbitq), 
to_sfixed(-244490544.0/4294967296.0,1,-nbitq), 
to_sfixed(46873486.0/4294967296.0,1,-nbitq), 
to_sfixed(68716734.0/4294967296.0,1,-nbitq), 
to_sfixed(-146553467.0/4294967296.0,1,-nbitq), 
to_sfixed(-96539009.0/4294967296.0,1,-nbitq), 
to_sfixed(542420652.0/4294967296.0,1,-nbitq), 
to_sfixed(-256425198.0/4294967296.0,1,-nbitq), 
to_sfixed(432071187.0/4294967296.0,1,-nbitq), 
to_sfixed(227006801.0/4294967296.0,1,-nbitq), 
to_sfixed(217158280.0/4294967296.0,1,-nbitq), 
to_sfixed(108744917.0/4294967296.0,1,-nbitq), 
to_sfixed(-435084308.0/4294967296.0,1,-nbitq), 
to_sfixed(284345237.0/4294967296.0,1,-nbitq), 
to_sfixed(-16088183.0/4294967296.0,1,-nbitq), 
to_sfixed(-194076631.0/4294967296.0,1,-nbitq), 
to_sfixed(-188029332.0/4294967296.0,1,-nbitq), 
to_sfixed(172215716.0/4294967296.0,1,-nbitq), 
to_sfixed(-329742039.0/4294967296.0,1,-nbitq), 
to_sfixed(375072020.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(165074960.0/4294967296.0,1,-nbitq), 
to_sfixed(-214773277.0/4294967296.0,1,-nbitq), 
to_sfixed(198974355.0/4294967296.0,1,-nbitq), 
to_sfixed(78409191.0/4294967296.0,1,-nbitq), 
to_sfixed(267426231.0/4294967296.0,1,-nbitq), 
to_sfixed(272750467.0/4294967296.0,1,-nbitq), 
to_sfixed(394577487.0/4294967296.0,1,-nbitq), 
to_sfixed(109024109.0/4294967296.0,1,-nbitq), 
to_sfixed(-16386638.0/4294967296.0,1,-nbitq), 
to_sfixed(-243152747.0/4294967296.0,1,-nbitq), 
to_sfixed(-214325033.0/4294967296.0,1,-nbitq), 
to_sfixed(171285860.0/4294967296.0,1,-nbitq), 
to_sfixed(-411690793.0/4294967296.0,1,-nbitq), 
to_sfixed(434580374.0/4294967296.0,1,-nbitq), 
to_sfixed(-227958949.0/4294967296.0,1,-nbitq), 
to_sfixed(-38855663.0/4294967296.0,1,-nbitq), 
to_sfixed(23072903.0/4294967296.0,1,-nbitq), 
to_sfixed(-244634842.0/4294967296.0,1,-nbitq), 
to_sfixed(-70886881.0/4294967296.0,1,-nbitq), 
to_sfixed(197600738.0/4294967296.0,1,-nbitq), 
to_sfixed(188763163.0/4294967296.0,1,-nbitq), 
to_sfixed(-228187837.0/4294967296.0,1,-nbitq), 
to_sfixed(6576402.0/4294967296.0,1,-nbitq), 
to_sfixed(-249715225.0/4294967296.0,1,-nbitq), 
to_sfixed(123212573.0/4294967296.0,1,-nbitq), 
to_sfixed(-222008715.0/4294967296.0,1,-nbitq), 
to_sfixed(-9408608.0/4294967296.0,1,-nbitq), 
to_sfixed(-630661197.0/4294967296.0,1,-nbitq), 
to_sfixed(228435762.0/4294967296.0,1,-nbitq), 
to_sfixed(-274255301.0/4294967296.0,1,-nbitq), 
to_sfixed(123695266.0/4294967296.0,1,-nbitq), 
to_sfixed(-357404734.0/4294967296.0,1,-nbitq), 
to_sfixed(-271482493.0/4294967296.0,1,-nbitq), 
to_sfixed(39942669.0/4294967296.0,1,-nbitq), 
to_sfixed(176328002.0/4294967296.0,1,-nbitq), 
to_sfixed(383396150.0/4294967296.0,1,-nbitq), 
to_sfixed(84210776.0/4294967296.0,1,-nbitq), 
to_sfixed(50724480.0/4294967296.0,1,-nbitq), 
to_sfixed(254015622.0/4294967296.0,1,-nbitq), 
to_sfixed(-76696742.0/4294967296.0,1,-nbitq), 
to_sfixed(-400699171.0/4294967296.0,1,-nbitq), 
to_sfixed(417835451.0/4294967296.0,1,-nbitq), 
to_sfixed(317450493.0/4294967296.0,1,-nbitq), 
to_sfixed(316083366.0/4294967296.0,1,-nbitq), 
to_sfixed(123716830.0/4294967296.0,1,-nbitq), 
to_sfixed(72294644.0/4294967296.0,1,-nbitq), 
to_sfixed(-56382557.0/4294967296.0,1,-nbitq), 
to_sfixed(-554603581.0/4294967296.0,1,-nbitq), 
to_sfixed(28646299.0/4294967296.0,1,-nbitq), 
to_sfixed(173031384.0/4294967296.0,1,-nbitq), 
to_sfixed(50437518.0/4294967296.0,1,-nbitq), 
to_sfixed(242491006.0/4294967296.0,1,-nbitq), 
to_sfixed(61414753.0/4294967296.0,1,-nbitq), 
to_sfixed(445686680.0/4294967296.0,1,-nbitq), 
to_sfixed(422453621.0/4294967296.0,1,-nbitq), 
to_sfixed(461502818.0/4294967296.0,1,-nbitq), 
to_sfixed(-152409043.0/4294967296.0,1,-nbitq), 
to_sfixed(-494225585.0/4294967296.0,1,-nbitq), 
to_sfixed(216136207.0/4294967296.0,1,-nbitq), 
to_sfixed(13802532.0/4294967296.0,1,-nbitq), 
to_sfixed(-166024208.0/4294967296.0,1,-nbitq), 
to_sfixed(578800363.0/4294967296.0,1,-nbitq), 
to_sfixed(-101583984.0/4294967296.0,1,-nbitq), 
to_sfixed(-182487095.0/4294967296.0,1,-nbitq), 
to_sfixed(32476480.0/4294967296.0,1,-nbitq), 
to_sfixed(-410172874.0/4294967296.0,1,-nbitq), 
to_sfixed(639120475.0/4294967296.0,1,-nbitq), 
to_sfixed(-4158898.0/4294967296.0,1,-nbitq), 
to_sfixed(89843174.0/4294967296.0,1,-nbitq), 
to_sfixed(-120506675.0/4294967296.0,1,-nbitq), 
to_sfixed(284871919.0/4294967296.0,1,-nbitq), 
to_sfixed(323194582.0/4294967296.0,1,-nbitq), 
to_sfixed(99977381.0/4294967296.0,1,-nbitq), 
to_sfixed(-235852914.0/4294967296.0,1,-nbitq), 
to_sfixed(6346906.0/4294967296.0,1,-nbitq), 
to_sfixed(-424961319.0/4294967296.0,1,-nbitq), 
to_sfixed(-237782302.0/4294967296.0,1,-nbitq), 
to_sfixed(77405655.0/4294967296.0,1,-nbitq), 
to_sfixed(-64066793.0/4294967296.0,1,-nbitq), 
to_sfixed(102170953.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(127680221.0/4294967296.0,1,-nbitq), 
to_sfixed(-4172808.0/4294967296.0,1,-nbitq), 
to_sfixed(198712528.0/4294967296.0,1,-nbitq), 
to_sfixed(-249568676.0/4294967296.0,1,-nbitq), 
to_sfixed(253275105.0/4294967296.0,1,-nbitq), 
to_sfixed(203293505.0/4294967296.0,1,-nbitq), 
to_sfixed(247109785.0/4294967296.0,1,-nbitq), 
to_sfixed(242088921.0/4294967296.0,1,-nbitq), 
to_sfixed(45327712.0/4294967296.0,1,-nbitq), 
to_sfixed(114925272.0/4294967296.0,1,-nbitq), 
to_sfixed(326218720.0/4294967296.0,1,-nbitq), 
to_sfixed(430944573.0/4294967296.0,1,-nbitq), 
to_sfixed(96212350.0/4294967296.0,1,-nbitq), 
to_sfixed(-43153651.0/4294967296.0,1,-nbitq), 
to_sfixed(-198497707.0/4294967296.0,1,-nbitq), 
to_sfixed(-380515804.0/4294967296.0,1,-nbitq), 
to_sfixed(49512706.0/4294967296.0,1,-nbitq), 
to_sfixed(360097349.0/4294967296.0,1,-nbitq), 
to_sfixed(139452663.0/4294967296.0,1,-nbitq), 
to_sfixed(36982738.0/4294967296.0,1,-nbitq), 
to_sfixed(89955486.0/4294967296.0,1,-nbitq), 
to_sfixed(292776270.0/4294967296.0,1,-nbitq), 
to_sfixed(479135506.0/4294967296.0,1,-nbitq), 
to_sfixed(-183516382.0/4294967296.0,1,-nbitq), 
to_sfixed(-265584107.0/4294967296.0,1,-nbitq), 
to_sfixed(195211842.0/4294967296.0,1,-nbitq), 
to_sfixed(344053755.0/4294967296.0,1,-nbitq), 
to_sfixed(-172863353.0/4294967296.0,1,-nbitq), 
to_sfixed(305153726.0/4294967296.0,1,-nbitq), 
to_sfixed(109016205.0/4294967296.0,1,-nbitq), 
to_sfixed(87057895.0/4294967296.0,1,-nbitq), 
to_sfixed(109708564.0/4294967296.0,1,-nbitq), 
to_sfixed(220908766.0/4294967296.0,1,-nbitq), 
to_sfixed(-100934350.0/4294967296.0,1,-nbitq), 
to_sfixed(447998669.0/4294967296.0,1,-nbitq), 
to_sfixed(-57272450.0/4294967296.0,1,-nbitq), 
to_sfixed(176384056.0/4294967296.0,1,-nbitq), 
to_sfixed(312923338.0/4294967296.0,1,-nbitq), 
to_sfixed(102475038.0/4294967296.0,1,-nbitq), 
to_sfixed(-263428362.0/4294967296.0,1,-nbitq), 
to_sfixed(219431906.0/4294967296.0,1,-nbitq), 
to_sfixed(468756353.0/4294967296.0,1,-nbitq), 
to_sfixed(74822827.0/4294967296.0,1,-nbitq), 
to_sfixed(233449690.0/4294967296.0,1,-nbitq), 
to_sfixed(276589902.0/4294967296.0,1,-nbitq), 
to_sfixed(319820756.0/4294967296.0,1,-nbitq), 
to_sfixed(-69604298.0/4294967296.0,1,-nbitq), 
to_sfixed(-53664752.0/4294967296.0,1,-nbitq), 
to_sfixed(-405622431.0/4294967296.0,1,-nbitq), 
to_sfixed(346160696.0/4294967296.0,1,-nbitq), 
to_sfixed(119589389.0/4294967296.0,1,-nbitq), 
to_sfixed(280081891.0/4294967296.0,1,-nbitq), 
to_sfixed(-337048206.0/4294967296.0,1,-nbitq), 
to_sfixed(-93215076.0/4294967296.0,1,-nbitq), 
to_sfixed(79565091.0/4294967296.0,1,-nbitq), 
to_sfixed(14111068.0/4294967296.0,1,-nbitq), 
to_sfixed(-227281720.0/4294967296.0,1,-nbitq), 
to_sfixed(93550736.0/4294967296.0,1,-nbitq), 
to_sfixed(258183260.0/4294967296.0,1,-nbitq), 
to_sfixed(-345175887.0/4294967296.0,1,-nbitq), 
to_sfixed(-38412260.0/4294967296.0,1,-nbitq), 
to_sfixed(333639250.0/4294967296.0,1,-nbitq), 
to_sfixed(98826756.0/4294967296.0,1,-nbitq), 
to_sfixed(240102591.0/4294967296.0,1,-nbitq), 
to_sfixed(-23421322.0/4294967296.0,1,-nbitq), 
to_sfixed(273943502.0/4294967296.0,1,-nbitq), 
to_sfixed(717020446.0/4294967296.0,1,-nbitq), 
to_sfixed(253392360.0/4294967296.0,1,-nbitq), 
to_sfixed(345381793.0/4294967296.0,1,-nbitq), 
to_sfixed(-60786455.0/4294967296.0,1,-nbitq), 
to_sfixed(148186694.0/4294967296.0,1,-nbitq), 
to_sfixed(-157619247.0/4294967296.0,1,-nbitq), 
to_sfixed(-437159003.0/4294967296.0,1,-nbitq), 
to_sfixed(344311905.0/4294967296.0,1,-nbitq), 
to_sfixed(365004588.0/4294967296.0,1,-nbitq), 
to_sfixed(-357014564.0/4294967296.0,1,-nbitq), 
to_sfixed(-306408377.0/4294967296.0,1,-nbitq), 
to_sfixed(32695097.0/4294967296.0,1,-nbitq), 
to_sfixed(-142918258.0/4294967296.0,1,-nbitq), 
to_sfixed(275747399.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(158958412.0/4294967296.0,1,-nbitq), 
to_sfixed(-392370528.0/4294967296.0,1,-nbitq), 
to_sfixed(202368289.0/4294967296.0,1,-nbitq), 
to_sfixed(382884119.0/4294967296.0,1,-nbitq), 
to_sfixed(151779186.0/4294967296.0,1,-nbitq), 
to_sfixed(-58055557.0/4294967296.0,1,-nbitq), 
to_sfixed(-5688970.0/4294967296.0,1,-nbitq), 
to_sfixed(104348162.0/4294967296.0,1,-nbitq), 
to_sfixed(559157820.0/4294967296.0,1,-nbitq), 
to_sfixed(-114737844.0/4294967296.0,1,-nbitq), 
to_sfixed(-17264533.0/4294967296.0,1,-nbitq), 
to_sfixed(383124163.0/4294967296.0,1,-nbitq), 
to_sfixed(-56546652.0/4294967296.0,1,-nbitq), 
to_sfixed(294849546.0/4294967296.0,1,-nbitq), 
to_sfixed(207628140.0/4294967296.0,1,-nbitq), 
to_sfixed(-364170320.0/4294967296.0,1,-nbitq), 
to_sfixed(269738710.0/4294967296.0,1,-nbitq), 
to_sfixed(-352466845.0/4294967296.0,1,-nbitq), 
to_sfixed(79872418.0/4294967296.0,1,-nbitq), 
to_sfixed(-231731418.0/4294967296.0,1,-nbitq), 
to_sfixed(-95800542.0/4294967296.0,1,-nbitq), 
to_sfixed(471474357.0/4294967296.0,1,-nbitq), 
to_sfixed(409631981.0/4294967296.0,1,-nbitq), 
to_sfixed(-264629376.0/4294967296.0,1,-nbitq), 
to_sfixed(304538513.0/4294967296.0,1,-nbitq), 
to_sfixed(360446361.0/4294967296.0,1,-nbitq), 
to_sfixed(369283287.0/4294967296.0,1,-nbitq), 
to_sfixed(-374828937.0/4294967296.0,1,-nbitq), 
to_sfixed(3294932.0/4294967296.0,1,-nbitq), 
to_sfixed(-94529431.0/4294967296.0,1,-nbitq), 
to_sfixed(-250933589.0/4294967296.0,1,-nbitq), 
to_sfixed(-223226234.0/4294967296.0,1,-nbitq), 
to_sfixed(361988738.0/4294967296.0,1,-nbitq), 
to_sfixed(-483721167.0/4294967296.0,1,-nbitq), 
to_sfixed(28041507.0/4294967296.0,1,-nbitq), 
to_sfixed(304332457.0/4294967296.0,1,-nbitq), 
to_sfixed(38556180.0/4294967296.0,1,-nbitq), 
to_sfixed(-154655205.0/4294967296.0,1,-nbitq), 
to_sfixed(-436418352.0/4294967296.0,1,-nbitq), 
to_sfixed(-227803695.0/4294967296.0,1,-nbitq), 
to_sfixed(-255682344.0/4294967296.0,1,-nbitq), 
to_sfixed(-8242737.0/4294967296.0,1,-nbitq), 
to_sfixed(-137705547.0/4294967296.0,1,-nbitq), 
to_sfixed(-332186122.0/4294967296.0,1,-nbitq), 
to_sfixed(848139.0/4294967296.0,1,-nbitq), 
to_sfixed(201801505.0/4294967296.0,1,-nbitq), 
to_sfixed(-275341044.0/4294967296.0,1,-nbitq), 
to_sfixed(158681762.0/4294967296.0,1,-nbitq), 
to_sfixed(102763327.0/4294967296.0,1,-nbitq), 
to_sfixed(-215586283.0/4294967296.0,1,-nbitq), 
to_sfixed(51652366.0/4294967296.0,1,-nbitq), 
to_sfixed(-156637953.0/4294967296.0,1,-nbitq), 
to_sfixed(-547931861.0/4294967296.0,1,-nbitq), 
to_sfixed(-25079602.0/4294967296.0,1,-nbitq), 
to_sfixed(82597053.0/4294967296.0,1,-nbitq), 
to_sfixed(-243955601.0/4294967296.0,1,-nbitq), 
to_sfixed(17492719.0/4294967296.0,1,-nbitq), 
to_sfixed(-59477997.0/4294967296.0,1,-nbitq), 
to_sfixed(-291824046.0/4294967296.0,1,-nbitq), 
to_sfixed(398285133.0/4294967296.0,1,-nbitq), 
to_sfixed(342659831.0/4294967296.0,1,-nbitq), 
to_sfixed(26646916.0/4294967296.0,1,-nbitq), 
to_sfixed(-607991487.0/4294967296.0,1,-nbitq), 
to_sfixed(-274631082.0/4294967296.0,1,-nbitq), 
to_sfixed(-358790752.0/4294967296.0,1,-nbitq), 
to_sfixed(-301325431.0/4294967296.0,1,-nbitq), 
to_sfixed(250124270.0/4294967296.0,1,-nbitq), 
to_sfixed(352369596.0/4294967296.0,1,-nbitq), 
to_sfixed(-220500790.0/4294967296.0,1,-nbitq), 
to_sfixed(-171789620.0/4294967296.0,1,-nbitq), 
to_sfixed(20892913.0/4294967296.0,1,-nbitq), 
to_sfixed(363045245.0/4294967296.0,1,-nbitq), 
to_sfixed(-343238050.0/4294967296.0,1,-nbitq), 
to_sfixed(234669734.0/4294967296.0,1,-nbitq), 
to_sfixed(111211814.0/4294967296.0,1,-nbitq), 
to_sfixed(-264005050.0/4294967296.0,1,-nbitq), 
to_sfixed(503299924.0/4294967296.0,1,-nbitq), 
to_sfixed(-324905048.0/4294967296.0,1,-nbitq), 
to_sfixed(-499989334.0/4294967296.0,1,-nbitq), 
to_sfixed(-366154221.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-58154254.0/4294967296.0,1,-nbitq), 
to_sfixed(-473940415.0/4294967296.0,1,-nbitq), 
to_sfixed(262326587.0/4294967296.0,1,-nbitq), 
to_sfixed(-279855148.0/4294967296.0,1,-nbitq), 
to_sfixed(-219346349.0/4294967296.0,1,-nbitq), 
to_sfixed(-374860110.0/4294967296.0,1,-nbitq), 
to_sfixed(8479771.0/4294967296.0,1,-nbitq), 
to_sfixed(-348612939.0/4294967296.0,1,-nbitq), 
to_sfixed(193237048.0/4294967296.0,1,-nbitq), 
to_sfixed(190598603.0/4294967296.0,1,-nbitq), 
to_sfixed(-173171434.0/4294967296.0,1,-nbitq), 
to_sfixed(-74962398.0/4294967296.0,1,-nbitq), 
to_sfixed(-477393407.0/4294967296.0,1,-nbitq), 
to_sfixed(-174946237.0/4294967296.0,1,-nbitq), 
to_sfixed(161672638.0/4294967296.0,1,-nbitq), 
to_sfixed(49753540.0/4294967296.0,1,-nbitq), 
to_sfixed(-410861425.0/4294967296.0,1,-nbitq), 
to_sfixed(354580259.0/4294967296.0,1,-nbitq), 
to_sfixed(90090508.0/4294967296.0,1,-nbitq), 
to_sfixed(-14074110.0/4294967296.0,1,-nbitq), 
to_sfixed(-287134345.0/4294967296.0,1,-nbitq), 
to_sfixed(-126791922.0/4294967296.0,1,-nbitq), 
to_sfixed(150126393.0/4294967296.0,1,-nbitq), 
to_sfixed(8720768.0/4294967296.0,1,-nbitq), 
to_sfixed(15670611.0/4294967296.0,1,-nbitq), 
to_sfixed(303245910.0/4294967296.0,1,-nbitq), 
to_sfixed(-220017584.0/4294967296.0,1,-nbitq), 
to_sfixed(-147466385.0/4294967296.0,1,-nbitq), 
to_sfixed(12597512.0/4294967296.0,1,-nbitq), 
to_sfixed(85346932.0/4294967296.0,1,-nbitq), 
to_sfixed(-82810442.0/4294967296.0,1,-nbitq), 
to_sfixed(-651524974.0/4294967296.0,1,-nbitq), 
to_sfixed(283518729.0/4294967296.0,1,-nbitq), 
to_sfixed(-257452892.0/4294967296.0,1,-nbitq), 
to_sfixed(-101800233.0/4294967296.0,1,-nbitq), 
to_sfixed(537933453.0/4294967296.0,1,-nbitq), 
to_sfixed(273186798.0/4294967296.0,1,-nbitq), 
to_sfixed(1309267.0/4294967296.0,1,-nbitq), 
to_sfixed(-514699722.0/4294967296.0,1,-nbitq), 
to_sfixed(289037796.0/4294967296.0,1,-nbitq), 
to_sfixed(-355247036.0/4294967296.0,1,-nbitq), 
to_sfixed(-52542631.0/4294967296.0,1,-nbitq), 
to_sfixed(-38309620.0/4294967296.0,1,-nbitq), 
to_sfixed(8379662.0/4294967296.0,1,-nbitq), 
to_sfixed(395387018.0/4294967296.0,1,-nbitq), 
to_sfixed(367787256.0/4294967296.0,1,-nbitq), 
to_sfixed(335144676.0/4294967296.0,1,-nbitq), 
to_sfixed(-325490065.0/4294967296.0,1,-nbitq), 
to_sfixed(279738467.0/4294967296.0,1,-nbitq), 
to_sfixed(162178863.0/4294967296.0,1,-nbitq), 
to_sfixed(-82590459.0/4294967296.0,1,-nbitq), 
to_sfixed(435658871.0/4294967296.0,1,-nbitq), 
to_sfixed(-633703787.0/4294967296.0,1,-nbitq), 
to_sfixed(-79687105.0/4294967296.0,1,-nbitq), 
to_sfixed(-172119946.0/4294967296.0,1,-nbitq), 
to_sfixed(498395408.0/4294967296.0,1,-nbitq), 
to_sfixed(-253513347.0/4294967296.0,1,-nbitq), 
to_sfixed(-312386558.0/4294967296.0,1,-nbitq), 
to_sfixed(357193020.0/4294967296.0,1,-nbitq), 
to_sfixed(409253958.0/4294967296.0,1,-nbitq), 
to_sfixed(240130982.0/4294967296.0,1,-nbitq), 
to_sfixed(378110290.0/4294967296.0,1,-nbitq), 
to_sfixed(-118616768.0/4294967296.0,1,-nbitq), 
to_sfixed(370302285.0/4294967296.0,1,-nbitq), 
to_sfixed(398632332.0/4294967296.0,1,-nbitq), 
to_sfixed(-418350558.0/4294967296.0,1,-nbitq), 
to_sfixed(57999714.0/4294967296.0,1,-nbitq), 
to_sfixed(-158680534.0/4294967296.0,1,-nbitq), 
to_sfixed(-295944457.0/4294967296.0,1,-nbitq), 
to_sfixed(202378234.0/4294967296.0,1,-nbitq), 
to_sfixed(173165063.0/4294967296.0,1,-nbitq), 
to_sfixed(214133738.0/4294967296.0,1,-nbitq), 
to_sfixed(-332502920.0/4294967296.0,1,-nbitq), 
to_sfixed(276297275.0/4294967296.0,1,-nbitq), 
to_sfixed(308865483.0/4294967296.0,1,-nbitq), 
to_sfixed(214154231.0/4294967296.0,1,-nbitq), 
to_sfixed(194893504.0/4294967296.0,1,-nbitq), 
to_sfixed(340733090.0/4294967296.0,1,-nbitq), 
to_sfixed(-371740472.0/4294967296.0,1,-nbitq), 
to_sfixed(-346761409.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(76330304.0/4294967296.0,1,-nbitq), 
to_sfixed(191716655.0/4294967296.0,1,-nbitq), 
to_sfixed(444460697.0/4294967296.0,1,-nbitq), 
to_sfixed(171133576.0/4294967296.0,1,-nbitq), 
to_sfixed(519020846.0/4294967296.0,1,-nbitq), 
to_sfixed(111690575.0/4294967296.0,1,-nbitq), 
to_sfixed(329718457.0/4294967296.0,1,-nbitq), 
to_sfixed(272346996.0/4294967296.0,1,-nbitq), 
to_sfixed(85945864.0/4294967296.0,1,-nbitq), 
to_sfixed(172898660.0/4294967296.0,1,-nbitq), 
to_sfixed(396578688.0/4294967296.0,1,-nbitq), 
to_sfixed(137534684.0/4294967296.0,1,-nbitq), 
to_sfixed(-159121943.0/4294967296.0,1,-nbitq), 
to_sfixed(544026734.0/4294967296.0,1,-nbitq), 
to_sfixed(27667792.0/4294967296.0,1,-nbitq), 
to_sfixed(-297116204.0/4294967296.0,1,-nbitq), 
to_sfixed(-312127860.0/4294967296.0,1,-nbitq), 
to_sfixed(-9612266.0/4294967296.0,1,-nbitq), 
to_sfixed(-316294305.0/4294967296.0,1,-nbitq), 
to_sfixed(58419117.0/4294967296.0,1,-nbitq), 
to_sfixed(-193776854.0/4294967296.0,1,-nbitq), 
to_sfixed(518814894.0/4294967296.0,1,-nbitq), 
to_sfixed(83605170.0/4294967296.0,1,-nbitq), 
to_sfixed(-428763273.0/4294967296.0,1,-nbitq), 
to_sfixed(809858.0/4294967296.0,1,-nbitq), 
to_sfixed(-155575317.0/4294967296.0,1,-nbitq), 
to_sfixed(132799916.0/4294967296.0,1,-nbitq), 
to_sfixed(-525723138.0/4294967296.0,1,-nbitq), 
to_sfixed(293688469.0/4294967296.0,1,-nbitq), 
to_sfixed(428732785.0/4294967296.0,1,-nbitq), 
to_sfixed(-36586033.0/4294967296.0,1,-nbitq), 
to_sfixed(-227959146.0/4294967296.0,1,-nbitq), 
to_sfixed(127551109.0/4294967296.0,1,-nbitq), 
to_sfixed(58398965.0/4294967296.0,1,-nbitq), 
to_sfixed(330183603.0/4294967296.0,1,-nbitq), 
to_sfixed(42587970.0/4294967296.0,1,-nbitq), 
to_sfixed(347593866.0/4294967296.0,1,-nbitq), 
to_sfixed(-55286834.0/4294967296.0,1,-nbitq), 
to_sfixed(-194220732.0/4294967296.0,1,-nbitq), 
to_sfixed(-168555568.0/4294967296.0,1,-nbitq), 
to_sfixed(108445466.0/4294967296.0,1,-nbitq), 
to_sfixed(141887791.0/4294967296.0,1,-nbitq), 
to_sfixed(370126304.0/4294967296.0,1,-nbitq), 
to_sfixed(511848326.0/4294967296.0,1,-nbitq), 
to_sfixed(-170941503.0/4294967296.0,1,-nbitq), 
to_sfixed(-173706455.0/4294967296.0,1,-nbitq), 
to_sfixed(223044479.0/4294967296.0,1,-nbitq), 
to_sfixed(-125220896.0/4294967296.0,1,-nbitq), 
to_sfixed(-40126342.0/4294967296.0,1,-nbitq), 
to_sfixed(-72222964.0/4294967296.0,1,-nbitq), 
to_sfixed(-593506849.0/4294967296.0,1,-nbitq), 
to_sfixed(-145499101.0/4294967296.0,1,-nbitq), 
to_sfixed(-708828804.0/4294967296.0,1,-nbitq), 
to_sfixed(-5660963.0/4294967296.0,1,-nbitq), 
to_sfixed(-155618271.0/4294967296.0,1,-nbitq), 
to_sfixed(-91942364.0/4294967296.0,1,-nbitq), 
to_sfixed(-252540353.0/4294967296.0,1,-nbitq), 
to_sfixed(-162088435.0/4294967296.0,1,-nbitq), 
to_sfixed(378747708.0/4294967296.0,1,-nbitq), 
to_sfixed(212874469.0/4294967296.0,1,-nbitq), 
to_sfixed(-325324284.0/4294967296.0,1,-nbitq), 
to_sfixed(-16592109.0/4294967296.0,1,-nbitq), 
to_sfixed(-400406007.0/4294967296.0,1,-nbitq), 
to_sfixed(-353514681.0/4294967296.0,1,-nbitq), 
to_sfixed(-316556854.0/4294967296.0,1,-nbitq), 
to_sfixed(-106176339.0/4294967296.0,1,-nbitq), 
to_sfixed(473385260.0/4294967296.0,1,-nbitq), 
to_sfixed(43584217.0/4294967296.0,1,-nbitq), 
to_sfixed(428012600.0/4294967296.0,1,-nbitq), 
to_sfixed(-426961976.0/4294967296.0,1,-nbitq), 
to_sfixed(-204682344.0/4294967296.0,1,-nbitq), 
to_sfixed(-108809171.0/4294967296.0,1,-nbitq), 
to_sfixed(120622490.0/4294967296.0,1,-nbitq), 
to_sfixed(-204899032.0/4294967296.0,1,-nbitq), 
to_sfixed(-140202846.0/4294967296.0,1,-nbitq), 
to_sfixed(329866014.0/4294967296.0,1,-nbitq), 
to_sfixed(372694814.0/4294967296.0,1,-nbitq), 
to_sfixed(336403379.0/4294967296.0,1,-nbitq), 
to_sfixed(-187879383.0/4294967296.0,1,-nbitq), 
to_sfixed(333680693.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(243734140.0/4294967296.0,1,-nbitq), 
to_sfixed(-403847272.0/4294967296.0,1,-nbitq), 
to_sfixed(-75099472.0/4294967296.0,1,-nbitq), 
to_sfixed(-239288726.0/4294967296.0,1,-nbitq), 
to_sfixed(-72454059.0/4294967296.0,1,-nbitq), 
to_sfixed(-216655039.0/4294967296.0,1,-nbitq), 
to_sfixed(-164917059.0/4294967296.0,1,-nbitq), 
to_sfixed(-391057708.0/4294967296.0,1,-nbitq), 
to_sfixed(275188767.0/4294967296.0,1,-nbitq), 
to_sfixed(407618427.0/4294967296.0,1,-nbitq), 
to_sfixed(518567656.0/4294967296.0,1,-nbitq), 
to_sfixed(687092376.0/4294967296.0,1,-nbitq), 
to_sfixed(-80804810.0/4294967296.0,1,-nbitq), 
to_sfixed(590044533.0/4294967296.0,1,-nbitq), 
to_sfixed(232641458.0/4294967296.0,1,-nbitq), 
to_sfixed(-257682166.0/4294967296.0,1,-nbitq), 
to_sfixed(-394642517.0/4294967296.0,1,-nbitq), 
to_sfixed(343947060.0/4294967296.0,1,-nbitq), 
to_sfixed(322809049.0/4294967296.0,1,-nbitq), 
to_sfixed(-110538164.0/4294967296.0,1,-nbitq), 
to_sfixed(42400844.0/4294967296.0,1,-nbitq), 
to_sfixed(-226107596.0/4294967296.0,1,-nbitq), 
to_sfixed(184945275.0/4294967296.0,1,-nbitq), 
to_sfixed(318815227.0/4294967296.0,1,-nbitq), 
to_sfixed(-237925144.0/4294967296.0,1,-nbitq), 
to_sfixed(-184567064.0/4294967296.0,1,-nbitq), 
to_sfixed(187852178.0/4294967296.0,1,-nbitq), 
to_sfixed(-252892974.0/4294967296.0,1,-nbitq), 
to_sfixed(-9152666.0/4294967296.0,1,-nbitq), 
to_sfixed(172640831.0/4294967296.0,1,-nbitq), 
to_sfixed(110231495.0/4294967296.0,1,-nbitq), 
to_sfixed(79216966.0/4294967296.0,1,-nbitq), 
to_sfixed(-214071782.0/4294967296.0,1,-nbitq), 
to_sfixed(9214365.0/4294967296.0,1,-nbitq), 
to_sfixed(-406373461.0/4294967296.0,1,-nbitq), 
to_sfixed(20138159.0/4294967296.0,1,-nbitq), 
to_sfixed(41230220.0/4294967296.0,1,-nbitq), 
to_sfixed(415397358.0/4294967296.0,1,-nbitq), 
to_sfixed(36601145.0/4294967296.0,1,-nbitq), 
to_sfixed(147519122.0/4294967296.0,1,-nbitq), 
to_sfixed(147769885.0/4294967296.0,1,-nbitq), 
to_sfixed(438825144.0/4294967296.0,1,-nbitq), 
to_sfixed(119171043.0/4294967296.0,1,-nbitq), 
to_sfixed(80748846.0/4294967296.0,1,-nbitq), 
to_sfixed(259042430.0/4294967296.0,1,-nbitq), 
to_sfixed(390021908.0/4294967296.0,1,-nbitq), 
to_sfixed(-96280444.0/4294967296.0,1,-nbitq), 
to_sfixed(73084719.0/4294967296.0,1,-nbitq), 
to_sfixed(360877521.0/4294967296.0,1,-nbitq), 
to_sfixed(147561090.0/4294967296.0,1,-nbitq), 
to_sfixed(55682715.0/4294967296.0,1,-nbitq), 
to_sfixed(-279179555.0/4294967296.0,1,-nbitq), 
to_sfixed(-667762481.0/4294967296.0,1,-nbitq), 
to_sfixed(411209736.0/4294967296.0,1,-nbitq), 
to_sfixed(-259533504.0/4294967296.0,1,-nbitq), 
to_sfixed(13372947.0/4294967296.0,1,-nbitq), 
to_sfixed(-99618782.0/4294967296.0,1,-nbitq), 
to_sfixed(-432901659.0/4294967296.0,1,-nbitq), 
to_sfixed(-3516859.0/4294967296.0,1,-nbitq), 
to_sfixed(-251691512.0/4294967296.0,1,-nbitq), 
to_sfixed(-16271869.0/4294967296.0,1,-nbitq), 
to_sfixed(-111389597.0/4294967296.0,1,-nbitq), 
to_sfixed(-313051164.0/4294967296.0,1,-nbitq), 
to_sfixed(-83059.0/4294967296.0,1,-nbitq), 
to_sfixed(23047049.0/4294967296.0,1,-nbitq), 
to_sfixed(41542582.0/4294967296.0,1,-nbitq), 
to_sfixed(134484826.0/4294967296.0,1,-nbitq), 
to_sfixed(-239690241.0/4294967296.0,1,-nbitq), 
to_sfixed(-9345757.0/4294967296.0,1,-nbitq), 
to_sfixed(118894810.0/4294967296.0,1,-nbitq), 
to_sfixed(-274048971.0/4294967296.0,1,-nbitq), 
to_sfixed(274034111.0/4294967296.0,1,-nbitq), 
to_sfixed(282017662.0/4294967296.0,1,-nbitq), 
to_sfixed(-305700739.0/4294967296.0,1,-nbitq), 
to_sfixed(330768946.0/4294967296.0,1,-nbitq), 
to_sfixed(-151484841.0/4294967296.0,1,-nbitq), 
to_sfixed(-77746131.0/4294967296.0,1,-nbitq), 
to_sfixed(-155587218.0/4294967296.0,1,-nbitq), 
to_sfixed(-49937308.0/4294967296.0,1,-nbitq), 
to_sfixed(182144298.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(444766278.0/4294967296.0,1,-nbitq), 
to_sfixed(-37093698.0/4294967296.0,1,-nbitq), 
to_sfixed(533522627.0/4294967296.0,1,-nbitq), 
to_sfixed(-243476687.0/4294967296.0,1,-nbitq), 
to_sfixed(183710210.0/4294967296.0,1,-nbitq), 
to_sfixed(48378474.0/4294967296.0,1,-nbitq), 
to_sfixed(319659650.0/4294967296.0,1,-nbitq), 
to_sfixed(-105597459.0/4294967296.0,1,-nbitq), 
to_sfixed(598077788.0/4294967296.0,1,-nbitq), 
to_sfixed(412000401.0/4294967296.0,1,-nbitq), 
to_sfixed(363405905.0/4294967296.0,1,-nbitq), 
to_sfixed(428830541.0/4294967296.0,1,-nbitq), 
to_sfixed(-336637445.0/4294967296.0,1,-nbitq), 
to_sfixed(-48590748.0/4294967296.0,1,-nbitq), 
to_sfixed(341282227.0/4294967296.0,1,-nbitq), 
to_sfixed(-273073199.0/4294967296.0,1,-nbitq), 
to_sfixed(-87329824.0/4294967296.0,1,-nbitq), 
to_sfixed(-159763514.0/4294967296.0,1,-nbitq), 
to_sfixed(45007991.0/4294967296.0,1,-nbitq), 
to_sfixed(85946367.0/4294967296.0,1,-nbitq), 
to_sfixed(-98626133.0/4294967296.0,1,-nbitq), 
to_sfixed(-113487164.0/4294967296.0,1,-nbitq), 
to_sfixed(488572604.0/4294967296.0,1,-nbitq), 
to_sfixed(-231465440.0/4294967296.0,1,-nbitq), 
to_sfixed(-189595604.0/4294967296.0,1,-nbitq), 
to_sfixed(-325174280.0/4294967296.0,1,-nbitq), 
to_sfixed(212865737.0/4294967296.0,1,-nbitq), 
to_sfixed(-343134113.0/4294967296.0,1,-nbitq), 
to_sfixed(133380995.0/4294967296.0,1,-nbitq), 
to_sfixed(277931171.0/4294967296.0,1,-nbitq), 
to_sfixed(208302528.0/4294967296.0,1,-nbitq), 
to_sfixed(196498816.0/4294967296.0,1,-nbitq), 
to_sfixed(34625397.0/4294967296.0,1,-nbitq), 
to_sfixed(721468.0/4294967296.0,1,-nbitq), 
to_sfixed(6876752.0/4294967296.0,1,-nbitq), 
to_sfixed(237693963.0/4294967296.0,1,-nbitq), 
to_sfixed(121915803.0/4294967296.0,1,-nbitq), 
to_sfixed(-6162101.0/4294967296.0,1,-nbitq), 
to_sfixed(-409937354.0/4294967296.0,1,-nbitq), 
to_sfixed(308095290.0/4294967296.0,1,-nbitq), 
to_sfixed(205898691.0/4294967296.0,1,-nbitq), 
to_sfixed(138456111.0/4294967296.0,1,-nbitq), 
to_sfixed(323880427.0/4294967296.0,1,-nbitq), 
to_sfixed(201447179.0/4294967296.0,1,-nbitq), 
to_sfixed(-313333080.0/4294967296.0,1,-nbitq), 
to_sfixed(235653383.0/4294967296.0,1,-nbitq), 
to_sfixed(-402290943.0/4294967296.0,1,-nbitq), 
to_sfixed(-24291302.0/4294967296.0,1,-nbitq), 
to_sfixed(55072196.0/4294967296.0,1,-nbitq), 
to_sfixed(280264523.0/4294967296.0,1,-nbitq), 
to_sfixed(-293911644.0/4294967296.0,1,-nbitq), 
to_sfixed(65273512.0/4294967296.0,1,-nbitq), 
to_sfixed(-465607135.0/4294967296.0,1,-nbitq), 
to_sfixed(373379929.0/4294967296.0,1,-nbitq), 
to_sfixed(-167671284.0/4294967296.0,1,-nbitq), 
to_sfixed(363131666.0/4294967296.0,1,-nbitq), 
to_sfixed(170320615.0/4294967296.0,1,-nbitq), 
to_sfixed(86685871.0/4294967296.0,1,-nbitq), 
to_sfixed(285496269.0/4294967296.0,1,-nbitq), 
to_sfixed(414892400.0/4294967296.0,1,-nbitq), 
to_sfixed(204071237.0/4294967296.0,1,-nbitq), 
to_sfixed(55720130.0/4294967296.0,1,-nbitq), 
to_sfixed(-450228719.0/4294967296.0,1,-nbitq), 
to_sfixed(166006289.0/4294967296.0,1,-nbitq), 
to_sfixed(-180106735.0/4294967296.0,1,-nbitq), 
to_sfixed(168723088.0/4294967296.0,1,-nbitq), 
to_sfixed(601961234.0/4294967296.0,1,-nbitq), 
to_sfixed(59384564.0/4294967296.0,1,-nbitq), 
to_sfixed(-353427111.0/4294967296.0,1,-nbitq), 
to_sfixed(-141186933.0/4294967296.0,1,-nbitq), 
to_sfixed(-127423883.0/4294967296.0,1,-nbitq), 
to_sfixed(-279734790.0/4294967296.0,1,-nbitq), 
to_sfixed(-14665016.0/4294967296.0,1,-nbitq), 
to_sfixed(88865357.0/4294967296.0,1,-nbitq), 
to_sfixed(199986736.0/4294967296.0,1,-nbitq), 
to_sfixed(-163822271.0/4294967296.0,1,-nbitq), 
to_sfixed(-28101653.0/4294967296.0,1,-nbitq), 
to_sfixed(-106524622.0/4294967296.0,1,-nbitq), 
to_sfixed(-118606458.0/4294967296.0,1,-nbitq), 
to_sfixed(-26771145.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(135194484.0/4294967296.0,1,-nbitq), 
to_sfixed(253279406.0/4294967296.0,1,-nbitq), 
to_sfixed(-228342447.0/4294967296.0,1,-nbitq), 
to_sfixed(-220355222.0/4294967296.0,1,-nbitq), 
to_sfixed(475394608.0/4294967296.0,1,-nbitq), 
to_sfixed(-199960252.0/4294967296.0,1,-nbitq), 
to_sfixed(-123263302.0/4294967296.0,1,-nbitq), 
to_sfixed(68722479.0/4294967296.0,1,-nbitq), 
to_sfixed(702863335.0/4294967296.0,1,-nbitq), 
to_sfixed(-281567802.0/4294967296.0,1,-nbitq), 
to_sfixed(390418059.0/4294967296.0,1,-nbitq), 
to_sfixed(121049219.0/4294967296.0,1,-nbitq), 
to_sfixed(-555294275.0/4294967296.0,1,-nbitq), 
to_sfixed(-224986734.0/4294967296.0,1,-nbitq), 
to_sfixed(41959521.0/4294967296.0,1,-nbitq), 
to_sfixed(276606466.0/4294967296.0,1,-nbitq), 
to_sfixed(-14913823.0/4294967296.0,1,-nbitq), 
to_sfixed(112242209.0/4294967296.0,1,-nbitq), 
to_sfixed(117332892.0/4294967296.0,1,-nbitq), 
to_sfixed(-233290117.0/4294967296.0,1,-nbitq), 
to_sfixed(-25335074.0/4294967296.0,1,-nbitq), 
to_sfixed(-280464528.0/4294967296.0,1,-nbitq), 
to_sfixed(279796930.0/4294967296.0,1,-nbitq), 
to_sfixed(55329422.0/4294967296.0,1,-nbitq), 
to_sfixed(254664422.0/4294967296.0,1,-nbitq), 
to_sfixed(-359144601.0/4294967296.0,1,-nbitq), 
to_sfixed(386210568.0/4294967296.0,1,-nbitq), 
to_sfixed(161906918.0/4294967296.0,1,-nbitq), 
to_sfixed(303679093.0/4294967296.0,1,-nbitq), 
to_sfixed(-378197913.0/4294967296.0,1,-nbitq), 
to_sfixed(175857167.0/4294967296.0,1,-nbitq), 
to_sfixed(330109083.0/4294967296.0,1,-nbitq), 
to_sfixed(149752287.0/4294967296.0,1,-nbitq), 
to_sfixed(3068701.0/4294967296.0,1,-nbitq), 
to_sfixed(-468445593.0/4294967296.0,1,-nbitq), 
to_sfixed(-304291717.0/4294967296.0,1,-nbitq), 
to_sfixed(-245995894.0/4294967296.0,1,-nbitq), 
to_sfixed(99373774.0/4294967296.0,1,-nbitq), 
to_sfixed(-494624014.0/4294967296.0,1,-nbitq), 
to_sfixed(100831114.0/4294967296.0,1,-nbitq), 
to_sfixed(390040938.0/4294967296.0,1,-nbitq), 
to_sfixed(-260890020.0/4294967296.0,1,-nbitq), 
to_sfixed(554710168.0/4294967296.0,1,-nbitq), 
to_sfixed(347945676.0/4294967296.0,1,-nbitq), 
to_sfixed(-252359877.0/4294967296.0,1,-nbitq), 
to_sfixed(-95705604.0/4294967296.0,1,-nbitq), 
to_sfixed(-4181494.0/4294967296.0,1,-nbitq), 
to_sfixed(-246579809.0/4294967296.0,1,-nbitq), 
to_sfixed(-111198980.0/4294967296.0,1,-nbitq), 
to_sfixed(19883212.0/4294967296.0,1,-nbitq), 
to_sfixed(-146886008.0/4294967296.0,1,-nbitq), 
to_sfixed(183858400.0/4294967296.0,1,-nbitq), 
to_sfixed(-505128012.0/4294967296.0,1,-nbitq), 
to_sfixed(274225154.0/4294967296.0,1,-nbitq), 
to_sfixed(112562850.0/4294967296.0,1,-nbitq), 
to_sfixed(-242948667.0/4294967296.0,1,-nbitq), 
to_sfixed(262813781.0/4294967296.0,1,-nbitq), 
to_sfixed(-325407726.0/4294967296.0,1,-nbitq), 
to_sfixed(-308484852.0/4294967296.0,1,-nbitq), 
to_sfixed(-358470131.0/4294967296.0,1,-nbitq), 
to_sfixed(-68281051.0/4294967296.0,1,-nbitq), 
to_sfixed(336245461.0/4294967296.0,1,-nbitq), 
to_sfixed(197149041.0/4294967296.0,1,-nbitq), 
to_sfixed(275031622.0/4294967296.0,1,-nbitq), 
to_sfixed(150154781.0/4294967296.0,1,-nbitq), 
to_sfixed(65271299.0/4294967296.0,1,-nbitq), 
to_sfixed(139350852.0/4294967296.0,1,-nbitq), 
to_sfixed(-300863553.0/4294967296.0,1,-nbitq), 
to_sfixed(43419593.0/4294967296.0,1,-nbitq), 
to_sfixed(-470402627.0/4294967296.0,1,-nbitq), 
to_sfixed(-436393218.0/4294967296.0,1,-nbitq), 
to_sfixed(180954395.0/4294967296.0,1,-nbitq), 
to_sfixed(-60603303.0/4294967296.0,1,-nbitq), 
to_sfixed(141773640.0/4294967296.0,1,-nbitq), 
to_sfixed(-203109970.0/4294967296.0,1,-nbitq), 
to_sfixed(-397821534.0/4294967296.0,1,-nbitq), 
to_sfixed(430316417.0/4294967296.0,1,-nbitq), 
to_sfixed(-553490412.0/4294967296.0,1,-nbitq), 
to_sfixed(256554825.0/4294967296.0,1,-nbitq), 
to_sfixed(150754628.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(340787913.0/4294967296.0,1,-nbitq), 
to_sfixed(259412211.0/4294967296.0,1,-nbitq), 
to_sfixed(-155631690.0/4294967296.0,1,-nbitq), 
to_sfixed(83718400.0/4294967296.0,1,-nbitq), 
to_sfixed(464332625.0/4294967296.0,1,-nbitq), 
to_sfixed(154216504.0/4294967296.0,1,-nbitq), 
to_sfixed(-175632374.0/4294967296.0,1,-nbitq), 
to_sfixed(139465257.0/4294967296.0,1,-nbitq), 
to_sfixed(298008594.0/4294967296.0,1,-nbitq), 
to_sfixed(86007801.0/4294967296.0,1,-nbitq), 
to_sfixed(415469698.0/4294967296.0,1,-nbitq), 
to_sfixed(356113123.0/4294967296.0,1,-nbitq), 
to_sfixed(-447417605.0/4294967296.0,1,-nbitq), 
to_sfixed(310383229.0/4294967296.0,1,-nbitq), 
to_sfixed(165386030.0/4294967296.0,1,-nbitq), 
to_sfixed(-153908994.0/4294967296.0,1,-nbitq), 
to_sfixed(-264796013.0/4294967296.0,1,-nbitq), 
to_sfixed(250612776.0/4294967296.0,1,-nbitq), 
to_sfixed(128208694.0/4294967296.0,1,-nbitq), 
to_sfixed(362260101.0/4294967296.0,1,-nbitq), 
to_sfixed(40667554.0/4294967296.0,1,-nbitq), 
to_sfixed(341426576.0/4294967296.0,1,-nbitq), 
to_sfixed(324646480.0/4294967296.0,1,-nbitq), 
to_sfixed(-185815085.0/4294967296.0,1,-nbitq), 
to_sfixed(220418269.0/4294967296.0,1,-nbitq), 
to_sfixed(47100413.0/4294967296.0,1,-nbitq), 
to_sfixed(47188603.0/4294967296.0,1,-nbitq), 
to_sfixed(-295731203.0/4294967296.0,1,-nbitq), 
to_sfixed(566382112.0/4294967296.0,1,-nbitq), 
to_sfixed(24375286.0/4294967296.0,1,-nbitq), 
to_sfixed(76309043.0/4294967296.0,1,-nbitq), 
to_sfixed(448071757.0/4294967296.0,1,-nbitq), 
to_sfixed(105099129.0/4294967296.0,1,-nbitq), 
to_sfixed(-320831742.0/4294967296.0,1,-nbitq), 
to_sfixed(-364226555.0/4294967296.0,1,-nbitq), 
to_sfixed(-481395933.0/4294967296.0,1,-nbitq), 
to_sfixed(-91307238.0/4294967296.0,1,-nbitq), 
to_sfixed(218345769.0/4294967296.0,1,-nbitq), 
to_sfixed(-307453252.0/4294967296.0,1,-nbitq), 
to_sfixed(-34586161.0/4294967296.0,1,-nbitq), 
to_sfixed(-284009894.0/4294967296.0,1,-nbitq), 
to_sfixed(-243020187.0/4294967296.0,1,-nbitq), 
to_sfixed(405662755.0/4294967296.0,1,-nbitq), 
to_sfixed(-42005615.0/4294967296.0,1,-nbitq), 
to_sfixed(-201901159.0/4294967296.0,1,-nbitq), 
to_sfixed(376301428.0/4294967296.0,1,-nbitq), 
to_sfixed(102862347.0/4294967296.0,1,-nbitq), 
to_sfixed(-417968032.0/4294967296.0,1,-nbitq), 
to_sfixed(-28844663.0/4294967296.0,1,-nbitq), 
to_sfixed(445407965.0/4294967296.0,1,-nbitq), 
to_sfixed(-46129551.0/4294967296.0,1,-nbitq), 
to_sfixed(-160531063.0/4294967296.0,1,-nbitq), 
to_sfixed(-293816114.0/4294967296.0,1,-nbitq), 
to_sfixed(83116798.0/4294967296.0,1,-nbitq), 
to_sfixed(-47965912.0/4294967296.0,1,-nbitq), 
to_sfixed(-105559923.0/4294967296.0,1,-nbitq), 
to_sfixed(-245856366.0/4294967296.0,1,-nbitq), 
to_sfixed(-534474514.0/4294967296.0,1,-nbitq), 
to_sfixed(-27153414.0/4294967296.0,1,-nbitq), 
to_sfixed(-285402520.0/4294967296.0,1,-nbitq), 
to_sfixed(172447588.0/4294967296.0,1,-nbitq), 
to_sfixed(-149288969.0/4294967296.0,1,-nbitq), 
to_sfixed(275342241.0/4294967296.0,1,-nbitq), 
to_sfixed(-418221428.0/4294967296.0,1,-nbitq), 
to_sfixed(297866847.0/4294967296.0,1,-nbitq), 
to_sfixed(-262223770.0/4294967296.0,1,-nbitq), 
to_sfixed(837434382.0/4294967296.0,1,-nbitq), 
to_sfixed(-52492180.0/4294967296.0,1,-nbitq), 
to_sfixed(291588787.0/4294967296.0,1,-nbitq), 
to_sfixed(26272143.0/4294967296.0,1,-nbitq), 
to_sfixed(251168876.0/4294967296.0,1,-nbitq), 
to_sfixed(470422133.0/4294967296.0,1,-nbitq), 
to_sfixed(529149140.0/4294967296.0,1,-nbitq), 
to_sfixed(-96868163.0/4294967296.0,1,-nbitq), 
to_sfixed(99352792.0/4294967296.0,1,-nbitq), 
to_sfixed(-163015725.0/4294967296.0,1,-nbitq), 
to_sfixed(317562238.0/4294967296.0,1,-nbitq), 
to_sfixed(-343673280.0/4294967296.0,1,-nbitq), 
to_sfixed(75252737.0/4294967296.0,1,-nbitq), 
to_sfixed(-58909360.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-96782204.0/4294967296.0,1,-nbitq), 
to_sfixed(310556812.0/4294967296.0,1,-nbitq), 
to_sfixed(478507137.0/4294967296.0,1,-nbitq), 
to_sfixed(-77782859.0/4294967296.0,1,-nbitq), 
to_sfixed(-644129.0/4294967296.0,1,-nbitq), 
to_sfixed(-454267958.0/4294967296.0,1,-nbitq), 
to_sfixed(-146358647.0/4294967296.0,1,-nbitq), 
to_sfixed(28482465.0/4294967296.0,1,-nbitq), 
to_sfixed(347734853.0/4294967296.0,1,-nbitq), 
to_sfixed(-353123728.0/4294967296.0,1,-nbitq), 
to_sfixed(338337290.0/4294967296.0,1,-nbitq), 
to_sfixed(691472772.0/4294967296.0,1,-nbitq), 
to_sfixed(-426183378.0/4294967296.0,1,-nbitq), 
to_sfixed(-104109369.0/4294967296.0,1,-nbitq), 
to_sfixed(-129578256.0/4294967296.0,1,-nbitq), 
to_sfixed(-115915696.0/4294967296.0,1,-nbitq), 
to_sfixed(-409301456.0/4294967296.0,1,-nbitq), 
to_sfixed(-26200202.0/4294967296.0,1,-nbitq), 
to_sfixed(94406429.0/4294967296.0,1,-nbitq), 
to_sfixed(-11443917.0/4294967296.0,1,-nbitq), 
to_sfixed(-316505315.0/4294967296.0,1,-nbitq), 
to_sfixed(128611867.0/4294967296.0,1,-nbitq), 
to_sfixed(215947031.0/4294967296.0,1,-nbitq), 
to_sfixed(132675296.0/4294967296.0,1,-nbitq), 
to_sfixed(178593241.0/4294967296.0,1,-nbitq), 
to_sfixed(-187258859.0/4294967296.0,1,-nbitq), 
to_sfixed(124382714.0/4294967296.0,1,-nbitq), 
to_sfixed(-401372607.0/4294967296.0,1,-nbitq), 
to_sfixed(284323008.0/4294967296.0,1,-nbitq), 
to_sfixed(144153600.0/4294967296.0,1,-nbitq), 
to_sfixed(-19047981.0/4294967296.0,1,-nbitq), 
to_sfixed(33498695.0/4294967296.0,1,-nbitq), 
to_sfixed(603300653.0/4294967296.0,1,-nbitq), 
to_sfixed(224116387.0/4294967296.0,1,-nbitq), 
to_sfixed(-220033251.0/4294967296.0,1,-nbitq), 
to_sfixed(-226238897.0/4294967296.0,1,-nbitq), 
to_sfixed(-83249549.0/4294967296.0,1,-nbitq), 
to_sfixed(321124.0/4294967296.0,1,-nbitq), 
to_sfixed(-467995742.0/4294967296.0,1,-nbitq), 
to_sfixed(143619130.0/4294967296.0,1,-nbitq), 
to_sfixed(312195652.0/4294967296.0,1,-nbitq), 
to_sfixed(-129752370.0/4294967296.0,1,-nbitq), 
to_sfixed(-110839108.0/4294967296.0,1,-nbitq), 
to_sfixed(143093818.0/4294967296.0,1,-nbitq), 
to_sfixed(-116299858.0/4294967296.0,1,-nbitq), 
to_sfixed(-89274637.0/4294967296.0,1,-nbitq), 
to_sfixed(-111983036.0/4294967296.0,1,-nbitq), 
to_sfixed(-59013258.0/4294967296.0,1,-nbitq), 
to_sfixed(61725992.0/4294967296.0,1,-nbitq), 
to_sfixed(87098401.0/4294967296.0,1,-nbitq), 
to_sfixed(-572166411.0/4294967296.0,1,-nbitq), 
to_sfixed(-193472002.0/4294967296.0,1,-nbitq), 
to_sfixed(-251138384.0/4294967296.0,1,-nbitq), 
to_sfixed(156492588.0/4294967296.0,1,-nbitq), 
to_sfixed(-14111541.0/4294967296.0,1,-nbitq), 
to_sfixed(-169848256.0/4294967296.0,1,-nbitq), 
to_sfixed(224562939.0/4294967296.0,1,-nbitq), 
to_sfixed(-522360987.0/4294967296.0,1,-nbitq), 
to_sfixed(-180044527.0/4294967296.0,1,-nbitq), 
to_sfixed(130178741.0/4294967296.0,1,-nbitq), 
to_sfixed(-295172115.0/4294967296.0,1,-nbitq), 
to_sfixed(-167923889.0/4294967296.0,1,-nbitq), 
to_sfixed(-101163822.0/4294967296.0,1,-nbitq), 
to_sfixed(-82379321.0/4294967296.0,1,-nbitq), 
to_sfixed(-45595370.0/4294967296.0,1,-nbitq), 
to_sfixed(-380303021.0/4294967296.0,1,-nbitq), 
to_sfixed(336437396.0/4294967296.0,1,-nbitq), 
to_sfixed(-163462866.0/4294967296.0,1,-nbitq), 
to_sfixed(388878402.0/4294967296.0,1,-nbitq), 
to_sfixed(72565467.0/4294967296.0,1,-nbitq), 
to_sfixed(-530532216.0/4294967296.0,1,-nbitq), 
to_sfixed(-244124174.0/4294967296.0,1,-nbitq), 
to_sfixed(69483455.0/4294967296.0,1,-nbitq), 
to_sfixed(354144303.0/4294967296.0,1,-nbitq), 
to_sfixed(42691298.0/4294967296.0,1,-nbitq), 
to_sfixed(97764567.0/4294967296.0,1,-nbitq), 
to_sfixed(-27209628.0/4294967296.0,1,-nbitq), 
to_sfixed(-62055771.0/4294967296.0,1,-nbitq), 
to_sfixed(3373107.0/4294967296.0,1,-nbitq), 
to_sfixed(-131533731.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-79351397.0/4294967296.0,1,-nbitq), 
to_sfixed(604832822.0/4294967296.0,1,-nbitq), 
to_sfixed(315382271.0/4294967296.0,1,-nbitq), 
to_sfixed(25067383.0/4294967296.0,1,-nbitq), 
to_sfixed(296017452.0/4294967296.0,1,-nbitq), 
to_sfixed(-505373747.0/4294967296.0,1,-nbitq), 
to_sfixed(249936900.0/4294967296.0,1,-nbitq), 
to_sfixed(-300110827.0/4294967296.0,1,-nbitq), 
to_sfixed(321059737.0/4294967296.0,1,-nbitq), 
to_sfixed(245791190.0/4294967296.0,1,-nbitq), 
to_sfixed(42926229.0/4294967296.0,1,-nbitq), 
to_sfixed(614502930.0/4294967296.0,1,-nbitq), 
to_sfixed(-323620284.0/4294967296.0,1,-nbitq), 
to_sfixed(36049358.0/4294967296.0,1,-nbitq), 
to_sfixed(-310694710.0/4294967296.0,1,-nbitq), 
to_sfixed(-212026189.0/4294967296.0,1,-nbitq), 
to_sfixed(-43261948.0/4294967296.0,1,-nbitq), 
to_sfixed(193944991.0/4294967296.0,1,-nbitq), 
to_sfixed(411091509.0/4294967296.0,1,-nbitq), 
to_sfixed(37656802.0/4294967296.0,1,-nbitq), 
to_sfixed(130682199.0/4294967296.0,1,-nbitq), 
to_sfixed(215920023.0/4294967296.0,1,-nbitq), 
to_sfixed(93470372.0/4294967296.0,1,-nbitq), 
to_sfixed(-69399529.0/4294967296.0,1,-nbitq), 
to_sfixed(-36890357.0/4294967296.0,1,-nbitq), 
to_sfixed(-206723086.0/4294967296.0,1,-nbitq), 
to_sfixed(-253089467.0/4294967296.0,1,-nbitq), 
to_sfixed(22560907.0/4294967296.0,1,-nbitq), 
to_sfixed(613364929.0/4294967296.0,1,-nbitq), 
to_sfixed(251096741.0/4294967296.0,1,-nbitq), 
to_sfixed(-312760642.0/4294967296.0,1,-nbitq), 
to_sfixed(259164211.0/4294967296.0,1,-nbitq), 
to_sfixed(396599411.0/4294967296.0,1,-nbitq), 
to_sfixed(117234849.0/4294967296.0,1,-nbitq), 
to_sfixed(-5183420.0/4294967296.0,1,-nbitq), 
to_sfixed(-668417515.0/4294967296.0,1,-nbitq), 
to_sfixed(-100105060.0/4294967296.0,1,-nbitq), 
to_sfixed(-285013178.0/4294967296.0,1,-nbitq), 
to_sfixed(73675324.0/4294967296.0,1,-nbitq), 
to_sfixed(-254051490.0/4294967296.0,1,-nbitq), 
to_sfixed(-74049279.0/4294967296.0,1,-nbitq), 
to_sfixed(162052663.0/4294967296.0,1,-nbitq), 
to_sfixed(-100037612.0/4294967296.0,1,-nbitq), 
to_sfixed(247187831.0/4294967296.0,1,-nbitq), 
to_sfixed(95579527.0/4294967296.0,1,-nbitq), 
to_sfixed(653803611.0/4294967296.0,1,-nbitq), 
to_sfixed(306693800.0/4294967296.0,1,-nbitq), 
to_sfixed(183464840.0/4294967296.0,1,-nbitq), 
to_sfixed(91106913.0/4294967296.0,1,-nbitq), 
to_sfixed(295590112.0/4294967296.0,1,-nbitq), 
to_sfixed(-515096879.0/4294967296.0,1,-nbitq), 
to_sfixed(54737056.0/4294967296.0,1,-nbitq), 
to_sfixed(77211478.0/4294967296.0,1,-nbitq), 
to_sfixed(430615203.0/4294967296.0,1,-nbitq), 
to_sfixed(256724124.0/4294967296.0,1,-nbitq), 
to_sfixed(-38403662.0/4294967296.0,1,-nbitq), 
to_sfixed(-298308675.0/4294967296.0,1,-nbitq), 
to_sfixed(-156254589.0/4294967296.0,1,-nbitq), 
to_sfixed(154958342.0/4294967296.0,1,-nbitq), 
to_sfixed(-190593100.0/4294967296.0,1,-nbitq), 
to_sfixed(-307344203.0/4294967296.0,1,-nbitq), 
to_sfixed(-215942566.0/4294967296.0,1,-nbitq), 
to_sfixed(-358514685.0/4294967296.0,1,-nbitq), 
to_sfixed(218122809.0/4294967296.0,1,-nbitq), 
to_sfixed(-69147945.0/4294967296.0,1,-nbitq), 
to_sfixed(46292066.0/4294967296.0,1,-nbitq), 
to_sfixed(108808943.0/4294967296.0,1,-nbitq), 
to_sfixed(-84722029.0/4294967296.0,1,-nbitq), 
to_sfixed(270343531.0/4294967296.0,1,-nbitq), 
to_sfixed(36723724.0/4294967296.0,1,-nbitq), 
to_sfixed(-268032201.0/4294967296.0,1,-nbitq), 
to_sfixed(175165020.0/4294967296.0,1,-nbitq), 
to_sfixed(-194904785.0/4294967296.0,1,-nbitq), 
to_sfixed(346985162.0/4294967296.0,1,-nbitq), 
to_sfixed(30313939.0/4294967296.0,1,-nbitq), 
to_sfixed(127944678.0/4294967296.0,1,-nbitq), 
to_sfixed(-168925964.0/4294967296.0,1,-nbitq), 
to_sfixed(-575069803.0/4294967296.0,1,-nbitq), 
to_sfixed(210891160.0/4294967296.0,1,-nbitq), 
to_sfixed(380477326.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(500907967.0/4294967296.0,1,-nbitq), 
to_sfixed(28869666.0/4294967296.0,1,-nbitq), 
to_sfixed(-199239227.0/4294967296.0,1,-nbitq), 
to_sfixed(196621320.0/4294967296.0,1,-nbitq), 
to_sfixed(-344543672.0/4294967296.0,1,-nbitq), 
to_sfixed(-211432223.0/4294967296.0,1,-nbitq), 
to_sfixed(-414184265.0/4294967296.0,1,-nbitq), 
to_sfixed(-195168704.0/4294967296.0,1,-nbitq), 
to_sfixed(-144504220.0/4294967296.0,1,-nbitq), 
to_sfixed(-330063132.0/4294967296.0,1,-nbitq), 
to_sfixed(-136815172.0/4294967296.0,1,-nbitq), 
to_sfixed(-231058711.0/4294967296.0,1,-nbitq), 
to_sfixed(-559262223.0/4294967296.0,1,-nbitq), 
to_sfixed(145636527.0/4294967296.0,1,-nbitq), 
to_sfixed(-188891471.0/4294967296.0,1,-nbitq), 
to_sfixed(-527812668.0/4294967296.0,1,-nbitq), 
to_sfixed(118987810.0/4294967296.0,1,-nbitq), 
to_sfixed(-252430546.0/4294967296.0,1,-nbitq), 
to_sfixed(150989066.0/4294967296.0,1,-nbitq), 
to_sfixed(-85820049.0/4294967296.0,1,-nbitq), 
to_sfixed(153050302.0/4294967296.0,1,-nbitq), 
to_sfixed(350748632.0/4294967296.0,1,-nbitq), 
to_sfixed(62244993.0/4294967296.0,1,-nbitq), 
to_sfixed(22589842.0/4294967296.0,1,-nbitq), 
to_sfixed(200166429.0/4294967296.0,1,-nbitq), 
to_sfixed(62524691.0/4294967296.0,1,-nbitq), 
to_sfixed(249342652.0/4294967296.0,1,-nbitq), 
to_sfixed(-196130443.0/4294967296.0,1,-nbitq), 
to_sfixed(385294374.0/4294967296.0,1,-nbitq), 
to_sfixed(155463425.0/4294967296.0,1,-nbitq), 
to_sfixed(-346049240.0/4294967296.0,1,-nbitq), 
to_sfixed(154979326.0/4294967296.0,1,-nbitq), 
to_sfixed(32006336.0/4294967296.0,1,-nbitq), 
to_sfixed(139837474.0/4294967296.0,1,-nbitq), 
to_sfixed(-174482165.0/4294967296.0,1,-nbitq), 
to_sfixed(-427144496.0/4294967296.0,1,-nbitq), 
to_sfixed(326996033.0/4294967296.0,1,-nbitq), 
to_sfixed(-16004482.0/4294967296.0,1,-nbitq), 
to_sfixed(-194693935.0/4294967296.0,1,-nbitq), 
to_sfixed(12026316.0/4294967296.0,1,-nbitq), 
to_sfixed(-148147496.0/4294967296.0,1,-nbitq), 
to_sfixed(-52496689.0/4294967296.0,1,-nbitq), 
to_sfixed(79040665.0/4294967296.0,1,-nbitq), 
to_sfixed(533826623.0/4294967296.0,1,-nbitq), 
to_sfixed(-312072529.0/4294967296.0,1,-nbitq), 
to_sfixed(29379301.0/4294967296.0,1,-nbitq), 
to_sfixed(-386653692.0/4294967296.0,1,-nbitq), 
to_sfixed(77978302.0/4294967296.0,1,-nbitq), 
to_sfixed(-201018974.0/4294967296.0,1,-nbitq), 
to_sfixed(312824784.0/4294967296.0,1,-nbitq), 
to_sfixed(-241247919.0/4294967296.0,1,-nbitq), 
to_sfixed(215776551.0/4294967296.0,1,-nbitq), 
to_sfixed(-370390476.0/4294967296.0,1,-nbitq), 
to_sfixed(-100418629.0/4294967296.0,1,-nbitq), 
to_sfixed(177655994.0/4294967296.0,1,-nbitq), 
to_sfixed(-135526884.0/4294967296.0,1,-nbitq), 
to_sfixed(-474628682.0/4294967296.0,1,-nbitq), 
to_sfixed(-91631968.0/4294967296.0,1,-nbitq), 
to_sfixed(228095628.0/4294967296.0,1,-nbitq), 
to_sfixed(124733592.0/4294967296.0,1,-nbitq), 
to_sfixed(-60013300.0/4294967296.0,1,-nbitq), 
to_sfixed(39217726.0/4294967296.0,1,-nbitq), 
to_sfixed(412409336.0/4294967296.0,1,-nbitq), 
to_sfixed(-477940073.0/4294967296.0,1,-nbitq), 
to_sfixed(165671241.0/4294967296.0,1,-nbitq), 
to_sfixed(-132493891.0/4294967296.0,1,-nbitq), 
to_sfixed(128872991.0/4294967296.0,1,-nbitq), 
to_sfixed(414376105.0/4294967296.0,1,-nbitq), 
to_sfixed(-13621031.0/4294967296.0,1,-nbitq), 
to_sfixed(-70519025.0/4294967296.0,1,-nbitq), 
to_sfixed(-370162637.0/4294967296.0,1,-nbitq), 
to_sfixed(397029229.0/4294967296.0,1,-nbitq), 
to_sfixed(71187583.0/4294967296.0,1,-nbitq), 
to_sfixed(357048480.0/4294967296.0,1,-nbitq), 
to_sfixed(124099462.0/4294967296.0,1,-nbitq), 
to_sfixed(-238217347.0/4294967296.0,1,-nbitq), 
to_sfixed(-66656071.0/4294967296.0,1,-nbitq), 
to_sfixed(-555417994.0/4294967296.0,1,-nbitq), 
to_sfixed(268268267.0/4294967296.0,1,-nbitq), 
to_sfixed(230153362.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-209980244.0/4294967296.0,1,-nbitq), 
to_sfixed(522423338.0/4294967296.0,1,-nbitq), 
to_sfixed(-289290462.0/4294967296.0,1,-nbitq), 
to_sfixed(211573610.0/4294967296.0,1,-nbitq), 
to_sfixed(-71849879.0/4294967296.0,1,-nbitq), 
to_sfixed(-115073304.0/4294967296.0,1,-nbitq), 
to_sfixed(351571430.0/4294967296.0,1,-nbitq), 
to_sfixed(107639248.0/4294967296.0,1,-nbitq), 
to_sfixed(271934094.0/4294967296.0,1,-nbitq), 
to_sfixed(348070944.0/4294967296.0,1,-nbitq), 
to_sfixed(-81264351.0/4294967296.0,1,-nbitq), 
to_sfixed(-252513262.0/4294967296.0,1,-nbitq), 
to_sfixed(-682821301.0/4294967296.0,1,-nbitq), 
to_sfixed(30815161.0/4294967296.0,1,-nbitq), 
to_sfixed(-8610531.0/4294967296.0,1,-nbitq), 
to_sfixed(-49637336.0/4294967296.0,1,-nbitq), 
to_sfixed(-48853420.0/4294967296.0,1,-nbitq), 
to_sfixed(386138127.0/4294967296.0,1,-nbitq), 
to_sfixed(192975783.0/4294967296.0,1,-nbitq), 
to_sfixed(183525737.0/4294967296.0,1,-nbitq), 
to_sfixed(-69371171.0/4294967296.0,1,-nbitq), 
to_sfixed(-96599965.0/4294967296.0,1,-nbitq), 
to_sfixed(-8077703.0/4294967296.0,1,-nbitq), 
to_sfixed(-8698537.0/4294967296.0,1,-nbitq), 
to_sfixed(-225935538.0/4294967296.0,1,-nbitq), 
to_sfixed(-195829958.0/4294967296.0,1,-nbitq), 
to_sfixed(119858301.0/4294967296.0,1,-nbitq), 
to_sfixed(-232874273.0/4294967296.0,1,-nbitq), 
to_sfixed(66432278.0/4294967296.0,1,-nbitq), 
to_sfixed(-107763491.0/4294967296.0,1,-nbitq), 
to_sfixed(-265919186.0/4294967296.0,1,-nbitq), 
to_sfixed(159715445.0/4294967296.0,1,-nbitq), 
to_sfixed(6668884.0/4294967296.0,1,-nbitq), 
to_sfixed(-191142705.0/4294967296.0,1,-nbitq), 
to_sfixed(114941169.0/4294967296.0,1,-nbitq), 
to_sfixed(-684956510.0/4294967296.0,1,-nbitq), 
to_sfixed(-215761445.0/4294967296.0,1,-nbitq), 
to_sfixed(-325997962.0/4294967296.0,1,-nbitq), 
to_sfixed(-202145183.0/4294967296.0,1,-nbitq), 
to_sfixed(286240370.0/4294967296.0,1,-nbitq), 
to_sfixed(-429794030.0/4294967296.0,1,-nbitq), 
to_sfixed(94375040.0/4294967296.0,1,-nbitq), 
to_sfixed(-80735095.0/4294967296.0,1,-nbitq), 
to_sfixed(497883403.0/4294967296.0,1,-nbitq), 
to_sfixed(339392425.0/4294967296.0,1,-nbitq), 
to_sfixed(33423030.0/4294967296.0,1,-nbitq), 
to_sfixed(65498404.0/4294967296.0,1,-nbitq), 
to_sfixed(168283393.0/4294967296.0,1,-nbitq), 
to_sfixed(98378278.0/4294967296.0,1,-nbitq), 
to_sfixed(101333620.0/4294967296.0,1,-nbitq), 
to_sfixed(-459463419.0/4294967296.0,1,-nbitq), 
to_sfixed(289138546.0/4294967296.0,1,-nbitq), 
to_sfixed(-162669563.0/4294967296.0,1,-nbitq), 
to_sfixed(-76743031.0/4294967296.0,1,-nbitq), 
to_sfixed(165279125.0/4294967296.0,1,-nbitq), 
to_sfixed(-350069112.0/4294967296.0,1,-nbitq), 
to_sfixed(-494953050.0/4294967296.0,1,-nbitq), 
to_sfixed(-278798726.0/4294967296.0,1,-nbitq), 
to_sfixed(-365899734.0/4294967296.0,1,-nbitq), 
to_sfixed(165790256.0/4294967296.0,1,-nbitq), 
to_sfixed(349082922.0/4294967296.0,1,-nbitq), 
to_sfixed(-179508954.0/4294967296.0,1,-nbitq), 
to_sfixed(297004384.0/4294967296.0,1,-nbitq), 
to_sfixed(267715302.0/4294967296.0,1,-nbitq), 
to_sfixed(-304097741.0/4294967296.0,1,-nbitq), 
to_sfixed(-39248136.0/4294967296.0,1,-nbitq), 
to_sfixed(176206150.0/4294967296.0,1,-nbitq), 
to_sfixed(-256877600.0/4294967296.0,1,-nbitq), 
to_sfixed(-180879621.0/4294967296.0,1,-nbitq), 
to_sfixed(-428841991.0/4294967296.0,1,-nbitq), 
to_sfixed(-283148195.0/4294967296.0,1,-nbitq), 
to_sfixed(-98904295.0/4294967296.0,1,-nbitq), 
to_sfixed(-17432275.0/4294967296.0,1,-nbitq), 
to_sfixed(39679987.0/4294967296.0,1,-nbitq), 
to_sfixed(523744964.0/4294967296.0,1,-nbitq), 
to_sfixed(305146797.0/4294967296.0,1,-nbitq), 
to_sfixed(12612963.0/4294967296.0,1,-nbitq), 
to_sfixed(-170658329.0/4294967296.0,1,-nbitq), 
to_sfixed(108640608.0/4294967296.0,1,-nbitq), 
to_sfixed(267925437.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(309358827.0/4294967296.0,1,-nbitq), 
to_sfixed(251311763.0/4294967296.0,1,-nbitq), 
to_sfixed(318762381.0/4294967296.0,1,-nbitq), 
to_sfixed(-7604732.0/4294967296.0,1,-nbitq), 
to_sfixed(-358106947.0/4294967296.0,1,-nbitq), 
to_sfixed(-300097134.0/4294967296.0,1,-nbitq), 
to_sfixed(-22034430.0/4294967296.0,1,-nbitq), 
to_sfixed(-344785150.0/4294967296.0,1,-nbitq), 
to_sfixed(103855072.0/4294967296.0,1,-nbitq), 
to_sfixed(-167986020.0/4294967296.0,1,-nbitq), 
to_sfixed(35907147.0/4294967296.0,1,-nbitq), 
to_sfixed(452710834.0/4294967296.0,1,-nbitq), 
to_sfixed(-513140090.0/4294967296.0,1,-nbitq), 
to_sfixed(527102692.0/4294967296.0,1,-nbitq), 
to_sfixed(-170214757.0/4294967296.0,1,-nbitq), 
to_sfixed(-481885894.0/4294967296.0,1,-nbitq), 
to_sfixed(218512611.0/4294967296.0,1,-nbitq), 
to_sfixed(-90784046.0/4294967296.0,1,-nbitq), 
to_sfixed(-169423301.0/4294967296.0,1,-nbitq), 
to_sfixed(324270643.0/4294967296.0,1,-nbitq), 
to_sfixed(343260597.0/4294967296.0,1,-nbitq), 
to_sfixed(-11362369.0/4294967296.0,1,-nbitq), 
to_sfixed(268186081.0/4294967296.0,1,-nbitq), 
to_sfixed(-1805492.0/4294967296.0,1,-nbitq), 
to_sfixed(-59412192.0/4294967296.0,1,-nbitq), 
to_sfixed(-176616774.0/4294967296.0,1,-nbitq), 
to_sfixed(-149287872.0/4294967296.0,1,-nbitq), 
to_sfixed(71748699.0/4294967296.0,1,-nbitq), 
to_sfixed(-250385969.0/4294967296.0,1,-nbitq), 
to_sfixed(-44740995.0/4294967296.0,1,-nbitq), 
to_sfixed(98337615.0/4294967296.0,1,-nbitq), 
to_sfixed(-239164775.0/4294967296.0,1,-nbitq), 
to_sfixed(242902954.0/4294967296.0,1,-nbitq), 
to_sfixed(-197551349.0/4294967296.0,1,-nbitq), 
to_sfixed(-39430422.0/4294967296.0,1,-nbitq), 
to_sfixed(-490129126.0/4294967296.0,1,-nbitq), 
to_sfixed(-114709785.0/4294967296.0,1,-nbitq), 
to_sfixed(88813851.0/4294967296.0,1,-nbitq), 
to_sfixed(354690816.0/4294967296.0,1,-nbitq), 
to_sfixed(-239658599.0/4294967296.0,1,-nbitq), 
to_sfixed(-363439016.0/4294967296.0,1,-nbitq), 
to_sfixed(-5649837.0/4294967296.0,1,-nbitq), 
to_sfixed(-151189868.0/4294967296.0,1,-nbitq), 
to_sfixed(164459955.0/4294967296.0,1,-nbitq), 
to_sfixed(54695097.0/4294967296.0,1,-nbitq), 
to_sfixed(6284884.0/4294967296.0,1,-nbitq), 
to_sfixed(328597296.0/4294967296.0,1,-nbitq), 
to_sfixed(-77828207.0/4294967296.0,1,-nbitq), 
to_sfixed(522029186.0/4294967296.0,1,-nbitq), 
to_sfixed(-210299838.0/4294967296.0,1,-nbitq), 
to_sfixed(-465365517.0/4294967296.0,1,-nbitq), 
to_sfixed(85606285.0/4294967296.0,1,-nbitq), 
to_sfixed(-221016018.0/4294967296.0,1,-nbitq), 
to_sfixed(133740862.0/4294967296.0,1,-nbitq), 
to_sfixed(127876308.0/4294967296.0,1,-nbitq), 
to_sfixed(72364618.0/4294967296.0,1,-nbitq), 
to_sfixed(107174862.0/4294967296.0,1,-nbitq), 
to_sfixed(-142404554.0/4294967296.0,1,-nbitq), 
to_sfixed(298469328.0/4294967296.0,1,-nbitq), 
to_sfixed(111702935.0/4294967296.0,1,-nbitq), 
to_sfixed(-410954221.0/4294967296.0,1,-nbitq), 
to_sfixed(375363770.0/4294967296.0,1,-nbitq), 
to_sfixed(107729484.0/4294967296.0,1,-nbitq), 
to_sfixed(-376984208.0/4294967296.0,1,-nbitq), 
to_sfixed(231719500.0/4294967296.0,1,-nbitq), 
to_sfixed(-460242927.0/4294967296.0,1,-nbitq), 
to_sfixed(573565743.0/4294967296.0,1,-nbitq), 
to_sfixed(80828605.0/4294967296.0,1,-nbitq), 
to_sfixed(-161103079.0/4294967296.0,1,-nbitq), 
to_sfixed(99421433.0/4294967296.0,1,-nbitq), 
to_sfixed(-290197362.0/4294967296.0,1,-nbitq), 
to_sfixed(-160925775.0/4294967296.0,1,-nbitq), 
to_sfixed(114211255.0/4294967296.0,1,-nbitq), 
to_sfixed(-41615517.0/4294967296.0,1,-nbitq), 
to_sfixed(281890285.0/4294967296.0,1,-nbitq), 
to_sfixed(-107377376.0/4294967296.0,1,-nbitq), 
to_sfixed(-407314178.0/4294967296.0,1,-nbitq), 
to_sfixed(220805486.0/4294967296.0,1,-nbitq), 
to_sfixed(237496351.0/4294967296.0,1,-nbitq), 
to_sfixed(305385520.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-5717611.0/4294967296.0,1,-nbitq), 
to_sfixed(323091227.0/4294967296.0,1,-nbitq), 
to_sfixed(208421153.0/4294967296.0,1,-nbitq), 
to_sfixed(-196219864.0/4294967296.0,1,-nbitq), 
to_sfixed(123196272.0/4294967296.0,1,-nbitq), 
to_sfixed(-72383765.0/4294967296.0,1,-nbitq), 
to_sfixed(280804141.0/4294967296.0,1,-nbitq), 
to_sfixed(-144364573.0/4294967296.0,1,-nbitq), 
to_sfixed(380940619.0/4294967296.0,1,-nbitq), 
to_sfixed(145190667.0/4294967296.0,1,-nbitq), 
to_sfixed(272925311.0/4294967296.0,1,-nbitq), 
to_sfixed(-162203361.0/4294967296.0,1,-nbitq), 
to_sfixed(-343772876.0/4294967296.0,1,-nbitq), 
to_sfixed(386095631.0/4294967296.0,1,-nbitq), 
to_sfixed(-95799449.0/4294967296.0,1,-nbitq), 
to_sfixed(-350671708.0/4294967296.0,1,-nbitq), 
to_sfixed(-284337653.0/4294967296.0,1,-nbitq), 
to_sfixed(264169067.0/4294967296.0,1,-nbitq), 
to_sfixed(135996615.0/4294967296.0,1,-nbitq), 
to_sfixed(230220281.0/4294967296.0,1,-nbitq), 
to_sfixed(371583904.0/4294967296.0,1,-nbitq), 
to_sfixed(269524523.0/4294967296.0,1,-nbitq), 
to_sfixed(292104883.0/4294967296.0,1,-nbitq), 
to_sfixed(-288460697.0/4294967296.0,1,-nbitq), 
to_sfixed(27384657.0/4294967296.0,1,-nbitq), 
to_sfixed(-130067815.0/4294967296.0,1,-nbitq), 
to_sfixed(-249478975.0/4294967296.0,1,-nbitq), 
to_sfixed(-623243257.0/4294967296.0,1,-nbitq), 
to_sfixed(-201694398.0/4294967296.0,1,-nbitq), 
to_sfixed(387125855.0/4294967296.0,1,-nbitq), 
to_sfixed(194311549.0/4294967296.0,1,-nbitq), 
to_sfixed(-514120202.0/4294967296.0,1,-nbitq), 
to_sfixed(153335012.0/4294967296.0,1,-nbitq), 
to_sfixed(52247026.0/4294967296.0,1,-nbitq), 
to_sfixed(558274271.0/4294967296.0,1,-nbitq), 
to_sfixed(-544354492.0/4294967296.0,1,-nbitq), 
to_sfixed(-273546812.0/4294967296.0,1,-nbitq), 
to_sfixed(-92933551.0/4294967296.0,1,-nbitq), 
to_sfixed(-221083909.0/4294967296.0,1,-nbitq), 
to_sfixed(329460469.0/4294967296.0,1,-nbitq), 
to_sfixed(137082095.0/4294967296.0,1,-nbitq), 
to_sfixed(-188206593.0/4294967296.0,1,-nbitq), 
to_sfixed(246344520.0/4294967296.0,1,-nbitq), 
to_sfixed(312335046.0/4294967296.0,1,-nbitq), 
to_sfixed(-204275702.0/4294967296.0,1,-nbitq), 
to_sfixed(-29325890.0/4294967296.0,1,-nbitq), 
to_sfixed(-333050556.0/4294967296.0,1,-nbitq), 
to_sfixed(-402797139.0/4294967296.0,1,-nbitq), 
to_sfixed(-296568751.0/4294967296.0,1,-nbitq), 
to_sfixed(372587467.0/4294967296.0,1,-nbitq), 
to_sfixed(-483973297.0/4294967296.0,1,-nbitq), 
to_sfixed(-246759077.0/4294967296.0,1,-nbitq), 
to_sfixed(-520588511.0/4294967296.0,1,-nbitq), 
to_sfixed(171707876.0/4294967296.0,1,-nbitq), 
to_sfixed(174750059.0/4294967296.0,1,-nbitq), 
to_sfixed(-91408342.0/4294967296.0,1,-nbitq), 
to_sfixed(-125307836.0/4294967296.0,1,-nbitq), 
to_sfixed(-361949230.0/4294967296.0,1,-nbitq), 
to_sfixed(224321672.0/4294967296.0,1,-nbitq), 
to_sfixed(292051775.0/4294967296.0,1,-nbitq), 
to_sfixed(-206631031.0/4294967296.0,1,-nbitq), 
to_sfixed(-211830849.0/4294967296.0,1,-nbitq), 
to_sfixed(-158984392.0/4294967296.0,1,-nbitq), 
to_sfixed(-83786899.0/4294967296.0,1,-nbitq), 
to_sfixed(-95088994.0/4294967296.0,1,-nbitq), 
to_sfixed(-394517777.0/4294967296.0,1,-nbitq), 
to_sfixed(334114102.0/4294967296.0,1,-nbitq), 
to_sfixed(377989771.0/4294967296.0,1,-nbitq), 
to_sfixed(146695093.0/4294967296.0,1,-nbitq), 
to_sfixed(-475971505.0/4294967296.0,1,-nbitq), 
to_sfixed(-184411157.0/4294967296.0,1,-nbitq), 
to_sfixed(-66567737.0/4294967296.0,1,-nbitq), 
to_sfixed(-302994283.0/4294967296.0,1,-nbitq), 
to_sfixed(-172714739.0/4294967296.0,1,-nbitq), 
to_sfixed(497556300.0/4294967296.0,1,-nbitq), 
to_sfixed(290583876.0/4294967296.0,1,-nbitq), 
to_sfixed(-94989894.0/4294967296.0,1,-nbitq), 
to_sfixed(191040346.0/4294967296.0,1,-nbitq), 
to_sfixed(-474970220.0/4294967296.0,1,-nbitq), 
to_sfixed(-105382563.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-38985429.0/4294967296.0,1,-nbitq), 
to_sfixed(-360598701.0/4294967296.0,1,-nbitq), 
to_sfixed(352007537.0/4294967296.0,1,-nbitq), 
to_sfixed(-289090253.0/4294967296.0,1,-nbitq), 
to_sfixed(-192897247.0/4294967296.0,1,-nbitq), 
to_sfixed(203698413.0/4294967296.0,1,-nbitq), 
to_sfixed(-327090962.0/4294967296.0,1,-nbitq), 
to_sfixed(-234714695.0/4294967296.0,1,-nbitq), 
to_sfixed(-186163989.0/4294967296.0,1,-nbitq), 
to_sfixed(-283907335.0/4294967296.0,1,-nbitq), 
to_sfixed(-405270541.0/4294967296.0,1,-nbitq), 
to_sfixed(302902349.0/4294967296.0,1,-nbitq), 
to_sfixed(-390395525.0/4294967296.0,1,-nbitq), 
to_sfixed(471326545.0/4294967296.0,1,-nbitq), 
to_sfixed(-132233865.0/4294967296.0,1,-nbitq), 
to_sfixed(194172332.0/4294967296.0,1,-nbitq), 
to_sfixed(-94176747.0/4294967296.0,1,-nbitq), 
to_sfixed(14411213.0/4294967296.0,1,-nbitq), 
to_sfixed(-186354546.0/4294967296.0,1,-nbitq), 
to_sfixed(-318766596.0/4294967296.0,1,-nbitq), 
to_sfixed(114200937.0/4294967296.0,1,-nbitq), 
to_sfixed(76854954.0/4294967296.0,1,-nbitq), 
to_sfixed(432205629.0/4294967296.0,1,-nbitq), 
to_sfixed(175032952.0/4294967296.0,1,-nbitq), 
to_sfixed(66123728.0/4294967296.0,1,-nbitq), 
to_sfixed(22543364.0/4294967296.0,1,-nbitq), 
to_sfixed(188293107.0/4294967296.0,1,-nbitq), 
to_sfixed(-272315202.0/4294967296.0,1,-nbitq), 
to_sfixed(96351036.0/4294967296.0,1,-nbitq), 
to_sfixed(-136451777.0/4294967296.0,1,-nbitq), 
to_sfixed(-374934459.0/4294967296.0,1,-nbitq), 
to_sfixed(-209825692.0/4294967296.0,1,-nbitq), 
to_sfixed(29262248.0/4294967296.0,1,-nbitq), 
to_sfixed(106531132.0/4294967296.0,1,-nbitq), 
to_sfixed(399807571.0/4294967296.0,1,-nbitq), 
to_sfixed(-448602788.0/4294967296.0,1,-nbitq), 
to_sfixed(-27735814.0/4294967296.0,1,-nbitq), 
to_sfixed(163382397.0/4294967296.0,1,-nbitq), 
to_sfixed(234112134.0/4294967296.0,1,-nbitq), 
to_sfixed(-16054077.0/4294967296.0,1,-nbitq), 
to_sfixed(-53626258.0/4294967296.0,1,-nbitq), 
to_sfixed(92024386.0/4294967296.0,1,-nbitq), 
to_sfixed(88839705.0/4294967296.0,1,-nbitq), 
to_sfixed(449387714.0/4294967296.0,1,-nbitq), 
to_sfixed(3613882.0/4294967296.0,1,-nbitq), 
to_sfixed(-201386859.0/4294967296.0,1,-nbitq), 
to_sfixed(-299724556.0/4294967296.0,1,-nbitq), 
to_sfixed(-342372043.0/4294967296.0,1,-nbitq), 
to_sfixed(-344689801.0/4294967296.0,1,-nbitq), 
to_sfixed(-237329963.0/4294967296.0,1,-nbitq), 
to_sfixed(-175431840.0/4294967296.0,1,-nbitq), 
to_sfixed(-206800307.0/4294967296.0,1,-nbitq), 
to_sfixed(17137711.0/4294967296.0,1,-nbitq), 
to_sfixed(27620817.0/4294967296.0,1,-nbitq), 
to_sfixed(484201358.0/4294967296.0,1,-nbitq), 
to_sfixed(-195510584.0/4294967296.0,1,-nbitq), 
to_sfixed(317015118.0/4294967296.0,1,-nbitq), 
to_sfixed(-70381410.0/4294967296.0,1,-nbitq), 
to_sfixed(-272326270.0/4294967296.0,1,-nbitq), 
to_sfixed(-306741285.0/4294967296.0,1,-nbitq), 
to_sfixed(-14533968.0/4294967296.0,1,-nbitq), 
to_sfixed(-226022366.0/4294967296.0,1,-nbitq), 
to_sfixed(-225461689.0/4294967296.0,1,-nbitq), 
to_sfixed(308644381.0/4294967296.0,1,-nbitq), 
to_sfixed(-218527143.0/4294967296.0,1,-nbitq), 
to_sfixed(68279813.0/4294967296.0,1,-nbitq), 
to_sfixed(371733246.0/4294967296.0,1,-nbitq), 
to_sfixed(9469020.0/4294967296.0,1,-nbitq), 
to_sfixed(119462682.0/4294967296.0,1,-nbitq), 
to_sfixed(-96080688.0/4294967296.0,1,-nbitq), 
to_sfixed(124208517.0/4294967296.0,1,-nbitq), 
to_sfixed(-212527376.0/4294967296.0,1,-nbitq), 
to_sfixed(35903479.0/4294967296.0,1,-nbitq), 
to_sfixed(-106368535.0/4294967296.0,1,-nbitq), 
to_sfixed(415722167.0/4294967296.0,1,-nbitq), 
to_sfixed(41039081.0/4294967296.0,1,-nbitq), 
to_sfixed(10496661.0/4294967296.0,1,-nbitq), 
to_sfixed(-397185890.0/4294967296.0,1,-nbitq), 
to_sfixed(-355286314.0/4294967296.0,1,-nbitq), 
to_sfixed(318611691.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-339522050.0/4294967296.0,1,-nbitq), 
to_sfixed(-563647694.0/4294967296.0,1,-nbitq), 
to_sfixed(61660309.0/4294967296.0,1,-nbitq), 
to_sfixed(-257463905.0/4294967296.0,1,-nbitq), 
to_sfixed(338750556.0/4294967296.0,1,-nbitq), 
to_sfixed(96643661.0/4294967296.0,1,-nbitq), 
to_sfixed(-275257444.0/4294967296.0,1,-nbitq), 
to_sfixed(-42936410.0/4294967296.0,1,-nbitq), 
to_sfixed(-180525422.0/4294967296.0,1,-nbitq), 
to_sfixed(54588264.0/4294967296.0,1,-nbitq), 
to_sfixed(167389607.0/4294967296.0,1,-nbitq), 
to_sfixed(192357991.0/4294967296.0,1,-nbitq), 
to_sfixed(-518291535.0/4294967296.0,1,-nbitq), 
to_sfixed(110370668.0/4294967296.0,1,-nbitq), 
to_sfixed(-234239300.0/4294967296.0,1,-nbitq), 
to_sfixed(-364484576.0/4294967296.0,1,-nbitq), 
to_sfixed(205828329.0/4294967296.0,1,-nbitq), 
to_sfixed(-46211122.0/4294967296.0,1,-nbitq), 
to_sfixed(-374262050.0/4294967296.0,1,-nbitq), 
to_sfixed(-290491877.0/4294967296.0,1,-nbitq), 
to_sfixed(223156134.0/4294967296.0,1,-nbitq), 
to_sfixed(-146611411.0/4294967296.0,1,-nbitq), 
to_sfixed(389025028.0/4294967296.0,1,-nbitq), 
to_sfixed(-391317517.0/4294967296.0,1,-nbitq), 
to_sfixed(397659605.0/4294967296.0,1,-nbitq), 
to_sfixed(188434892.0/4294967296.0,1,-nbitq), 
to_sfixed(346827861.0/4294967296.0,1,-nbitq), 
to_sfixed(-142835089.0/4294967296.0,1,-nbitq), 
to_sfixed(-74626285.0/4294967296.0,1,-nbitq), 
to_sfixed(22332905.0/4294967296.0,1,-nbitq), 
to_sfixed(-260781660.0/4294967296.0,1,-nbitq), 
to_sfixed(156079249.0/4294967296.0,1,-nbitq), 
to_sfixed(213824753.0/4294967296.0,1,-nbitq), 
to_sfixed(-102107271.0/4294967296.0,1,-nbitq), 
to_sfixed(464591115.0/4294967296.0,1,-nbitq), 
to_sfixed(-367719664.0/4294967296.0,1,-nbitq), 
to_sfixed(-17125558.0/4294967296.0,1,-nbitq), 
to_sfixed(-270952327.0/4294967296.0,1,-nbitq), 
to_sfixed(-140502211.0/4294967296.0,1,-nbitq), 
to_sfixed(275426133.0/4294967296.0,1,-nbitq), 
to_sfixed(-143769559.0/4294967296.0,1,-nbitq), 
to_sfixed(41780209.0/4294967296.0,1,-nbitq), 
to_sfixed(107403982.0/4294967296.0,1,-nbitq), 
to_sfixed(371048386.0/4294967296.0,1,-nbitq), 
to_sfixed(-144197597.0/4294967296.0,1,-nbitq), 
to_sfixed(360021405.0/4294967296.0,1,-nbitq), 
to_sfixed(2565663.0/4294967296.0,1,-nbitq), 
to_sfixed(-148283982.0/4294967296.0,1,-nbitq), 
to_sfixed(155408699.0/4294967296.0,1,-nbitq), 
to_sfixed(-84780832.0/4294967296.0,1,-nbitq), 
to_sfixed(391969499.0/4294967296.0,1,-nbitq), 
to_sfixed(139450365.0/4294967296.0,1,-nbitq), 
to_sfixed(-203220863.0/4294967296.0,1,-nbitq), 
to_sfixed(342831768.0/4294967296.0,1,-nbitq), 
to_sfixed(344789881.0/4294967296.0,1,-nbitq), 
to_sfixed(62945826.0/4294967296.0,1,-nbitq), 
to_sfixed(-148753544.0/4294967296.0,1,-nbitq), 
to_sfixed(53783882.0/4294967296.0,1,-nbitq), 
to_sfixed(-100546498.0/4294967296.0,1,-nbitq), 
to_sfixed(364640400.0/4294967296.0,1,-nbitq), 
to_sfixed(-269006860.0/4294967296.0,1,-nbitq), 
to_sfixed(391094021.0/4294967296.0,1,-nbitq), 
to_sfixed(-25489221.0/4294967296.0,1,-nbitq), 
to_sfixed(93885796.0/4294967296.0,1,-nbitq), 
to_sfixed(-23058964.0/4294967296.0,1,-nbitq), 
to_sfixed(-33095603.0/4294967296.0,1,-nbitq), 
to_sfixed(72647530.0/4294967296.0,1,-nbitq), 
to_sfixed(-317243556.0/4294967296.0,1,-nbitq), 
to_sfixed(417093223.0/4294967296.0,1,-nbitq), 
to_sfixed(510881199.0/4294967296.0,1,-nbitq), 
to_sfixed(128348996.0/4294967296.0,1,-nbitq), 
to_sfixed(-71826158.0/4294967296.0,1,-nbitq), 
to_sfixed(-25885487.0/4294967296.0,1,-nbitq), 
to_sfixed(-198051701.0/4294967296.0,1,-nbitq), 
to_sfixed(-112018225.0/4294967296.0,1,-nbitq), 
to_sfixed(89563105.0/4294967296.0,1,-nbitq), 
to_sfixed(444172255.0/4294967296.0,1,-nbitq), 
to_sfixed(250350430.0/4294967296.0,1,-nbitq), 
to_sfixed(-505373078.0/4294967296.0,1,-nbitq), 
to_sfixed(20055071.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-176988216.0/4294967296.0,1,-nbitq), 
to_sfixed(-379984375.0/4294967296.0,1,-nbitq), 
to_sfixed(-36304716.0/4294967296.0,1,-nbitq), 
to_sfixed(395975340.0/4294967296.0,1,-nbitq), 
to_sfixed(-204614446.0/4294967296.0,1,-nbitq), 
to_sfixed(394484436.0/4294967296.0,1,-nbitq), 
to_sfixed(166938109.0/4294967296.0,1,-nbitq), 
to_sfixed(14493202.0/4294967296.0,1,-nbitq), 
to_sfixed(245565650.0/4294967296.0,1,-nbitq), 
to_sfixed(143263104.0/4294967296.0,1,-nbitq), 
to_sfixed(334881409.0/4294967296.0,1,-nbitq), 
to_sfixed(271589995.0/4294967296.0,1,-nbitq), 
to_sfixed(-301176464.0/4294967296.0,1,-nbitq), 
to_sfixed(-285991268.0/4294967296.0,1,-nbitq), 
to_sfixed(342487402.0/4294967296.0,1,-nbitq), 
to_sfixed(-263871625.0/4294967296.0,1,-nbitq), 
to_sfixed(-93837683.0/4294967296.0,1,-nbitq), 
to_sfixed(-34678697.0/4294967296.0,1,-nbitq), 
to_sfixed(112205709.0/4294967296.0,1,-nbitq), 
to_sfixed(226543011.0/4294967296.0,1,-nbitq), 
to_sfixed(-72547922.0/4294967296.0,1,-nbitq), 
to_sfixed(438085860.0/4294967296.0,1,-nbitq), 
to_sfixed(167392314.0/4294967296.0,1,-nbitq), 
to_sfixed(58024030.0/4294967296.0,1,-nbitq), 
to_sfixed(48411055.0/4294967296.0,1,-nbitq), 
to_sfixed(313587114.0/4294967296.0,1,-nbitq), 
to_sfixed(-96724084.0/4294967296.0,1,-nbitq), 
to_sfixed(-487680040.0/4294967296.0,1,-nbitq), 
to_sfixed(-147690787.0/4294967296.0,1,-nbitq), 
to_sfixed(-57979765.0/4294967296.0,1,-nbitq), 
to_sfixed(-191979459.0/4294967296.0,1,-nbitq), 
to_sfixed(-389525365.0/4294967296.0,1,-nbitq), 
to_sfixed(113572592.0/4294967296.0,1,-nbitq), 
to_sfixed(83372039.0/4294967296.0,1,-nbitq), 
to_sfixed(19268366.0/4294967296.0,1,-nbitq), 
to_sfixed(340569352.0/4294967296.0,1,-nbitq), 
to_sfixed(374235527.0/4294967296.0,1,-nbitq), 
to_sfixed(44049598.0/4294967296.0,1,-nbitq), 
to_sfixed(286269631.0/4294967296.0,1,-nbitq), 
to_sfixed(134382859.0/4294967296.0,1,-nbitq), 
to_sfixed(-133121129.0/4294967296.0,1,-nbitq), 
to_sfixed(335585227.0/4294967296.0,1,-nbitq), 
to_sfixed(10837507.0/4294967296.0,1,-nbitq), 
to_sfixed(-131629110.0/4294967296.0,1,-nbitq), 
to_sfixed(364804457.0/4294967296.0,1,-nbitq), 
to_sfixed(305887276.0/4294967296.0,1,-nbitq), 
to_sfixed(292915928.0/4294967296.0,1,-nbitq), 
to_sfixed(-208591893.0/4294967296.0,1,-nbitq), 
to_sfixed(330285330.0/4294967296.0,1,-nbitq), 
to_sfixed(-231452476.0/4294967296.0,1,-nbitq), 
to_sfixed(-343487525.0/4294967296.0,1,-nbitq), 
to_sfixed(10380474.0/4294967296.0,1,-nbitq), 
to_sfixed(-31068586.0/4294967296.0,1,-nbitq), 
to_sfixed(-14830416.0/4294967296.0,1,-nbitq), 
to_sfixed(-157257373.0/4294967296.0,1,-nbitq), 
to_sfixed(-200097677.0/4294967296.0,1,-nbitq), 
to_sfixed(-106857097.0/4294967296.0,1,-nbitq), 
to_sfixed(-409392174.0/4294967296.0,1,-nbitq), 
to_sfixed(-35746562.0/4294967296.0,1,-nbitq), 
to_sfixed(142866254.0/4294967296.0,1,-nbitq), 
to_sfixed(292248711.0/4294967296.0,1,-nbitq), 
to_sfixed(304089892.0/4294967296.0,1,-nbitq), 
to_sfixed(-95915327.0/4294967296.0,1,-nbitq), 
to_sfixed(-311663320.0/4294967296.0,1,-nbitq), 
to_sfixed(397713037.0/4294967296.0,1,-nbitq), 
to_sfixed(-162023888.0/4294967296.0,1,-nbitq), 
to_sfixed(-26649412.0/4294967296.0,1,-nbitq), 
to_sfixed(-255355046.0/4294967296.0,1,-nbitq), 
to_sfixed(-282557928.0/4294967296.0,1,-nbitq), 
to_sfixed(-85676526.0/4294967296.0,1,-nbitq), 
to_sfixed(58158618.0/4294967296.0,1,-nbitq), 
to_sfixed(170481674.0/4294967296.0,1,-nbitq), 
to_sfixed(-138523383.0/4294967296.0,1,-nbitq), 
to_sfixed(360133550.0/4294967296.0,1,-nbitq), 
to_sfixed(-170618892.0/4294967296.0,1,-nbitq), 
to_sfixed(-36624031.0/4294967296.0,1,-nbitq), 
to_sfixed(28523304.0/4294967296.0,1,-nbitq), 
to_sfixed(-141908507.0/4294967296.0,1,-nbitq), 
to_sfixed(-370095786.0/4294967296.0,1,-nbitq), 
to_sfixed(129973037.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-213329832.0/4294967296.0,1,-nbitq), 
to_sfixed(-213446823.0/4294967296.0,1,-nbitq), 
to_sfixed(80678527.0/4294967296.0,1,-nbitq), 
to_sfixed(124685848.0/4294967296.0,1,-nbitq), 
to_sfixed(111162376.0/4294967296.0,1,-nbitq), 
to_sfixed(289148794.0/4294967296.0,1,-nbitq), 
to_sfixed(313391804.0/4294967296.0,1,-nbitq), 
to_sfixed(-23936608.0/4294967296.0,1,-nbitq), 
to_sfixed(-356304205.0/4294967296.0,1,-nbitq), 
to_sfixed(262038116.0/4294967296.0,1,-nbitq), 
to_sfixed(-400757076.0/4294967296.0,1,-nbitq), 
to_sfixed(243031947.0/4294967296.0,1,-nbitq), 
to_sfixed(-346979689.0/4294967296.0,1,-nbitq), 
to_sfixed(184783344.0/4294967296.0,1,-nbitq), 
to_sfixed(-26144435.0/4294967296.0,1,-nbitq), 
to_sfixed(-109344590.0/4294967296.0,1,-nbitq), 
to_sfixed(-392450619.0/4294967296.0,1,-nbitq), 
to_sfixed(121509628.0/4294967296.0,1,-nbitq), 
to_sfixed(25243656.0/4294967296.0,1,-nbitq), 
to_sfixed(-209475237.0/4294967296.0,1,-nbitq), 
to_sfixed(217150305.0/4294967296.0,1,-nbitq), 
to_sfixed(266863824.0/4294967296.0,1,-nbitq), 
to_sfixed(496630778.0/4294967296.0,1,-nbitq), 
to_sfixed(195712607.0/4294967296.0,1,-nbitq), 
to_sfixed(-13637486.0/4294967296.0,1,-nbitq), 
to_sfixed(342504328.0/4294967296.0,1,-nbitq), 
to_sfixed(98589649.0/4294967296.0,1,-nbitq), 
to_sfixed(-351622101.0/4294967296.0,1,-nbitq), 
to_sfixed(331019412.0/4294967296.0,1,-nbitq), 
to_sfixed(229302533.0/4294967296.0,1,-nbitq), 
to_sfixed(-451093262.0/4294967296.0,1,-nbitq), 
to_sfixed(-157152654.0/4294967296.0,1,-nbitq), 
to_sfixed(-61298593.0/4294967296.0,1,-nbitq), 
to_sfixed(-511805749.0/4294967296.0,1,-nbitq), 
to_sfixed(159929401.0/4294967296.0,1,-nbitq), 
to_sfixed(62272626.0/4294967296.0,1,-nbitq), 
to_sfixed(241114347.0/4294967296.0,1,-nbitq), 
to_sfixed(100780710.0/4294967296.0,1,-nbitq), 
to_sfixed(-21188700.0/4294967296.0,1,-nbitq), 
to_sfixed(-155076669.0/4294967296.0,1,-nbitq), 
to_sfixed(6407538.0/4294967296.0,1,-nbitq), 
to_sfixed(-249221479.0/4294967296.0,1,-nbitq), 
to_sfixed(-115191212.0/4294967296.0,1,-nbitq), 
to_sfixed(-329536717.0/4294967296.0,1,-nbitq), 
to_sfixed(322037385.0/4294967296.0,1,-nbitq), 
to_sfixed(416175193.0/4294967296.0,1,-nbitq), 
to_sfixed(-339272392.0/4294967296.0,1,-nbitq), 
to_sfixed(224419245.0/4294967296.0,1,-nbitq), 
to_sfixed(-383420093.0/4294967296.0,1,-nbitq), 
to_sfixed(-72383115.0/4294967296.0,1,-nbitq), 
to_sfixed(-291290518.0/4294967296.0,1,-nbitq), 
to_sfixed(177449946.0/4294967296.0,1,-nbitq), 
to_sfixed(-92704256.0/4294967296.0,1,-nbitq), 
to_sfixed(14256606.0/4294967296.0,1,-nbitq), 
to_sfixed(288933255.0/4294967296.0,1,-nbitq), 
to_sfixed(-406336.0/4294967296.0,1,-nbitq), 
to_sfixed(427008458.0/4294967296.0,1,-nbitq), 
to_sfixed(39142122.0/4294967296.0,1,-nbitq), 
to_sfixed(-286787120.0/4294967296.0,1,-nbitq), 
to_sfixed(1163323.0/4294967296.0,1,-nbitq), 
to_sfixed(232089616.0/4294967296.0,1,-nbitq), 
to_sfixed(375985896.0/4294967296.0,1,-nbitq), 
to_sfixed(152439399.0/4294967296.0,1,-nbitq), 
to_sfixed(122790985.0/4294967296.0,1,-nbitq), 
to_sfixed(-35429066.0/4294967296.0,1,-nbitq), 
to_sfixed(-407868165.0/4294967296.0,1,-nbitq), 
to_sfixed(455388503.0/4294967296.0,1,-nbitq), 
to_sfixed(-360262795.0/4294967296.0,1,-nbitq), 
to_sfixed(43867582.0/4294967296.0,1,-nbitq), 
to_sfixed(10025517.0/4294967296.0,1,-nbitq), 
to_sfixed(-425075027.0/4294967296.0,1,-nbitq), 
to_sfixed(-323447715.0/4294967296.0,1,-nbitq), 
to_sfixed(-304925261.0/4294967296.0,1,-nbitq), 
to_sfixed(376455214.0/4294967296.0,1,-nbitq), 
to_sfixed(408976509.0/4294967296.0,1,-nbitq), 
to_sfixed(-461389640.0/4294967296.0,1,-nbitq), 
to_sfixed(-231908117.0/4294967296.0,1,-nbitq), 
to_sfixed(-187698793.0/4294967296.0,1,-nbitq), 
to_sfixed(-487853651.0/4294967296.0,1,-nbitq), 
to_sfixed(-372007032.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-39863313.0/4294967296.0,1,-nbitq), 
to_sfixed(-270738990.0/4294967296.0,1,-nbitq), 
to_sfixed(27163388.0/4294967296.0,1,-nbitq), 
to_sfixed(-9438293.0/4294967296.0,1,-nbitq), 
to_sfixed(65775378.0/4294967296.0,1,-nbitq), 
to_sfixed(237112028.0/4294967296.0,1,-nbitq), 
to_sfixed(115682533.0/4294967296.0,1,-nbitq), 
to_sfixed(-410817185.0/4294967296.0,1,-nbitq), 
to_sfixed(126663775.0/4294967296.0,1,-nbitq), 
to_sfixed(-220582365.0/4294967296.0,1,-nbitq), 
to_sfixed(-341655313.0/4294967296.0,1,-nbitq), 
to_sfixed(151214938.0/4294967296.0,1,-nbitq), 
to_sfixed(146226771.0/4294967296.0,1,-nbitq), 
to_sfixed(340873600.0/4294967296.0,1,-nbitq), 
to_sfixed(-230286500.0/4294967296.0,1,-nbitq), 
to_sfixed(-214588041.0/4294967296.0,1,-nbitq), 
to_sfixed(24834017.0/4294967296.0,1,-nbitq), 
to_sfixed(251239366.0/4294967296.0,1,-nbitq), 
to_sfixed(27349301.0/4294967296.0,1,-nbitq), 
to_sfixed(-359963088.0/4294967296.0,1,-nbitq), 
to_sfixed(-370232724.0/4294967296.0,1,-nbitq), 
to_sfixed(230163225.0/4294967296.0,1,-nbitq), 
to_sfixed(266595266.0/4294967296.0,1,-nbitq), 
to_sfixed(278697658.0/4294967296.0,1,-nbitq), 
to_sfixed(-311624788.0/4294967296.0,1,-nbitq), 
to_sfixed(-158155598.0/4294967296.0,1,-nbitq), 
to_sfixed(204374416.0/4294967296.0,1,-nbitq), 
to_sfixed(15200013.0/4294967296.0,1,-nbitq), 
to_sfixed(12189261.0/4294967296.0,1,-nbitq), 
to_sfixed(126066332.0/4294967296.0,1,-nbitq), 
to_sfixed(-302314308.0/4294967296.0,1,-nbitq), 
to_sfixed(-543232031.0/4294967296.0,1,-nbitq), 
to_sfixed(-9890943.0/4294967296.0,1,-nbitq), 
to_sfixed(-195430335.0/4294967296.0,1,-nbitq), 
to_sfixed(281823022.0/4294967296.0,1,-nbitq), 
to_sfixed(-7363503.0/4294967296.0,1,-nbitq), 
to_sfixed(-291168840.0/4294967296.0,1,-nbitq), 
to_sfixed(71660383.0/4294967296.0,1,-nbitq), 
to_sfixed(274729147.0/4294967296.0,1,-nbitq), 
to_sfixed(348346842.0/4294967296.0,1,-nbitq), 
to_sfixed(-43011052.0/4294967296.0,1,-nbitq), 
to_sfixed(304945599.0/4294967296.0,1,-nbitq), 
to_sfixed(5797925.0/4294967296.0,1,-nbitq), 
to_sfixed(227032028.0/4294967296.0,1,-nbitq), 
to_sfixed(130237877.0/4294967296.0,1,-nbitq), 
to_sfixed(354750537.0/4294967296.0,1,-nbitq), 
to_sfixed(-259446161.0/4294967296.0,1,-nbitq), 
to_sfixed(-468679878.0/4294967296.0,1,-nbitq), 
to_sfixed(-88465012.0/4294967296.0,1,-nbitq), 
to_sfixed(13639661.0/4294967296.0,1,-nbitq), 
to_sfixed(-23082561.0/4294967296.0,1,-nbitq), 
to_sfixed(76394068.0/4294967296.0,1,-nbitq), 
to_sfixed(-424483158.0/4294967296.0,1,-nbitq), 
to_sfixed(-251296152.0/4294967296.0,1,-nbitq), 
to_sfixed(71158644.0/4294967296.0,1,-nbitq), 
to_sfixed(180988009.0/4294967296.0,1,-nbitq), 
to_sfixed(111220346.0/4294967296.0,1,-nbitq), 
to_sfixed(-266781687.0/4294967296.0,1,-nbitq), 
to_sfixed(327597690.0/4294967296.0,1,-nbitq), 
to_sfixed(311855704.0/4294967296.0,1,-nbitq), 
to_sfixed(-258908843.0/4294967296.0,1,-nbitq), 
to_sfixed(72758793.0/4294967296.0,1,-nbitq), 
to_sfixed(267716948.0/4294967296.0,1,-nbitq), 
to_sfixed(-242647825.0/4294967296.0,1,-nbitq), 
to_sfixed(-147866069.0/4294967296.0,1,-nbitq), 
to_sfixed(232356611.0/4294967296.0,1,-nbitq), 
to_sfixed(373526931.0/4294967296.0,1,-nbitq), 
to_sfixed(350146860.0/4294967296.0,1,-nbitq), 
to_sfixed(-242708907.0/4294967296.0,1,-nbitq), 
to_sfixed(238888430.0/4294967296.0,1,-nbitq), 
to_sfixed(-444320588.0/4294967296.0,1,-nbitq), 
to_sfixed(-221471721.0/4294967296.0,1,-nbitq), 
to_sfixed(-139970501.0/4294967296.0,1,-nbitq), 
to_sfixed(-329485054.0/4294967296.0,1,-nbitq), 
to_sfixed(142877824.0/4294967296.0,1,-nbitq), 
to_sfixed(110408951.0/4294967296.0,1,-nbitq), 
to_sfixed(263422824.0/4294967296.0,1,-nbitq), 
to_sfixed(223774856.0/4294967296.0,1,-nbitq), 
to_sfixed(-90985024.0/4294967296.0,1,-nbitq), 
to_sfixed(-40836446.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-48263626.0/4294967296.0,1,-nbitq), 
to_sfixed(191292592.0/4294967296.0,1,-nbitq), 
to_sfixed(98377745.0/4294967296.0,1,-nbitq), 
to_sfixed(-357442878.0/4294967296.0,1,-nbitq), 
to_sfixed(-178254571.0/4294967296.0,1,-nbitq), 
to_sfixed(320057372.0/4294967296.0,1,-nbitq), 
to_sfixed(-323373892.0/4294967296.0,1,-nbitq), 
to_sfixed(-143862935.0/4294967296.0,1,-nbitq), 
to_sfixed(215339009.0/4294967296.0,1,-nbitq), 
to_sfixed(109078452.0/4294967296.0,1,-nbitq), 
to_sfixed(-86345587.0/4294967296.0,1,-nbitq), 
to_sfixed(85169727.0/4294967296.0,1,-nbitq), 
to_sfixed(286978752.0/4294967296.0,1,-nbitq), 
to_sfixed(20084313.0/4294967296.0,1,-nbitq), 
to_sfixed(-385091.0/4294967296.0,1,-nbitq), 
to_sfixed(337181372.0/4294967296.0,1,-nbitq), 
to_sfixed(-221843984.0/4294967296.0,1,-nbitq), 
to_sfixed(416924200.0/4294967296.0,1,-nbitq), 
to_sfixed(149625744.0/4294967296.0,1,-nbitq), 
to_sfixed(-397974459.0/4294967296.0,1,-nbitq), 
to_sfixed(315403532.0/4294967296.0,1,-nbitq), 
to_sfixed(-253316844.0/4294967296.0,1,-nbitq), 
to_sfixed(181321370.0/4294967296.0,1,-nbitq), 
to_sfixed(315013208.0/4294967296.0,1,-nbitq), 
to_sfixed(54282372.0/4294967296.0,1,-nbitq), 
to_sfixed(-68554868.0/4294967296.0,1,-nbitq), 
to_sfixed(-355301902.0/4294967296.0,1,-nbitq), 
to_sfixed(-262354193.0/4294967296.0,1,-nbitq), 
to_sfixed(400803929.0/4294967296.0,1,-nbitq), 
to_sfixed(336442559.0/4294967296.0,1,-nbitq), 
to_sfixed(-398577139.0/4294967296.0,1,-nbitq), 
to_sfixed(-210177722.0/4294967296.0,1,-nbitq), 
to_sfixed(-178079764.0/4294967296.0,1,-nbitq), 
to_sfixed(150695436.0/4294967296.0,1,-nbitq), 
to_sfixed(7750378.0/4294967296.0,1,-nbitq), 
to_sfixed(282256184.0/4294967296.0,1,-nbitq), 
to_sfixed(366689116.0/4294967296.0,1,-nbitq), 
to_sfixed(274356311.0/4294967296.0,1,-nbitq), 
to_sfixed(-263025960.0/4294967296.0,1,-nbitq), 
to_sfixed(-157424104.0/4294967296.0,1,-nbitq), 
to_sfixed(287510258.0/4294967296.0,1,-nbitq), 
to_sfixed(435756920.0/4294967296.0,1,-nbitq), 
to_sfixed(-399290839.0/4294967296.0,1,-nbitq), 
to_sfixed(157062098.0/4294967296.0,1,-nbitq), 
to_sfixed(106224116.0/4294967296.0,1,-nbitq), 
to_sfixed(-175572334.0/4294967296.0,1,-nbitq), 
to_sfixed(-431608546.0/4294967296.0,1,-nbitq), 
to_sfixed(-473895336.0/4294967296.0,1,-nbitq), 
to_sfixed(28463041.0/4294967296.0,1,-nbitq), 
to_sfixed(-191660608.0/4294967296.0,1,-nbitq), 
to_sfixed(-281088569.0/4294967296.0,1,-nbitq), 
to_sfixed(202205780.0/4294967296.0,1,-nbitq), 
to_sfixed(89184599.0/4294967296.0,1,-nbitq), 
to_sfixed(103063472.0/4294967296.0,1,-nbitq), 
to_sfixed(-165046175.0/4294967296.0,1,-nbitq), 
to_sfixed(-329688814.0/4294967296.0,1,-nbitq), 
to_sfixed(444016831.0/4294967296.0,1,-nbitq), 
to_sfixed(114645463.0/4294967296.0,1,-nbitq), 
to_sfixed(-332667204.0/4294967296.0,1,-nbitq), 
to_sfixed(120584559.0/4294967296.0,1,-nbitq), 
to_sfixed(-183305142.0/4294967296.0,1,-nbitq), 
to_sfixed(74500681.0/4294967296.0,1,-nbitq), 
to_sfixed(-174123626.0/4294967296.0,1,-nbitq), 
to_sfixed(52703409.0/4294967296.0,1,-nbitq), 
to_sfixed(443938522.0/4294967296.0,1,-nbitq), 
to_sfixed(188932989.0/4294967296.0,1,-nbitq), 
to_sfixed(292889927.0/4294967296.0,1,-nbitq), 
to_sfixed(217791985.0/4294967296.0,1,-nbitq), 
to_sfixed(435373749.0/4294967296.0,1,-nbitq), 
to_sfixed(175072644.0/4294967296.0,1,-nbitq), 
to_sfixed(101064655.0/4294967296.0,1,-nbitq), 
to_sfixed(334319260.0/4294967296.0,1,-nbitq), 
to_sfixed(-366325243.0/4294967296.0,1,-nbitq), 
to_sfixed(448176583.0/4294967296.0,1,-nbitq), 
to_sfixed(366602548.0/4294967296.0,1,-nbitq), 
to_sfixed(-193277146.0/4294967296.0,1,-nbitq), 
to_sfixed(292173169.0/4294967296.0,1,-nbitq), 
to_sfixed(200081988.0/4294967296.0,1,-nbitq), 
to_sfixed(44370004.0/4294967296.0,1,-nbitq), 
to_sfixed(290663661.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-102273549.0/4294967296.0,1,-nbitq), 
to_sfixed(-140098597.0/4294967296.0,1,-nbitq), 
to_sfixed(-11068568.0/4294967296.0,1,-nbitq), 
to_sfixed(-322236199.0/4294967296.0,1,-nbitq), 
to_sfixed(393490198.0/4294967296.0,1,-nbitq), 
to_sfixed(213384505.0/4294967296.0,1,-nbitq), 
to_sfixed(194847043.0/4294967296.0,1,-nbitq), 
to_sfixed(366491015.0/4294967296.0,1,-nbitq), 
to_sfixed(349727268.0/4294967296.0,1,-nbitq), 
to_sfixed(-128609364.0/4294967296.0,1,-nbitq), 
to_sfixed(317270949.0/4294967296.0,1,-nbitq), 
to_sfixed(212243703.0/4294967296.0,1,-nbitq), 
to_sfixed(33081476.0/4294967296.0,1,-nbitq), 
to_sfixed(449183748.0/4294967296.0,1,-nbitq), 
to_sfixed(-371235605.0/4294967296.0,1,-nbitq), 
to_sfixed(-321496144.0/4294967296.0,1,-nbitq), 
to_sfixed(206828072.0/4294967296.0,1,-nbitq), 
to_sfixed(320663693.0/4294967296.0,1,-nbitq), 
to_sfixed(132211408.0/4294967296.0,1,-nbitq), 
to_sfixed(-311599487.0/4294967296.0,1,-nbitq), 
to_sfixed(-344605861.0/4294967296.0,1,-nbitq), 
to_sfixed(-1126322.0/4294967296.0,1,-nbitq), 
to_sfixed(27879550.0/4294967296.0,1,-nbitq), 
to_sfixed(-141555008.0/4294967296.0,1,-nbitq), 
to_sfixed(-213499394.0/4294967296.0,1,-nbitq), 
to_sfixed(-147143001.0/4294967296.0,1,-nbitq), 
to_sfixed(316485140.0/4294967296.0,1,-nbitq), 
to_sfixed(-453412483.0/4294967296.0,1,-nbitq), 
to_sfixed(160554841.0/4294967296.0,1,-nbitq), 
to_sfixed(243178344.0/4294967296.0,1,-nbitq), 
to_sfixed(27932531.0/4294967296.0,1,-nbitq), 
to_sfixed(-345711343.0/4294967296.0,1,-nbitq), 
to_sfixed(324234587.0/4294967296.0,1,-nbitq), 
to_sfixed(216205739.0/4294967296.0,1,-nbitq), 
to_sfixed(-100023303.0/4294967296.0,1,-nbitq), 
to_sfixed(38599085.0/4294967296.0,1,-nbitq), 
to_sfixed(399201502.0/4294967296.0,1,-nbitq), 
to_sfixed(450568138.0/4294967296.0,1,-nbitq), 
to_sfixed(-20747389.0/4294967296.0,1,-nbitq), 
to_sfixed(-203771594.0/4294967296.0,1,-nbitq), 
to_sfixed(129887661.0/4294967296.0,1,-nbitq), 
to_sfixed(194917078.0/4294967296.0,1,-nbitq), 
to_sfixed(89698087.0/4294967296.0,1,-nbitq), 
to_sfixed(271212831.0/4294967296.0,1,-nbitq), 
to_sfixed(423957429.0/4294967296.0,1,-nbitq), 
to_sfixed(-10027328.0/4294967296.0,1,-nbitq), 
to_sfixed(84284089.0/4294967296.0,1,-nbitq), 
to_sfixed(-406559337.0/4294967296.0,1,-nbitq), 
to_sfixed(238838852.0/4294967296.0,1,-nbitq), 
to_sfixed(8616844.0/4294967296.0,1,-nbitq), 
to_sfixed(327822228.0/4294967296.0,1,-nbitq), 
to_sfixed(-91898956.0/4294967296.0,1,-nbitq), 
to_sfixed(-324558963.0/4294967296.0,1,-nbitq), 
to_sfixed(-128188384.0/4294967296.0,1,-nbitq), 
to_sfixed(100582671.0/4294967296.0,1,-nbitq), 
to_sfixed(536131788.0/4294967296.0,1,-nbitq), 
to_sfixed(387012159.0/4294967296.0,1,-nbitq), 
to_sfixed(-168754279.0/4294967296.0,1,-nbitq), 
to_sfixed(241540280.0/4294967296.0,1,-nbitq), 
to_sfixed(322068345.0/4294967296.0,1,-nbitq), 
to_sfixed(-66205281.0/4294967296.0,1,-nbitq), 
to_sfixed(-195786607.0/4294967296.0,1,-nbitq), 
to_sfixed(-362956101.0/4294967296.0,1,-nbitq), 
to_sfixed(-280376481.0/4294967296.0,1,-nbitq), 
to_sfixed(155862495.0/4294967296.0,1,-nbitq), 
to_sfixed(52747114.0/4294967296.0,1,-nbitq), 
to_sfixed(597504103.0/4294967296.0,1,-nbitq), 
to_sfixed(-227348176.0/4294967296.0,1,-nbitq), 
to_sfixed(385543662.0/4294967296.0,1,-nbitq), 
to_sfixed(109394971.0/4294967296.0,1,-nbitq), 
to_sfixed(256016202.0/4294967296.0,1,-nbitq), 
to_sfixed(-21456696.0/4294967296.0,1,-nbitq), 
to_sfixed(-71867367.0/4294967296.0,1,-nbitq), 
to_sfixed(-314542822.0/4294967296.0,1,-nbitq), 
to_sfixed(306476838.0/4294967296.0,1,-nbitq), 
to_sfixed(-293534748.0/4294967296.0,1,-nbitq), 
to_sfixed(-19361745.0/4294967296.0,1,-nbitq), 
to_sfixed(38315997.0/4294967296.0,1,-nbitq), 
to_sfixed(14916181.0/4294967296.0,1,-nbitq), 
to_sfixed(-236362436.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(330796707.0/4294967296.0,1,-nbitq), 
to_sfixed(-52454186.0/4294967296.0,1,-nbitq), 
to_sfixed(-218461157.0/4294967296.0,1,-nbitq), 
to_sfixed(-319040320.0/4294967296.0,1,-nbitq), 
to_sfixed(-69228243.0/4294967296.0,1,-nbitq), 
to_sfixed(322487613.0/4294967296.0,1,-nbitq), 
to_sfixed(196119398.0/4294967296.0,1,-nbitq), 
to_sfixed(68778981.0/4294967296.0,1,-nbitq), 
to_sfixed(101647985.0/4294967296.0,1,-nbitq), 
to_sfixed(196148090.0/4294967296.0,1,-nbitq), 
to_sfixed(-8420728.0/4294967296.0,1,-nbitq), 
to_sfixed(249153625.0/4294967296.0,1,-nbitq), 
to_sfixed(-231809167.0/4294967296.0,1,-nbitq), 
to_sfixed(225636881.0/4294967296.0,1,-nbitq), 
to_sfixed(226235119.0/4294967296.0,1,-nbitq), 
to_sfixed(-235958734.0/4294967296.0,1,-nbitq), 
to_sfixed(333306453.0/4294967296.0,1,-nbitq), 
to_sfixed(-59277254.0/4294967296.0,1,-nbitq), 
to_sfixed(503545313.0/4294967296.0,1,-nbitq), 
to_sfixed(-298626363.0/4294967296.0,1,-nbitq), 
to_sfixed(49503439.0/4294967296.0,1,-nbitq), 
to_sfixed(171412611.0/4294967296.0,1,-nbitq), 
to_sfixed(556854455.0/4294967296.0,1,-nbitq), 
to_sfixed(408663784.0/4294967296.0,1,-nbitq), 
to_sfixed(248861524.0/4294967296.0,1,-nbitq), 
to_sfixed(365089148.0/4294967296.0,1,-nbitq), 
to_sfixed(-66902936.0/4294967296.0,1,-nbitq), 
to_sfixed(51120878.0/4294967296.0,1,-nbitq), 
to_sfixed(321911225.0/4294967296.0,1,-nbitq), 
to_sfixed(192288815.0/4294967296.0,1,-nbitq), 
to_sfixed(124223461.0/4294967296.0,1,-nbitq), 
to_sfixed(-176151057.0/4294967296.0,1,-nbitq), 
to_sfixed(-109909486.0/4294967296.0,1,-nbitq), 
to_sfixed(243267664.0/4294967296.0,1,-nbitq), 
to_sfixed(556773339.0/4294967296.0,1,-nbitq), 
to_sfixed(483675724.0/4294967296.0,1,-nbitq), 
to_sfixed(316046112.0/4294967296.0,1,-nbitq), 
to_sfixed(185114305.0/4294967296.0,1,-nbitq), 
to_sfixed(334708843.0/4294967296.0,1,-nbitq), 
to_sfixed(462197029.0/4294967296.0,1,-nbitq), 
to_sfixed(-287204970.0/4294967296.0,1,-nbitq), 
to_sfixed(446991279.0/4294967296.0,1,-nbitq), 
to_sfixed(227926223.0/4294967296.0,1,-nbitq), 
to_sfixed(51096862.0/4294967296.0,1,-nbitq), 
to_sfixed(231317847.0/4294967296.0,1,-nbitq), 
to_sfixed(-285842154.0/4294967296.0,1,-nbitq), 
to_sfixed(92754101.0/4294967296.0,1,-nbitq), 
to_sfixed(116012604.0/4294967296.0,1,-nbitq), 
to_sfixed(131015125.0/4294967296.0,1,-nbitq), 
to_sfixed(-211876664.0/4294967296.0,1,-nbitq), 
to_sfixed(-138193043.0/4294967296.0,1,-nbitq), 
to_sfixed(-149985299.0/4294967296.0,1,-nbitq), 
to_sfixed(-452840245.0/4294967296.0,1,-nbitq), 
to_sfixed(-219799196.0/4294967296.0,1,-nbitq), 
to_sfixed(-149633696.0/4294967296.0,1,-nbitq), 
to_sfixed(43331977.0/4294967296.0,1,-nbitq), 
to_sfixed(418792835.0/4294967296.0,1,-nbitq), 
to_sfixed(-96000460.0/4294967296.0,1,-nbitq), 
to_sfixed(6864213.0/4294967296.0,1,-nbitq), 
to_sfixed(-126634007.0/4294967296.0,1,-nbitq), 
to_sfixed(203946764.0/4294967296.0,1,-nbitq), 
to_sfixed(-201620077.0/4294967296.0,1,-nbitq), 
to_sfixed(-374952067.0/4294967296.0,1,-nbitq), 
to_sfixed(-318221906.0/4294967296.0,1,-nbitq), 
to_sfixed(12930302.0/4294967296.0,1,-nbitq), 
to_sfixed(-273339613.0/4294967296.0,1,-nbitq), 
to_sfixed(693877446.0/4294967296.0,1,-nbitq), 
to_sfixed(-359364173.0/4294967296.0,1,-nbitq), 
to_sfixed(-301820012.0/4294967296.0,1,-nbitq), 
to_sfixed(171661588.0/4294967296.0,1,-nbitq), 
to_sfixed(1890586.0/4294967296.0,1,-nbitq), 
to_sfixed(19195991.0/4294967296.0,1,-nbitq), 
to_sfixed(-223961293.0/4294967296.0,1,-nbitq), 
to_sfixed(291628025.0/4294967296.0,1,-nbitq), 
to_sfixed(227991811.0/4294967296.0,1,-nbitq), 
to_sfixed(-449996557.0/4294967296.0,1,-nbitq), 
to_sfixed(-266666497.0/4294967296.0,1,-nbitq), 
to_sfixed(-37848513.0/4294967296.0,1,-nbitq), 
to_sfixed(-244999595.0/4294967296.0,1,-nbitq), 
to_sfixed(399415335.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-323759358.0/4294967296.0,1,-nbitq), 
to_sfixed(-107211985.0/4294967296.0,1,-nbitq), 
to_sfixed(111301681.0/4294967296.0,1,-nbitq), 
to_sfixed(-68307635.0/4294967296.0,1,-nbitq), 
to_sfixed(384138032.0/4294967296.0,1,-nbitq), 
to_sfixed(173486682.0/4294967296.0,1,-nbitq), 
to_sfixed(117670663.0/4294967296.0,1,-nbitq), 
to_sfixed(55897032.0/4294967296.0,1,-nbitq), 
to_sfixed(145633474.0/4294967296.0,1,-nbitq), 
to_sfixed(-28069131.0/4294967296.0,1,-nbitq), 
to_sfixed(-209038226.0/4294967296.0,1,-nbitq), 
to_sfixed(314139142.0/4294967296.0,1,-nbitq), 
to_sfixed(-444057291.0/4294967296.0,1,-nbitq), 
to_sfixed(-175255903.0/4294967296.0,1,-nbitq), 
to_sfixed(-230250361.0/4294967296.0,1,-nbitq), 
to_sfixed(50411497.0/4294967296.0,1,-nbitq), 
to_sfixed(282941355.0/4294967296.0,1,-nbitq), 
to_sfixed(-274944561.0/4294967296.0,1,-nbitq), 
to_sfixed(334970008.0/4294967296.0,1,-nbitq), 
to_sfixed(66175012.0/4294967296.0,1,-nbitq), 
to_sfixed(-63820329.0/4294967296.0,1,-nbitq), 
to_sfixed(-260806083.0/4294967296.0,1,-nbitq), 
to_sfixed(-142811843.0/4294967296.0,1,-nbitq), 
to_sfixed(-396340074.0/4294967296.0,1,-nbitq), 
to_sfixed(333605426.0/4294967296.0,1,-nbitq), 
to_sfixed(-266283403.0/4294967296.0,1,-nbitq), 
to_sfixed(323711655.0/4294967296.0,1,-nbitq), 
to_sfixed(180821843.0/4294967296.0,1,-nbitq), 
to_sfixed(171782108.0/4294967296.0,1,-nbitq), 
to_sfixed(559026058.0/4294967296.0,1,-nbitq), 
to_sfixed(-185272111.0/4294967296.0,1,-nbitq), 
to_sfixed(-431678398.0/4294967296.0,1,-nbitq), 
to_sfixed(393434784.0/4294967296.0,1,-nbitq), 
to_sfixed(-475719315.0/4294967296.0,1,-nbitq), 
to_sfixed(-267157794.0/4294967296.0,1,-nbitq), 
to_sfixed(-10617780.0/4294967296.0,1,-nbitq), 
to_sfixed(477944399.0/4294967296.0,1,-nbitq), 
to_sfixed(266329841.0/4294967296.0,1,-nbitq), 
to_sfixed(-505909714.0/4294967296.0,1,-nbitq), 
to_sfixed(475523287.0/4294967296.0,1,-nbitq), 
to_sfixed(-220198793.0/4294967296.0,1,-nbitq), 
to_sfixed(-212780410.0/4294967296.0,1,-nbitq), 
to_sfixed(214269969.0/4294967296.0,1,-nbitq), 
to_sfixed(-97140791.0/4294967296.0,1,-nbitq), 
to_sfixed(271844356.0/4294967296.0,1,-nbitq), 
to_sfixed(28948591.0/4294967296.0,1,-nbitq), 
to_sfixed(33128331.0/4294967296.0,1,-nbitq), 
to_sfixed(-181375017.0/4294967296.0,1,-nbitq), 
to_sfixed(-360290720.0/4294967296.0,1,-nbitq), 
to_sfixed(319749332.0/4294967296.0,1,-nbitq), 
to_sfixed(220055272.0/4294967296.0,1,-nbitq), 
to_sfixed(-76012486.0/4294967296.0,1,-nbitq), 
to_sfixed(-384823872.0/4294967296.0,1,-nbitq), 
to_sfixed(420169486.0/4294967296.0,1,-nbitq), 
to_sfixed(155077950.0/4294967296.0,1,-nbitq), 
to_sfixed(359958316.0/4294967296.0,1,-nbitq), 
to_sfixed(-77805181.0/4294967296.0,1,-nbitq), 
to_sfixed(-27516474.0/4294967296.0,1,-nbitq), 
to_sfixed(-53503036.0/4294967296.0,1,-nbitq), 
to_sfixed(115593281.0/4294967296.0,1,-nbitq), 
to_sfixed(55195881.0/4294967296.0,1,-nbitq), 
to_sfixed(-255494697.0/4294967296.0,1,-nbitq), 
to_sfixed(-44704963.0/4294967296.0,1,-nbitq), 
to_sfixed(420119424.0/4294967296.0,1,-nbitq), 
to_sfixed(410365463.0/4294967296.0,1,-nbitq), 
to_sfixed(-369117959.0/4294967296.0,1,-nbitq), 
to_sfixed(331136980.0/4294967296.0,1,-nbitq), 
to_sfixed(234647612.0/4294967296.0,1,-nbitq), 
to_sfixed(298406578.0/4294967296.0,1,-nbitq), 
to_sfixed(-52679819.0/4294967296.0,1,-nbitq), 
to_sfixed(77311072.0/4294967296.0,1,-nbitq), 
to_sfixed(-19128916.0/4294967296.0,1,-nbitq), 
to_sfixed(-533652844.0/4294967296.0,1,-nbitq), 
to_sfixed(211300999.0/4294967296.0,1,-nbitq), 
to_sfixed(522687154.0/4294967296.0,1,-nbitq), 
to_sfixed(-431940634.0/4294967296.0,1,-nbitq), 
to_sfixed(-116439465.0/4294967296.0,1,-nbitq), 
to_sfixed(432573556.0/4294967296.0,1,-nbitq), 
to_sfixed(-424553018.0/4294967296.0,1,-nbitq), 
to_sfixed(349822773.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-135062708.0/4294967296.0,1,-nbitq), 
to_sfixed(-231059740.0/4294967296.0,1,-nbitq), 
to_sfixed(-194776007.0/4294967296.0,1,-nbitq), 
to_sfixed(-250530563.0/4294967296.0,1,-nbitq), 
to_sfixed(108009325.0/4294967296.0,1,-nbitq), 
to_sfixed(427454558.0/4294967296.0,1,-nbitq), 
to_sfixed(68231471.0/4294967296.0,1,-nbitq), 
to_sfixed(-245634271.0/4294967296.0,1,-nbitq), 
to_sfixed(705326718.0/4294967296.0,1,-nbitq), 
to_sfixed(195880012.0/4294967296.0,1,-nbitq), 
to_sfixed(-222348833.0/4294967296.0,1,-nbitq), 
to_sfixed(465344702.0/4294967296.0,1,-nbitq), 
to_sfixed(-628304380.0/4294967296.0,1,-nbitq), 
to_sfixed(189675191.0/4294967296.0,1,-nbitq), 
to_sfixed(148437834.0/4294967296.0,1,-nbitq), 
to_sfixed(-115881949.0/4294967296.0,1,-nbitq), 
to_sfixed(248843071.0/4294967296.0,1,-nbitq), 
to_sfixed(-204819639.0/4294967296.0,1,-nbitq), 
to_sfixed(-347268394.0/4294967296.0,1,-nbitq), 
to_sfixed(-164704400.0/4294967296.0,1,-nbitq), 
to_sfixed(-408558394.0/4294967296.0,1,-nbitq), 
to_sfixed(223441267.0/4294967296.0,1,-nbitq), 
to_sfixed(346925040.0/4294967296.0,1,-nbitq), 
to_sfixed(-579427029.0/4294967296.0,1,-nbitq), 
to_sfixed(332415196.0/4294967296.0,1,-nbitq), 
to_sfixed(-218966730.0/4294967296.0,1,-nbitq), 
to_sfixed(396116289.0/4294967296.0,1,-nbitq), 
to_sfixed(-26544438.0/4294967296.0,1,-nbitq), 
to_sfixed(-116246702.0/4294967296.0,1,-nbitq), 
to_sfixed(21199388.0/4294967296.0,1,-nbitq), 
to_sfixed(89277321.0/4294967296.0,1,-nbitq), 
to_sfixed(-595221214.0/4294967296.0,1,-nbitq), 
to_sfixed(-152436495.0/4294967296.0,1,-nbitq), 
to_sfixed(-34976361.0/4294967296.0,1,-nbitq), 
to_sfixed(-223112529.0/4294967296.0,1,-nbitq), 
to_sfixed(-250743113.0/4294967296.0,1,-nbitq), 
to_sfixed(780677295.0/4294967296.0,1,-nbitq), 
to_sfixed(98209029.0/4294967296.0,1,-nbitq), 
to_sfixed(-206324588.0/4294967296.0,1,-nbitq), 
to_sfixed(391305806.0/4294967296.0,1,-nbitq), 
to_sfixed(-402717578.0/4294967296.0,1,-nbitq), 
to_sfixed(205429211.0/4294967296.0,1,-nbitq), 
to_sfixed(-236687992.0/4294967296.0,1,-nbitq), 
to_sfixed(487436672.0/4294967296.0,1,-nbitq), 
to_sfixed(-420960013.0/4294967296.0,1,-nbitq), 
to_sfixed(85720230.0/4294967296.0,1,-nbitq), 
to_sfixed(-188788274.0/4294967296.0,1,-nbitq), 
to_sfixed(-364940723.0/4294967296.0,1,-nbitq), 
to_sfixed(-354208220.0/4294967296.0,1,-nbitq), 
to_sfixed(607980304.0/4294967296.0,1,-nbitq), 
to_sfixed(-195721496.0/4294967296.0,1,-nbitq), 
to_sfixed(-249848438.0/4294967296.0,1,-nbitq), 
to_sfixed(-521709315.0/4294967296.0,1,-nbitq), 
to_sfixed(360674541.0/4294967296.0,1,-nbitq), 
to_sfixed(-256063861.0/4294967296.0,1,-nbitq), 
to_sfixed(-95890609.0/4294967296.0,1,-nbitq), 
to_sfixed(-11409209.0/4294967296.0,1,-nbitq), 
to_sfixed(-252301578.0/4294967296.0,1,-nbitq), 
to_sfixed(74186950.0/4294967296.0,1,-nbitq), 
to_sfixed(369297706.0/4294967296.0,1,-nbitq), 
to_sfixed(-173540621.0/4294967296.0,1,-nbitq), 
to_sfixed(219158323.0/4294967296.0,1,-nbitq), 
to_sfixed(-154146918.0/4294967296.0,1,-nbitq), 
to_sfixed(-269289036.0/4294967296.0,1,-nbitq), 
to_sfixed(-188926080.0/4294967296.0,1,-nbitq), 
to_sfixed(-177147291.0/4294967296.0,1,-nbitq), 
to_sfixed(648426434.0/4294967296.0,1,-nbitq), 
to_sfixed(85732363.0/4294967296.0,1,-nbitq), 
to_sfixed(-132277053.0/4294967296.0,1,-nbitq), 
to_sfixed(320020367.0/4294967296.0,1,-nbitq), 
to_sfixed(-272013152.0/4294967296.0,1,-nbitq), 
to_sfixed(291207479.0/4294967296.0,1,-nbitq), 
to_sfixed(-70081910.0/4294967296.0,1,-nbitq), 
to_sfixed(-323494302.0/4294967296.0,1,-nbitq), 
to_sfixed(-235134254.0/4294967296.0,1,-nbitq), 
to_sfixed(170778387.0/4294967296.0,1,-nbitq), 
to_sfixed(585692070.0/4294967296.0,1,-nbitq), 
to_sfixed(364768412.0/4294967296.0,1,-nbitq), 
to_sfixed(-393119607.0/4294967296.0,1,-nbitq), 
to_sfixed(227236912.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(368268949.0/4294967296.0,1,-nbitq), 
to_sfixed(-520445861.0/4294967296.0,1,-nbitq), 
to_sfixed(-61517331.0/4294967296.0,1,-nbitq), 
to_sfixed(-70510078.0/4294967296.0,1,-nbitq), 
to_sfixed(604850199.0/4294967296.0,1,-nbitq), 
to_sfixed(-38640522.0/4294967296.0,1,-nbitq), 
to_sfixed(-315875208.0/4294967296.0,1,-nbitq), 
to_sfixed(-270990664.0/4294967296.0,1,-nbitq), 
to_sfixed(795786996.0/4294967296.0,1,-nbitq), 
to_sfixed(-219511285.0/4294967296.0,1,-nbitq), 
to_sfixed(85008203.0/4294967296.0,1,-nbitq), 
to_sfixed(689673486.0/4294967296.0,1,-nbitq), 
to_sfixed(-476277251.0/4294967296.0,1,-nbitq), 
to_sfixed(90969691.0/4294967296.0,1,-nbitq), 
to_sfixed(-243430065.0/4294967296.0,1,-nbitq), 
to_sfixed(-23698309.0/4294967296.0,1,-nbitq), 
to_sfixed(-21018010.0/4294967296.0,1,-nbitq), 
to_sfixed(-230442720.0/4294967296.0,1,-nbitq), 
to_sfixed(138202216.0/4294967296.0,1,-nbitq), 
to_sfixed(116513031.0/4294967296.0,1,-nbitq), 
to_sfixed(-161383357.0/4294967296.0,1,-nbitq), 
to_sfixed(-39370425.0/4294967296.0,1,-nbitq), 
to_sfixed(284701349.0/4294967296.0,1,-nbitq), 
to_sfixed(240875575.0/4294967296.0,1,-nbitq), 
to_sfixed(-73853435.0/4294967296.0,1,-nbitq), 
to_sfixed(-418121957.0/4294967296.0,1,-nbitq), 
to_sfixed(385398230.0/4294967296.0,1,-nbitq), 
to_sfixed(-236587445.0/4294967296.0,1,-nbitq), 
to_sfixed(184922548.0/4294967296.0,1,-nbitq), 
to_sfixed(257993234.0/4294967296.0,1,-nbitq), 
to_sfixed(-263059404.0/4294967296.0,1,-nbitq), 
to_sfixed(-229964036.0/4294967296.0,1,-nbitq), 
to_sfixed(328969826.0/4294967296.0,1,-nbitq), 
to_sfixed(44310039.0/4294967296.0,1,-nbitq), 
to_sfixed(-261395809.0/4294967296.0,1,-nbitq), 
to_sfixed(24023574.0/4294967296.0,1,-nbitq), 
to_sfixed(70309865.0/4294967296.0,1,-nbitq), 
to_sfixed(-260130889.0/4294967296.0,1,-nbitq), 
to_sfixed(-167672096.0/4294967296.0,1,-nbitq), 
to_sfixed(-101185289.0/4294967296.0,1,-nbitq), 
to_sfixed(-347579769.0/4294967296.0,1,-nbitq), 
to_sfixed(266305266.0/4294967296.0,1,-nbitq), 
to_sfixed(-185149114.0/4294967296.0,1,-nbitq), 
to_sfixed(395938203.0/4294967296.0,1,-nbitq), 
to_sfixed(130616992.0/4294967296.0,1,-nbitq), 
to_sfixed(-55141100.0/4294967296.0,1,-nbitq), 
to_sfixed(204663135.0/4294967296.0,1,-nbitq), 
to_sfixed(-262530392.0/4294967296.0,1,-nbitq), 
to_sfixed(-383462987.0/4294967296.0,1,-nbitq), 
to_sfixed(424280075.0/4294967296.0,1,-nbitq), 
to_sfixed(-399227225.0/4294967296.0,1,-nbitq), 
to_sfixed(381821570.0/4294967296.0,1,-nbitq), 
to_sfixed(-24237453.0/4294967296.0,1,-nbitq), 
to_sfixed(377700446.0/4294967296.0,1,-nbitq), 
to_sfixed(-342146919.0/4294967296.0,1,-nbitq), 
to_sfixed(-46798066.0/4294967296.0,1,-nbitq), 
to_sfixed(326464815.0/4294967296.0,1,-nbitq), 
to_sfixed(45762934.0/4294967296.0,1,-nbitq), 
to_sfixed(-34351649.0/4294967296.0,1,-nbitq), 
to_sfixed(96116764.0/4294967296.0,1,-nbitq), 
to_sfixed(-209312620.0/4294967296.0,1,-nbitq), 
to_sfixed(-103972607.0/4294967296.0,1,-nbitq), 
to_sfixed(-370403953.0/4294967296.0,1,-nbitq), 
to_sfixed(272632324.0/4294967296.0,1,-nbitq), 
to_sfixed(-175269121.0/4294967296.0,1,-nbitq), 
to_sfixed(-73979321.0/4294967296.0,1,-nbitq), 
to_sfixed(124485199.0/4294967296.0,1,-nbitq), 
to_sfixed(-239081374.0/4294967296.0,1,-nbitq), 
to_sfixed(351518896.0/4294967296.0,1,-nbitq), 
to_sfixed(45156820.0/4294967296.0,1,-nbitq), 
to_sfixed(-672607876.0/4294967296.0,1,-nbitq), 
to_sfixed(-355149172.0/4294967296.0,1,-nbitq), 
to_sfixed(-168310060.0/4294967296.0,1,-nbitq), 
to_sfixed(124153398.0/4294967296.0,1,-nbitq), 
to_sfixed(-218055261.0/4294967296.0,1,-nbitq), 
to_sfixed(-198563632.0/4294967296.0,1,-nbitq), 
to_sfixed(251298820.0/4294967296.0,1,-nbitq), 
to_sfixed(-248458039.0/4294967296.0,1,-nbitq), 
to_sfixed(72449072.0/4294967296.0,1,-nbitq), 
to_sfixed(186423450.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-63580660.0/4294967296.0,1,-nbitq), 
to_sfixed(-420473653.0/4294967296.0,1,-nbitq), 
to_sfixed(435320720.0/4294967296.0,1,-nbitq), 
to_sfixed(-57438616.0/4294967296.0,1,-nbitq), 
to_sfixed(89447549.0/4294967296.0,1,-nbitq), 
to_sfixed(140635904.0/4294967296.0,1,-nbitq), 
to_sfixed(325160899.0/4294967296.0,1,-nbitq), 
to_sfixed(220505230.0/4294967296.0,1,-nbitq), 
to_sfixed(813602103.0/4294967296.0,1,-nbitq), 
to_sfixed(133689714.0/4294967296.0,1,-nbitq), 
to_sfixed(288519452.0/4294967296.0,1,-nbitq), 
to_sfixed(490436712.0/4294967296.0,1,-nbitq), 
to_sfixed(-812409967.0/4294967296.0,1,-nbitq), 
to_sfixed(195547840.0/4294967296.0,1,-nbitq), 
to_sfixed(-25847465.0/4294967296.0,1,-nbitq), 
to_sfixed(-143575066.0/4294967296.0,1,-nbitq), 
to_sfixed(88471839.0/4294967296.0,1,-nbitq), 
to_sfixed(416911290.0/4294967296.0,1,-nbitq), 
to_sfixed(287843912.0/4294967296.0,1,-nbitq), 
to_sfixed(-235437125.0/4294967296.0,1,-nbitq), 
to_sfixed(-356857783.0/4294967296.0,1,-nbitq), 
to_sfixed(-136216111.0/4294967296.0,1,-nbitq), 
to_sfixed(548450902.0/4294967296.0,1,-nbitq), 
to_sfixed(66397689.0/4294967296.0,1,-nbitq), 
to_sfixed(193858830.0/4294967296.0,1,-nbitq), 
to_sfixed(-214659364.0/4294967296.0,1,-nbitq), 
to_sfixed(-134635474.0/4294967296.0,1,-nbitq), 
to_sfixed(-349040587.0/4294967296.0,1,-nbitq), 
to_sfixed(223835716.0/4294967296.0,1,-nbitq), 
to_sfixed(197327252.0/4294967296.0,1,-nbitq), 
to_sfixed(-630863220.0/4294967296.0,1,-nbitq), 
to_sfixed(429197455.0/4294967296.0,1,-nbitq), 
to_sfixed(298872740.0/4294967296.0,1,-nbitq), 
to_sfixed(-3371026.0/4294967296.0,1,-nbitq), 
to_sfixed(-416276930.0/4294967296.0,1,-nbitq), 
to_sfixed(-70752703.0/4294967296.0,1,-nbitq), 
to_sfixed(564231424.0/4294967296.0,1,-nbitq), 
to_sfixed(-132030184.0/4294967296.0,1,-nbitq), 
to_sfixed(-58263216.0/4294967296.0,1,-nbitq), 
to_sfixed(308188727.0/4294967296.0,1,-nbitq), 
to_sfixed(348455120.0/4294967296.0,1,-nbitq), 
to_sfixed(12234507.0/4294967296.0,1,-nbitq), 
to_sfixed(-204569240.0/4294967296.0,1,-nbitq), 
to_sfixed(207084442.0/4294967296.0,1,-nbitq), 
to_sfixed(359445926.0/4294967296.0,1,-nbitq), 
to_sfixed(191115264.0/4294967296.0,1,-nbitq), 
to_sfixed(55116078.0/4294967296.0,1,-nbitq), 
to_sfixed(103664719.0/4294967296.0,1,-nbitq), 
to_sfixed(-277595284.0/4294967296.0,1,-nbitq), 
to_sfixed(422518641.0/4294967296.0,1,-nbitq), 
to_sfixed(143893691.0/4294967296.0,1,-nbitq), 
to_sfixed(-361268495.0/4294967296.0,1,-nbitq), 
to_sfixed(-103428512.0/4294967296.0,1,-nbitq), 
to_sfixed(-153050065.0/4294967296.0,1,-nbitq), 
to_sfixed(-32682894.0/4294967296.0,1,-nbitq), 
to_sfixed(630090198.0/4294967296.0,1,-nbitq), 
to_sfixed(5040077.0/4294967296.0,1,-nbitq), 
to_sfixed(-361436373.0/4294967296.0,1,-nbitq), 
to_sfixed(-179475607.0/4294967296.0,1,-nbitq), 
to_sfixed(380753141.0/4294967296.0,1,-nbitq), 
to_sfixed(54189796.0/4294967296.0,1,-nbitq), 
to_sfixed(17889704.0/4294967296.0,1,-nbitq), 
to_sfixed(-588754685.0/4294967296.0,1,-nbitq), 
to_sfixed(-297564158.0/4294967296.0,1,-nbitq), 
to_sfixed(245854491.0/4294967296.0,1,-nbitq), 
to_sfixed(-482919562.0/4294967296.0,1,-nbitq), 
to_sfixed(165076174.0/4294967296.0,1,-nbitq), 
to_sfixed(337339202.0/4294967296.0,1,-nbitq), 
to_sfixed(-35658276.0/4294967296.0,1,-nbitq), 
to_sfixed(-215927072.0/4294967296.0,1,-nbitq), 
to_sfixed(-330607302.0/4294967296.0,1,-nbitq), 
to_sfixed(27166807.0/4294967296.0,1,-nbitq), 
to_sfixed(319214940.0/4294967296.0,1,-nbitq), 
to_sfixed(-175486173.0/4294967296.0,1,-nbitq), 
to_sfixed(64261456.0/4294967296.0,1,-nbitq), 
to_sfixed(37792663.0/4294967296.0,1,-nbitq), 
to_sfixed(-31772406.0/4294967296.0,1,-nbitq), 
to_sfixed(207503708.0/4294967296.0,1,-nbitq), 
to_sfixed(50166479.0/4294967296.0,1,-nbitq), 
to_sfixed(-360993498.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(472452608.0/4294967296.0,1,-nbitq), 
to_sfixed(155582148.0/4294967296.0,1,-nbitq), 
to_sfixed(-139798514.0/4294967296.0,1,-nbitq), 
to_sfixed(-76332197.0/4294967296.0,1,-nbitq), 
to_sfixed(-144890439.0/4294967296.0,1,-nbitq), 
to_sfixed(-162268499.0/4294967296.0,1,-nbitq), 
to_sfixed(86521317.0/4294967296.0,1,-nbitq), 
to_sfixed(74243917.0/4294967296.0,1,-nbitq), 
to_sfixed(802374369.0/4294967296.0,1,-nbitq), 
to_sfixed(39568961.0/4294967296.0,1,-nbitq), 
to_sfixed(4174691.0/4294967296.0,1,-nbitq), 
to_sfixed(316336605.0/4294967296.0,1,-nbitq), 
to_sfixed(-255801858.0/4294967296.0,1,-nbitq), 
to_sfixed(-274068320.0/4294967296.0,1,-nbitq), 
to_sfixed(162018981.0/4294967296.0,1,-nbitq), 
to_sfixed(147086460.0/4294967296.0,1,-nbitq), 
to_sfixed(-48316868.0/4294967296.0,1,-nbitq), 
to_sfixed(-52556493.0/4294967296.0,1,-nbitq), 
to_sfixed(378367064.0/4294967296.0,1,-nbitq), 
to_sfixed(40974146.0/4294967296.0,1,-nbitq), 
to_sfixed(5158678.0/4294967296.0,1,-nbitq), 
to_sfixed(403268380.0/4294967296.0,1,-nbitq), 
to_sfixed(177315681.0/4294967296.0,1,-nbitq), 
to_sfixed(-25103475.0/4294967296.0,1,-nbitq), 
to_sfixed(-199162894.0/4294967296.0,1,-nbitq), 
to_sfixed(387766505.0/4294967296.0,1,-nbitq), 
to_sfixed(-18520047.0/4294967296.0,1,-nbitq), 
to_sfixed(173532854.0/4294967296.0,1,-nbitq), 
to_sfixed(4507095.0/4294967296.0,1,-nbitq), 
to_sfixed(197064293.0/4294967296.0,1,-nbitq), 
to_sfixed(-414723659.0/4294967296.0,1,-nbitq), 
to_sfixed(-255716786.0/4294967296.0,1,-nbitq), 
to_sfixed(-211064327.0/4294967296.0,1,-nbitq), 
to_sfixed(-200095664.0/4294967296.0,1,-nbitq), 
to_sfixed(-121391287.0/4294967296.0,1,-nbitq), 
to_sfixed(-497958320.0/4294967296.0,1,-nbitq), 
to_sfixed(108437118.0/4294967296.0,1,-nbitq), 
to_sfixed(-217679339.0/4294967296.0,1,-nbitq), 
to_sfixed(-112746994.0/4294967296.0,1,-nbitq), 
to_sfixed(-110526083.0/4294967296.0,1,-nbitq), 
to_sfixed(-287125074.0/4294967296.0,1,-nbitq), 
to_sfixed(-57258851.0/4294967296.0,1,-nbitq), 
to_sfixed(84673364.0/4294967296.0,1,-nbitq), 
to_sfixed(680135318.0/4294967296.0,1,-nbitq), 
to_sfixed(-5065795.0/4294967296.0,1,-nbitq), 
to_sfixed(139276171.0/4294967296.0,1,-nbitq), 
to_sfixed(312698562.0/4294967296.0,1,-nbitq), 
to_sfixed(-365692218.0/4294967296.0,1,-nbitq), 
to_sfixed(199532017.0/4294967296.0,1,-nbitq), 
to_sfixed(318900333.0/4294967296.0,1,-nbitq), 
to_sfixed(-362411280.0/4294967296.0,1,-nbitq), 
to_sfixed(228930656.0/4294967296.0,1,-nbitq), 
to_sfixed(-654354513.0/4294967296.0,1,-nbitq), 
to_sfixed(-506769688.0/4294967296.0,1,-nbitq), 
to_sfixed(204672880.0/4294967296.0,1,-nbitq), 
to_sfixed(189382949.0/4294967296.0,1,-nbitq), 
to_sfixed(340279087.0/4294967296.0,1,-nbitq), 
to_sfixed(-117403885.0/4294967296.0,1,-nbitq), 
to_sfixed(277460587.0/4294967296.0,1,-nbitq), 
to_sfixed(194494323.0/4294967296.0,1,-nbitq), 
to_sfixed(-203722242.0/4294967296.0,1,-nbitq), 
to_sfixed(-147239815.0/4294967296.0,1,-nbitq), 
to_sfixed(168754594.0/4294967296.0,1,-nbitq), 
to_sfixed(-166455374.0/4294967296.0,1,-nbitq), 
to_sfixed(-335001058.0/4294967296.0,1,-nbitq), 
to_sfixed(282641958.0/4294967296.0,1,-nbitq), 
to_sfixed(556496291.0/4294967296.0,1,-nbitq), 
to_sfixed(114587532.0/4294967296.0,1,-nbitq), 
to_sfixed(-253727643.0/4294967296.0,1,-nbitq), 
to_sfixed(260090372.0/4294967296.0,1,-nbitq), 
to_sfixed(-155509137.0/4294967296.0,1,-nbitq), 
to_sfixed(-110931756.0/4294967296.0,1,-nbitq), 
to_sfixed(-4885444.0/4294967296.0,1,-nbitq), 
to_sfixed(55420096.0/4294967296.0,1,-nbitq), 
to_sfixed(279146743.0/4294967296.0,1,-nbitq), 
to_sfixed(-271501402.0/4294967296.0,1,-nbitq), 
to_sfixed(-116100381.0/4294967296.0,1,-nbitq), 
to_sfixed(-515684377.0/4294967296.0,1,-nbitq), 
to_sfixed(-321899718.0/4294967296.0,1,-nbitq), 
to_sfixed(211303821.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(394285858.0/4294967296.0,1,-nbitq), 
to_sfixed(318058196.0/4294967296.0,1,-nbitq), 
to_sfixed(147515678.0/4294967296.0,1,-nbitq), 
to_sfixed(244437733.0/4294967296.0,1,-nbitq), 
to_sfixed(-310799909.0/4294967296.0,1,-nbitq), 
to_sfixed(-76213692.0/4294967296.0,1,-nbitq), 
to_sfixed(-127933758.0/4294967296.0,1,-nbitq), 
to_sfixed(31748635.0/4294967296.0,1,-nbitq), 
to_sfixed(290309593.0/4294967296.0,1,-nbitq), 
to_sfixed(121516850.0/4294967296.0,1,-nbitq), 
to_sfixed(213237148.0/4294967296.0,1,-nbitq), 
to_sfixed(674776983.0/4294967296.0,1,-nbitq), 
to_sfixed(-535837310.0/4294967296.0,1,-nbitq), 
to_sfixed(-386383053.0/4294967296.0,1,-nbitq), 
to_sfixed(-25027499.0/4294967296.0,1,-nbitq), 
to_sfixed(-153277077.0/4294967296.0,1,-nbitq), 
to_sfixed(27609860.0/4294967296.0,1,-nbitq), 
to_sfixed(-96396501.0/4294967296.0,1,-nbitq), 
to_sfixed(-6863458.0/4294967296.0,1,-nbitq), 
to_sfixed(-88568322.0/4294967296.0,1,-nbitq), 
to_sfixed(-220135638.0/4294967296.0,1,-nbitq), 
to_sfixed(-220867213.0/4294967296.0,1,-nbitq), 
to_sfixed(-105430816.0/4294967296.0,1,-nbitq), 
to_sfixed(-35809251.0/4294967296.0,1,-nbitq), 
to_sfixed(41356462.0/4294967296.0,1,-nbitq), 
to_sfixed(-326077402.0/4294967296.0,1,-nbitq), 
to_sfixed(-383023619.0/4294967296.0,1,-nbitq), 
to_sfixed(-215680778.0/4294967296.0,1,-nbitq), 
to_sfixed(423939374.0/4294967296.0,1,-nbitq), 
to_sfixed(132043125.0/4294967296.0,1,-nbitq), 
to_sfixed(-50921851.0/4294967296.0,1,-nbitq), 
to_sfixed(-104608857.0/4294967296.0,1,-nbitq), 
to_sfixed(25081646.0/4294967296.0,1,-nbitq), 
to_sfixed(-155655058.0/4294967296.0,1,-nbitq), 
to_sfixed(-240111522.0/4294967296.0,1,-nbitq), 
to_sfixed(-496965643.0/4294967296.0,1,-nbitq), 
to_sfixed(-40644483.0/4294967296.0,1,-nbitq), 
to_sfixed(-257320282.0/4294967296.0,1,-nbitq), 
to_sfixed(97785188.0/4294967296.0,1,-nbitq), 
to_sfixed(31581151.0/4294967296.0,1,-nbitq), 
to_sfixed(260051971.0/4294967296.0,1,-nbitq), 
to_sfixed(-344559049.0/4294967296.0,1,-nbitq), 
to_sfixed(180861341.0/4294967296.0,1,-nbitq), 
to_sfixed(-67946237.0/4294967296.0,1,-nbitq), 
to_sfixed(-423663057.0/4294967296.0,1,-nbitq), 
to_sfixed(525913462.0/4294967296.0,1,-nbitq), 
to_sfixed(-10838128.0/4294967296.0,1,-nbitq), 
to_sfixed(-72032077.0/4294967296.0,1,-nbitq), 
to_sfixed(26754306.0/4294967296.0,1,-nbitq), 
to_sfixed(250527605.0/4294967296.0,1,-nbitq), 
to_sfixed(-283897065.0/4294967296.0,1,-nbitq), 
to_sfixed(-42752568.0/4294967296.0,1,-nbitq), 
to_sfixed(-291321725.0/4294967296.0,1,-nbitq), 
to_sfixed(117595372.0/4294967296.0,1,-nbitq), 
to_sfixed(64307431.0/4294967296.0,1,-nbitq), 
to_sfixed(746873365.0/4294967296.0,1,-nbitq), 
to_sfixed(59251142.0/4294967296.0,1,-nbitq), 
to_sfixed(273290399.0/4294967296.0,1,-nbitq), 
to_sfixed(92459360.0/4294967296.0,1,-nbitq), 
to_sfixed(20230043.0/4294967296.0,1,-nbitq), 
to_sfixed(-277821259.0/4294967296.0,1,-nbitq), 
to_sfixed(200947036.0/4294967296.0,1,-nbitq), 
to_sfixed(-620990543.0/4294967296.0,1,-nbitq), 
to_sfixed(330710699.0/4294967296.0,1,-nbitq), 
to_sfixed(-131774617.0/4294967296.0,1,-nbitq), 
to_sfixed(22466953.0/4294967296.0,1,-nbitq), 
to_sfixed(753329954.0/4294967296.0,1,-nbitq), 
to_sfixed(-324419347.0/4294967296.0,1,-nbitq), 
to_sfixed(182146856.0/4294967296.0,1,-nbitq), 
to_sfixed(368614022.0/4294967296.0,1,-nbitq), 
to_sfixed(-130266498.0/4294967296.0,1,-nbitq), 
to_sfixed(-527461739.0/4294967296.0,1,-nbitq), 
to_sfixed(134814310.0/4294967296.0,1,-nbitq), 
to_sfixed(201410799.0/4294967296.0,1,-nbitq), 
to_sfixed(58256013.0/4294967296.0,1,-nbitq), 
to_sfixed(53665800.0/4294967296.0,1,-nbitq), 
to_sfixed(306534163.0/4294967296.0,1,-nbitq), 
to_sfixed(-35304932.0/4294967296.0,1,-nbitq), 
to_sfixed(-460405792.0/4294967296.0,1,-nbitq), 
to_sfixed(357307474.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(389119753.0/4294967296.0,1,-nbitq), 
to_sfixed(590726917.0/4294967296.0,1,-nbitq), 
to_sfixed(54959533.0/4294967296.0,1,-nbitq), 
to_sfixed(412881591.0/4294967296.0,1,-nbitq), 
to_sfixed(-335096362.0/4294967296.0,1,-nbitq), 
to_sfixed(-6630227.0/4294967296.0,1,-nbitq), 
to_sfixed(-236803256.0/4294967296.0,1,-nbitq), 
to_sfixed(-298434457.0/4294967296.0,1,-nbitq), 
to_sfixed(419113089.0/4294967296.0,1,-nbitq), 
to_sfixed(228657734.0/4294967296.0,1,-nbitq), 
to_sfixed(153324020.0/4294967296.0,1,-nbitq), 
to_sfixed(355980094.0/4294967296.0,1,-nbitq), 
to_sfixed(-169420230.0/4294967296.0,1,-nbitq), 
to_sfixed(-634247108.0/4294967296.0,1,-nbitq), 
to_sfixed(225919425.0/4294967296.0,1,-nbitq), 
to_sfixed(-127211007.0/4294967296.0,1,-nbitq), 
to_sfixed(315520839.0/4294967296.0,1,-nbitq), 
to_sfixed(394995143.0/4294967296.0,1,-nbitq), 
to_sfixed(274072113.0/4294967296.0,1,-nbitq), 
to_sfixed(-199537069.0/4294967296.0,1,-nbitq), 
to_sfixed(-368023034.0/4294967296.0,1,-nbitq), 
to_sfixed(250181291.0/4294967296.0,1,-nbitq), 
to_sfixed(-126982218.0/4294967296.0,1,-nbitq), 
to_sfixed(-111244253.0/4294967296.0,1,-nbitq), 
to_sfixed(134287375.0/4294967296.0,1,-nbitq), 
to_sfixed(-75724434.0/4294967296.0,1,-nbitq), 
to_sfixed(-178794765.0/4294967296.0,1,-nbitq), 
to_sfixed(-285344502.0/4294967296.0,1,-nbitq), 
to_sfixed(484608329.0/4294967296.0,1,-nbitq), 
to_sfixed(-331871065.0/4294967296.0,1,-nbitq), 
to_sfixed(146052042.0/4294967296.0,1,-nbitq), 
to_sfixed(2339099.0/4294967296.0,1,-nbitq), 
to_sfixed(-424318189.0/4294967296.0,1,-nbitq), 
to_sfixed(241347429.0/4294967296.0,1,-nbitq), 
to_sfixed(-382280703.0/4294967296.0,1,-nbitq), 
to_sfixed(-362684281.0/4294967296.0,1,-nbitq), 
to_sfixed(202270485.0/4294967296.0,1,-nbitq), 
to_sfixed(-64258323.0/4294967296.0,1,-nbitq), 
to_sfixed(275328443.0/4294967296.0,1,-nbitq), 
to_sfixed(-141517968.0/4294967296.0,1,-nbitq), 
to_sfixed(521132215.0/4294967296.0,1,-nbitq), 
to_sfixed(72770706.0/4294967296.0,1,-nbitq), 
to_sfixed(480483775.0/4294967296.0,1,-nbitq), 
to_sfixed(376206926.0/4294967296.0,1,-nbitq), 
to_sfixed(402040756.0/4294967296.0,1,-nbitq), 
to_sfixed(341914481.0/4294967296.0,1,-nbitq), 
to_sfixed(106307151.0/4294967296.0,1,-nbitq), 
to_sfixed(507061296.0/4294967296.0,1,-nbitq), 
to_sfixed(-225399795.0/4294967296.0,1,-nbitq), 
to_sfixed(169247207.0/4294967296.0,1,-nbitq), 
to_sfixed(-127056041.0/4294967296.0,1,-nbitq), 
to_sfixed(420427114.0/4294967296.0,1,-nbitq), 
to_sfixed(-238884162.0/4294967296.0,1,-nbitq), 
to_sfixed(-482035891.0/4294967296.0,1,-nbitq), 
to_sfixed(-544023645.0/4294967296.0,1,-nbitq), 
to_sfixed(92783787.0/4294967296.0,1,-nbitq), 
to_sfixed(220718013.0/4294967296.0,1,-nbitq), 
to_sfixed(239783258.0/4294967296.0,1,-nbitq), 
to_sfixed(-143056482.0/4294967296.0,1,-nbitq), 
to_sfixed(-158616555.0/4294967296.0,1,-nbitq), 
to_sfixed(74736605.0/4294967296.0,1,-nbitq), 
to_sfixed(-347576269.0/4294967296.0,1,-nbitq), 
to_sfixed(-142982091.0/4294967296.0,1,-nbitq), 
to_sfixed(33114158.0/4294967296.0,1,-nbitq), 
to_sfixed(329808318.0/4294967296.0,1,-nbitq), 
to_sfixed(-441511512.0/4294967296.0,1,-nbitq), 
to_sfixed(371478509.0/4294967296.0,1,-nbitq), 
to_sfixed(-140525488.0/4294967296.0,1,-nbitq), 
to_sfixed(324269422.0/4294967296.0,1,-nbitq), 
to_sfixed(123095975.0/4294967296.0,1,-nbitq), 
to_sfixed(258649331.0/4294967296.0,1,-nbitq), 
to_sfixed(-337916567.0/4294967296.0,1,-nbitq), 
to_sfixed(-89398411.0/4294967296.0,1,-nbitq), 
to_sfixed(1900974.0/4294967296.0,1,-nbitq), 
to_sfixed(219611013.0/4294967296.0,1,-nbitq), 
to_sfixed(-219924388.0/4294967296.0,1,-nbitq), 
to_sfixed(311048720.0/4294967296.0,1,-nbitq), 
to_sfixed(-543993328.0/4294967296.0,1,-nbitq), 
to_sfixed(-121712829.0/4294967296.0,1,-nbitq), 
to_sfixed(-108106408.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-74160468.0/4294967296.0,1,-nbitq), 
to_sfixed(364607007.0/4294967296.0,1,-nbitq), 
to_sfixed(-319778860.0/4294967296.0,1,-nbitq), 
to_sfixed(-31831774.0/4294967296.0,1,-nbitq), 
to_sfixed(-502417430.0/4294967296.0,1,-nbitq), 
to_sfixed(-59012279.0/4294967296.0,1,-nbitq), 
to_sfixed(-10307126.0/4294967296.0,1,-nbitq), 
to_sfixed(87106536.0/4294967296.0,1,-nbitq), 
to_sfixed(526022882.0/4294967296.0,1,-nbitq), 
to_sfixed(430787839.0/4294967296.0,1,-nbitq), 
to_sfixed(480993082.0/4294967296.0,1,-nbitq), 
to_sfixed(525325296.0/4294967296.0,1,-nbitq), 
to_sfixed(164405179.0/4294967296.0,1,-nbitq), 
to_sfixed(-322077074.0/4294967296.0,1,-nbitq), 
to_sfixed(62378511.0/4294967296.0,1,-nbitq), 
to_sfixed(-241869669.0/4294967296.0,1,-nbitq), 
to_sfixed(122071676.0/4294967296.0,1,-nbitq), 
to_sfixed(140033346.0/4294967296.0,1,-nbitq), 
to_sfixed(-231048962.0/4294967296.0,1,-nbitq), 
to_sfixed(-261530163.0/4294967296.0,1,-nbitq), 
to_sfixed(356901157.0/4294967296.0,1,-nbitq), 
to_sfixed(72657562.0/4294967296.0,1,-nbitq), 
to_sfixed(345979935.0/4294967296.0,1,-nbitq), 
to_sfixed(28891581.0/4294967296.0,1,-nbitq), 
to_sfixed(-173935807.0/4294967296.0,1,-nbitq), 
to_sfixed(347120896.0/4294967296.0,1,-nbitq), 
to_sfixed(-229629380.0/4294967296.0,1,-nbitq), 
to_sfixed(66225805.0/4294967296.0,1,-nbitq), 
to_sfixed(-131789433.0/4294967296.0,1,-nbitq), 
to_sfixed(135663655.0/4294967296.0,1,-nbitq), 
to_sfixed(145555684.0/4294967296.0,1,-nbitq), 
to_sfixed(-332464769.0/4294967296.0,1,-nbitq), 
to_sfixed(390151631.0/4294967296.0,1,-nbitq), 
to_sfixed(248644883.0/4294967296.0,1,-nbitq), 
to_sfixed(-616465526.0/4294967296.0,1,-nbitq), 
to_sfixed(-223618730.0/4294967296.0,1,-nbitq), 
to_sfixed(-63213641.0/4294967296.0,1,-nbitq), 
to_sfixed(-187335077.0/4294967296.0,1,-nbitq), 
to_sfixed(-414539390.0/4294967296.0,1,-nbitq), 
to_sfixed(141664930.0/4294967296.0,1,-nbitq), 
to_sfixed(-105714092.0/4294967296.0,1,-nbitq), 
to_sfixed(313693600.0/4294967296.0,1,-nbitq), 
to_sfixed(520900862.0/4294967296.0,1,-nbitq), 
to_sfixed(192511550.0/4294967296.0,1,-nbitq), 
to_sfixed(332893558.0/4294967296.0,1,-nbitq), 
to_sfixed(-100037939.0/4294967296.0,1,-nbitq), 
to_sfixed(129396228.0/4294967296.0,1,-nbitq), 
to_sfixed(70924429.0/4294967296.0,1,-nbitq), 
to_sfixed(485323267.0/4294967296.0,1,-nbitq), 
to_sfixed(301810597.0/4294967296.0,1,-nbitq), 
to_sfixed(-45154102.0/4294967296.0,1,-nbitq), 
to_sfixed(168651532.0/4294967296.0,1,-nbitq), 
to_sfixed(-364720088.0/4294967296.0,1,-nbitq), 
to_sfixed(413487993.0/4294967296.0,1,-nbitq), 
to_sfixed(-234833994.0/4294967296.0,1,-nbitq), 
to_sfixed(145736061.0/4294967296.0,1,-nbitq), 
to_sfixed(195956042.0/4294967296.0,1,-nbitq), 
to_sfixed(-381154840.0/4294967296.0,1,-nbitq), 
to_sfixed(-211312753.0/4294967296.0,1,-nbitq), 
to_sfixed(-127040472.0/4294967296.0,1,-nbitq), 
to_sfixed(260004446.0/4294967296.0,1,-nbitq), 
to_sfixed(-24064952.0/4294967296.0,1,-nbitq), 
to_sfixed(-401381336.0/4294967296.0,1,-nbitq), 
to_sfixed(358250711.0/4294967296.0,1,-nbitq), 
to_sfixed(-401740675.0/4294967296.0,1,-nbitq), 
to_sfixed(-330042222.0/4294967296.0,1,-nbitq), 
to_sfixed(805105037.0/4294967296.0,1,-nbitq), 
to_sfixed(319962380.0/4294967296.0,1,-nbitq), 
to_sfixed(250483600.0/4294967296.0,1,-nbitq), 
to_sfixed(-317942274.0/4294967296.0,1,-nbitq), 
to_sfixed(-2096317.0/4294967296.0,1,-nbitq), 
to_sfixed(-187522943.0/4294967296.0,1,-nbitq), 
to_sfixed(-254799394.0/4294967296.0,1,-nbitq), 
to_sfixed(306857513.0/4294967296.0,1,-nbitq), 
to_sfixed(22768658.0/4294967296.0,1,-nbitq), 
to_sfixed(358879648.0/4294967296.0,1,-nbitq), 
to_sfixed(608623701.0/4294967296.0,1,-nbitq), 
to_sfixed(-420516755.0/4294967296.0,1,-nbitq), 
to_sfixed(264835934.0/4294967296.0,1,-nbitq), 
to_sfixed(-189420756.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-190417024.0/4294967296.0,1,-nbitq), 
to_sfixed(602424322.0/4294967296.0,1,-nbitq), 
to_sfixed(-314395201.0/4294967296.0,1,-nbitq), 
to_sfixed(111447353.0/4294967296.0,1,-nbitq), 
to_sfixed(-105080360.0/4294967296.0,1,-nbitq), 
to_sfixed(-205869404.0/4294967296.0,1,-nbitq), 
to_sfixed(-394597497.0/4294967296.0,1,-nbitq), 
to_sfixed(36085338.0/4294967296.0,1,-nbitq), 
to_sfixed(895171473.0/4294967296.0,1,-nbitq), 
to_sfixed(-22394926.0/4294967296.0,1,-nbitq), 
to_sfixed(95003462.0/4294967296.0,1,-nbitq), 
to_sfixed(178006321.0/4294967296.0,1,-nbitq), 
to_sfixed(330838915.0/4294967296.0,1,-nbitq), 
to_sfixed(-188420174.0/4294967296.0,1,-nbitq), 
to_sfixed(-408584545.0/4294967296.0,1,-nbitq), 
to_sfixed(-409878460.0/4294967296.0,1,-nbitq), 
to_sfixed(34968989.0/4294967296.0,1,-nbitq), 
to_sfixed(318923691.0/4294967296.0,1,-nbitq), 
to_sfixed(72456456.0/4294967296.0,1,-nbitq), 
to_sfixed(-276239976.0/4294967296.0,1,-nbitq), 
to_sfixed(-67815849.0/4294967296.0,1,-nbitq), 
to_sfixed(-233902661.0/4294967296.0,1,-nbitq), 
to_sfixed(-267521677.0/4294967296.0,1,-nbitq), 
to_sfixed(-485483902.0/4294967296.0,1,-nbitq), 
to_sfixed(108668127.0/4294967296.0,1,-nbitq), 
to_sfixed(229029216.0/4294967296.0,1,-nbitq), 
to_sfixed(-244638551.0/4294967296.0,1,-nbitq), 
to_sfixed(-538797155.0/4294967296.0,1,-nbitq), 
to_sfixed(412893109.0/4294967296.0,1,-nbitq), 
to_sfixed(-148390414.0/4294967296.0,1,-nbitq), 
to_sfixed(237207403.0/4294967296.0,1,-nbitq), 
to_sfixed(267791420.0/4294967296.0,1,-nbitq), 
to_sfixed(133132675.0/4294967296.0,1,-nbitq), 
to_sfixed(-60265315.0/4294967296.0,1,-nbitq), 
to_sfixed(-122209910.0/4294967296.0,1,-nbitq), 
to_sfixed(80630274.0/4294967296.0,1,-nbitq), 
to_sfixed(-57764738.0/4294967296.0,1,-nbitq), 
to_sfixed(216847693.0/4294967296.0,1,-nbitq), 
to_sfixed(104862167.0/4294967296.0,1,-nbitq), 
to_sfixed(202999980.0/4294967296.0,1,-nbitq), 
to_sfixed(-230060821.0/4294967296.0,1,-nbitq), 
to_sfixed(492349875.0/4294967296.0,1,-nbitq), 
to_sfixed(610923462.0/4294967296.0,1,-nbitq), 
to_sfixed(861113083.0/4294967296.0,1,-nbitq), 
to_sfixed(-338623264.0/4294967296.0,1,-nbitq), 
to_sfixed(238127223.0/4294967296.0,1,-nbitq), 
to_sfixed(-100008483.0/4294967296.0,1,-nbitq), 
to_sfixed(236189876.0/4294967296.0,1,-nbitq), 
to_sfixed(400248156.0/4294967296.0,1,-nbitq), 
to_sfixed(715833446.0/4294967296.0,1,-nbitq), 
to_sfixed(73983581.0/4294967296.0,1,-nbitq), 
to_sfixed(-311032719.0/4294967296.0,1,-nbitq), 
to_sfixed(-260725654.0/4294967296.0,1,-nbitq), 
to_sfixed(-178392476.0/4294967296.0,1,-nbitq), 
to_sfixed(-111213305.0/4294967296.0,1,-nbitq), 
to_sfixed(464854898.0/4294967296.0,1,-nbitq), 
to_sfixed(-385411846.0/4294967296.0,1,-nbitq), 
to_sfixed(-31537605.0/4294967296.0,1,-nbitq), 
to_sfixed(-329571009.0/4294967296.0,1,-nbitq), 
to_sfixed(253636958.0/4294967296.0,1,-nbitq), 
to_sfixed(-120938794.0/4294967296.0,1,-nbitq), 
to_sfixed(277520231.0/4294967296.0,1,-nbitq), 
to_sfixed(-381166620.0/4294967296.0,1,-nbitq), 
to_sfixed(-440137828.0/4294967296.0,1,-nbitq), 
to_sfixed(339721259.0/4294967296.0,1,-nbitq), 
to_sfixed(-266741309.0/4294967296.0,1,-nbitq), 
to_sfixed(-77855154.0/4294967296.0,1,-nbitq), 
to_sfixed(106850433.0/4294967296.0,1,-nbitq), 
to_sfixed(-73324486.0/4294967296.0,1,-nbitq), 
to_sfixed(260899379.0/4294967296.0,1,-nbitq), 
to_sfixed(25923315.0/4294967296.0,1,-nbitq), 
to_sfixed(151540531.0/4294967296.0,1,-nbitq), 
to_sfixed(299736724.0/4294967296.0,1,-nbitq), 
to_sfixed(195286653.0/4294967296.0,1,-nbitq), 
to_sfixed(-135665234.0/4294967296.0,1,-nbitq), 
to_sfixed(266799422.0/4294967296.0,1,-nbitq), 
to_sfixed(-67800163.0/4294967296.0,1,-nbitq), 
to_sfixed(-452373891.0/4294967296.0,1,-nbitq), 
to_sfixed(477535009.0/4294967296.0,1,-nbitq), 
to_sfixed(-224820535.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-228855306.0/4294967296.0,1,-nbitq), 
to_sfixed(541994652.0/4294967296.0,1,-nbitq), 
to_sfixed(8488573.0/4294967296.0,1,-nbitq), 
to_sfixed(424441355.0/4294967296.0,1,-nbitq), 
to_sfixed(-766223875.0/4294967296.0,1,-nbitq), 
to_sfixed(-292518333.0/4294967296.0,1,-nbitq), 
to_sfixed(-405234513.0/4294967296.0,1,-nbitq), 
to_sfixed(-426801453.0/4294967296.0,1,-nbitq), 
to_sfixed(400674932.0/4294967296.0,1,-nbitq), 
to_sfixed(205613898.0/4294967296.0,1,-nbitq), 
to_sfixed(85408810.0/4294967296.0,1,-nbitq), 
to_sfixed(335827145.0/4294967296.0,1,-nbitq), 
to_sfixed(234939314.0/4294967296.0,1,-nbitq), 
to_sfixed(51398321.0/4294967296.0,1,-nbitq), 
to_sfixed(-230242715.0/4294967296.0,1,-nbitq), 
to_sfixed(240526991.0/4294967296.0,1,-nbitq), 
to_sfixed(249923230.0/4294967296.0,1,-nbitq), 
to_sfixed(265797846.0/4294967296.0,1,-nbitq), 
to_sfixed(125159801.0/4294967296.0,1,-nbitq), 
to_sfixed(-345629875.0/4294967296.0,1,-nbitq), 
to_sfixed(207025233.0/4294967296.0,1,-nbitq), 
to_sfixed(58939409.0/4294967296.0,1,-nbitq), 
to_sfixed(-171105799.0/4294967296.0,1,-nbitq), 
to_sfixed(197866694.0/4294967296.0,1,-nbitq), 
to_sfixed(376648068.0/4294967296.0,1,-nbitq), 
to_sfixed(387657970.0/4294967296.0,1,-nbitq), 
to_sfixed(-338869308.0/4294967296.0,1,-nbitq), 
to_sfixed(82183275.0/4294967296.0,1,-nbitq), 
to_sfixed(203430827.0/4294967296.0,1,-nbitq), 
to_sfixed(409973729.0/4294967296.0,1,-nbitq), 
to_sfixed(-223329878.0/4294967296.0,1,-nbitq), 
to_sfixed(175408089.0/4294967296.0,1,-nbitq), 
to_sfixed(431190451.0/4294967296.0,1,-nbitq), 
to_sfixed(-640792526.0/4294967296.0,1,-nbitq), 
to_sfixed(312699891.0/4294967296.0,1,-nbitq), 
to_sfixed(100894259.0/4294967296.0,1,-nbitq), 
to_sfixed(174936903.0/4294967296.0,1,-nbitq), 
to_sfixed(441716946.0/4294967296.0,1,-nbitq), 
to_sfixed(-480985119.0/4294967296.0,1,-nbitq), 
to_sfixed(-291044250.0/4294967296.0,1,-nbitq), 
to_sfixed(234776759.0/4294967296.0,1,-nbitq), 
to_sfixed(218592025.0/4294967296.0,1,-nbitq), 
to_sfixed(296464987.0/4294967296.0,1,-nbitq), 
to_sfixed(622627881.0/4294967296.0,1,-nbitq), 
to_sfixed(219029278.0/4294967296.0,1,-nbitq), 
to_sfixed(45858146.0/4294967296.0,1,-nbitq), 
to_sfixed(100702171.0/4294967296.0,1,-nbitq), 
to_sfixed(-201162969.0/4294967296.0,1,-nbitq), 
to_sfixed(187281108.0/4294967296.0,1,-nbitq), 
to_sfixed(79080342.0/4294967296.0,1,-nbitq), 
to_sfixed(-202723865.0/4294967296.0,1,-nbitq), 
to_sfixed(-451712301.0/4294967296.0,1,-nbitq), 
to_sfixed(42804877.0/4294967296.0,1,-nbitq), 
to_sfixed(146964857.0/4294967296.0,1,-nbitq), 
to_sfixed(-105821919.0/4294967296.0,1,-nbitq), 
to_sfixed(-238640049.0/4294967296.0,1,-nbitq), 
to_sfixed(-421577593.0/4294967296.0,1,-nbitq), 
to_sfixed(-194793536.0/4294967296.0,1,-nbitq), 
to_sfixed(-154433362.0/4294967296.0,1,-nbitq), 
to_sfixed(-86728899.0/4294967296.0,1,-nbitq), 
to_sfixed(-116385518.0/4294967296.0,1,-nbitq), 
to_sfixed(-302815025.0/4294967296.0,1,-nbitq), 
to_sfixed(182228039.0/4294967296.0,1,-nbitq), 
to_sfixed(312920044.0/4294967296.0,1,-nbitq), 
to_sfixed(-186641802.0/4294967296.0,1,-nbitq), 
to_sfixed(-371867085.0/4294967296.0,1,-nbitq), 
to_sfixed(574414812.0/4294967296.0,1,-nbitq), 
to_sfixed(638452681.0/4294967296.0,1,-nbitq), 
to_sfixed(-271998054.0/4294967296.0,1,-nbitq), 
to_sfixed(-434673529.0/4294967296.0,1,-nbitq), 
to_sfixed(76462131.0/4294967296.0,1,-nbitq), 
to_sfixed(-336566917.0/4294967296.0,1,-nbitq), 
to_sfixed(-245280683.0/4294967296.0,1,-nbitq), 
to_sfixed(122120638.0/4294967296.0,1,-nbitq), 
to_sfixed(-45215767.0/4294967296.0,1,-nbitq), 
to_sfixed(36632673.0/4294967296.0,1,-nbitq), 
to_sfixed(-390415588.0/4294967296.0,1,-nbitq), 
to_sfixed(88779387.0/4294967296.0,1,-nbitq), 
to_sfixed(557907093.0/4294967296.0,1,-nbitq), 
to_sfixed(116056024.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-204873076.0/4294967296.0,1,-nbitq), 
to_sfixed(257033046.0/4294967296.0,1,-nbitq), 
to_sfixed(24717491.0/4294967296.0,1,-nbitq), 
to_sfixed(-137960490.0/4294967296.0,1,-nbitq), 
to_sfixed(-345813707.0/4294967296.0,1,-nbitq), 
to_sfixed(-387234474.0/4294967296.0,1,-nbitq), 
to_sfixed(354305506.0/4294967296.0,1,-nbitq), 
to_sfixed(-14676811.0/4294967296.0,1,-nbitq), 
to_sfixed(607412473.0/4294967296.0,1,-nbitq), 
to_sfixed(318147184.0/4294967296.0,1,-nbitq), 
to_sfixed(-61670062.0/4294967296.0,1,-nbitq), 
to_sfixed(-46740469.0/4294967296.0,1,-nbitq), 
to_sfixed(10953807.0/4294967296.0,1,-nbitq), 
to_sfixed(34050037.0/4294967296.0,1,-nbitq), 
to_sfixed(-410221663.0/4294967296.0,1,-nbitq), 
to_sfixed(-371161654.0/4294967296.0,1,-nbitq), 
to_sfixed(-82756388.0/4294967296.0,1,-nbitq), 
to_sfixed(-35844977.0/4294967296.0,1,-nbitq), 
to_sfixed(-84201349.0/4294967296.0,1,-nbitq), 
to_sfixed(-34117677.0/4294967296.0,1,-nbitq), 
to_sfixed(166079561.0/4294967296.0,1,-nbitq), 
to_sfixed(337607105.0/4294967296.0,1,-nbitq), 
to_sfixed(333695389.0/4294967296.0,1,-nbitq), 
to_sfixed(171119066.0/4294967296.0,1,-nbitq), 
to_sfixed(418362007.0/4294967296.0,1,-nbitq), 
to_sfixed(-94216015.0/4294967296.0,1,-nbitq), 
to_sfixed(-390217815.0/4294967296.0,1,-nbitq), 
to_sfixed(-34507155.0/4294967296.0,1,-nbitq), 
to_sfixed(165157855.0/4294967296.0,1,-nbitq), 
to_sfixed(-349642394.0/4294967296.0,1,-nbitq), 
to_sfixed(-372882054.0/4294967296.0,1,-nbitq), 
to_sfixed(219242117.0/4294967296.0,1,-nbitq), 
to_sfixed(101096388.0/4294967296.0,1,-nbitq), 
to_sfixed(-578590025.0/4294967296.0,1,-nbitq), 
to_sfixed(-2770893.0/4294967296.0,1,-nbitq), 
to_sfixed(-55315201.0/4294967296.0,1,-nbitq), 
to_sfixed(361320851.0/4294967296.0,1,-nbitq), 
to_sfixed(386590665.0/4294967296.0,1,-nbitq), 
to_sfixed(-52551689.0/4294967296.0,1,-nbitq), 
to_sfixed(322613571.0/4294967296.0,1,-nbitq), 
to_sfixed(79320443.0/4294967296.0,1,-nbitq), 
to_sfixed(352343733.0/4294967296.0,1,-nbitq), 
to_sfixed(664684157.0/4294967296.0,1,-nbitq), 
to_sfixed(509263602.0/4294967296.0,1,-nbitq), 
to_sfixed(-39510231.0/4294967296.0,1,-nbitq), 
to_sfixed(342487007.0/4294967296.0,1,-nbitq), 
to_sfixed(195488567.0/4294967296.0,1,-nbitq), 
to_sfixed(327179351.0/4294967296.0,1,-nbitq), 
to_sfixed(-136364199.0/4294967296.0,1,-nbitq), 
to_sfixed(-128392792.0/4294967296.0,1,-nbitq), 
to_sfixed(386498985.0/4294967296.0,1,-nbitq), 
to_sfixed(-266181175.0/4294967296.0,1,-nbitq), 
to_sfixed(81579192.0/4294967296.0,1,-nbitq), 
to_sfixed(361047387.0/4294967296.0,1,-nbitq), 
to_sfixed(428645998.0/4294967296.0,1,-nbitq), 
to_sfixed(-259107581.0/4294967296.0,1,-nbitq), 
to_sfixed(-371008203.0/4294967296.0,1,-nbitq), 
to_sfixed(-499596026.0/4294967296.0,1,-nbitq), 
to_sfixed(3938086.0/4294967296.0,1,-nbitq), 
to_sfixed(-87908154.0/4294967296.0,1,-nbitq), 
to_sfixed(100758148.0/4294967296.0,1,-nbitq), 
to_sfixed(-149602372.0/4294967296.0,1,-nbitq), 
to_sfixed(-190693140.0/4294967296.0,1,-nbitq), 
to_sfixed(-404910254.0/4294967296.0,1,-nbitq), 
to_sfixed(-124379412.0/4294967296.0,1,-nbitq), 
to_sfixed(30688558.0/4294967296.0,1,-nbitq), 
to_sfixed(128246392.0/4294967296.0,1,-nbitq), 
to_sfixed(773230171.0/4294967296.0,1,-nbitq), 
to_sfixed(-181738054.0/4294967296.0,1,-nbitq), 
to_sfixed(-31441435.0/4294967296.0,1,-nbitq), 
to_sfixed(408039625.0/4294967296.0,1,-nbitq), 
to_sfixed(357399033.0/4294967296.0,1,-nbitq), 
to_sfixed(46712475.0/4294967296.0,1,-nbitq), 
to_sfixed(-334347434.0/4294967296.0,1,-nbitq), 
to_sfixed(220427937.0/4294967296.0,1,-nbitq), 
to_sfixed(54444788.0/4294967296.0,1,-nbitq), 
to_sfixed(116423086.0/4294967296.0,1,-nbitq), 
to_sfixed(-381378420.0/4294967296.0,1,-nbitq), 
to_sfixed(243868853.0/4294967296.0,1,-nbitq), 
to_sfixed(94217164.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-293200795.0/4294967296.0,1,-nbitq), 
to_sfixed(493225906.0/4294967296.0,1,-nbitq), 
to_sfixed(96176657.0/4294967296.0,1,-nbitq), 
to_sfixed(-37972887.0/4294967296.0,1,-nbitq), 
to_sfixed(-89406096.0/4294967296.0,1,-nbitq), 
to_sfixed(-167695676.0/4294967296.0,1,-nbitq), 
to_sfixed(-60572902.0/4294967296.0,1,-nbitq), 
to_sfixed(233036584.0/4294967296.0,1,-nbitq), 
to_sfixed(349074522.0/4294967296.0,1,-nbitq), 
to_sfixed(375811966.0/4294967296.0,1,-nbitq), 
to_sfixed(-405435318.0/4294967296.0,1,-nbitq), 
to_sfixed(-312708715.0/4294967296.0,1,-nbitq), 
to_sfixed(-523744321.0/4294967296.0,1,-nbitq), 
to_sfixed(138955601.0/4294967296.0,1,-nbitq), 
to_sfixed(-352716668.0/4294967296.0,1,-nbitq), 
to_sfixed(220738421.0/4294967296.0,1,-nbitq), 
to_sfixed(-415773325.0/4294967296.0,1,-nbitq), 
to_sfixed(129153373.0/4294967296.0,1,-nbitq), 
to_sfixed(190567649.0/4294967296.0,1,-nbitq), 
to_sfixed(215351593.0/4294967296.0,1,-nbitq), 
to_sfixed(373212891.0/4294967296.0,1,-nbitq), 
to_sfixed(-337544288.0/4294967296.0,1,-nbitq), 
to_sfixed(-208187070.0/4294967296.0,1,-nbitq), 
to_sfixed(331830733.0/4294967296.0,1,-nbitq), 
to_sfixed(-103047682.0/4294967296.0,1,-nbitq), 
to_sfixed(68968267.0/4294967296.0,1,-nbitq), 
to_sfixed(39099115.0/4294967296.0,1,-nbitq), 
to_sfixed(-351907981.0/4294967296.0,1,-nbitq), 
to_sfixed(-113082577.0/4294967296.0,1,-nbitq), 
to_sfixed(207794198.0/4294967296.0,1,-nbitq), 
to_sfixed(301226903.0/4294967296.0,1,-nbitq), 
to_sfixed(-523573410.0/4294967296.0,1,-nbitq), 
to_sfixed(503214772.0/4294967296.0,1,-nbitq), 
to_sfixed(-141513379.0/4294967296.0,1,-nbitq), 
to_sfixed(686369085.0/4294967296.0,1,-nbitq), 
to_sfixed(-251541794.0/4294967296.0,1,-nbitq), 
to_sfixed(552048851.0/4294967296.0,1,-nbitq), 
to_sfixed(-11501350.0/4294967296.0,1,-nbitq), 
to_sfixed(-451677629.0/4294967296.0,1,-nbitq), 
to_sfixed(417583853.0/4294967296.0,1,-nbitq), 
to_sfixed(111640293.0/4294967296.0,1,-nbitq), 
to_sfixed(156550342.0/4294967296.0,1,-nbitq), 
to_sfixed(381861965.0/4294967296.0,1,-nbitq), 
to_sfixed(782940242.0/4294967296.0,1,-nbitq), 
to_sfixed(-266153180.0/4294967296.0,1,-nbitq), 
to_sfixed(508030284.0/4294967296.0,1,-nbitq), 
to_sfixed(182464982.0/4294967296.0,1,-nbitq), 
to_sfixed(-382742581.0/4294967296.0,1,-nbitq), 
to_sfixed(44450677.0/4294967296.0,1,-nbitq), 
to_sfixed(348692888.0/4294967296.0,1,-nbitq), 
to_sfixed(445005068.0/4294967296.0,1,-nbitq), 
to_sfixed(38501115.0/4294967296.0,1,-nbitq), 
to_sfixed(8949011.0/4294967296.0,1,-nbitq), 
to_sfixed(734098893.0/4294967296.0,1,-nbitq), 
to_sfixed(191131447.0/4294967296.0,1,-nbitq), 
to_sfixed(-146516076.0/4294967296.0,1,-nbitq), 
to_sfixed(-153768422.0/4294967296.0,1,-nbitq), 
to_sfixed(23821107.0/4294967296.0,1,-nbitq), 
to_sfixed(8940485.0/4294967296.0,1,-nbitq), 
to_sfixed(-190991418.0/4294967296.0,1,-nbitq), 
to_sfixed(-337251091.0/4294967296.0,1,-nbitq), 
to_sfixed(-421079657.0/4294967296.0,1,-nbitq), 
to_sfixed(62199759.0/4294967296.0,1,-nbitq), 
to_sfixed(-83858134.0/4294967296.0,1,-nbitq), 
to_sfixed(563870645.0/4294967296.0,1,-nbitq), 
to_sfixed(-354333803.0/4294967296.0,1,-nbitq), 
to_sfixed(293655995.0/4294967296.0,1,-nbitq), 
to_sfixed(716644918.0/4294967296.0,1,-nbitq), 
to_sfixed(-98120780.0/4294967296.0,1,-nbitq), 
to_sfixed(165991814.0/4294967296.0,1,-nbitq), 
to_sfixed(225896014.0/4294967296.0,1,-nbitq), 
to_sfixed(184398132.0/4294967296.0,1,-nbitq), 
to_sfixed(2205348.0/4294967296.0,1,-nbitq), 
to_sfixed(-32339126.0/4294967296.0,1,-nbitq), 
to_sfixed(-156491698.0/4294967296.0,1,-nbitq), 
to_sfixed(-144925680.0/4294967296.0,1,-nbitq), 
to_sfixed(204806241.0/4294967296.0,1,-nbitq), 
to_sfixed(-445801951.0/4294967296.0,1,-nbitq), 
to_sfixed(65606578.0/4294967296.0,1,-nbitq), 
to_sfixed(-13844900.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(55480654.0/4294967296.0,1,-nbitq), 
to_sfixed(156282874.0/4294967296.0,1,-nbitq), 
to_sfixed(328446336.0/4294967296.0,1,-nbitq), 
to_sfixed(245330487.0/4294967296.0,1,-nbitq), 
to_sfixed(-544717223.0/4294967296.0,1,-nbitq), 
to_sfixed(61173106.0/4294967296.0,1,-nbitq), 
to_sfixed(-101553116.0/4294967296.0,1,-nbitq), 
to_sfixed(-192152401.0/4294967296.0,1,-nbitq), 
to_sfixed(423973277.0/4294967296.0,1,-nbitq), 
to_sfixed(73706488.0/4294967296.0,1,-nbitq), 
to_sfixed(-9206449.0/4294967296.0,1,-nbitq), 
to_sfixed(-173710050.0/4294967296.0,1,-nbitq), 
to_sfixed(-519073377.0/4294967296.0,1,-nbitq), 
to_sfixed(23292706.0/4294967296.0,1,-nbitq), 
to_sfixed(71602609.0/4294967296.0,1,-nbitq), 
to_sfixed(-150596540.0/4294967296.0,1,-nbitq), 
to_sfixed(-282554831.0/4294967296.0,1,-nbitq), 
to_sfixed(69828832.0/4294967296.0,1,-nbitq), 
to_sfixed(524387001.0/4294967296.0,1,-nbitq), 
to_sfixed(-298265305.0/4294967296.0,1,-nbitq), 
to_sfixed(-361589113.0/4294967296.0,1,-nbitq), 
to_sfixed(-255842126.0/4294967296.0,1,-nbitq), 
to_sfixed(-50348109.0/4294967296.0,1,-nbitq), 
to_sfixed(-119742053.0/4294967296.0,1,-nbitq), 
to_sfixed(268306673.0/4294967296.0,1,-nbitq), 
to_sfixed(-45486130.0/4294967296.0,1,-nbitq), 
to_sfixed(130692179.0/4294967296.0,1,-nbitq), 
to_sfixed(-47813212.0/4294967296.0,1,-nbitq), 
to_sfixed(381922811.0/4294967296.0,1,-nbitq), 
to_sfixed(-24679033.0/4294967296.0,1,-nbitq), 
to_sfixed(-291393768.0/4294967296.0,1,-nbitq), 
to_sfixed(-335275501.0/4294967296.0,1,-nbitq), 
to_sfixed(-185088.0/4294967296.0,1,-nbitq), 
to_sfixed(-218233436.0/4294967296.0,1,-nbitq), 
to_sfixed(550796727.0/4294967296.0,1,-nbitq), 
to_sfixed(-187819538.0/4294967296.0,1,-nbitq), 
to_sfixed(265864882.0/4294967296.0,1,-nbitq), 
to_sfixed(390597863.0/4294967296.0,1,-nbitq), 
to_sfixed(265371896.0/4294967296.0,1,-nbitq), 
to_sfixed(66575684.0/4294967296.0,1,-nbitq), 
to_sfixed(-8872333.0/4294967296.0,1,-nbitq), 
to_sfixed(-116165593.0/4294967296.0,1,-nbitq), 
to_sfixed(384391441.0/4294967296.0,1,-nbitq), 
to_sfixed(136219904.0/4294967296.0,1,-nbitq), 
to_sfixed(67574185.0/4294967296.0,1,-nbitq), 
to_sfixed(-133150575.0/4294967296.0,1,-nbitq), 
to_sfixed(-125560689.0/4294967296.0,1,-nbitq), 
to_sfixed(304626175.0/4294967296.0,1,-nbitq), 
to_sfixed(273078634.0/4294967296.0,1,-nbitq), 
to_sfixed(370276698.0/4294967296.0,1,-nbitq), 
to_sfixed(-99638181.0/4294967296.0,1,-nbitq), 
to_sfixed(97074657.0/4294967296.0,1,-nbitq), 
to_sfixed(-347374536.0/4294967296.0,1,-nbitq), 
to_sfixed(458177.0/4294967296.0,1,-nbitq), 
to_sfixed(329690085.0/4294967296.0,1,-nbitq), 
to_sfixed(367539413.0/4294967296.0,1,-nbitq), 
to_sfixed(-681428656.0/4294967296.0,1,-nbitq), 
to_sfixed(-277404626.0/4294967296.0,1,-nbitq), 
to_sfixed(286451213.0/4294967296.0,1,-nbitq), 
to_sfixed(136417745.0/4294967296.0,1,-nbitq), 
to_sfixed(151185795.0/4294967296.0,1,-nbitq), 
to_sfixed(-398911408.0/4294967296.0,1,-nbitq), 
to_sfixed(-36001326.0/4294967296.0,1,-nbitq), 
to_sfixed(-321517105.0/4294967296.0,1,-nbitq), 
to_sfixed(-67787749.0/4294967296.0,1,-nbitq), 
to_sfixed(-60388305.0/4294967296.0,1,-nbitq), 
to_sfixed(-312012292.0/4294967296.0,1,-nbitq), 
to_sfixed(809414417.0/4294967296.0,1,-nbitq), 
to_sfixed(259843567.0/4294967296.0,1,-nbitq), 
to_sfixed(-262882476.0/4294967296.0,1,-nbitq), 
to_sfixed(526238491.0/4294967296.0,1,-nbitq), 
to_sfixed(-59913314.0/4294967296.0,1,-nbitq), 
to_sfixed(-184251892.0/4294967296.0,1,-nbitq), 
to_sfixed(-162059752.0/4294967296.0,1,-nbitq), 
to_sfixed(-153185843.0/4294967296.0,1,-nbitq), 
to_sfixed(54775789.0/4294967296.0,1,-nbitq), 
to_sfixed(228322904.0/4294967296.0,1,-nbitq), 
to_sfixed(-49793846.0/4294967296.0,1,-nbitq), 
to_sfixed(579406393.0/4294967296.0,1,-nbitq), 
to_sfixed(340389186.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(178294717.0/4294967296.0,1,-nbitq), 
to_sfixed(695001734.0/4294967296.0,1,-nbitq), 
to_sfixed(-367247236.0/4294967296.0,1,-nbitq), 
to_sfixed(-167909079.0/4294967296.0,1,-nbitq), 
to_sfixed(81059694.0/4294967296.0,1,-nbitq), 
to_sfixed(331410996.0/4294967296.0,1,-nbitq), 
to_sfixed(-247069955.0/4294967296.0,1,-nbitq), 
to_sfixed(156904825.0/4294967296.0,1,-nbitq), 
to_sfixed(485226361.0/4294967296.0,1,-nbitq), 
to_sfixed(-42506065.0/4294967296.0,1,-nbitq), 
to_sfixed(-528169681.0/4294967296.0,1,-nbitq), 
to_sfixed(-329582555.0/4294967296.0,1,-nbitq), 
to_sfixed(-928245659.0/4294967296.0,1,-nbitq), 
to_sfixed(335912118.0/4294967296.0,1,-nbitq), 
to_sfixed(-113874686.0/4294967296.0,1,-nbitq), 
to_sfixed(-9931346.0/4294967296.0,1,-nbitq), 
to_sfixed(-242636201.0/4294967296.0,1,-nbitq), 
to_sfixed(239787501.0/4294967296.0,1,-nbitq), 
to_sfixed(-30533499.0/4294967296.0,1,-nbitq), 
to_sfixed(-212223415.0/4294967296.0,1,-nbitq), 
to_sfixed(63969296.0/4294967296.0,1,-nbitq), 
to_sfixed(3364565.0/4294967296.0,1,-nbitq), 
to_sfixed(550274169.0/4294967296.0,1,-nbitq), 
to_sfixed(108475349.0/4294967296.0,1,-nbitq), 
to_sfixed(273084248.0/4294967296.0,1,-nbitq), 
to_sfixed(-257454387.0/4294967296.0,1,-nbitq), 
to_sfixed(-161399122.0/4294967296.0,1,-nbitq), 
to_sfixed(-55679237.0/4294967296.0,1,-nbitq), 
to_sfixed(-101768756.0/4294967296.0,1,-nbitq), 
to_sfixed(428237518.0/4294967296.0,1,-nbitq), 
to_sfixed(-623791963.0/4294967296.0,1,-nbitq), 
to_sfixed(-402218363.0/4294967296.0,1,-nbitq), 
to_sfixed(-48261936.0/4294967296.0,1,-nbitq), 
to_sfixed(-92320152.0/4294967296.0,1,-nbitq), 
to_sfixed(506037365.0/4294967296.0,1,-nbitq), 
to_sfixed(95843020.0/4294967296.0,1,-nbitq), 
to_sfixed(373480864.0/4294967296.0,1,-nbitq), 
to_sfixed(-291207512.0/4294967296.0,1,-nbitq), 
to_sfixed(-37757729.0/4294967296.0,1,-nbitq), 
to_sfixed(-268860285.0/4294967296.0,1,-nbitq), 
to_sfixed(-372942148.0/4294967296.0,1,-nbitq), 
to_sfixed(225357492.0/4294967296.0,1,-nbitq), 
to_sfixed(-46399394.0/4294967296.0,1,-nbitq), 
to_sfixed(-34167711.0/4294967296.0,1,-nbitq), 
to_sfixed(123513071.0/4294967296.0,1,-nbitq), 
to_sfixed(-124532927.0/4294967296.0,1,-nbitq), 
to_sfixed(124177007.0/4294967296.0,1,-nbitq), 
to_sfixed(191210.0/4294967296.0,1,-nbitq), 
to_sfixed(546171379.0/4294967296.0,1,-nbitq), 
to_sfixed(-14433852.0/4294967296.0,1,-nbitq), 
to_sfixed(136891404.0/4294967296.0,1,-nbitq), 
to_sfixed(-156985486.0/4294967296.0,1,-nbitq), 
to_sfixed(-335654215.0/4294967296.0,1,-nbitq), 
to_sfixed(337064865.0/4294967296.0,1,-nbitq), 
to_sfixed(-278155299.0/4294967296.0,1,-nbitq), 
to_sfixed(-182473567.0/4294967296.0,1,-nbitq), 
to_sfixed(200032755.0/4294967296.0,1,-nbitq), 
to_sfixed(220013754.0/4294967296.0,1,-nbitq), 
to_sfixed(267662896.0/4294967296.0,1,-nbitq), 
to_sfixed(163099800.0/4294967296.0,1,-nbitq), 
to_sfixed(-110856385.0/4294967296.0,1,-nbitq), 
to_sfixed(158299175.0/4294967296.0,1,-nbitq), 
to_sfixed(114870536.0/4294967296.0,1,-nbitq), 
to_sfixed(290006693.0/4294967296.0,1,-nbitq), 
to_sfixed(349987957.0/4294967296.0,1,-nbitq), 
to_sfixed(-49340857.0/4294967296.0,1,-nbitq), 
to_sfixed(-225572767.0/4294967296.0,1,-nbitq), 
to_sfixed(-28308470.0/4294967296.0,1,-nbitq), 
to_sfixed(-313931244.0/4294967296.0,1,-nbitq), 
to_sfixed(99391168.0/4294967296.0,1,-nbitq), 
to_sfixed(386656470.0/4294967296.0,1,-nbitq), 
to_sfixed(-2134850.0/4294967296.0,1,-nbitq), 
to_sfixed(-651265735.0/4294967296.0,1,-nbitq), 
to_sfixed(-42809322.0/4294967296.0,1,-nbitq), 
to_sfixed(-206302436.0/4294967296.0,1,-nbitq), 
to_sfixed(266707828.0/4294967296.0,1,-nbitq), 
to_sfixed(265090971.0/4294967296.0,1,-nbitq), 
to_sfixed(-235061194.0/4294967296.0,1,-nbitq), 
to_sfixed(462912970.0/4294967296.0,1,-nbitq), 
to_sfixed(267247396.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-129900761.0/4294967296.0,1,-nbitq), 
to_sfixed(227852094.0/4294967296.0,1,-nbitq), 
to_sfixed(319960911.0/4294967296.0,1,-nbitq), 
to_sfixed(-6733330.0/4294967296.0,1,-nbitq), 
to_sfixed(-110178235.0/4294967296.0,1,-nbitq), 
to_sfixed(-8317114.0/4294967296.0,1,-nbitq), 
to_sfixed(72430988.0/4294967296.0,1,-nbitq), 
to_sfixed(-373271768.0/4294967296.0,1,-nbitq), 
to_sfixed(-222992665.0/4294967296.0,1,-nbitq), 
to_sfixed(210003144.0/4294967296.0,1,-nbitq), 
to_sfixed(194819330.0/4294967296.0,1,-nbitq), 
to_sfixed(533449503.0/4294967296.0,1,-nbitq), 
to_sfixed(-660502586.0/4294967296.0,1,-nbitq), 
to_sfixed(576954374.0/4294967296.0,1,-nbitq), 
to_sfixed(-171393316.0/4294967296.0,1,-nbitq), 
to_sfixed(-143542561.0/4294967296.0,1,-nbitq), 
to_sfixed(-393192970.0/4294967296.0,1,-nbitq), 
to_sfixed(429666339.0/4294967296.0,1,-nbitq), 
to_sfixed(257856006.0/4294967296.0,1,-nbitq), 
to_sfixed(-321308701.0/4294967296.0,1,-nbitq), 
to_sfixed(327071387.0/4294967296.0,1,-nbitq), 
to_sfixed(-169560423.0/4294967296.0,1,-nbitq), 
to_sfixed(447859879.0/4294967296.0,1,-nbitq), 
to_sfixed(130934999.0/4294967296.0,1,-nbitq), 
to_sfixed(384024743.0/4294967296.0,1,-nbitq), 
to_sfixed(149128400.0/4294967296.0,1,-nbitq), 
to_sfixed(-405793527.0/4294967296.0,1,-nbitq), 
to_sfixed(-113218499.0/4294967296.0,1,-nbitq), 
to_sfixed(10481691.0/4294967296.0,1,-nbitq), 
to_sfixed(359802728.0/4294967296.0,1,-nbitq), 
to_sfixed(-372383141.0/4294967296.0,1,-nbitq), 
to_sfixed(-722990913.0/4294967296.0,1,-nbitq), 
to_sfixed(-27934426.0/4294967296.0,1,-nbitq), 
to_sfixed(-64465613.0/4294967296.0,1,-nbitq), 
to_sfixed(264590510.0/4294967296.0,1,-nbitq), 
to_sfixed(-146569678.0/4294967296.0,1,-nbitq), 
to_sfixed(427326411.0/4294967296.0,1,-nbitq), 
to_sfixed(-126612459.0/4294967296.0,1,-nbitq), 
to_sfixed(16963379.0/4294967296.0,1,-nbitq), 
to_sfixed(-136695414.0/4294967296.0,1,-nbitq), 
to_sfixed(-225944433.0/4294967296.0,1,-nbitq), 
to_sfixed(61642009.0/4294967296.0,1,-nbitq), 
to_sfixed(543458856.0/4294967296.0,1,-nbitq), 
to_sfixed(175149455.0/4294967296.0,1,-nbitq), 
to_sfixed(-273512601.0/4294967296.0,1,-nbitq), 
to_sfixed(-136125777.0/4294967296.0,1,-nbitq), 
to_sfixed(169464637.0/4294967296.0,1,-nbitq), 
to_sfixed(114992376.0/4294967296.0,1,-nbitq), 
to_sfixed(339611646.0/4294967296.0,1,-nbitq), 
to_sfixed(-128344981.0/4294967296.0,1,-nbitq), 
to_sfixed(-349763426.0/4294967296.0,1,-nbitq), 
to_sfixed(117880117.0/4294967296.0,1,-nbitq), 
to_sfixed(-92648237.0/4294967296.0,1,-nbitq), 
to_sfixed(-353028794.0/4294967296.0,1,-nbitq), 
to_sfixed(76598870.0/4294967296.0,1,-nbitq), 
to_sfixed(-124060517.0/4294967296.0,1,-nbitq), 
to_sfixed(90942248.0/4294967296.0,1,-nbitq), 
to_sfixed(-136865665.0/4294967296.0,1,-nbitq), 
to_sfixed(158349492.0/4294967296.0,1,-nbitq), 
to_sfixed(-264571119.0/4294967296.0,1,-nbitq), 
to_sfixed(-175417669.0/4294967296.0,1,-nbitq), 
to_sfixed(145958902.0/4294967296.0,1,-nbitq), 
to_sfixed(197308539.0/4294967296.0,1,-nbitq), 
to_sfixed(89366831.0/4294967296.0,1,-nbitq), 
to_sfixed(17712188.0/4294967296.0,1,-nbitq), 
to_sfixed(-430686463.0/4294967296.0,1,-nbitq), 
to_sfixed(-99638412.0/4294967296.0,1,-nbitq), 
to_sfixed(-348993602.0/4294967296.0,1,-nbitq), 
to_sfixed(-234733137.0/4294967296.0,1,-nbitq), 
to_sfixed(192866837.0/4294967296.0,1,-nbitq), 
to_sfixed(-315767205.0/4294967296.0,1,-nbitq), 
to_sfixed(327130745.0/4294967296.0,1,-nbitq), 
to_sfixed(107002367.0/4294967296.0,1,-nbitq), 
to_sfixed(112857602.0/4294967296.0,1,-nbitq), 
to_sfixed(444408867.0/4294967296.0,1,-nbitq), 
to_sfixed(-341216115.0/4294967296.0,1,-nbitq), 
to_sfixed(176394030.0/4294967296.0,1,-nbitq), 
to_sfixed(182874006.0/4294967296.0,1,-nbitq), 
to_sfixed(84349749.0/4294967296.0,1,-nbitq), 
to_sfixed(-148599849.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-401348452.0/4294967296.0,1,-nbitq), 
to_sfixed(74882396.0/4294967296.0,1,-nbitq), 
to_sfixed(-125507871.0/4294967296.0,1,-nbitq), 
to_sfixed(-485011228.0/4294967296.0,1,-nbitq), 
to_sfixed(-17489104.0/4294967296.0,1,-nbitq), 
to_sfixed(158524646.0/4294967296.0,1,-nbitq), 
to_sfixed(-347980263.0/4294967296.0,1,-nbitq), 
to_sfixed(89407106.0/4294967296.0,1,-nbitq), 
to_sfixed(-42062602.0/4294967296.0,1,-nbitq), 
to_sfixed(-321872921.0/4294967296.0,1,-nbitq), 
to_sfixed(107354487.0/4294967296.0,1,-nbitq), 
to_sfixed(348525857.0/4294967296.0,1,-nbitq), 
to_sfixed(-405739949.0/4294967296.0,1,-nbitq), 
to_sfixed(282520203.0/4294967296.0,1,-nbitq), 
to_sfixed(-204454498.0/4294967296.0,1,-nbitq), 
to_sfixed(-79970413.0/4294967296.0,1,-nbitq), 
to_sfixed(-343916711.0/4294967296.0,1,-nbitq), 
to_sfixed(163707895.0/4294967296.0,1,-nbitq), 
to_sfixed(93608188.0/4294967296.0,1,-nbitq), 
to_sfixed(-192527081.0/4294967296.0,1,-nbitq), 
to_sfixed(-179506493.0/4294967296.0,1,-nbitq), 
to_sfixed(243830826.0/4294967296.0,1,-nbitq), 
to_sfixed(235730553.0/4294967296.0,1,-nbitq), 
to_sfixed(261024462.0/4294967296.0,1,-nbitq), 
to_sfixed(-264438042.0/4294967296.0,1,-nbitq), 
to_sfixed(-215145942.0/4294967296.0,1,-nbitq), 
to_sfixed(-172405401.0/4294967296.0,1,-nbitq), 
to_sfixed(-469041222.0/4294967296.0,1,-nbitq), 
to_sfixed(-71777409.0/4294967296.0,1,-nbitq), 
to_sfixed(161630341.0/4294967296.0,1,-nbitq), 
to_sfixed(122890512.0/4294967296.0,1,-nbitq), 
to_sfixed(-271742398.0/4294967296.0,1,-nbitq), 
to_sfixed(-21139763.0/4294967296.0,1,-nbitq), 
to_sfixed(-327661378.0/4294967296.0,1,-nbitq), 
to_sfixed(339148121.0/4294967296.0,1,-nbitq), 
to_sfixed(117899727.0/4294967296.0,1,-nbitq), 
to_sfixed(-50809240.0/4294967296.0,1,-nbitq), 
to_sfixed(-291158967.0/4294967296.0,1,-nbitq), 
to_sfixed(368613721.0/4294967296.0,1,-nbitq), 
to_sfixed(-32160904.0/4294967296.0,1,-nbitq), 
to_sfixed(44350692.0/4294967296.0,1,-nbitq), 
to_sfixed(-64457171.0/4294967296.0,1,-nbitq), 
to_sfixed(-74026311.0/4294967296.0,1,-nbitq), 
to_sfixed(139301241.0/4294967296.0,1,-nbitq), 
to_sfixed(242097561.0/4294967296.0,1,-nbitq), 
to_sfixed(64569115.0/4294967296.0,1,-nbitq), 
to_sfixed(-94979594.0/4294967296.0,1,-nbitq), 
to_sfixed(-220451209.0/4294967296.0,1,-nbitq), 
to_sfixed(-94944124.0/4294967296.0,1,-nbitq), 
to_sfixed(-263799125.0/4294967296.0,1,-nbitq), 
to_sfixed(163217996.0/4294967296.0,1,-nbitq), 
to_sfixed(-7842130.0/4294967296.0,1,-nbitq), 
to_sfixed(-215857602.0/4294967296.0,1,-nbitq), 
to_sfixed(-193389615.0/4294967296.0,1,-nbitq), 
to_sfixed(432446048.0/4294967296.0,1,-nbitq), 
to_sfixed(-81530069.0/4294967296.0,1,-nbitq), 
to_sfixed(-161462331.0/4294967296.0,1,-nbitq), 
to_sfixed(208392514.0/4294967296.0,1,-nbitq), 
to_sfixed(-265335146.0/4294967296.0,1,-nbitq), 
to_sfixed(389321805.0/4294967296.0,1,-nbitq), 
to_sfixed(358918948.0/4294967296.0,1,-nbitq), 
to_sfixed(192719460.0/4294967296.0,1,-nbitq), 
to_sfixed(-314734684.0/4294967296.0,1,-nbitq), 
to_sfixed(-236843573.0/4294967296.0,1,-nbitq), 
to_sfixed(-238067859.0/4294967296.0,1,-nbitq), 
to_sfixed(262229344.0/4294967296.0,1,-nbitq), 
to_sfixed(-11201634.0/4294967296.0,1,-nbitq), 
to_sfixed(-124744969.0/4294967296.0,1,-nbitq), 
to_sfixed(-278096826.0/4294967296.0,1,-nbitq), 
to_sfixed(303166596.0/4294967296.0,1,-nbitq), 
to_sfixed(-58795954.0/4294967296.0,1,-nbitq), 
to_sfixed(136790005.0/4294967296.0,1,-nbitq), 
to_sfixed(-361389575.0/4294967296.0,1,-nbitq), 
to_sfixed(150335768.0/4294967296.0,1,-nbitq), 
to_sfixed(179371980.0/4294967296.0,1,-nbitq), 
to_sfixed(164015051.0/4294967296.0,1,-nbitq), 
to_sfixed(-91224939.0/4294967296.0,1,-nbitq), 
to_sfixed(-189423572.0/4294967296.0,1,-nbitq), 
to_sfixed(-345724112.0/4294967296.0,1,-nbitq), 
to_sfixed(334131220.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(249683452.0/4294967296.0,1,-nbitq), 
to_sfixed(182259148.0/4294967296.0,1,-nbitq), 
to_sfixed(232493193.0/4294967296.0,1,-nbitq), 
to_sfixed(-356394540.0/4294967296.0,1,-nbitq), 
to_sfixed(-90639214.0/4294967296.0,1,-nbitq), 
to_sfixed(11265390.0/4294967296.0,1,-nbitq), 
to_sfixed(-110895537.0/4294967296.0,1,-nbitq), 
to_sfixed(-305544937.0/4294967296.0,1,-nbitq), 
to_sfixed(-381975205.0/4294967296.0,1,-nbitq), 
to_sfixed(-173094275.0/4294967296.0,1,-nbitq), 
to_sfixed(-225403978.0/4294967296.0,1,-nbitq), 
to_sfixed(111775595.0/4294967296.0,1,-nbitq), 
to_sfixed(278168422.0/4294967296.0,1,-nbitq), 
to_sfixed(459225059.0/4294967296.0,1,-nbitq), 
to_sfixed(-329756479.0/4294967296.0,1,-nbitq), 
to_sfixed(-269873316.0/4294967296.0,1,-nbitq), 
to_sfixed(230226570.0/4294967296.0,1,-nbitq), 
to_sfixed(-63273677.0/4294967296.0,1,-nbitq), 
to_sfixed(294459279.0/4294967296.0,1,-nbitq), 
to_sfixed(-44049156.0/4294967296.0,1,-nbitq), 
to_sfixed(-323160679.0/4294967296.0,1,-nbitq), 
to_sfixed(114576742.0/4294967296.0,1,-nbitq), 
to_sfixed(580331686.0/4294967296.0,1,-nbitq), 
to_sfixed(354173187.0/4294967296.0,1,-nbitq), 
to_sfixed(235523222.0/4294967296.0,1,-nbitq), 
to_sfixed(573708725.0/4294967296.0,1,-nbitq), 
to_sfixed(-4135355.0/4294967296.0,1,-nbitq), 
to_sfixed(-7314436.0/4294967296.0,1,-nbitq), 
to_sfixed(85710800.0/4294967296.0,1,-nbitq), 
to_sfixed(-92746044.0/4294967296.0,1,-nbitq), 
to_sfixed(-477462742.0/4294967296.0,1,-nbitq), 
to_sfixed(-202876275.0/4294967296.0,1,-nbitq), 
to_sfixed(-129680003.0/4294967296.0,1,-nbitq), 
to_sfixed(-150790546.0/4294967296.0,1,-nbitq), 
to_sfixed(68930884.0/4294967296.0,1,-nbitq), 
to_sfixed(-277500813.0/4294967296.0,1,-nbitq), 
to_sfixed(-74806521.0/4294967296.0,1,-nbitq), 
to_sfixed(-1517240.0/4294967296.0,1,-nbitq), 
to_sfixed(61126957.0/4294967296.0,1,-nbitq), 
to_sfixed(89059974.0/4294967296.0,1,-nbitq), 
to_sfixed(220817808.0/4294967296.0,1,-nbitq), 
to_sfixed(133403713.0/4294967296.0,1,-nbitq), 
to_sfixed(29475657.0/4294967296.0,1,-nbitq), 
to_sfixed(-349052521.0/4294967296.0,1,-nbitq), 
to_sfixed(276037226.0/4294967296.0,1,-nbitq), 
to_sfixed(435887215.0/4294967296.0,1,-nbitq), 
to_sfixed(-269212496.0/4294967296.0,1,-nbitq), 
to_sfixed(-377805582.0/4294967296.0,1,-nbitq), 
to_sfixed(13033389.0/4294967296.0,1,-nbitq), 
to_sfixed(206879149.0/4294967296.0,1,-nbitq), 
to_sfixed(-54058483.0/4294967296.0,1,-nbitq), 
to_sfixed(83804284.0/4294967296.0,1,-nbitq), 
to_sfixed(98995869.0/4294967296.0,1,-nbitq), 
to_sfixed(285789010.0/4294967296.0,1,-nbitq), 
to_sfixed(325028999.0/4294967296.0,1,-nbitq), 
to_sfixed(360265280.0/4294967296.0,1,-nbitq), 
to_sfixed(95937284.0/4294967296.0,1,-nbitq), 
to_sfixed(147308814.0/4294967296.0,1,-nbitq), 
to_sfixed(142066279.0/4294967296.0,1,-nbitq), 
to_sfixed(170161168.0/4294967296.0,1,-nbitq), 
to_sfixed(-108859391.0/4294967296.0,1,-nbitq), 
to_sfixed(-172317667.0/4294967296.0,1,-nbitq), 
to_sfixed(-318097627.0/4294967296.0,1,-nbitq), 
to_sfixed(281992969.0/4294967296.0,1,-nbitq), 
to_sfixed(-266325068.0/4294967296.0,1,-nbitq), 
to_sfixed(203813628.0/4294967296.0,1,-nbitq), 
to_sfixed(666676298.0/4294967296.0,1,-nbitq), 
to_sfixed(7118464.0/4294967296.0,1,-nbitq), 
to_sfixed(-338181098.0/4294967296.0,1,-nbitq), 
to_sfixed(-191148239.0/4294967296.0,1,-nbitq), 
to_sfixed(105452076.0/4294967296.0,1,-nbitq), 
to_sfixed(-284864193.0/4294967296.0,1,-nbitq), 
to_sfixed(-276661459.0/4294967296.0,1,-nbitq), 
to_sfixed(461962592.0/4294967296.0,1,-nbitq), 
to_sfixed(-7015784.0/4294967296.0,1,-nbitq), 
to_sfixed(-318149385.0/4294967296.0,1,-nbitq), 
to_sfixed(-142747181.0/4294967296.0,1,-nbitq), 
to_sfixed(-458516785.0/4294967296.0,1,-nbitq), 
to_sfixed(-310314338.0/4294967296.0,1,-nbitq), 
to_sfixed(-362507433.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(262069422.0/4294967296.0,1,-nbitq), 
to_sfixed(330084732.0/4294967296.0,1,-nbitq), 
to_sfixed(201641480.0/4294967296.0,1,-nbitq), 
to_sfixed(-275763895.0/4294967296.0,1,-nbitq), 
to_sfixed(91177715.0/4294967296.0,1,-nbitq), 
to_sfixed(-23542500.0/4294967296.0,1,-nbitq), 
to_sfixed(-260575894.0/4294967296.0,1,-nbitq), 
to_sfixed(6127105.0/4294967296.0,1,-nbitq), 
to_sfixed(-178834423.0/4294967296.0,1,-nbitq), 
to_sfixed(52827679.0/4294967296.0,1,-nbitq), 
to_sfixed(-65446578.0/4294967296.0,1,-nbitq), 
to_sfixed(366036427.0/4294967296.0,1,-nbitq), 
to_sfixed(-31091853.0/4294967296.0,1,-nbitq), 
to_sfixed(437815553.0/4294967296.0,1,-nbitq), 
to_sfixed(-388913210.0/4294967296.0,1,-nbitq), 
to_sfixed(-48326727.0/4294967296.0,1,-nbitq), 
to_sfixed(295504226.0/4294967296.0,1,-nbitq), 
to_sfixed(-310743147.0/4294967296.0,1,-nbitq), 
to_sfixed(-155115196.0/4294967296.0,1,-nbitq), 
to_sfixed(-316487697.0/4294967296.0,1,-nbitq), 
to_sfixed(-182336382.0/4294967296.0,1,-nbitq), 
to_sfixed(243360410.0/4294967296.0,1,-nbitq), 
to_sfixed(425484972.0/4294967296.0,1,-nbitq), 
to_sfixed(-135469249.0/4294967296.0,1,-nbitq), 
to_sfixed(-254491230.0/4294967296.0,1,-nbitq), 
to_sfixed(-62182158.0/4294967296.0,1,-nbitq), 
to_sfixed(-305508232.0/4294967296.0,1,-nbitq), 
to_sfixed(20702505.0/4294967296.0,1,-nbitq), 
to_sfixed(-249793138.0/4294967296.0,1,-nbitq), 
to_sfixed(50039482.0/4294967296.0,1,-nbitq), 
to_sfixed(-5069270.0/4294967296.0,1,-nbitq), 
to_sfixed(-274343707.0/4294967296.0,1,-nbitq), 
to_sfixed(16052532.0/4294967296.0,1,-nbitq), 
to_sfixed(40945586.0/4294967296.0,1,-nbitq), 
to_sfixed(-113168209.0/4294967296.0,1,-nbitq), 
to_sfixed(161196955.0/4294967296.0,1,-nbitq), 
to_sfixed(325311111.0/4294967296.0,1,-nbitq), 
to_sfixed(86735412.0/4294967296.0,1,-nbitq), 
to_sfixed(21111455.0/4294967296.0,1,-nbitq), 
to_sfixed(161306571.0/4294967296.0,1,-nbitq), 
to_sfixed(125049319.0/4294967296.0,1,-nbitq), 
to_sfixed(33539705.0/4294967296.0,1,-nbitq), 
to_sfixed(-107832814.0/4294967296.0,1,-nbitq), 
to_sfixed(-349200590.0/4294967296.0,1,-nbitq), 
to_sfixed(-375680450.0/4294967296.0,1,-nbitq), 
to_sfixed(-78707458.0/4294967296.0,1,-nbitq), 
to_sfixed(235579353.0/4294967296.0,1,-nbitq), 
to_sfixed(-40074653.0/4294967296.0,1,-nbitq), 
to_sfixed(-252792745.0/4294967296.0,1,-nbitq), 
to_sfixed(-106539327.0/4294967296.0,1,-nbitq), 
to_sfixed(-71616652.0/4294967296.0,1,-nbitq), 
to_sfixed(-297872569.0/4294967296.0,1,-nbitq), 
to_sfixed(-515998382.0/4294967296.0,1,-nbitq), 
to_sfixed(-227889192.0/4294967296.0,1,-nbitq), 
to_sfixed(-154652922.0/4294967296.0,1,-nbitq), 
to_sfixed(-133706187.0/4294967296.0,1,-nbitq), 
to_sfixed(-129760176.0/4294967296.0,1,-nbitq), 
to_sfixed(-191273765.0/4294967296.0,1,-nbitq), 
to_sfixed(364169129.0/4294967296.0,1,-nbitq), 
to_sfixed(-240063537.0/4294967296.0,1,-nbitq), 
to_sfixed(-189479710.0/4294967296.0,1,-nbitq), 
to_sfixed(158790887.0/4294967296.0,1,-nbitq), 
to_sfixed(285019074.0/4294967296.0,1,-nbitq), 
to_sfixed(-304967678.0/4294967296.0,1,-nbitq), 
to_sfixed(-303255578.0/4294967296.0,1,-nbitq), 
to_sfixed(239011984.0/4294967296.0,1,-nbitq), 
to_sfixed(668485871.0/4294967296.0,1,-nbitq), 
to_sfixed(114253517.0/4294967296.0,1,-nbitq), 
to_sfixed(159976452.0/4294967296.0,1,-nbitq), 
to_sfixed(-66676005.0/4294967296.0,1,-nbitq), 
to_sfixed(192528911.0/4294967296.0,1,-nbitq), 
to_sfixed(-138456858.0/4294967296.0,1,-nbitq), 
to_sfixed(-307632713.0/4294967296.0,1,-nbitq), 
to_sfixed(11391341.0/4294967296.0,1,-nbitq), 
to_sfixed(-202342737.0/4294967296.0,1,-nbitq), 
to_sfixed(-450145988.0/4294967296.0,1,-nbitq), 
to_sfixed(-118361870.0/4294967296.0,1,-nbitq), 
to_sfixed(249604540.0/4294967296.0,1,-nbitq), 
to_sfixed(-321388889.0/4294967296.0,1,-nbitq), 
to_sfixed(22261640.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(273910299.0/4294967296.0,1,-nbitq), 
to_sfixed(30682340.0/4294967296.0,1,-nbitq), 
to_sfixed(-245361305.0/4294967296.0,1,-nbitq), 
to_sfixed(-99465752.0/4294967296.0,1,-nbitq), 
to_sfixed(197736512.0/4294967296.0,1,-nbitq), 
to_sfixed(198744166.0/4294967296.0,1,-nbitq), 
to_sfixed(179213474.0/4294967296.0,1,-nbitq), 
to_sfixed(-290236133.0/4294967296.0,1,-nbitq), 
to_sfixed(-272104026.0/4294967296.0,1,-nbitq), 
to_sfixed(-164279853.0/4294967296.0,1,-nbitq), 
to_sfixed(254207588.0/4294967296.0,1,-nbitq), 
to_sfixed(-223918380.0/4294967296.0,1,-nbitq), 
to_sfixed(213643703.0/4294967296.0,1,-nbitq), 
to_sfixed(-50932731.0/4294967296.0,1,-nbitq), 
to_sfixed(-304437439.0/4294967296.0,1,-nbitq), 
to_sfixed(-278705720.0/4294967296.0,1,-nbitq), 
to_sfixed(-382783587.0/4294967296.0,1,-nbitq), 
to_sfixed(240276429.0/4294967296.0,1,-nbitq), 
to_sfixed(-28497532.0/4294967296.0,1,-nbitq), 
to_sfixed(224272764.0/4294967296.0,1,-nbitq), 
to_sfixed(-132701838.0/4294967296.0,1,-nbitq), 
to_sfixed(-220435481.0/4294967296.0,1,-nbitq), 
to_sfixed(-46708849.0/4294967296.0,1,-nbitq), 
to_sfixed(258337000.0/4294967296.0,1,-nbitq), 
to_sfixed(63518062.0/4294967296.0,1,-nbitq), 
to_sfixed(-202771917.0/4294967296.0,1,-nbitq), 
to_sfixed(-99623895.0/4294967296.0,1,-nbitq), 
to_sfixed(-404052025.0/4294967296.0,1,-nbitq), 
to_sfixed(-213323000.0/4294967296.0,1,-nbitq), 
to_sfixed(282799436.0/4294967296.0,1,-nbitq), 
to_sfixed(-85503878.0/4294967296.0,1,-nbitq), 
to_sfixed(-292134247.0/4294967296.0,1,-nbitq), 
to_sfixed(417436367.0/4294967296.0,1,-nbitq), 
to_sfixed(-230196386.0/4294967296.0,1,-nbitq), 
to_sfixed(31983390.0/4294967296.0,1,-nbitq), 
to_sfixed(278011025.0/4294967296.0,1,-nbitq), 
to_sfixed(359048739.0/4294967296.0,1,-nbitq), 
to_sfixed(-234673525.0/4294967296.0,1,-nbitq), 
to_sfixed(-375004753.0/4294967296.0,1,-nbitq), 
to_sfixed(-131310715.0/4294967296.0,1,-nbitq), 
to_sfixed(22144316.0/4294967296.0,1,-nbitq), 
to_sfixed(191018945.0/4294967296.0,1,-nbitq), 
to_sfixed(102973470.0/4294967296.0,1,-nbitq), 
to_sfixed(204288213.0/4294967296.0,1,-nbitq), 
to_sfixed(-234953016.0/4294967296.0,1,-nbitq), 
to_sfixed(458611086.0/4294967296.0,1,-nbitq), 
to_sfixed(-246628111.0/4294967296.0,1,-nbitq), 
to_sfixed(-39947087.0/4294967296.0,1,-nbitq), 
to_sfixed(-156633993.0/4294967296.0,1,-nbitq), 
to_sfixed(-19625237.0/4294967296.0,1,-nbitq), 
to_sfixed(-226845264.0/4294967296.0,1,-nbitq), 
to_sfixed(177587633.0/4294967296.0,1,-nbitq), 
to_sfixed(-386529042.0/4294967296.0,1,-nbitq), 
to_sfixed(458921491.0/4294967296.0,1,-nbitq), 
to_sfixed(269527167.0/4294967296.0,1,-nbitq), 
to_sfixed(-196001209.0/4294967296.0,1,-nbitq), 
to_sfixed(-303312883.0/4294967296.0,1,-nbitq), 
to_sfixed(-449221754.0/4294967296.0,1,-nbitq), 
to_sfixed(346414228.0/4294967296.0,1,-nbitq), 
to_sfixed(367707791.0/4294967296.0,1,-nbitq), 
to_sfixed(-68873282.0/4294967296.0,1,-nbitq), 
to_sfixed(83916298.0/4294967296.0,1,-nbitq), 
to_sfixed(27582385.0/4294967296.0,1,-nbitq), 
to_sfixed(3318817.0/4294967296.0,1,-nbitq), 
to_sfixed(45732511.0/4294967296.0,1,-nbitq), 
to_sfixed(-7810793.0/4294967296.0,1,-nbitq), 
to_sfixed(46099895.0/4294967296.0,1,-nbitq), 
to_sfixed(-87414393.0/4294967296.0,1,-nbitq), 
to_sfixed(161980993.0/4294967296.0,1,-nbitq), 
to_sfixed(-241663888.0/4294967296.0,1,-nbitq), 
to_sfixed(-49340286.0/4294967296.0,1,-nbitq), 
to_sfixed(-184033363.0/4294967296.0,1,-nbitq), 
to_sfixed(134471039.0/4294967296.0,1,-nbitq), 
to_sfixed(-227037363.0/4294967296.0,1,-nbitq), 
to_sfixed(-119484173.0/4294967296.0,1,-nbitq), 
to_sfixed(-573612535.0/4294967296.0,1,-nbitq), 
to_sfixed(305319114.0/4294967296.0,1,-nbitq), 
to_sfixed(-425873494.0/4294967296.0,1,-nbitq), 
to_sfixed(-590057333.0/4294967296.0,1,-nbitq), 
to_sfixed(325770173.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(106273100.0/4294967296.0,1,-nbitq), 
to_sfixed(-182182218.0/4294967296.0,1,-nbitq), 
to_sfixed(21049735.0/4294967296.0,1,-nbitq), 
to_sfixed(-63728060.0/4294967296.0,1,-nbitq), 
to_sfixed(292076871.0/4294967296.0,1,-nbitq), 
to_sfixed(93175023.0/4294967296.0,1,-nbitq), 
to_sfixed(-86547953.0/4294967296.0,1,-nbitq), 
to_sfixed(-23458892.0/4294967296.0,1,-nbitq), 
to_sfixed(-118446216.0/4294967296.0,1,-nbitq), 
to_sfixed(312359620.0/4294967296.0,1,-nbitq), 
to_sfixed(-265182261.0/4294967296.0,1,-nbitq), 
to_sfixed(212115771.0/4294967296.0,1,-nbitq), 
to_sfixed(138166460.0/4294967296.0,1,-nbitq), 
to_sfixed(-322403420.0/4294967296.0,1,-nbitq), 
to_sfixed(161575260.0/4294967296.0,1,-nbitq), 
to_sfixed(138651852.0/4294967296.0,1,-nbitq), 
to_sfixed(-151752776.0/4294967296.0,1,-nbitq), 
to_sfixed(-192870541.0/4294967296.0,1,-nbitq), 
to_sfixed(-112752173.0/4294967296.0,1,-nbitq), 
to_sfixed(-203522660.0/4294967296.0,1,-nbitq), 
to_sfixed(-344824034.0/4294967296.0,1,-nbitq), 
to_sfixed(177641121.0/4294967296.0,1,-nbitq), 
to_sfixed(518756482.0/4294967296.0,1,-nbitq), 
to_sfixed(-144624937.0/4294967296.0,1,-nbitq), 
to_sfixed(57670150.0/4294967296.0,1,-nbitq), 
to_sfixed(-9865157.0/4294967296.0,1,-nbitq), 
to_sfixed(357247873.0/4294967296.0,1,-nbitq), 
to_sfixed(-308443837.0/4294967296.0,1,-nbitq), 
to_sfixed(14057575.0/4294967296.0,1,-nbitq), 
to_sfixed(-210586893.0/4294967296.0,1,-nbitq), 
to_sfixed(-245394561.0/4294967296.0,1,-nbitq), 
to_sfixed(-102291539.0/4294967296.0,1,-nbitq), 
to_sfixed(115475167.0/4294967296.0,1,-nbitq), 
to_sfixed(-77099951.0/4294967296.0,1,-nbitq), 
to_sfixed(459195294.0/4294967296.0,1,-nbitq), 
to_sfixed(225426794.0/4294967296.0,1,-nbitq), 
to_sfixed(93509649.0/4294967296.0,1,-nbitq), 
to_sfixed(144071273.0/4294967296.0,1,-nbitq), 
to_sfixed(-248118940.0/4294967296.0,1,-nbitq), 
to_sfixed(201271232.0/4294967296.0,1,-nbitq), 
to_sfixed(-297333246.0/4294967296.0,1,-nbitq), 
to_sfixed(466747263.0/4294967296.0,1,-nbitq), 
to_sfixed(204351634.0/4294967296.0,1,-nbitq), 
to_sfixed(233291878.0/4294967296.0,1,-nbitq), 
to_sfixed(-144075145.0/4294967296.0,1,-nbitq), 
to_sfixed(86510980.0/4294967296.0,1,-nbitq), 
to_sfixed(-59160912.0/4294967296.0,1,-nbitq), 
to_sfixed(-362557054.0/4294967296.0,1,-nbitq), 
to_sfixed(-293328145.0/4294967296.0,1,-nbitq), 
to_sfixed(-73280571.0/4294967296.0,1,-nbitq), 
to_sfixed(132473146.0/4294967296.0,1,-nbitq), 
to_sfixed(-2655383.0/4294967296.0,1,-nbitq), 
to_sfixed(-308916144.0/4294967296.0,1,-nbitq), 
to_sfixed(246914625.0/4294967296.0,1,-nbitq), 
to_sfixed(-144669001.0/4294967296.0,1,-nbitq), 
to_sfixed(54852801.0/4294967296.0,1,-nbitq), 
to_sfixed(-276415024.0/4294967296.0,1,-nbitq), 
to_sfixed(205592588.0/4294967296.0,1,-nbitq), 
to_sfixed(376524253.0/4294967296.0,1,-nbitq), 
to_sfixed(310253331.0/4294967296.0,1,-nbitq), 
to_sfixed(232939192.0/4294967296.0,1,-nbitq), 
to_sfixed(578010673.0/4294967296.0,1,-nbitq), 
to_sfixed(-344437079.0/4294967296.0,1,-nbitq), 
to_sfixed(402582635.0/4294967296.0,1,-nbitq), 
to_sfixed(-92255954.0/4294967296.0,1,-nbitq), 
to_sfixed(-117423392.0/4294967296.0,1,-nbitq), 
to_sfixed(554771305.0/4294967296.0,1,-nbitq), 
to_sfixed(49808860.0/4294967296.0,1,-nbitq), 
to_sfixed(-167644448.0/4294967296.0,1,-nbitq), 
to_sfixed(-112210318.0/4294967296.0,1,-nbitq), 
to_sfixed(7138352.0/4294967296.0,1,-nbitq), 
to_sfixed(44683512.0/4294967296.0,1,-nbitq), 
to_sfixed(101775783.0/4294967296.0,1,-nbitq), 
to_sfixed(141456603.0/4294967296.0,1,-nbitq), 
to_sfixed(480309053.0/4294967296.0,1,-nbitq), 
to_sfixed(16509428.0/4294967296.0,1,-nbitq), 
to_sfixed(62004123.0/4294967296.0,1,-nbitq), 
to_sfixed(26143753.0/4294967296.0,1,-nbitq), 
to_sfixed(-559332841.0/4294967296.0,1,-nbitq), 
to_sfixed(93633766.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(260285667.0/4294967296.0,1,-nbitq), 
to_sfixed(-217095719.0/4294967296.0,1,-nbitq), 
to_sfixed(-36533023.0/4294967296.0,1,-nbitq), 
to_sfixed(23919992.0/4294967296.0,1,-nbitq), 
to_sfixed(395875086.0/4294967296.0,1,-nbitq), 
to_sfixed(-85178505.0/4294967296.0,1,-nbitq), 
to_sfixed(409254581.0/4294967296.0,1,-nbitq), 
to_sfixed(411471537.0/4294967296.0,1,-nbitq), 
to_sfixed(153142856.0/4294967296.0,1,-nbitq), 
to_sfixed(3131740.0/4294967296.0,1,-nbitq), 
to_sfixed(21416196.0/4294967296.0,1,-nbitq), 
to_sfixed(163058463.0/4294967296.0,1,-nbitq), 
to_sfixed(-315488382.0/4294967296.0,1,-nbitq), 
to_sfixed(-102037263.0/4294967296.0,1,-nbitq), 
to_sfixed(170033018.0/4294967296.0,1,-nbitq), 
to_sfixed(-364324267.0/4294967296.0,1,-nbitq), 
to_sfixed(-111774379.0/4294967296.0,1,-nbitq), 
to_sfixed(16118404.0/4294967296.0,1,-nbitq), 
to_sfixed(-201881033.0/4294967296.0,1,-nbitq), 
to_sfixed(157681003.0/4294967296.0,1,-nbitq), 
to_sfixed(-191884958.0/4294967296.0,1,-nbitq), 
to_sfixed(181378720.0/4294967296.0,1,-nbitq), 
to_sfixed(680536553.0/4294967296.0,1,-nbitq), 
to_sfixed(359376839.0/4294967296.0,1,-nbitq), 
to_sfixed(-11071740.0/4294967296.0,1,-nbitq), 
to_sfixed(-434170452.0/4294967296.0,1,-nbitq), 
to_sfixed(-170641760.0/4294967296.0,1,-nbitq), 
to_sfixed(-623781537.0/4294967296.0,1,-nbitq), 
to_sfixed(-3418662.0/4294967296.0,1,-nbitq), 
to_sfixed(-252161248.0/4294967296.0,1,-nbitq), 
to_sfixed(-613790857.0/4294967296.0,1,-nbitq), 
to_sfixed(-411516040.0/4294967296.0,1,-nbitq), 
to_sfixed(-159113679.0/4294967296.0,1,-nbitq), 
to_sfixed(229151549.0/4294967296.0,1,-nbitq), 
to_sfixed(365513265.0/4294967296.0,1,-nbitq), 
to_sfixed(40515806.0/4294967296.0,1,-nbitq), 
to_sfixed(149785108.0/4294967296.0,1,-nbitq), 
to_sfixed(536180172.0/4294967296.0,1,-nbitq), 
to_sfixed(145203943.0/4294967296.0,1,-nbitq), 
to_sfixed(504873146.0/4294967296.0,1,-nbitq), 
to_sfixed(8452567.0/4294967296.0,1,-nbitq), 
to_sfixed(-56689803.0/4294967296.0,1,-nbitq), 
to_sfixed(-77584346.0/4294967296.0,1,-nbitq), 
to_sfixed(117435732.0/4294967296.0,1,-nbitq), 
to_sfixed(-72700596.0/4294967296.0,1,-nbitq), 
to_sfixed(14934495.0/4294967296.0,1,-nbitq), 
to_sfixed(-109796871.0/4294967296.0,1,-nbitq), 
to_sfixed(-62911825.0/4294967296.0,1,-nbitq), 
to_sfixed(-327537956.0/4294967296.0,1,-nbitq), 
to_sfixed(8610147.0/4294967296.0,1,-nbitq), 
to_sfixed(53348853.0/4294967296.0,1,-nbitq), 
to_sfixed(233119588.0/4294967296.0,1,-nbitq), 
to_sfixed(-36503465.0/4294967296.0,1,-nbitq), 
to_sfixed(209752649.0/4294967296.0,1,-nbitq), 
to_sfixed(363501625.0/4294967296.0,1,-nbitq), 
to_sfixed(98958864.0/4294967296.0,1,-nbitq), 
to_sfixed(330877926.0/4294967296.0,1,-nbitq), 
to_sfixed(-220139618.0/4294967296.0,1,-nbitq), 
to_sfixed(-222104578.0/4294967296.0,1,-nbitq), 
to_sfixed(162707488.0/4294967296.0,1,-nbitq), 
to_sfixed(325679613.0/4294967296.0,1,-nbitq), 
to_sfixed(-35903155.0/4294967296.0,1,-nbitq), 
to_sfixed(7514025.0/4294967296.0,1,-nbitq), 
to_sfixed(69496982.0/4294967296.0,1,-nbitq), 
to_sfixed(-193314467.0/4294967296.0,1,-nbitq), 
to_sfixed(-186645271.0/4294967296.0,1,-nbitq), 
to_sfixed(447004394.0/4294967296.0,1,-nbitq), 
to_sfixed(-68663530.0/4294967296.0,1,-nbitq), 
to_sfixed(-100605213.0/4294967296.0,1,-nbitq), 
to_sfixed(188303664.0/4294967296.0,1,-nbitq), 
to_sfixed(-232671768.0/4294967296.0,1,-nbitq), 
to_sfixed(-42739198.0/4294967296.0,1,-nbitq), 
to_sfixed(-60979508.0/4294967296.0,1,-nbitq), 
to_sfixed(418805914.0/4294967296.0,1,-nbitq), 
to_sfixed(15661829.0/4294967296.0,1,-nbitq), 
to_sfixed(-85324240.0/4294967296.0,1,-nbitq), 
to_sfixed(423949124.0/4294967296.0,1,-nbitq), 
to_sfixed(-21337022.0/4294967296.0,1,-nbitq), 
to_sfixed(-344523040.0/4294967296.0,1,-nbitq), 
to_sfixed(385067472.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-245841750.0/4294967296.0,1,-nbitq), 
to_sfixed(109119515.0/4294967296.0,1,-nbitq), 
to_sfixed(82244183.0/4294967296.0,1,-nbitq), 
to_sfixed(214565929.0/4294967296.0,1,-nbitq), 
to_sfixed(567261014.0/4294967296.0,1,-nbitq), 
to_sfixed(-168358743.0/4294967296.0,1,-nbitq), 
to_sfixed(441765238.0/4294967296.0,1,-nbitq), 
to_sfixed(-248857135.0/4294967296.0,1,-nbitq), 
to_sfixed(466407465.0/4294967296.0,1,-nbitq), 
to_sfixed(326738686.0/4294967296.0,1,-nbitq), 
to_sfixed(-259655939.0/4294967296.0,1,-nbitq), 
to_sfixed(650528804.0/4294967296.0,1,-nbitq), 
to_sfixed(45626353.0/4294967296.0,1,-nbitq), 
to_sfixed(156614527.0/4294967296.0,1,-nbitq), 
to_sfixed(-304041248.0/4294967296.0,1,-nbitq), 
to_sfixed(31686075.0/4294967296.0,1,-nbitq), 
to_sfixed(-414824829.0/4294967296.0,1,-nbitq), 
to_sfixed(-45486554.0/4294967296.0,1,-nbitq), 
to_sfixed(-441328110.0/4294967296.0,1,-nbitq), 
to_sfixed(-318829253.0/4294967296.0,1,-nbitq), 
to_sfixed(-33415813.0/4294967296.0,1,-nbitq), 
to_sfixed(14654023.0/4294967296.0,1,-nbitq), 
to_sfixed(-25751780.0/4294967296.0,1,-nbitq), 
to_sfixed(195525460.0/4294967296.0,1,-nbitq), 
to_sfixed(-233984358.0/4294967296.0,1,-nbitq), 
to_sfixed(135682396.0/4294967296.0,1,-nbitq), 
to_sfixed(-342246733.0/4294967296.0,1,-nbitq), 
to_sfixed(4310426.0/4294967296.0,1,-nbitq), 
to_sfixed(-238979311.0/4294967296.0,1,-nbitq), 
to_sfixed(-93719751.0/4294967296.0,1,-nbitq), 
to_sfixed(-361145905.0/4294967296.0,1,-nbitq), 
to_sfixed(-627420161.0/4294967296.0,1,-nbitq), 
to_sfixed(5462281.0/4294967296.0,1,-nbitq), 
to_sfixed(100455154.0/4294967296.0,1,-nbitq), 
to_sfixed(485187638.0/4294967296.0,1,-nbitq), 
to_sfixed(458091489.0/4294967296.0,1,-nbitq), 
to_sfixed(-194300214.0/4294967296.0,1,-nbitq), 
to_sfixed(263580768.0/4294967296.0,1,-nbitq), 
to_sfixed(-283947110.0/4294967296.0,1,-nbitq), 
to_sfixed(-50681470.0/4294967296.0,1,-nbitq), 
to_sfixed(-197485776.0/4294967296.0,1,-nbitq), 
to_sfixed(-92804308.0/4294967296.0,1,-nbitq), 
to_sfixed(-380573940.0/4294967296.0,1,-nbitq), 
to_sfixed(-358057640.0/4294967296.0,1,-nbitq), 
to_sfixed(306544310.0/4294967296.0,1,-nbitq), 
to_sfixed(-281651483.0/4294967296.0,1,-nbitq), 
to_sfixed(-175236794.0/4294967296.0,1,-nbitq), 
to_sfixed(-6226501.0/4294967296.0,1,-nbitq), 
to_sfixed(-162333905.0/4294967296.0,1,-nbitq), 
to_sfixed(512193002.0/4294967296.0,1,-nbitq), 
to_sfixed(-136783615.0/4294967296.0,1,-nbitq), 
to_sfixed(-123808456.0/4294967296.0,1,-nbitq), 
to_sfixed(-323891691.0/4294967296.0,1,-nbitq), 
to_sfixed(-72073618.0/4294967296.0,1,-nbitq), 
to_sfixed(192752474.0/4294967296.0,1,-nbitq), 
to_sfixed(-47992999.0/4294967296.0,1,-nbitq), 
to_sfixed(333739906.0/4294967296.0,1,-nbitq), 
to_sfixed(-495443289.0/4294967296.0,1,-nbitq), 
to_sfixed(-186940189.0/4294967296.0,1,-nbitq), 
to_sfixed(317909063.0/4294967296.0,1,-nbitq), 
to_sfixed(-220631623.0/4294967296.0,1,-nbitq), 
to_sfixed(126314203.0/4294967296.0,1,-nbitq), 
to_sfixed(-472494983.0/4294967296.0,1,-nbitq), 
to_sfixed(200915719.0/4294967296.0,1,-nbitq), 
to_sfixed(-113578162.0/4294967296.0,1,-nbitq), 
to_sfixed(48266346.0/4294967296.0,1,-nbitq), 
to_sfixed(-17130514.0/4294967296.0,1,-nbitq), 
to_sfixed(-127555874.0/4294967296.0,1,-nbitq), 
to_sfixed(-350640069.0/4294967296.0,1,-nbitq), 
to_sfixed(222693556.0/4294967296.0,1,-nbitq), 
to_sfixed(-89070097.0/4294967296.0,1,-nbitq), 
to_sfixed(-129179659.0/4294967296.0,1,-nbitq), 
to_sfixed(-342663228.0/4294967296.0,1,-nbitq), 
to_sfixed(443545147.0/4294967296.0,1,-nbitq), 
to_sfixed(-216556919.0/4294967296.0,1,-nbitq), 
to_sfixed(-288463728.0/4294967296.0,1,-nbitq), 
to_sfixed(385740256.0/4294967296.0,1,-nbitq), 
to_sfixed(-340256132.0/4294967296.0,1,-nbitq), 
to_sfixed(-285076877.0/4294967296.0,1,-nbitq), 
to_sfixed(-133123145.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(71580881.0/4294967296.0,1,-nbitq), 
to_sfixed(-137230142.0/4294967296.0,1,-nbitq), 
to_sfixed(206715877.0/4294967296.0,1,-nbitq), 
to_sfixed(-284198233.0/4294967296.0,1,-nbitq), 
to_sfixed(225215437.0/4294967296.0,1,-nbitq), 
to_sfixed(98153740.0/4294967296.0,1,-nbitq), 
to_sfixed(384314847.0/4294967296.0,1,-nbitq), 
to_sfixed(226609319.0/4294967296.0,1,-nbitq), 
to_sfixed(469968398.0/4294967296.0,1,-nbitq), 
to_sfixed(242896938.0/4294967296.0,1,-nbitq), 
to_sfixed(-265448945.0/4294967296.0,1,-nbitq), 
to_sfixed(350819794.0/4294967296.0,1,-nbitq), 
to_sfixed(-58310508.0/4294967296.0,1,-nbitq), 
to_sfixed(-324878789.0/4294967296.0,1,-nbitq), 
to_sfixed(244235713.0/4294967296.0,1,-nbitq), 
to_sfixed(-169844716.0/4294967296.0,1,-nbitq), 
to_sfixed(337097450.0/4294967296.0,1,-nbitq), 
to_sfixed(-196666028.0/4294967296.0,1,-nbitq), 
to_sfixed(110410649.0/4294967296.0,1,-nbitq), 
to_sfixed(-197833960.0/4294967296.0,1,-nbitq), 
to_sfixed(-339728474.0/4294967296.0,1,-nbitq), 
to_sfixed(-150980003.0/4294967296.0,1,-nbitq), 
to_sfixed(194235978.0/4294967296.0,1,-nbitq), 
to_sfixed(58424584.0/4294967296.0,1,-nbitq), 
to_sfixed(324393711.0/4294967296.0,1,-nbitq), 
to_sfixed(-532817189.0/4294967296.0,1,-nbitq), 
to_sfixed(-322338334.0/4294967296.0,1,-nbitq), 
to_sfixed(-366865609.0/4294967296.0,1,-nbitq), 
to_sfixed(-151180762.0/4294967296.0,1,-nbitq), 
to_sfixed(-137193723.0/4294967296.0,1,-nbitq), 
to_sfixed(14311588.0/4294967296.0,1,-nbitq), 
to_sfixed(-97087273.0/4294967296.0,1,-nbitq), 
to_sfixed(60643061.0/4294967296.0,1,-nbitq), 
to_sfixed(-347465631.0/4294967296.0,1,-nbitq), 
to_sfixed(81190543.0/4294967296.0,1,-nbitq), 
to_sfixed(-84692812.0/4294967296.0,1,-nbitq), 
to_sfixed(238078952.0/4294967296.0,1,-nbitq), 
to_sfixed(148267722.0/4294967296.0,1,-nbitq), 
to_sfixed(-562191093.0/4294967296.0,1,-nbitq), 
to_sfixed(359846742.0/4294967296.0,1,-nbitq), 
to_sfixed(-285617261.0/4294967296.0,1,-nbitq), 
to_sfixed(431871182.0/4294967296.0,1,-nbitq), 
to_sfixed(357303818.0/4294967296.0,1,-nbitq), 
to_sfixed(-158781546.0/4294967296.0,1,-nbitq), 
to_sfixed(-10617215.0/4294967296.0,1,-nbitq), 
to_sfixed(428956471.0/4294967296.0,1,-nbitq), 
to_sfixed(22798009.0/4294967296.0,1,-nbitq), 
to_sfixed(-197289886.0/4294967296.0,1,-nbitq), 
to_sfixed(-271772123.0/4294967296.0,1,-nbitq), 
to_sfixed(209793409.0/4294967296.0,1,-nbitq), 
to_sfixed(-292368390.0/4294967296.0,1,-nbitq), 
to_sfixed(-142441307.0/4294967296.0,1,-nbitq), 
to_sfixed(96670290.0/4294967296.0,1,-nbitq), 
to_sfixed(-103177700.0/4294967296.0,1,-nbitq), 
to_sfixed(312720231.0/4294967296.0,1,-nbitq), 
to_sfixed(-56860919.0/4294967296.0,1,-nbitq), 
to_sfixed(508141211.0/4294967296.0,1,-nbitq), 
to_sfixed(-177428897.0/4294967296.0,1,-nbitq), 
to_sfixed(22403900.0/4294967296.0,1,-nbitq), 
to_sfixed(251515405.0/4294967296.0,1,-nbitq), 
to_sfixed(377434292.0/4294967296.0,1,-nbitq), 
to_sfixed(-115795534.0/4294967296.0,1,-nbitq), 
to_sfixed(19769192.0/4294967296.0,1,-nbitq), 
to_sfixed(351234191.0/4294967296.0,1,-nbitq), 
to_sfixed(387709164.0/4294967296.0,1,-nbitq), 
to_sfixed(-167187398.0/4294967296.0,1,-nbitq), 
to_sfixed(582183916.0/4294967296.0,1,-nbitq), 
to_sfixed(-26238565.0/4294967296.0,1,-nbitq), 
to_sfixed(369717743.0/4294967296.0,1,-nbitq), 
to_sfixed(424216568.0/4294967296.0,1,-nbitq), 
to_sfixed(-241353143.0/4294967296.0,1,-nbitq), 
to_sfixed(260963862.0/4294967296.0,1,-nbitq), 
to_sfixed(356622209.0/4294967296.0,1,-nbitq), 
to_sfixed(334615657.0/4294967296.0,1,-nbitq), 
to_sfixed(123880905.0/4294967296.0,1,-nbitq), 
to_sfixed(344866721.0/4294967296.0,1,-nbitq), 
to_sfixed(-81463360.0/4294967296.0,1,-nbitq), 
to_sfixed(-73866778.0/4294967296.0,1,-nbitq), 
to_sfixed(-400768870.0/4294967296.0,1,-nbitq), 
to_sfixed(293534050.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(243741212.0/4294967296.0,1,-nbitq), 
to_sfixed(-12990857.0/4294967296.0,1,-nbitq), 
to_sfixed(607977968.0/4294967296.0,1,-nbitq), 
to_sfixed(-390532201.0/4294967296.0,1,-nbitq), 
to_sfixed(201710584.0/4294967296.0,1,-nbitq), 
to_sfixed(-277537884.0/4294967296.0,1,-nbitq), 
to_sfixed(-222030796.0/4294967296.0,1,-nbitq), 
to_sfixed(317764089.0/4294967296.0,1,-nbitq), 
to_sfixed(1087219910.0/4294967296.0,1,-nbitq), 
to_sfixed(464769934.0/4294967296.0,1,-nbitq), 
to_sfixed(144276980.0/4294967296.0,1,-nbitq), 
to_sfixed(870359392.0/4294967296.0,1,-nbitq), 
to_sfixed(-849892104.0/4294967296.0,1,-nbitq), 
to_sfixed(-155134597.0/4294967296.0,1,-nbitq), 
to_sfixed(-227679058.0/4294967296.0,1,-nbitq), 
to_sfixed(268312627.0/4294967296.0,1,-nbitq), 
to_sfixed(3547398.0/4294967296.0,1,-nbitq), 
to_sfixed(308677635.0/4294967296.0,1,-nbitq), 
to_sfixed(-26110775.0/4294967296.0,1,-nbitq), 
to_sfixed(297668453.0/4294967296.0,1,-nbitq), 
to_sfixed(29514530.0/4294967296.0,1,-nbitq), 
to_sfixed(242621036.0/4294967296.0,1,-nbitq), 
to_sfixed(550117099.0/4294967296.0,1,-nbitq), 
to_sfixed(165346780.0/4294967296.0,1,-nbitq), 
to_sfixed(350068842.0/4294967296.0,1,-nbitq), 
to_sfixed(155544855.0/4294967296.0,1,-nbitq), 
to_sfixed(-22712045.0/4294967296.0,1,-nbitq), 
to_sfixed(1075786.0/4294967296.0,1,-nbitq), 
to_sfixed(-320934266.0/4294967296.0,1,-nbitq), 
to_sfixed(152528044.0/4294967296.0,1,-nbitq), 
to_sfixed(-701428982.0/4294967296.0,1,-nbitq), 
to_sfixed(-834471.0/4294967296.0,1,-nbitq), 
to_sfixed(-80216285.0/4294967296.0,1,-nbitq), 
to_sfixed(-82176278.0/4294967296.0,1,-nbitq), 
to_sfixed(-237423773.0/4294967296.0,1,-nbitq), 
to_sfixed(-144931054.0/4294967296.0,1,-nbitq), 
to_sfixed(454121434.0/4294967296.0,1,-nbitq), 
to_sfixed(-219153070.0/4294967296.0,1,-nbitq), 
to_sfixed(-393910430.0/4294967296.0,1,-nbitq), 
to_sfixed(189594120.0/4294967296.0,1,-nbitq), 
to_sfixed(404746836.0/4294967296.0,1,-nbitq), 
to_sfixed(-268352454.0/4294967296.0,1,-nbitq), 
to_sfixed(301156019.0/4294967296.0,1,-nbitq), 
to_sfixed(34796058.0/4294967296.0,1,-nbitq), 
to_sfixed(112012551.0/4294967296.0,1,-nbitq), 
to_sfixed(690071212.0/4294967296.0,1,-nbitq), 
to_sfixed(-301841265.0/4294967296.0,1,-nbitq), 
to_sfixed(343560181.0/4294967296.0,1,-nbitq), 
to_sfixed(89791603.0/4294967296.0,1,-nbitq), 
to_sfixed(286793263.0/4294967296.0,1,-nbitq), 
to_sfixed(-369729739.0/4294967296.0,1,-nbitq), 
to_sfixed(361566037.0/4294967296.0,1,-nbitq), 
to_sfixed(-697458697.0/4294967296.0,1,-nbitq), 
to_sfixed(-224936707.0/4294967296.0,1,-nbitq), 
to_sfixed(687202.0/4294967296.0,1,-nbitq), 
to_sfixed(127882117.0/4294967296.0,1,-nbitq), 
to_sfixed(-143902109.0/4294967296.0,1,-nbitq), 
to_sfixed(-50798748.0/4294967296.0,1,-nbitq), 
to_sfixed(347937297.0/4294967296.0,1,-nbitq), 
to_sfixed(149394534.0/4294967296.0,1,-nbitq), 
to_sfixed(347082549.0/4294967296.0,1,-nbitq), 
to_sfixed(271165518.0/4294967296.0,1,-nbitq), 
to_sfixed(-732845515.0/4294967296.0,1,-nbitq), 
to_sfixed(-193626187.0/4294967296.0,1,-nbitq), 
to_sfixed(181740683.0/4294967296.0,1,-nbitq), 
to_sfixed(-185781236.0/4294967296.0,1,-nbitq), 
to_sfixed(227125467.0/4294967296.0,1,-nbitq), 
to_sfixed(149294745.0/4294967296.0,1,-nbitq), 
to_sfixed(426934908.0/4294967296.0,1,-nbitq), 
to_sfixed(-115470957.0/4294967296.0,1,-nbitq), 
to_sfixed(42456025.0/4294967296.0,1,-nbitq), 
to_sfixed(-165022718.0/4294967296.0,1,-nbitq), 
to_sfixed(233055553.0/4294967296.0,1,-nbitq), 
to_sfixed(205354261.0/4294967296.0,1,-nbitq), 
to_sfixed(-18371722.0/4294967296.0,1,-nbitq), 
to_sfixed(117055872.0/4294967296.0,1,-nbitq), 
to_sfixed(128414423.0/4294967296.0,1,-nbitq), 
to_sfixed(-373834679.0/4294967296.0,1,-nbitq), 
to_sfixed(-568715705.0/4294967296.0,1,-nbitq), 
to_sfixed(106904370.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(82825510.0/4294967296.0,1,-nbitq), 
to_sfixed(-661717561.0/4294967296.0,1,-nbitq), 
to_sfixed(731640739.0/4294967296.0,1,-nbitq), 
to_sfixed(115097163.0/4294967296.0,1,-nbitq), 
to_sfixed(354659672.0/4294967296.0,1,-nbitq), 
to_sfixed(398794638.0/4294967296.0,1,-nbitq), 
to_sfixed(386563438.0/4294967296.0,1,-nbitq), 
to_sfixed(-128633757.0/4294967296.0,1,-nbitq), 
to_sfixed(505639583.0/4294967296.0,1,-nbitq), 
to_sfixed(18092092.0/4294967296.0,1,-nbitq), 
to_sfixed(278373426.0/4294967296.0,1,-nbitq), 
to_sfixed(631460751.0/4294967296.0,1,-nbitq), 
to_sfixed(-740029178.0/4294967296.0,1,-nbitq), 
to_sfixed(-559497675.0/4294967296.0,1,-nbitq), 
to_sfixed(346709891.0/4294967296.0,1,-nbitq), 
to_sfixed(285237979.0/4294967296.0,1,-nbitq), 
to_sfixed(353423657.0/4294967296.0,1,-nbitq), 
to_sfixed(-301393825.0/4294967296.0,1,-nbitq), 
to_sfixed(-252815243.0/4294967296.0,1,-nbitq), 
to_sfixed(-102554020.0/4294967296.0,1,-nbitq), 
to_sfixed(96789525.0/4294967296.0,1,-nbitq), 
to_sfixed(-133921349.0/4294967296.0,1,-nbitq), 
to_sfixed(660919651.0/4294967296.0,1,-nbitq), 
to_sfixed(-48373943.0/4294967296.0,1,-nbitq), 
to_sfixed(410997506.0/4294967296.0,1,-nbitq), 
to_sfixed(-184589159.0/4294967296.0,1,-nbitq), 
to_sfixed(-514704699.0/4294967296.0,1,-nbitq), 
to_sfixed(107685535.0/4294967296.0,1,-nbitq), 
to_sfixed(265584928.0/4294967296.0,1,-nbitq), 
to_sfixed(-129605352.0/4294967296.0,1,-nbitq), 
to_sfixed(-203401238.0/4294967296.0,1,-nbitq), 
to_sfixed(-261568007.0/4294967296.0,1,-nbitq), 
to_sfixed(-234588255.0/4294967296.0,1,-nbitq), 
to_sfixed(57714516.0/4294967296.0,1,-nbitq), 
to_sfixed(81917319.0/4294967296.0,1,-nbitq), 
to_sfixed(-64699328.0/4294967296.0,1,-nbitq), 
to_sfixed(103156975.0/4294967296.0,1,-nbitq), 
to_sfixed(-513499371.0/4294967296.0,1,-nbitq), 
to_sfixed(-351705927.0/4294967296.0,1,-nbitq), 
to_sfixed(-126675802.0/4294967296.0,1,-nbitq), 
to_sfixed(406425000.0/4294967296.0,1,-nbitq), 
to_sfixed(-89693033.0/4294967296.0,1,-nbitq), 
to_sfixed(357878098.0/4294967296.0,1,-nbitq), 
to_sfixed(125351274.0/4294967296.0,1,-nbitq), 
to_sfixed(268522443.0/4294967296.0,1,-nbitq), 
to_sfixed(706044440.0/4294967296.0,1,-nbitq), 
to_sfixed(-278335395.0/4294967296.0,1,-nbitq), 
to_sfixed(196252198.0/4294967296.0,1,-nbitq), 
to_sfixed(-403934962.0/4294967296.0,1,-nbitq), 
to_sfixed(334835932.0/4294967296.0,1,-nbitq), 
to_sfixed(-305120427.0/4294967296.0,1,-nbitq), 
to_sfixed(512596512.0/4294967296.0,1,-nbitq), 
to_sfixed(-337814553.0/4294967296.0,1,-nbitq), 
to_sfixed(-310992696.0/4294967296.0,1,-nbitq), 
to_sfixed(165014303.0/4294967296.0,1,-nbitq), 
to_sfixed(554388407.0/4294967296.0,1,-nbitq), 
to_sfixed(384862232.0/4294967296.0,1,-nbitq), 
to_sfixed(-369227373.0/4294967296.0,1,-nbitq), 
to_sfixed(-23453719.0/4294967296.0,1,-nbitq), 
to_sfixed(416439931.0/4294967296.0,1,-nbitq), 
to_sfixed(-36224656.0/4294967296.0,1,-nbitq), 
to_sfixed(-327122388.0/4294967296.0,1,-nbitq), 
to_sfixed(-436918035.0/4294967296.0,1,-nbitq), 
to_sfixed(173000635.0/4294967296.0,1,-nbitq), 
to_sfixed(-30607723.0/4294967296.0,1,-nbitq), 
to_sfixed(109319724.0/4294967296.0,1,-nbitq), 
to_sfixed(163288559.0/4294967296.0,1,-nbitq), 
to_sfixed(-125726763.0/4294967296.0,1,-nbitq), 
to_sfixed(178390160.0/4294967296.0,1,-nbitq), 
to_sfixed(-21712793.0/4294967296.0,1,-nbitq), 
to_sfixed(-363133246.0/4294967296.0,1,-nbitq), 
to_sfixed(-112761807.0/4294967296.0,1,-nbitq), 
to_sfixed(333047251.0/4294967296.0,1,-nbitq), 
to_sfixed(-284297819.0/4294967296.0,1,-nbitq), 
to_sfixed(351009382.0/4294967296.0,1,-nbitq), 
to_sfixed(63182810.0/4294967296.0,1,-nbitq), 
to_sfixed(742917029.0/4294967296.0,1,-nbitq), 
to_sfixed(234615212.0/4294967296.0,1,-nbitq), 
to_sfixed(198558668.0/4294967296.0,1,-nbitq), 
to_sfixed(-111602541.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(307421566.0/4294967296.0,1,-nbitq), 
to_sfixed(-359984967.0/4294967296.0,1,-nbitq), 
to_sfixed(-29530703.0/4294967296.0,1,-nbitq), 
to_sfixed(-56804265.0/4294967296.0,1,-nbitq), 
to_sfixed(351924183.0/4294967296.0,1,-nbitq), 
to_sfixed(4790390.0/4294967296.0,1,-nbitq), 
to_sfixed(109995488.0/4294967296.0,1,-nbitq), 
to_sfixed(-197853165.0/4294967296.0,1,-nbitq), 
to_sfixed(348115750.0/4294967296.0,1,-nbitq), 
to_sfixed(65565820.0/4294967296.0,1,-nbitq), 
to_sfixed(439474881.0/4294967296.0,1,-nbitq), 
to_sfixed(586497086.0/4294967296.0,1,-nbitq), 
to_sfixed(-559193423.0/4294967296.0,1,-nbitq), 
to_sfixed(-644900778.0/4294967296.0,1,-nbitq), 
to_sfixed(-154954551.0/4294967296.0,1,-nbitq), 
to_sfixed(-157271894.0/4294967296.0,1,-nbitq), 
to_sfixed(31750860.0/4294967296.0,1,-nbitq), 
to_sfixed(-152920639.0/4294967296.0,1,-nbitq), 
to_sfixed(-198014439.0/4294967296.0,1,-nbitq), 
to_sfixed(-2768633.0/4294967296.0,1,-nbitq), 
to_sfixed(256660543.0/4294967296.0,1,-nbitq), 
to_sfixed(-368662364.0/4294967296.0,1,-nbitq), 
to_sfixed(304184199.0/4294967296.0,1,-nbitq), 
to_sfixed(-241738815.0/4294967296.0,1,-nbitq), 
to_sfixed(272801763.0/4294967296.0,1,-nbitq), 
to_sfixed(-217305201.0/4294967296.0,1,-nbitq), 
to_sfixed(-542448236.0/4294967296.0,1,-nbitq), 
to_sfixed(-129249640.0/4294967296.0,1,-nbitq), 
to_sfixed(-146422149.0/4294967296.0,1,-nbitq), 
to_sfixed(302675396.0/4294967296.0,1,-nbitq), 
to_sfixed(287938712.0/4294967296.0,1,-nbitq), 
to_sfixed(-321875366.0/4294967296.0,1,-nbitq), 
to_sfixed(237960638.0/4294967296.0,1,-nbitq), 
to_sfixed(393018396.0/4294967296.0,1,-nbitq), 
to_sfixed(-144765836.0/4294967296.0,1,-nbitq), 
to_sfixed(-398004222.0/4294967296.0,1,-nbitq), 
to_sfixed(467648421.0/4294967296.0,1,-nbitq), 
to_sfixed(52416823.0/4294967296.0,1,-nbitq), 
to_sfixed(-365305011.0/4294967296.0,1,-nbitq), 
to_sfixed(-157336397.0/4294967296.0,1,-nbitq), 
to_sfixed(335333771.0/4294967296.0,1,-nbitq), 
to_sfixed(-202361244.0/4294967296.0,1,-nbitq), 
to_sfixed(182883976.0/4294967296.0,1,-nbitq), 
to_sfixed(180366832.0/4294967296.0,1,-nbitq), 
to_sfixed(-116209924.0/4294967296.0,1,-nbitq), 
to_sfixed(467736120.0/4294967296.0,1,-nbitq), 
to_sfixed(209322499.0/4294967296.0,1,-nbitq), 
to_sfixed(470876441.0/4294967296.0,1,-nbitq), 
to_sfixed(-197454353.0/4294967296.0,1,-nbitq), 
to_sfixed(-217462862.0/4294967296.0,1,-nbitq), 
to_sfixed(-368914962.0/4294967296.0,1,-nbitq), 
to_sfixed(478438167.0/4294967296.0,1,-nbitq), 
to_sfixed(-141079610.0/4294967296.0,1,-nbitq), 
to_sfixed(-178448168.0/4294967296.0,1,-nbitq), 
to_sfixed(-403718668.0/4294967296.0,1,-nbitq), 
to_sfixed(211475084.0/4294967296.0,1,-nbitq), 
to_sfixed(158710354.0/4294967296.0,1,-nbitq), 
to_sfixed(-216536117.0/4294967296.0,1,-nbitq), 
to_sfixed(-172458640.0/4294967296.0,1,-nbitq), 
to_sfixed(-66780721.0/4294967296.0,1,-nbitq), 
to_sfixed(-366944658.0/4294967296.0,1,-nbitq), 
to_sfixed(-16316966.0/4294967296.0,1,-nbitq), 
to_sfixed(-96297443.0/4294967296.0,1,-nbitq), 
to_sfixed(-256660171.0/4294967296.0,1,-nbitq), 
to_sfixed(-432512290.0/4294967296.0,1,-nbitq), 
to_sfixed(181092359.0/4294967296.0,1,-nbitq), 
to_sfixed(289560049.0/4294967296.0,1,-nbitq), 
to_sfixed(-182879293.0/4294967296.0,1,-nbitq), 
to_sfixed(287114084.0/4294967296.0,1,-nbitq), 
to_sfixed(-18161199.0/4294967296.0,1,-nbitq), 
to_sfixed(141410087.0/4294967296.0,1,-nbitq), 
to_sfixed(-261896267.0/4294967296.0,1,-nbitq), 
to_sfixed(402176496.0/4294967296.0,1,-nbitq), 
to_sfixed(18311963.0/4294967296.0,1,-nbitq), 
to_sfixed(351545261.0/4294967296.0,1,-nbitq), 
to_sfixed(105848969.0/4294967296.0,1,-nbitq), 
to_sfixed(-220237154.0/4294967296.0,1,-nbitq), 
to_sfixed(-205817212.0/4294967296.0,1,-nbitq), 
to_sfixed(12170770.0/4294967296.0,1,-nbitq), 
to_sfixed(-268625976.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-7718171.0/4294967296.0,1,-nbitq), 
to_sfixed(-351217890.0/4294967296.0,1,-nbitq), 
to_sfixed(60277192.0/4294967296.0,1,-nbitq), 
to_sfixed(-171517126.0/4294967296.0,1,-nbitq), 
to_sfixed(-492619432.0/4294967296.0,1,-nbitq), 
to_sfixed(339144808.0/4294967296.0,1,-nbitq), 
to_sfixed(138871210.0/4294967296.0,1,-nbitq), 
to_sfixed(28212162.0/4294967296.0,1,-nbitq), 
to_sfixed(845175387.0/4294967296.0,1,-nbitq), 
to_sfixed(318073930.0/4294967296.0,1,-nbitq), 
to_sfixed(109171986.0/4294967296.0,1,-nbitq), 
to_sfixed(820012189.0/4294967296.0,1,-nbitq), 
to_sfixed(-339201452.0/4294967296.0,1,-nbitq), 
to_sfixed(-500166904.0/4294967296.0,1,-nbitq), 
to_sfixed(191911990.0/4294967296.0,1,-nbitq), 
to_sfixed(-395711784.0/4294967296.0,1,-nbitq), 
to_sfixed(-255206381.0/4294967296.0,1,-nbitq), 
to_sfixed(352859011.0/4294967296.0,1,-nbitq), 
to_sfixed(26391866.0/4294967296.0,1,-nbitq), 
to_sfixed(-37015012.0/4294967296.0,1,-nbitq), 
to_sfixed(-284584735.0/4294967296.0,1,-nbitq), 
to_sfixed(230928802.0/4294967296.0,1,-nbitq), 
to_sfixed(500333179.0/4294967296.0,1,-nbitq), 
to_sfixed(-517725898.0/4294967296.0,1,-nbitq), 
to_sfixed(-58884319.0/4294967296.0,1,-nbitq), 
to_sfixed(527381282.0/4294967296.0,1,-nbitq), 
to_sfixed(-284364390.0/4294967296.0,1,-nbitq), 
to_sfixed(-136626509.0/4294967296.0,1,-nbitq), 
to_sfixed(-116636151.0/4294967296.0,1,-nbitq), 
to_sfixed(111233863.0/4294967296.0,1,-nbitq), 
to_sfixed(31666549.0/4294967296.0,1,-nbitq), 
to_sfixed(-617347908.0/4294967296.0,1,-nbitq), 
to_sfixed(-381526344.0/4294967296.0,1,-nbitq), 
to_sfixed(863106479.0/4294967296.0,1,-nbitq), 
to_sfixed(-394851759.0/4294967296.0,1,-nbitq), 
to_sfixed(-487766293.0/4294967296.0,1,-nbitq), 
to_sfixed(424442441.0/4294967296.0,1,-nbitq), 
to_sfixed(11602039.0/4294967296.0,1,-nbitq), 
to_sfixed(-58588654.0/4294967296.0,1,-nbitq), 
to_sfixed(73442987.0/4294967296.0,1,-nbitq), 
to_sfixed(5837169.0/4294967296.0,1,-nbitq), 
to_sfixed(-429772289.0/4294967296.0,1,-nbitq), 
to_sfixed(224962060.0/4294967296.0,1,-nbitq), 
to_sfixed(449828925.0/4294967296.0,1,-nbitq), 
to_sfixed(-88157609.0/4294967296.0,1,-nbitq), 
to_sfixed(-197375424.0/4294967296.0,1,-nbitq), 
to_sfixed(-359052773.0/4294967296.0,1,-nbitq), 
to_sfixed(45550151.0/4294967296.0,1,-nbitq), 
to_sfixed(10681851.0/4294967296.0,1,-nbitq), 
to_sfixed(-17315304.0/4294967296.0,1,-nbitq), 
to_sfixed(273519349.0/4294967296.0,1,-nbitq), 
to_sfixed(-24861763.0/4294967296.0,1,-nbitq), 
to_sfixed(-71676114.0/4294967296.0,1,-nbitq), 
to_sfixed(-527657961.0/4294967296.0,1,-nbitq), 
to_sfixed(-517761473.0/4294967296.0,1,-nbitq), 
to_sfixed(779945711.0/4294967296.0,1,-nbitq), 
to_sfixed(255838934.0/4294967296.0,1,-nbitq), 
to_sfixed(371194580.0/4294967296.0,1,-nbitq), 
to_sfixed(166124863.0/4294967296.0,1,-nbitq), 
to_sfixed(30604086.0/4294967296.0,1,-nbitq), 
to_sfixed(61941718.0/4294967296.0,1,-nbitq), 
to_sfixed(-90115638.0/4294967296.0,1,-nbitq), 
to_sfixed(31430346.0/4294967296.0,1,-nbitq), 
to_sfixed(545974380.0/4294967296.0,1,-nbitq), 
to_sfixed(122549422.0/4294967296.0,1,-nbitq), 
to_sfixed(-187549084.0/4294967296.0,1,-nbitq), 
to_sfixed(-165867949.0/4294967296.0,1,-nbitq), 
to_sfixed(-580693952.0/4294967296.0,1,-nbitq), 
to_sfixed(-230996714.0/4294967296.0,1,-nbitq), 
to_sfixed(-161927589.0/4294967296.0,1,-nbitq), 
to_sfixed(-164154264.0/4294967296.0,1,-nbitq), 
to_sfixed(-523435083.0/4294967296.0,1,-nbitq), 
to_sfixed(542921749.0/4294967296.0,1,-nbitq), 
to_sfixed(294530079.0/4294967296.0,1,-nbitq), 
to_sfixed(435850964.0/4294967296.0,1,-nbitq), 
to_sfixed(21741302.0/4294967296.0,1,-nbitq), 
to_sfixed(414259206.0/4294967296.0,1,-nbitq), 
to_sfixed(-584854401.0/4294967296.0,1,-nbitq), 
to_sfixed(116484436.0/4294967296.0,1,-nbitq), 
to_sfixed(338497071.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(428656686.0/4294967296.0,1,-nbitq), 
to_sfixed(392588955.0/4294967296.0,1,-nbitq), 
to_sfixed(61736507.0/4294967296.0,1,-nbitq), 
to_sfixed(207806440.0/4294967296.0,1,-nbitq), 
to_sfixed(-408874034.0/4294967296.0,1,-nbitq), 
to_sfixed(158249981.0/4294967296.0,1,-nbitq), 
to_sfixed(-38649035.0/4294967296.0,1,-nbitq), 
to_sfixed(288531650.0/4294967296.0,1,-nbitq), 
to_sfixed(335799664.0/4294967296.0,1,-nbitq), 
to_sfixed(171604812.0/4294967296.0,1,-nbitq), 
to_sfixed(106559718.0/4294967296.0,1,-nbitq), 
to_sfixed(208153870.0/4294967296.0,1,-nbitq), 
to_sfixed(-141612981.0/4294967296.0,1,-nbitq), 
to_sfixed(-530985754.0/4294967296.0,1,-nbitq), 
to_sfixed(-46997496.0/4294967296.0,1,-nbitq), 
to_sfixed(-174810939.0/4294967296.0,1,-nbitq), 
to_sfixed(-39740491.0/4294967296.0,1,-nbitq), 
to_sfixed(-106947416.0/4294967296.0,1,-nbitq), 
to_sfixed(-89918933.0/4294967296.0,1,-nbitq), 
to_sfixed(-118413323.0/4294967296.0,1,-nbitq), 
to_sfixed(17955874.0/4294967296.0,1,-nbitq), 
to_sfixed(-265247392.0/4294967296.0,1,-nbitq), 
to_sfixed(270946376.0/4294967296.0,1,-nbitq), 
to_sfixed(88539443.0/4294967296.0,1,-nbitq), 
to_sfixed(-37668358.0/4294967296.0,1,-nbitq), 
to_sfixed(458347662.0/4294967296.0,1,-nbitq), 
to_sfixed(-236829590.0/4294967296.0,1,-nbitq), 
to_sfixed(-18418434.0/4294967296.0,1,-nbitq), 
to_sfixed(236214761.0/4294967296.0,1,-nbitq), 
to_sfixed(-474667761.0/4294967296.0,1,-nbitq), 
to_sfixed(474688076.0/4294967296.0,1,-nbitq), 
to_sfixed(-523580968.0/4294967296.0,1,-nbitq), 
to_sfixed(-161215725.0/4294967296.0,1,-nbitq), 
to_sfixed(-101107569.0/4294967296.0,1,-nbitq), 
to_sfixed(-82330471.0/4294967296.0,1,-nbitq), 
to_sfixed(-413580334.0/4294967296.0,1,-nbitq), 
to_sfixed(526877599.0/4294967296.0,1,-nbitq), 
to_sfixed(344371059.0/4294967296.0,1,-nbitq), 
to_sfixed(-390995875.0/4294967296.0,1,-nbitq), 
to_sfixed(462153046.0/4294967296.0,1,-nbitq), 
to_sfixed(127202886.0/4294967296.0,1,-nbitq), 
to_sfixed(84675551.0/4294967296.0,1,-nbitq), 
to_sfixed(88458605.0/4294967296.0,1,-nbitq), 
to_sfixed(732624196.0/4294967296.0,1,-nbitq), 
to_sfixed(62257196.0/4294967296.0,1,-nbitq), 
to_sfixed(-101666253.0/4294967296.0,1,-nbitq), 
to_sfixed(111363472.0/4294967296.0,1,-nbitq), 
to_sfixed(521032623.0/4294967296.0,1,-nbitq), 
to_sfixed(-243656611.0/4294967296.0,1,-nbitq), 
to_sfixed(513278121.0/4294967296.0,1,-nbitq), 
to_sfixed(202702465.0/4294967296.0,1,-nbitq), 
to_sfixed(243123408.0/4294967296.0,1,-nbitq), 
to_sfixed(-373682302.0/4294967296.0,1,-nbitq), 
to_sfixed(110358304.0/4294967296.0,1,-nbitq), 
to_sfixed(-558573811.0/4294967296.0,1,-nbitq), 
to_sfixed(283728600.0/4294967296.0,1,-nbitq), 
to_sfixed(-299322396.0/4294967296.0,1,-nbitq), 
to_sfixed(13513510.0/4294967296.0,1,-nbitq), 
to_sfixed(-161003736.0/4294967296.0,1,-nbitq), 
to_sfixed(-273668258.0/4294967296.0,1,-nbitq), 
to_sfixed(-262732490.0/4294967296.0,1,-nbitq), 
to_sfixed(-420261480.0/4294967296.0,1,-nbitq), 
to_sfixed(-548009792.0/4294967296.0,1,-nbitq), 
to_sfixed(90348499.0/4294967296.0,1,-nbitq), 
to_sfixed(-201511202.0/4294967296.0,1,-nbitq), 
to_sfixed(-95891183.0/4294967296.0,1,-nbitq), 
to_sfixed(295046559.0/4294967296.0,1,-nbitq), 
to_sfixed(225154089.0/4294967296.0,1,-nbitq), 
to_sfixed(286059832.0/4294967296.0,1,-nbitq), 
to_sfixed(284003085.0/4294967296.0,1,-nbitq), 
to_sfixed(681578055.0/4294967296.0,1,-nbitq), 
to_sfixed(-459997090.0/4294967296.0,1,-nbitq), 
to_sfixed(494098821.0/4294967296.0,1,-nbitq), 
to_sfixed(-49925062.0/4294967296.0,1,-nbitq), 
to_sfixed(383920926.0/4294967296.0,1,-nbitq), 
to_sfixed(-42678993.0/4294967296.0,1,-nbitq), 
to_sfixed(157578449.0/4294967296.0,1,-nbitq), 
to_sfixed(-213610851.0/4294967296.0,1,-nbitq), 
to_sfixed(-160077450.0/4294967296.0,1,-nbitq), 
to_sfixed(-341360243.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(441720079.0/4294967296.0,1,-nbitq), 
to_sfixed(482399921.0/4294967296.0,1,-nbitq), 
to_sfixed(-166199576.0/4294967296.0,1,-nbitq), 
to_sfixed(-209860967.0/4294967296.0,1,-nbitq), 
to_sfixed(-363649012.0/4294967296.0,1,-nbitq), 
to_sfixed(272176283.0/4294967296.0,1,-nbitq), 
to_sfixed(-99391338.0/4294967296.0,1,-nbitq), 
to_sfixed(183014431.0/4294967296.0,1,-nbitq), 
to_sfixed(685586102.0/4294967296.0,1,-nbitq), 
to_sfixed(-77017422.0/4294967296.0,1,-nbitq), 
to_sfixed(21038121.0/4294967296.0,1,-nbitq), 
to_sfixed(493006181.0/4294967296.0,1,-nbitq), 
to_sfixed(25740334.0/4294967296.0,1,-nbitq), 
to_sfixed(-502293033.0/4294967296.0,1,-nbitq), 
to_sfixed(-87959454.0/4294967296.0,1,-nbitq), 
to_sfixed(-212149072.0/4294967296.0,1,-nbitq), 
to_sfixed(-76014314.0/4294967296.0,1,-nbitq), 
to_sfixed(-184606112.0/4294967296.0,1,-nbitq), 
to_sfixed(-171878311.0/4294967296.0,1,-nbitq), 
to_sfixed(-45897845.0/4294967296.0,1,-nbitq), 
to_sfixed(227798796.0/4294967296.0,1,-nbitq), 
to_sfixed(-324165074.0/4294967296.0,1,-nbitq), 
to_sfixed(-189202764.0/4294967296.0,1,-nbitq), 
to_sfixed(-17648687.0/4294967296.0,1,-nbitq), 
to_sfixed(-244223340.0/4294967296.0,1,-nbitq), 
to_sfixed(1259605707.0/4294967296.0,1,-nbitq), 
to_sfixed(-522562789.0/4294967296.0,1,-nbitq), 
to_sfixed(-38123074.0/4294967296.0,1,-nbitq), 
to_sfixed(325424924.0/4294967296.0,1,-nbitq), 
to_sfixed(120208729.0/4294967296.0,1,-nbitq), 
to_sfixed(551029097.0/4294967296.0,1,-nbitq), 
to_sfixed(-35444089.0/4294967296.0,1,-nbitq), 
to_sfixed(-99257717.0/4294967296.0,1,-nbitq), 
to_sfixed(415590891.0/4294967296.0,1,-nbitq), 
to_sfixed(-457148815.0/4294967296.0,1,-nbitq), 
to_sfixed(250033921.0/4294967296.0,1,-nbitq), 
to_sfixed(446588021.0/4294967296.0,1,-nbitq), 
to_sfixed(457683300.0/4294967296.0,1,-nbitq), 
to_sfixed(172538139.0/4294967296.0,1,-nbitq), 
to_sfixed(34599644.0/4294967296.0,1,-nbitq), 
to_sfixed(683925999.0/4294967296.0,1,-nbitq), 
to_sfixed(490368680.0/4294967296.0,1,-nbitq), 
to_sfixed(606183574.0/4294967296.0,1,-nbitq), 
to_sfixed(814037126.0/4294967296.0,1,-nbitq), 
to_sfixed(-321645519.0/4294967296.0,1,-nbitq), 
to_sfixed(341924577.0/4294967296.0,1,-nbitq), 
to_sfixed(120566243.0/4294967296.0,1,-nbitq), 
to_sfixed(-79115171.0/4294967296.0,1,-nbitq), 
to_sfixed(-166326123.0/4294967296.0,1,-nbitq), 
to_sfixed(-110925677.0/4294967296.0,1,-nbitq), 
to_sfixed(333174147.0/4294967296.0,1,-nbitq), 
to_sfixed(378653648.0/4294967296.0,1,-nbitq), 
to_sfixed(-807750987.0/4294967296.0,1,-nbitq), 
to_sfixed(246581867.0/4294967296.0,1,-nbitq), 
to_sfixed(196925362.0/4294967296.0,1,-nbitq), 
to_sfixed(202777887.0/4294967296.0,1,-nbitq), 
to_sfixed(-240913248.0/4294967296.0,1,-nbitq), 
to_sfixed(259399240.0/4294967296.0,1,-nbitq), 
to_sfixed(-69942493.0/4294967296.0,1,-nbitq), 
to_sfixed(265785595.0/4294967296.0,1,-nbitq), 
to_sfixed(276266250.0/4294967296.0,1,-nbitq), 
to_sfixed(-121308179.0/4294967296.0,1,-nbitq), 
to_sfixed(-992789708.0/4294967296.0,1,-nbitq), 
to_sfixed(264551511.0/4294967296.0,1,-nbitq), 
to_sfixed(-111148345.0/4294967296.0,1,-nbitq), 
to_sfixed(-437618993.0/4294967296.0,1,-nbitq), 
to_sfixed(311577283.0/4294967296.0,1,-nbitq), 
to_sfixed(-170654940.0/4294967296.0,1,-nbitq), 
to_sfixed(-363064950.0/4294967296.0,1,-nbitq), 
to_sfixed(-331654244.0/4294967296.0,1,-nbitq), 
to_sfixed(124847452.0/4294967296.0,1,-nbitq), 
to_sfixed(-362890246.0/4294967296.0,1,-nbitq), 
to_sfixed(102673257.0/4294967296.0,1,-nbitq), 
to_sfixed(-71454415.0/4294967296.0,1,-nbitq), 
to_sfixed(-285783883.0/4294967296.0,1,-nbitq), 
to_sfixed(-195646416.0/4294967296.0,1,-nbitq), 
to_sfixed(272047527.0/4294967296.0,1,-nbitq), 
to_sfixed(161374235.0/4294967296.0,1,-nbitq), 
to_sfixed(50218124.0/4294967296.0,1,-nbitq), 
to_sfixed(-282205241.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(549944756.0/4294967296.0,1,-nbitq), 
to_sfixed(1035993861.0/4294967296.0,1,-nbitq), 
to_sfixed(-146569196.0/4294967296.0,1,-nbitq), 
to_sfixed(188708832.0/4294967296.0,1,-nbitq), 
to_sfixed(-140297206.0/4294967296.0,1,-nbitq), 
to_sfixed(-578363115.0/4294967296.0,1,-nbitq), 
to_sfixed(328518531.0/4294967296.0,1,-nbitq), 
to_sfixed(80649739.0/4294967296.0,1,-nbitq), 
to_sfixed(289757555.0/4294967296.0,1,-nbitq), 
to_sfixed(-343850146.0/4294967296.0,1,-nbitq), 
to_sfixed(-506352033.0/4294967296.0,1,-nbitq), 
to_sfixed(212446773.0/4294967296.0,1,-nbitq), 
to_sfixed(-52930206.0/4294967296.0,1,-nbitq), 
to_sfixed(-113360612.0/4294967296.0,1,-nbitq), 
to_sfixed(135284565.0/4294967296.0,1,-nbitq), 
to_sfixed(-509725691.0/4294967296.0,1,-nbitq), 
to_sfixed(373770268.0/4294967296.0,1,-nbitq), 
to_sfixed(-125374401.0/4294967296.0,1,-nbitq), 
to_sfixed(-689233947.0/4294967296.0,1,-nbitq), 
to_sfixed(-221190948.0/4294967296.0,1,-nbitq), 
to_sfixed(229334963.0/4294967296.0,1,-nbitq), 
to_sfixed(215816453.0/4294967296.0,1,-nbitq), 
to_sfixed(56386659.0/4294967296.0,1,-nbitq), 
to_sfixed(408178444.0/4294967296.0,1,-nbitq), 
to_sfixed(-237808111.0/4294967296.0,1,-nbitq), 
to_sfixed(1178173896.0/4294967296.0,1,-nbitq), 
to_sfixed(-114675519.0/4294967296.0,1,-nbitq), 
to_sfixed(-418143835.0/4294967296.0,1,-nbitq), 
to_sfixed(186976926.0/4294967296.0,1,-nbitq), 
to_sfixed(-538765410.0/4294967296.0,1,-nbitq), 
to_sfixed(167195253.0/4294967296.0,1,-nbitq), 
to_sfixed(-428269078.0/4294967296.0,1,-nbitq), 
to_sfixed(235949309.0/4294967296.0,1,-nbitq), 
to_sfixed(-433925342.0/4294967296.0,1,-nbitq), 
to_sfixed(-195845014.0/4294967296.0,1,-nbitq), 
to_sfixed(24345839.0/4294967296.0,1,-nbitq), 
to_sfixed(-355271913.0/4294967296.0,1,-nbitq), 
to_sfixed(-214392303.0/4294967296.0,1,-nbitq), 
to_sfixed(-375486354.0/4294967296.0,1,-nbitq), 
to_sfixed(-230453057.0/4294967296.0,1,-nbitq), 
to_sfixed(281972926.0/4294967296.0,1,-nbitq), 
to_sfixed(-37032287.0/4294967296.0,1,-nbitq), 
to_sfixed(1324887060.0/4294967296.0,1,-nbitq), 
to_sfixed(1128549840.0/4294967296.0,1,-nbitq), 
to_sfixed(-25626026.0/4294967296.0,1,-nbitq), 
to_sfixed(462155988.0/4294967296.0,1,-nbitq), 
to_sfixed(-119980860.0/4294967296.0,1,-nbitq), 
to_sfixed(29436545.0/4294967296.0,1,-nbitq), 
to_sfixed(28959241.0/4294967296.0,1,-nbitq), 
to_sfixed(275442133.0/4294967296.0,1,-nbitq), 
to_sfixed(297703173.0/4294967296.0,1,-nbitq), 
to_sfixed(96367511.0/4294967296.0,1,-nbitq), 
to_sfixed(-740227294.0/4294967296.0,1,-nbitq), 
to_sfixed(169823179.0/4294967296.0,1,-nbitq), 
to_sfixed(1170015479.0/4294967296.0,1,-nbitq), 
to_sfixed(-80842327.0/4294967296.0,1,-nbitq), 
to_sfixed(19907640.0/4294967296.0,1,-nbitq), 
to_sfixed(496606183.0/4294967296.0,1,-nbitq), 
to_sfixed(106210527.0/4294967296.0,1,-nbitq), 
to_sfixed(112322873.0/4294967296.0,1,-nbitq), 
to_sfixed(-151280987.0/4294967296.0,1,-nbitq), 
to_sfixed(-546453249.0/4294967296.0,1,-nbitq), 
to_sfixed(-884333221.0/4294967296.0,1,-nbitq), 
to_sfixed(518004889.0/4294967296.0,1,-nbitq), 
to_sfixed(155950120.0/4294967296.0,1,-nbitq), 
to_sfixed(-173628267.0/4294967296.0,1,-nbitq), 
to_sfixed(30350772.0/4294967296.0,1,-nbitq), 
to_sfixed(962887250.0/4294967296.0,1,-nbitq), 
to_sfixed(385953302.0/4294967296.0,1,-nbitq), 
to_sfixed(-731521958.0/4294967296.0,1,-nbitq), 
to_sfixed(531785440.0/4294967296.0,1,-nbitq), 
to_sfixed(-4723725.0/4294967296.0,1,-nbitq), 
to_sfixed(-79177319.0/4294967296.0,1,-nbitq), 
to_sfixed(-123686254.0/4294967296.0,1,-nbitq), 
to_sfixed(267092094.0/4294967296.0,1,-nbitq), 
to_sfixed(150133928.0/4294967296.0,1,-nbitq), 
to_sfixed(328543989.0/4294967296.0,1,-nbitq), 
to_sfixed(-298882198.0/4294967296.0,1,-nbitq), 
to_sfixed(224774631.0/4294967296.0,1,-nbitq), 
to_sfixed(343201584.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-103125331.0/4294967296.0,1,-nbitq), 
to_sfixed(325908704.0/4294967296.0,1,-nbitq), 
to_sfixed(85439254.0/4294967296.0,1,-nbitq), 
to_sfixed(182485023.0/4294967296.0,1,-nbitq), 
to_sfixed(-436056076.0/4294967296.0,1,-nbitq), 
to_sfixed(-316461075.0/4294967296.0,1,-nbitq), 
to_sfixed(-489396209.0/4294967296.0,1,-nbitq), 
to_sfixed(-534640595.0/4294967296.0,1,-nbitq), 
to_sfixed(314845918.0/4294967296.0,1,-nbitq), 
to_sfixed(417078349.0/4294967296.0,1,-nbitq), 
to_sfixed(-445193224.0/4294967296.0,1,-nbitq), 
to_sfixed(-58603320.0/4294967296.0,1,-nbitq), 
to_sfixed(147854638.0/4294967296.0,1,-nbitq), 
to_sfixed(227477833.0/4294967296.0,1,-nbitq), 
to_sfixed(16278515.0/4294967296.0,1,-nbitq), 
to_sfixed(15437972.0/4294967296.0,1,-nbitq), 
to_sfixed(31373628.0/4294967296.0,1,-nbitq), 
to_sfixed(-42317854.0/4294967296.0,1,-nbitq), 
to_sfixed(-790996985.0/4294967296.0,1,-nbitq), 
to_sfixed(-399365617.0/4294967296.0,1,-nbitq), 
to_sfixed(32411551.0/4294967296.0,1,-nbitq), 
to_sfixed(-206830871.0/4294967296.0,1,-nbitq), 
to_sfixed(-152250661.0/4294967296.0,1,-nbitq), 
to_sfixed(163291205.0/4294967296.0,1,-nbitq), 
to_sfixed(28953622.0/4294967296.0,1,-nbitq), 
to_sfixed(331765546.0/4294967296.0,1,-nbitq), 
to_sfixed(-99091600.0/4294967296.0,1,-nbitq), 
to_sfixed(78024683.0/4294967296.0,1,-nbitq), 
to_sfixed(152891525.0/4294967296.0,1,-nbitq), 
to_sfixed(-161491964.0/4294967296.0,1,-nbitq), 
to_sfixed(360690508.0/4294967296.0,1,-nbitq), 
to_sfixed(-330289427.0/4294967296.0,1,-nbitq), 
to_sfixed(83114506.0/4294967296.0,1,-nbitq), 
to_sfixed(142323855.0/4294967296.0,1,-nbitq), 
to_sfixed(71578086.0/4294967296.0,1,-nbitq), 
to_sfixed(-286983845.0/4294967296.0,1,-nbitq), 
to_sfixed(-194947328.0/4294967296.0,1,-nbitq), 
to_sfixed(-162384769.0/4294967296.0,1,-nbitq), 
to_sfixed(106185767.0/4294967296.0,1,-nbitq), 
to_sfixed(-392565174.0/4294967296.0,1,-nbitq), 
to_sfixed(575605512.0/4294967296.0,1,-nbitq), 
to_sfixed(417341251.0/4294967296.0,1,-nbitq), 
to_sfixed(1426486181.0/4294967296.0,1,-nbitq), 
to_sfixed(1099952173.0/4294967296.0,1,-nbitq), 
to_sfixed(44818939.0/4294967296.0,1,-nbitq), 
to_sfixed(1067895349.0/4294967296.0,1,-nbitq), 
to_sfixed(18619681.0/4294967296.0,1,-nbitq), 
to_sfixed(463384322.0/4294967296.0,1,-nbitq), 
to_sfixed(25467131.0/4294967296.0,1,-nbitq), 
to_sfixed(-82740426.0/4294967296.0,1,-nbitq), 
to_sfixed(22825550.0/4294967296.0,1,-nbitq), 
to_sfixed(-426918202.0/4294967296.0,1,-nbitq), 
to_sfixed(-271663457.0/4294967296.0,1,-nbitq), 
to_sfixed(645875964.0/4294967296.0,1,-nbitq), 
to_sfixed(1268939229.0/4294967296.0,1,-nbitq), 
to_sfixed(-259461621.0/4294967296.0,1,-nbitq), 
to_sfixed(204519038.0/4294967296.0,1,-nbitq), 
to_sfixed(19439102.0/4294967296.0,1,-nbitq), 
to_sfixed(291085519.0/4294967296.0,1,-nbitq), 
to_sfixed(174317340.0/4294967296.0,1,-nbitq), 
to_sfixed(29066524.0/4294967296.0,1,-nbitq), 
to_sfixed(-261179016.0/4294967296.0,1,-nbitq), 
to_sfixed(66250354.0/4294967296.0,1,-nbitq), 
to_sfixed(180787358.0/4294967296.0,1,-nbitq), 
to_sfixed(163128860.0/4294967296.0,1,-nbitq), 
to_sfixed(-318714520.0/4294967296.0,1,-nbitq), 
to_sfixed(175376172.0/4294967296.0,1,-nbitq), 
to_sfixed(972640657.0/4294967296.0,1,-nbitq), 
to_sfixed(317077792.0/4294967296.0,1,-nbitq), 
to_sfixed(-1130143159.0/4294967296.0,1,-nbitq), 
to_sfixed(-53116534.0/4294967296.0,1,-nbitq), 
to_sfixed(-404996917.0/4294967296.0,1,-nbitq), 
to_sfixed(152452461.0/4294967296.0,1,-nbitq), 
to_sfixed(-78172163.0/4294967296.0,1,-nbitq), 
to_sfixed(-55296903.0/4294967296.0,1,-nbitq), 
to_sfixed(-84080713.0/4294967296.0,1,-nbitq), 
to_sfixed(-595644182.0/4294967296.0,1,-nbitq), 
to_sfixed(77914922.0/4294967296.0,1,-nbitq), 
to_sfixed(548037886.0/4294967296.0,1,-nbitq), 
to_sfixed(111385800.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-6627646.0/4294967296.0,1,-nbitq), 
to_sfixed(621639323.0/4294967296.0,1,-nbitq), 
to_sfixed(-284519645.0/4294967296.0,1,-nbitq), 
to_sfixed(70378271.0/4294967296.0,1,-nbitq), 
to_sfixed(-816788536.0/4294967296.0,1,-nbitq), 
to_sfixed(-128764439.0/4294967296.0,1,-nbitq), 
to_sfixed(-69632335.0/4294967296.0,1,-nbitq), 
to_sfixed(-643214902.0/4294967296.0,1,-nbitq), 
to_sfixed(154080057.0/4294967296.0,1,-nbitq), 
to_sfixed(330160464.0/4294967296.0,1,-nbitq), 
to_sfixed(-136117653.0/4294967296.0,1,-nbitq), 
to_sfixed(-336754168.0/4294967296.0,1,-nbitq), 
to_sfixed(250933341.0/4294967296.0,1,-nbitq), 
to_sfixed(-29229292.0/4294967296.0,1,-nbitq), 
to_sfixed(-147979116.0/4294967296.0,1,-nbitq), 
to_sfixed(-354433369.0/4294967296.0,1,-nbitq), 
to_sfixed(104909266.0/4294967296.0,1,-nbitq), 
to_sfixed(-152649201.0/4294967296.0,1,-nbitq), 
to_sfixed(-478643177.0/4294967296.0,1,-nbitq), 
to_sfixed(-372681374.0/4294967296.0,1,-nbitq), 
to_sfixed(23458719.0/4294967296.0,1,-nbitq), 
to_sfixed(-118629089.0/4294967296.0,1,-nbitq), 
to_sfixed(-6892606.0/4294967296.0,1,-nbitq), 
to_sfixed(-331599677.0/4294967296.0,1,-nbitq), 
to_sfixed(-149899699.0/4294967296.0,1,-nbitq), 
to_sfixed(321855965.0/4294967296.0,1,-nbitq), 
to_sfixed(364705002.0/4294967296.0,1,-nbitq), 
to_sfixed(101650.0/4294967296.0,1,-nbitq), 
to_sfixed(275990643.0/4294967296.0,1,-nbitq), 
to_sfixed(-551008028.0/4294967296.0,1,-nbitq), 
to_sfixed(347019304.0/4294967296.0,1,-nbitq), 
to_sfixed(273181713.0/4294967296.0,1,-nbitq), 
to_sfixed(462951182.0/4294967296.0,1,-nbitq), 
to_sfixed(-233071374.0/4294967296.0,1,-nbitq), 
to_sfixed(-7493068.0/4294967296.0,1,-nbitq), 
to_sfixed(-544360831.0/4294967296.0,1,-nbitq), 
to_sfixed(148603398.0/4294967296.0,1,-nbitq), 
to_sfixed(14204593.0/4294967296.0,1,-nbitq), 
to_sfixed(-400935763.0/4294967296.0,1,-nbitq), 
to_sfixed(203906776.0/4294967296.0,1,-nbitq), 
to_sfixed(-241247264.0/4294967296.0,1,-nbitq), 
to_sfixed(292107068.0/4294967296.0,1,-nbitq), 
to_sfixed(1174458796.0/4294967296.0,1,-nbitq), 
to_sfixed(702822067.0/4294967296.0,1,-nbitq), 
to_sfixed(225792485.0/4294967296.0,1,-nbitq), 
to_sfixed(297449634.0/4294967296.0,1,-nbitq), 
to_sfixed(-232999416.0/4294967296.0,1,-nbitq), 
to_sfixed(688343034.0/4294967296.0,1,-nbitq), 
to_sfixed(-161948814.0/4294967296.0,1,-nbitq), 
to_sfixed(530510641.0/4294967296.0,1,-nbitq), 
to_sfixed(484657936.0/4294967296.0,1,-nbitq), 
to_sfixed(-657041439.0/4294967296.0,1,-nbitq), 
to_sfixed(61218543.0/4294967296.0,1,-nbitq), 
to_sfixed(488909565.0/4294967296.0,1,-nbitq), 
to_sfixed(947493563.0/4294967296.0,1,-nbitq), 
to_sfixed(-182845.0/4294967296.0,1,-nbitq), 
to_sfixed(138906444.0/4294967296.0,1,-nbitq), 
to_sfixed(-398606316.0/4294967296.0,1,-nbitq), 
to_sfixed(125515555.0/4294967296.0,1,-nbitq), 
to_sfixed(-38351924.0/4294967296.0,1,-nbitq), 
to_sfixed(132583521.0/4294967296.0,1,-nbitq), 
to_sfixed(-622353913.0/4294967296.0,1,-nbitq), 
to_sfixed(148528896.0/4294967296.0,1,-nbitq), 
to_sfixed(-143387053.0/4294967296.0,1,-nbitq), 
to_sfixed(-52061282.0/4294967296.0,1,-nbitq), 
to_sfixed(-211324164.0/4294967296.0,1,-nbitq), 
to_sfixed(-371855957.0/4294967296.0,1,-nbitq), 
to_sfixed(1200148685.0/4294967296.0,1,-nbitq), 
to_sfixed(205953104.0/4294967296.0,1,-nbitq), 
to_sfixed(-440637247.0/4294967296.0,1,-nbitq), 
to_sfixed(336640025.0/4294967296.0,1,-nbitq), 
to_sfixed(-148876577.0/4294967296.0,1,-nbitq), 
to_sfixed(44476189.0/4294967296.0,1,-nbitq), 
to_sfixed(-35160248.0/4294967296.0,1,-nbitq), 
to_sfixed(-326310327.0/4294967296.0,1,-nbitq), 
to_sfixed(-233176616.0/4294967296.0,1,-nbitq), 
to_sfixed(-344297152.0/4294967296.0,1,-nbitq), 
to_sfixed(-324919060.0/4294967296.0,1,-nbitq), 
to_sfixed(227442092.0/4294967296.0,1,-nbitq), 
to_sfixed(47108465.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-71687975.0/4294967296.0,1,-nbitq), 
to_sfixed(831424971.0/4294967296.0,1,-nbitq), 
to_sfixed(33615188.0/4294967296.0,1,-nbitq), 
to_sfixed(-20563036.0/4294967296.0,1,-nbitq), 
to_sfixed(-290593076.0/4294967296.0,1,-nbitq), 
to_sfixed(-356764365.0/4294967296.0,1,-nbitq), 
to_sfixed(-481613933.0/4294967296.0,1,-nbitq), 
to_sfixed(-220202807.0/4294967296.0,1,-nbitq), 
to_sfixed(445763662.0/4294967296.0,1,-nbitq), 
to_sfixed(347055438.0/4294967296.0,1,-nbitq), 
to_sfixed(300013122.0/4294967296.0,1,-nbitq), 
to_sfixed(-25899377.0/4294967296.0,1,-nbitq), 
to_sfixed(408579494.0/4294967296.0,1,-nbitq), 
to_sfixed(-269847991.0/4294967296.0,1,-nbitq), 
to_sfixed(-458073582.0/4294967296.0,1,-nbitq), 
to_sfixed(141000329.0/4294967296.0,1,-nbitq), 
to_sfixed(-335422413.0/4294967296.0,1,-nbitq), 
to_sfixed(-267540640.0/4294967296.0,1,-nbitq), 
to_sfixed(-695621557.0/4294967296.0,1,-nbitq), 
to_sfixed(-327440162.0/4294967296.0,1,-nbitq), 
to_sfixed(-109352886.0/4294967296.0,1,-nbitq), 
to_sfixed(-416435794.0/4294967296.0,1,-nbitq), 
to_sfixed(-288666646.0/4294967296.0,1,-nbitq), 
to_sfixed(541572604.0/4294967296.0,1,-nbitq), 
to_sfixed(58213548.0/4294967296.0,1,-nbitq), 
to_sfixed(237504960.0/4294967296.0,1,-nbitq), 
to_sfixed(-243646384.0/4294967296.0,1,-nbitq), 
to_sfixed(-171205940.0/4294967296.0,1,-nbitq), 
to_sfixed(109120506.0/4294967296.0,1,-nbitq), 
to_sfixed(-31929158.0/4294967296.0,1,-nbitq), 
to_sfixed(-137437453.0/4294967296.0,1,-nbitq), 
to_sfixed(213706545.0/4294967296.0,1,-nbitq), 
to_sfixed(310511685.0/4294967296.0,1,-nbitq), 
to_sfixed(-630128330.0/4294967296.0,1,-nbitq), 
to_sfixed(289477570.0/4294967296.0,1,-nbitq), 
to_sfixed(22545820.0/4294967296.0,1,-nbitq), 
to_sfixed(205140803.0/4294967296.0,1,-nbitq), 
to_sfixed(-86024209.0/4294967296.0,1,-nbitq), 
to_sfixed(-128146291.0/4294967296.0,1,-nbitq), 
to_sfixed(-124751765.0/4294967296.0,1,-nbitq), 
to_sfixed(-96876908.0/4294967296.0,1,-nbitq), 
to_sfixed(-38136231.0/4294967296.0,1,-nbitq), 
to_sfixed(1080668064.0/4294967296.0,1,-nbitq), 
to_sfixed(1155358908.0/4294967296.0,1,-nbitq), 
to_sfixed(112085378.0/4294967296.0,1,-nbitq), 
to_sfixed(579460457.0/4294967296.0,1,-nbitq), 
to_sfixed(-376354080.0/4294967296.0,1,-nbitq), 
to_sfixed(284236635.0/4294967296.0,1,-nbitq), 
to_sfixed(220690655.0/4294967296.0,1,-nbitq), 
to_sfixed(258224608.0/4294967296.0,1,-nbitq), 
to_sfixed(508363657.0/4294967296.0,1,-nbitq), 
to_sfixed(-150001694.0/4294967296.0,1,-nbitq), 
to_sfixed(626704418.0/4294967296.0,1,-nbitq), 
to_sfixed(143250590.0/4294967296.0,1,-nbitq), 
to_sfixed(1023225346.0/4294967296.0,1,-nbitq), 
to_sfixed(-182849444.0/4294967296.0,1,-nbitq), 
to_sfixed(136681266.0/4294967296.0,1,-nbitq), 
to_sfixed(313227.0/4294967296.0,1,-nbitq), 
to_sfixed(220076510.0/4294967296.0,1,-nbitq), 
to_sfixed(-2237376.0/4294967296.0,1,-nbitq), 
to_sfixed(17010668.0/4294967296.0,1,-nbitq), 
to_sfixed(-788491630.0/4294967296.0,1,-nbitq), 
to_sfixed(48400685.0/4294967296.0,1,-nbitq), 
to_sfixed(157286835.0/4294967296.0,1,-nbitq), 
to_sfixed(71113307.0/4294967296.0,1,-nbitq), 
to_sfixed(126763015.0/4294967296.0,1,-nbitq), 
to_sfixed(-466823245.0/4294967296.0,1,-nbitq), 
to_sfixed(1408162747.0/4294967296.0,1,-nbitq), 
to_sfixed(272645694.0/4294967296.0,1,-nbitq), 
to_sfixed(-283278645.0/4294967296.0,1,-nbitq), 
to_sfixed(326260498.0/4294967296.0,1,-nbitq), 
to_sfixed(108996679.0/4294967296.0,1,-nbitq), 
to_sfixed(370848010.0/4294967296.0,1,-nbitq), 
to_sfixed(173492929.0/4294967296.0,1,-nbitq), 
to_sfixed(-83208619.0/4294967296.0,1,-nbitq), 
to_sfixed(576765502.0/4294967296.0,1,-nbitq), 
to_sfixed(-1197202972.0/4294967296.0,1,-nbitq), 
to_sfixed(355161117.0/4294967296.0,1,-nbitq), 
to_sfixed(641937713.0/4294967296.0,1,-nbitq), 
to_sfixed(13247402.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-19855366.0/4294967296.0,1,-nbitq), 
to_sfixed(1467334128.0/4294967296.0,1,-nbitq), 
to_sfixed(-146218021.0/4294967296.0,1,-nbitq), 
to_sfixed(288297933.0/4294967296.0,1,-nbitq), 
to_sfixed(-262857472.0/4294967296.0,1,-nbitq), 
to_sfixed(-31792986.0/4294967296.0,1,-nbitq), 
to_sfixed(-132524306.0/4294967296.0,1,-nbitq), 
to_sfixed(31941515.0/4294967296.0,1,-nbitq), 
to_sfixed(542767834.0/4294967296.0,1,-nbitq), 
to_sfixed(-300533387.0/4294967296.0,1,-nbitq), 
to_sfixed(319832792.0/4294967296.0,1,-nbitq), 
to_sfixed(152461097.0/4294967296.0,1,-nbitq), 
to_sfixed(303866725.0/4294967296.0,1,-nbitq), 
to_sfixed(-256624156.0/4294967296.0,1,-nbitq), 
to_sfixed(-421702550.0/4294967296.0,1,-nbitq), 
to_sfixed(297441832.0/4294967296.0,1,-nbitq), 
to_sfixed(342108800.0/4294967296.0,1,-nbitq), 
to_sfixed(221938285.0/4294967296.0,1,-nbitq), 
to_sfixed(172823384.0/4294967296.0,1,-nbitq), 
to_sfixed(45206177.0/4294967296.0,1,-nbitq), 
to_sfixed(35727594.0/4294967296.0,1,-nbitq), 
to_sfixed(440035746.0/4294967296.0,1,-nbitq), 
to_sfixed(130031417.0/4294967296.0,1,-nbitq), 
to_sfixed(586784895.0/4294967296.0,1,-nbitq), 
to_sfixed(258309786.0/4294967296.0,1,-nbitq), 
to_sfixed(260760567.0/4294967296.0,1,-nbitq), 
to_sfixed(-248084579.0/4294967296.0,1,-nbitq), 
to_sfixed(6280564.0/4294967296.0,1,-nbitq), 
to_sfixed(387991418.0/4294967296.0,1,-nbitq), 
to_sfixed(-198254000.0/4294967296.0,1,-nbitq), 
to_sfixed(261469946.0/4294967296.0,1,-nbitq), 
to_sfixed(-100402754.0/4294967296.0,1,-nbitq), 
to_sfixed(802522663.0/4294967296.0,1,-nbitq), 
to_sfixed(-769262484.0/4294967296.0,1,-nbitq), 
to_sfixed(1428012.0/4294967296.0,1,-nbitq), 
to_sfixed(-416085771.0/4294967296.0,1,-nbitq), 
to_sfixed(36999020.0/4294967296.0,1,-nbitq), 
to_sfixed(240355179.0/4294967296.0,1,-nbitq), 
to_sfixed(-360840221.0/4294967296.0,1,-nbitq), 
to_sfixed(35081710.0/4294967296.0,1,-nbitq), 
to_sfixed(-47943817.0/4294967296.0,1,-nbitq), 
to_sfixed(295294860.0/4294967296.0,1,-nbitq), 
to_sfixed(630336817.0/4294967296.0,1,-nbitq), 
to_sfixed(828670224.0/4294967296.0,1,-nbitq), 
to_sfixed(449127570.0/4294967296.0,1,-nbitq), 
to_sfixed(1044294454.0/4294967296.0,1,-nbitq), 
to_sfixed(174872530.0/4294967296.0,1,-nbitq), 
to_sfixed(-152013458.0/4294967296.0,1,-nbitq), 
to_sfixed(-39042424.0/4294967296.0,1,-nbitq), 
to_sfixed(-168638525.0/4294967296.0,1,-nbitq), 
to_sfixed(59461937.0/4294967296.0,1,-nbitq), 
to_sfixed(-634973788.0/4294967296.0,1,-nbitq), 
to_sfixed(608935418.0/4294967296.0,1,-nbitq), 
to_sfixed(36771665.0/4294967296.0,1,-nbitq), 
to_sfixed(587777892.0/4294967296.0,1,-nbitq), 
to_sfixed(-32384365.0/4294967296.0,1,-nbitq), 
to_sfixed(-430242883.0/4294967296.0,1,-nbitq), 
to_sfixed(119429948.0/4294967296.0,1,-nbitq), 
to_sfixed(-17216112.0/4294967296.0,1,-nbitq), 
to_sfixed(-89928467.0/4294967296.0,1,-nbitq), 
to_sfixed(119831570.0/4294967296.0,1,-nbitq), 
to_sfixed(-340003544.0/4294967296.0,1,-nbitq), 
to_sfixed(110670803.0/4294967296.0,1,-nbitq), 
to_sfixed(-243596748.0/4294967296.0,1,-nbitq), 
to_sfixed(207280614.0/4294967296.0,1,-nbitq), 
to_sfixed(-328786502.0/4294967296.0,1,-nbitq), 
to_sfixed(-550031333.0/4294967296.0,1,-nbitq), 
to_sfixed(2166480694.0/4294967296.0,1,-nbitq), 
to_sfixed(68711143.0/4294967296.0,1,-nbitq), 
to_sfixed(-333159490.0/4294967296.0,1,-nbitq), 
to_sfixed(286643791.0/4294967296.0,1,-nbitq), 
to_sfixed(305206232.0/4294967296.0,1,-nbitq), 
to_sfixed(197612480.0/4294967296.0,1,-nbitq), 
to_sfixed(-27861872.0/4294967296.0,1,-nbitq), 
to_sfixed(-229355320.0/4294967296.0,1,-nbitq), 
to_sfixed(646945710.0/4294967296.0,1,-nbitq), 
to_sfixed(-1058553750.0/4294967296.0,1,-nbitq), 
to_sfixed(-248160809.0/4294967296.0,1,-nbitq), 
to_sfixed(737340113.0/4294967296.0,1,-nbitq), 
to_sfixed(-165264744.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(101375284.0/4294967296.0,1,-nbitq), 
to_sfixed(978236189.0/4294967296.0,1,-nbitq), 
to_sfixed(-16449627.0/4294967296.0,1,-nbitq), 
to_sfixed(-130939256.0/4294967296.0,1,-nbitq), 
to_sfixed(-155178680.0/4294967296.0,1,-nbitq), 
to_sfixed(259204714.0/4294967296.0,1,-nbitq), 
to_sfixed(58790616.0/4294967296.0,1,-nbitq), 
to_sfixed(-46310186.0/4294967296.0,1,-nbitq), 
to_sfixed(774424944.0/4294967296.0,1,-nbitq), 
to_sfixed(106221281.0/4294967296.0,1,-nbitq), 
to_sfixed(373960917.0/4294967296.0,1,-nbitq), 
to_sfixed(337601713.0/4294967296.0,1,-nbitq), 
to_sfixed(52811482.0/4294967296.0,1,-nbitq), 
to_sfixed(-278848898.0/4294967296.0,1,-nbitq), 
to_sfixed(-120953869.0/4294967296.0,1,-nbitq), 
to_sfixed(-187638346.0/4294967296.0,1,-nbitq), 
to_sfixed(-367966111.0/4294967296.0,1,-nbitq), 
to_sfixed(303906652.0/4294967296.0,1,-nbitq), 
to_sfixed(532511091.0/4294967296.0,1,-nbitq), 
to_sfixed(-104247580.0/4294967296.0,1,-nbitq), 
to_sfixed(376673629.0/4294967296.0,1,-nbitq), 
to_sfixed(-13064396.0/4294967296.0,1,-nbitq), 
to_sfixed(208660416.0/4294967296.0,1,-nbitq), 
to_sfixed(219789675.0/4294967296.0,1,-nbitq), 
to_sfixed(368885270.0/4294967296.0,1,-nbitq), 
to_sfixed(223530474.0/4294967296.0,1,-nbitq), 
to_sfixed(-21381929.0/4294967296.0,1,-nbitq), 
to_sfixed(281716146.0/4294967296.0,1,-nbitq), 
to_sfixed(178199600.0/4294967296.0,1,-nbitq), 
to_sfixed(444698061.0/4294967296.0,1,-nbitq), 
to_sfixed(164653765.0/4294967296.0,1,-nbitq), 
to_sfixed(-348344104.0/4294967296.0,1,-nbitq), 
to_sfixed(413321493.0/4294967296.0,1,-nbitq), 
to_sfixed(-375802211.0/4294967296.0,1,-nbitq), 
to_sfixed(710858124.0/4294967296.0,1,-nbitq), 
to_sfixed(568122167.0/4294967296.0,1,-nbitq), 
to_sfixed(351591976.0/4294967296.0,1,-nbitq), 
to_sfixed(145651581.0/4294967296.0,1,-nbitq), 
to_sfixed(44111674.0/4294967296.0,1,-nbitq), 
to_sfixed(-293412447.0/4294967296.0,1,-nbitq), 
to_sfixed(-107247600.0/4294967296.0,1,-nbitq), 
to_sfixed(763190557.0/4294967296.0,1,-nbitq), 
to_sfixed(619620125.0/4294967296.0,1,-nbitq), 
to_sfixed(468494595.0/4294967296.0,1,-nbitq), 
to_sfixed(190096594.0/4294967296.0,1,-nbitq), 
to_sfixed(742840215.0/4294967296.0,1,-nbitq), 
to_sfixed(201844675.0/4294967296.0,1,-nbitq), 
to_sfixed(-8716735.0/4294967296.0,1,-nbitq), 
to_sfixed(-212437249.0/4294967296.0,1,-nbitq), 
to_sfixed(-201222100.0/4294967296.0,1,-nbitq), 
to_sfixed(-222069373.0/4294967296.0,1,-nbitq), 
to_sfixed(-512219734.0/4294967296.0,1,-nbitq), 
to_sfixed(-176173652.0/4294967296.0,1,-nbitq), 
to_sfixed(140356557.0/4294967296.0,1,-nbitq), 
to_sfixed(837336468.0/4294967296.0,1,-nbitq), 
to_sfixed(-598941277.0/4294967296.0,1,-nbitq), 
to_sfixed(-589978130.0/4294967296.0,1,-nbitq), 
to_sfixed(63464943.0/4294967296.0,1,-nbitq), 
to_sfixed(378214895.0/4294967296.0,1,-nbitq), 
to_sfixed(-245962091.0/4294967296.0,1,-nbitq), 
to_sfixed(-329077361.0/4294967296.0,1,-nbitq), 
to_sfixed(147814427.0/4294967296.0,1,-nbitq), 
to_sfixed(124313423.0/4294967296.0,1,-nbitq), 
to_sfixed(-212036002.0/4294967296.0,1,-nbitq), 
to_sfixed(200570472.0/4294967296.0,1,-nbitq), 
to_sfixed(-130922100.0/4294967296.0,1,-nbitq), 
to_sfixed(-564165581.0/4294967296.0,1,-nbitq), 
to_sfixed(1670610797.0/4294967296.0,1,-nbitq), 
to_sfixed(-351989786.0/4294967296.0,1,-nbitq), 
to_sfixed(-756108083.0/4294967296.0,1,-nbitq), 
to_sfixed(145801346.0/4294967296.0,1,-nbitq), 
to_sfixed(-96892485.0/4294967296.0,1,-nbitq), 
to_sfixed(-396502033.0/4294967296.0,1,-nbitq), 
to_sfixed(-160151367.0/4294967296.0,1,-nbitq), 
to_sfixed(-77504207.0/4294967296.0,1,-nbitq), 
to_sfixed(901102301.0/4294967296.0,1,-nbitq), 
to_sfixed(-424634793.0/4294967296.0,1,-nbitq), 
to_sfixed(119538923.0/4294967296.0,1,-nbitq), 
to_sfixed(455506078.0/4294967296.0,1,-nbitq), 
to_sfixed(322175532.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(17985000.0/4294967296.0,1,-nbitq), 
to_sfixed(428111666.0/4294967296.0,1,-nbitq), 
to_sfixed(375057129.0/4294967296.0,1,-nbitq), 
to_sfixed(429526693.0/4294967296.0,1,-nbitq), 
to_sfixed(-294524216.0/4294967296.0,1,-nbitq), 
to_sfixed(952582913.0/4294967296.0,1,-nbitq), 
to_sfixed(173043371.0/4294967296.0,1,-nbitq), 
to_sfixed(38776152.0/4294967296.0,1,-nbitq), 
to_sfixed(200997375.0/4294967296.0,1,-nbitq), 
to_sfixed(134761013.0/4294967296.0,1,-nbitq), 
to_sfixed(29400199.0/4294967296.0,1,-nbitq), 
to_sfixed(-110511136.0/4294967296.0,1,-nbitq), 
to_sfixed(-452141837.0/4294967296.0,1,-nbitq), 
to_sfixed(-200839300.0/4294967296.0,1,-nbitq), 
to_sfixed(-122113266.0/4294967296.0,1,-nbitq), 
to_sfixed(109081334.0/4294967296.0,1,-nbitq), 
to_sfixed(186308425.0/4294967296.0,1,-nbitq), 
to_sfixed(12770438.0/4294967296.0,1,-nbitq), 
to_sfixed(616932797.0/4294967296.0,1,-nbitq), 
to_sfixed(333263788.0/4294967296.0,1,-nbitq), 
to_sfixed(1986320.0/4294967296.0,1,-nbitq), 
to_sfixed(494512311.0/4294967296.0,1,-nbitq), 
to_sfixed(72758358.0/4294967296.0,1,-nbitq), 
to_sfixed(588162128.0/4294967296.0,1,-nbitq), 
to_sfixed(158834570.0/4294967296.0,1,-nbitq), 
to_sfixed(348662679.0/4294967296.0,1,-nbitq), 
to_sfixed(-5707258.0/4294967296.0,1,-nbitq), 
to_sfixed(168948861.0/4294967296.0,1,-nbitq), 
to_sfixed(-427268302.0/4294967296.0,1,-nbitq), 
to_sfixed(223253656.0/4294967296.0,1,-nbitq), 
to_sfixed(-433496380.0/4294967296.0,1,-nbitq), 
to_sfixed(-385414110.0/4294967296.0,1,-nbitq), 
to_sfixed(205527640.0/4294967296.0,1,-nbitq), 
to_sfixed(-714148174.0/4294967296.0,1,-nbitq), 
to_sfixed(843185559.0/4294967296.0,1,-nbitq), 
to_sfixed(443319288.0/4294967296.0,1,-nbitq), 
to_sfixed(278627106.0/4294967296.0,1,-nbitq), 
to_sfixed(101793804.0/4294967296.0,1,-nbitq), 
to_sfixed(-482828296.0/4294967296.0,1,-nbitq), 
to_sfixed(-102291329.0/4294967296.0,1,-nbitq), 
to_sfixed(-254748857.0/4294967296.0,1,-nbitq), 
to_sfixed(628150726.0/4294967296.0,1,-nbitq), 
to_sfixed(826143003.0/4294967296.0,1,-nbitq), 
to_sfixed(269336001.0/4294967296.0,1,-nbitq), 
to_sfixed(556792153.0/4294967296.0,1,-nbitq), 
to_sfixed(755986487.0/4294967296.0,1,-nbitq), 
to_sfixed(-28529326.0/4294967296.0,1,-nbitq), 
to_sfixed(-431298283.0/4294967296.0,1,-nbitq), 
to_sfixed(330556508.0/4294967296.0,1,-nbitq), 
to_sfixed(-111703647.0/4294967296.0,1,-nbitq), 
to_sfixed(-273844708.0/4294967296.0,1,-nbitq), 
to_sfixed(-122312941.0/4294967296.0,1,-nbitq), 
to_sfixed(23533733.0/4294967296.0,1,-nbitq), 
to_sfixed(120760974.0/4294967296.0,1,-nbitq), 
to_sfixed(434239508.0/4294967296.0,1,-nbitq), 
to_sfixed(165551552.0/4294967296.0,1,-nbitq), 
to_sfixed(-612034565.0/4294967296.0,1,-nbitq), 
to_sfixed(329897942.0/4294967296.0,1,-nbitq), 
to_sfixed(237790916.0/4294967296.0,1,-nbitq), 
to_sfixed(413113929.0/4294967296.0,1,-nbitq), 
to_sfixed(-213324737.0/4294967296.0,1,-nbitq), 
to_sfixed(511072297.0/4294967296.0,1,-nbitq), 
to_sfixed(-325204857.0/4294967296.0,1,-nbitq), 
to_sfixed(262318876.0/4294967296.0,1,-nbitq), 
to_sfixed(90931156.0/4294967296.0,1,-nbitq), 
to_sfixed(-95667007.0/4294967296.0,1,-nbitq), 
to_sfixed(-119875150.0/4294967296.0,1,-nbitq), 
to_sfixed(608991031.0/4294967296.0,1,-nbitq), 
to_sfixed(-145428016.0/4294967296.0,1,-nbitq), 
to_sfixed(-651226165.0/4294967296.0,1,-nbitq), 
to_sfixed(238593046.0/4294967296.0,1,-nbitq), 
to_sfixed(428150688.0/4294967296.0,1,-nbitq), 
to_sfixed(-275638113.0/4294967296.0,1,-nbitq), 
to_sfixed(309774270.0/4294967296.0,1,-nbitq), 
to_sfixed(283242270.0/4294967296.0,1,-nbitq), 
to_sfixed(388159930.0/4294967296.0,1,-nbitq), 
to_sfixed(-351130730.0/4294967296.0,1,-nbitq), 
to_sfixed(208625840.0/4294967296.0,1,-nbitq), 
to_sfixed(596010865.0/4294967296.0,1,-nbitq), 
to_sfixed(-133713357.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-125423125.0/4294967296.0,1,-nbitq), 
to_sfixed(686924811.0/4294967296.0,1,-nbitq), 
to_sfixed(-163370718.0/4294967296.0,1,-nbitq), 
to_sfixed(-162008711.0/4294967296.0,1,-nbitq), 
to_sfixed(217741359.0/4294967296.0,1,-nbitq), 
to_sfixed(633929395.0/4294967296.0,1,-nbitq), 
to_sfixed(274060336.0/4294967296.0,1,-nbitq), 
to_sfixed(-130745696.0/4294967296.0,1,-nbitq), 
to_sfixed(28125108.0/4294967296.0,1,-nbitq), 
to_sfixed(252204321.0/4294967296.0,1,-nbitq), 
to_sfixed(291748963.0/4294967296.0,1,-nbitq), 
to_sfixed(-232427780.0/4294967296.0,1,-nbitq), 
to_sfixed(-259821501.0/4294967296.0,1,-nbitq), 
to_sfixed(314952669.0/4294967296.0,1,-nbitq), 
to_sfixed(67536555.0/4294967296.0,1,-nbitq), 
to_sfixed(354465347.0/4294967296.0,1,-nbitq), 
to_sfixed(-95956959.0/4294967296.0,1,-nbitq), 
to_sfixed(348637839.0/4294967296.0,1,-nbitq), 
to_sfixed(300825252.0/4294967296.0,1,-nbitq), 
to_sfixed(-292021332.0/4294967296.0,1,-nbitq), 
to_sfixed(-343251532.0/4294967296.0,1,-nbitq), 
to_sfixed(628470618.0/4294967296.0,1,-nbitq), 
to_sfixed(208290812.0/4294967296.0,1,-nbitq), 
to_sfixed(-276882842.0/4294967296.0,1,-nbitq), 
to_sfixed(-263208858.0/4294967296.0,1,-nbitq), 
to_sfixed(214189966.0/4294967296.0,1,-nbitq), 
to_sfixed(18767978.0/4294967296.0,1,-nbitq), 
to_sfixed(465721073.0/4294967296.0,1,-nbitq), 
to_sfixed(19797547.0/4294967296.0,1,-nbitq), 
to_sfixed(-214147130.0/4294967296.0,1,-nbitq), 
to_sfixed(18902397.0/4294967296.0,1,-nbitq), 
to_sfixed(-56593468.0/4294967296.0,1,-nbitq), 
to_sfixed(669149274.0/4294967296.0,1,-nbitq), 
to_sfixed(32896130.0/4294967296.0,1,-nbitq), 
to_sfixed(630632695.0/4294967296.0,1,-nbitq), 
to_sfixed(213365655.0/4294967296.0,1,-nbitq), 
to_sfixed(567525816.0/4294967296.0,1,-nbitq), 
to_sfixed(-220043033.0/4294967296.0,1,-nbitq), 
to_sfixed(-407476298.0/4294967296.0,1,-nbitq), 
to_sfixed(-62262455.0/4294967296.0,1,-nbitq), 
to_sfixed(133262199.0/4294967296.0,1,-nbitq), 
to_sfixed(-145973142.0/4294967296.0,1,-nbitq), 
to_sfixed(459904049.0/4294967296.0,1,-nbitq), 
to_sfixed(70136662.0/4294967296.0,1,-nbitq), 
to_sfixed(354747961.0/4294967296.0,1,-nbitq), 
to_sfixed(386234419.0/4294967296.0,1,-nbitq), 
to_sfixed(228945139.0/4294967296.0,1,-nbitq), 
to_sfixed(-171925121.0/4294967296.0,1,-nbitq), 
to_sfixed(83970876.0/4294967296.0,1,-nbitq), 
to_sfixed(60361994.0/4294967296.0,1,-nbitq), 
to_sfixed(323713795.0/4294967296.0,1,-nbitq), 
to_sfixed(-5577126.0/4294967296.0,1,-nbitq), 
to_sfixed(59174400.0/4294967296.0,1,-nbitq), 
to_sfixed(-46273055.0/4294967296.0,1,-nbitq), 
to_sfixed(431465758.0/4294967296.0,1,-nbitq), 
to_sfixed(136165671.0/4294967296.0,1,-nbitq), 
to_sfixed(-505560688.0/4294967296.0,1,-nbitq), 
to_sfixed(311203692.0/4294967296.0,1,-nbitq), 
to_sfixed(-170415298.0/4294967296.0,1,-nbitq), 
to_sfixed(394422187.0/4294967296.0,1,-nbitq), 
to_sfixed(63938982.0/4294967296.0,1,-nbitq), 
to_sfixed(134508128.0/4294967296.0,1,-nbitq), 
to_sfixed(437437108.0/4294967296.0,1,-nbitq), 
to_sfixed(47009815.0/4294967296.0,1,-nbitq), 
to_sfixed(-302737335.0/4294967296.0,1,-nbitq), 
to_sfixed(-344358570.0/4294967296.0,1,-nbitq), 
to_sfixed(-367950665.0/4294967296.0,1,-nbitq), 
to_sfixed(694199585.0/4294967296.0,1,-nbitq), 
to_sfixed(156890664.0/4294967296.0,1,-nbitq), 
to_sfixed(-232728621.0/4294967296.0,1,-nbitq), 
to_sfixed(264023118.0/4294967296.0,1,-nbitq), 
to_sfixed(-142566489.0/4294967296.0,1,-nbitq), 
to_sfixed(-358466138.0/4294967296.0,1,-nbitq), 
to_sfixed(219242753.0/4294967296.0,1,-nbitq), 
to_sfixed(84433239.0/4294967296.0,1,-nbitq), 
to_sfixed(363191732.0/4294967296.0,1,-nbitq), 
to_sfixed(-322129694.0/4294967296.0,1,-nbitq), 
to_sfixed(-641648086.0/4294967296.0,1,-nbitq), 
to_sfixed(-19084983.0/4294967296.0,1,-nbitq), 
to_sfixed(-306879841.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(374007806.0/4294967296.0,1,-nbitq), 
to_sfixed(546197477.0/4294967296.0,1,-nbitq), 
to_sfixed(-125960027.0/4294967296.0,1,-nbitq), 
to_sfixed(47777921.0/4294967296.0,1,-nbitq), 
to_sfixed(389335615.0/4294967296.0,1,-nbitq), 
to_sfixed(409804168.0/4294967296.0,1,-nbitq), 
to_sfixed(144177939.0/4294967296.0,1,-nbitq), 
to_sfixed(-141732522.0/4294967296.0,1,-nbitq), 
to_sfixed(-171967287.0/4294967296.0,1,-nbitq), 
to_sfixed(-95796413.0/4294967296.0,1,-nbitq), 
to_sfixed(67463205.0/4294967296.0,1,-nbitq), 
to_sfixed(219847555.0/4294967296.0,1,-nbitq), 
to_sfixed(-435789094.0/4294967296.0,1,-nbitq), 
to_sfixed(427081825.0/4294967296.0,1,-nbitq), 
to_sfixed(-358637438.0/4294967296.0,1,-nbitq), 
to_sfixed(422927424.0/4294967296.0,1,-nbitq), 
to_sfixed(110117687.0/4294967296.0,1,-nbitq), 
to_sfixed(42756255.0/4294967296.0,1,-nbitq), 
to_sfixed(619768665.0/4294967296.0,1,-nbitq), 
to_sfixed(114444615.0/4294967296.0,1,-nbitq), 
to_sfixed(294725010.0/4294967296.0,1,-nbitq), 
to_sfixed(-171736866.0/4294967296.0,1,-nbitq), 
to_sfixed(498990441.0/4294967296.0,1,-nbitq), 
to_sfixed(114124505.0/4294967296.0,1,-nbitq), 
to_sfixed(-59040761.0/4294967296.0,1,-nbitq), 
to_sfixed(445800411.0/4294967296.0,1,-nbitq), 
to_sfixed(-316170136.0/4294967296.0,1,-nbitq), 
to_sfixed(-313814225.0/4294967296.0,1,-nbitq), 
to_sfixed(-1571539.0/4294967296.0,1,-nbitq), 
to_sfixed(388379447.0/4294967296.0,1,-nbitq), 
to_sfixed(188332784.0/4294967296.0,1,-nbitq), 
to_sfixed(-350777179.0/4294967296.0,1,-nbitq), 
to_sfixed(319200055.0/4294967296.0,1,-nbitq), 
to_sfixed(9734942.0/4294967296.0,1,-nbitq), 
to_sfixed(-71546027.0/4294967296.0,1,-nbitq), 
to_sfixed(-436130091.0/4294967296.0,1,-nbitq), 
to_sfixed(-84054127.0/4294967296.0,1,-nbitq), 
to_sfixed(246164457.0/4294967296.0,1,-nbitq), 
to_sfixed(-356893861.0/4294967296.0,1,-nbitq), 
to_sfixed(335760866.0/4294967296.0,1,-nbitq), 
to_sfixed(-302442819.0/4294967296.0,1,-nbitq), 
to_sfixed(-60354847.0/4294967296.0,1,-nbitq), 
to_sfixed(31622467.0/4294967296.0,1,-nbitq), 
to_sfixed(321457356.0/4294967296.0,1,-nbitq), 
to_sfixed(-308752769.0/4294967296.0,1,-nbitq), 
to_sfixed(210568041.0/4294967296.0,1,-nbitq), 
to_sfixed(-229853876.0/4294967296.0,1,-nbitq), 
to_sfixed(-2031990.0/4294967296.0,1,-nbitq), 
to_sfixed(-125297315.0/4294967296.0,1,-nbitq), 
to_sfixed(145245875.0/4294967296.0,1,-nbitq), 
to_sfixed(-105258198.0/4294967296.0,1,-nbitq), 
to_sfixed(-315028168.0/4294967296.0,1,-nbitq), 
to_sfixed(-22867693.0/4294967296.0,1,-nbitq), 
to_sfixed(380657914.0/4294967296.0,1,-nbitq), 
to_sfixed(48803394.0/4294967296.0,1,-nbitq), 
to_sfixed(106631049.0/4294967296.0,1,-nbitq), 
to_sfixed(372458643.0/4294967296.0,1,-nbitq), 
to_sfixed(73903745.0/4294967296.0,1,-nbitq), 
to_sfixed(172291685.0/4294967296.0,1,-nbitq), 
to_sfixed(410149438.0/4294967296.0,1,-nbitq), 
to_sfixed(260858155.0/4294967296.0,1,-nbitq), 
to_sfixed(-4692202.0/4294967296.0,1,-nbitq), 
to_sfixed(310231601.0/4294967296.0,1,-nbitq), 
to_sfixed(-87453505.0/4294967296.0,1,-nbitq), 
to_sfixed(208525412.0/4294967296.0,1,-nbitq), 
to_sfixed(-423488113.0/4294967296.0,1,-nbitq), 
to_sfixed(7653564.0/4294967296.0,1,-nbitq), 
to_sfixed(-300985764.0/4294967296.0,1,-nbitq), 
to_sfixed(-153919132.0/4294967296.0,1,-nbitq), 
to_sfixed(224662176.0/4294967296.0,1,-nbitq), 
to_sfixed(-347329396.0/4294967296.0,1,-nbitq), 
to_sfixed(276103588.0/4294967296.0,1,-nbitq), 
to_sfixed(-454967059.0/4294967296.0,1,-nbitq), 
to_sfixed(-128288505.0/4294967296.0,1,-nbitq), 
to_sfixed(438605344.0/4294967296.0,1,-nbitq), 
to_sfixed(116856671.0/4294967296.0,1,-nbitq), 
to_sfixed(-18830489.0/4294967296.0,1,-nbitq), 
to_sfixed(-569294686.0/4294967296.0,1,-nbitq), 
to_sfixed(214554299.0/4294967296.0,1,-nbitq), 
to_sfixed(-122544151.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(103413102.0/4294967296.0,1,-nbitq), 
to_sfixed(-41730293.0/4294967296.0,1,-nbitq), 
to_sfixed(135405551.0/4294967296.0,1,-nbitq), 
to_sfixed(45116814.0/4294967296.0,1,-nbitq), 
to_sfixed(66228513.0/4294967296.0,1,-nbitq), 
to_sfixed(277019958.0/4294967296.0,1,-nbitq), 
to_sfixed(-265641696.0/4294967296.0,1,-nbitq), 
to_sfixed(-376416653.0/4294967296.0,1,-nbitq), 
to_sfixed(-366011494.0/4294967296.0,1,-nbitq), 
to_sfixed(275723148.0/4294967296.0,1,-nbitq), 
to_sfixed(238813561.0/4294967296.0,1,-nbitq), 
to_sfixed(65578309.0/4294967296.0,1,-nbitq), 
to_sfixed(-308150192.0/4294967296.0,1,-nbitq), 
to_sfixed(-160521248.0/4294967296.0,1,-nbitq), 
to_sfixed(140491600.0/4294967296.0,1,-nbitq), 
to_sfixed(-34406050.0/4294967296.0,1,-nbitq), 
to_sfixed(-101741213.0/4294967296.0,1,-nbitq), 
to_sfixed(-402845780.0/4294967296.0,1,-nbitq), 
to_sfixed(324149087.0/4294967296.0,1,-nbitq), 
to_sfixed(-168484145.0/4294967296.0,1,-nbitq), 
to_sfixed(-406040275.0/4294967296.0,1,-nbitq), 
to_sfixed(-130479593.0/4294967296.0,1,-nbitq), 
to_sfixed(244777825.0/4294967296.0,1,-nbitq), 
to_sfixed(166530092.0/4294967296.0,1,-nbitq), 
to_sfixed(-87594697.0/4294967296.0,1,-nbitq), 
to_sfixed(-99968690.0/4294967296.0,1,-nbitq), 
to_sfixed(95531237.0/4294967296.0,1,-nbitq), 
to_sfixed(-413774395.0/4294967296.0,1,-nbitq), 
to_sfixed(-281909333.0/4294967296.0,1,-nbitq), 
to_sfixed(-161904236.0/4294967296.0,1,-nbitq), 
to_sfixed(121490228.0/4294967296.0,1,-nbitq), 
to_sfixed(74138512.0/4294967296.0,1,-nbitq), 
to_sfixed(359977356.0/4294967296.0,1,-nbitq), 
to_sfixed(222584933.0/4294967296.0,1,-nbitq), 
to_sfixed(302254966.0/4294967296.0,1,-nbitq), 
to_sfixed(-16664543.0/4294967296.0,1,-nbitq), 
to_sfixed(-105400069.0/4294967296.0,1,-nbitq), 
to_sfixed(-121375101.0/4294967296.0,1,-nbitq), 
to_sfixed(235670900.0/4294967296.0,1,-nbitq), 
to_sfixed(32165623.0/4294967296.0,1,-nbitq), 
to_sfixed(189991415.0/4294967296.0,1,-nbitq), 
to_sfixed(468620594.0/4294967296.0,1,-nbitq), 
to_sfixed(267112454.0/4294967296.0,1,-nbitq), 
to_sfixed(210859490.0/4294967296.0,1,-nbitq), 
to_sfixed(18408767.0/4294967296.0,1,-nbitq), 
to_sfixed(297642025.0/4294967296.0,1,-nbitq), 
to_sfixed(-148994955.0/4294967296.0,1,-nbitq), 
to_sfixed(3634557.0/4294967296.0,1,-nbitq), 
to_sfixed(-275092739.0/4294967296.0,1,-nbitq), 
to_sfixed(201098600.0/4294967296.0,1,-nbitq), 
to_sfixed(47755070.0/4294967296.0,1,-nbitq), 
to_sfixed(-56681169.0/4294967296.0,1,-nbitq), 
to_sfixed(-31065957.0/4294967296.0,1,-nbitq), 
to_sfixed(72397753.0/4294967296.0,1,-nbitq), 
to_sfixed(-218294025.0/4294967296.0,1,-nbitq), 
to_sfixed(-296396301.0/4294967296.0,1,-nbitq), 
to_sfixed(425647302.0/4294967296.0,1,-nbitq), 
to_sfixed(-286036979.0/4294967296.0,1,-nbitq), 
to_sfixed(-20892477.0/4294967296.0,1,-nbitq), 
to_sfixed(164796811.0/4294967296.0,1,-nbitq), 
to_sfixed(-224104912.0/4294967296.0,1,-nbitq), 
to_sfixed(294166644.0/4294967296.0,1,-nbitq), 
to_sfixed(-287218054.0/4294967296.0,1,-nbitq), 
to_sfixed(-65608899.0/4294967296.0,1,-nbitq), 
to_sfixed(167753055.0/4294967296.0,1,-nbitq), 
to_sfixed(90896986.0/4294967296.0,1,-nbitq), 
to_sfixed(397902229.0/4294967296.0,1,-nbitq), 
to_sfixed(38832588.0/4294967296.0,1,-nbitq), 
to_sfixed(-300970894.0/4294967296.0,1,-nbitq), 
to_sfixed(196820087.0/4294967296.0,1,-nbitq), 
to_sfixed(-428476169.0/4294967296.0,1,-nbitq), 
to_sfixed(102833576.0/4294967296.0,1,-nbitq), 
to_sfixed(-286078952.0/4294967296.0,1,-nbitq), 
to_sfixed(-327732894.0/4294967296.0,1,-nbitq), 
to_sfixed(388555172.0/4294967296.0,1,-nbitq), 
to_sfixed(-491986573.0/4294967296.0,1,-nbitq), 
to_sfixed(37809213.0/4294967296.0,1,-nbitq), 
to_sfixed(-274585610.0/4294967296.0,1,-nbitq), 
to_sfixed(247400719.0/4294967296.0,1,-nbitq), 
to_sfixed(-319255971.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-52726986.0/4294967296.0,1,-nbitq), 
to_sfixed(200894586.0/4294967296.0,1,-nbitq), 
to_sfixed(-206938156.0/4294967296.0,1,-nbitq), 
to_sfixed(249203101.0/4294967296.0,1,-nbitq), 
to_sfixed(-260392355.0/4294967296.0,1,-nbitq), 
to_sfixed(253198755.0/4294967296.0,1,-nbitq), 
to_sfixed(-130413331.0/4294967296.0,1,-nbitq), 
to_sfixed(-299564325.0/4294967296.0,1,-nbitq), 
to_sfixed(-289814569.0/4294967296.0,1,-nbitq), 
to_sfixed(-315191602.0/4294967296.0,1,-nbitq), 
to_sfixed(-228423567.0/4294967296.0,1,-nbitq), 
to_sfixed(135471921.0/4294967296.0,1,-nbitq), 
to_sfixed(94276303.0/4294967296.0,1,-nbitq), 
to_sfixed(-158217971.0/4294967296.0,1,-nbitq), 
to_sfixed(-382136856.0/4294967296.0,1,-nbitq), 
to_sfixed(228341411.0/4294967296.0,1,-nbitq), 
to_sfixed(234920669.0/4294967296.0,1,-nbitq), 
to_sfixed(193162999.0/4294967296.0,1,-nbitq), 
to_sfixed(339508273.0/4294967296.0,1,-nbitq), 
to_sfixed(-296354248.0/4294967296.0,1,-nbitq), 
to_sfixed(10459058.0/4294967296.0,1,-nbitq), 
to_sfixed(52569816.0/4294967296.0,1,-nbitq), 
to_sfixed(543843942.0/4294967296.0,1,-nbitq), 
to_sfixed(-23606366.0/4294967296.0,1,-nbitq), 
to_sfixed(14543387.0/4294967296.0,1,-nbitq), 
to_sfixed(71201320.0/4294967296.0,1,-nbitq), 
to_sfixed(17851845.0/4294967296.0,1,-nbitq), 
to_sfixed(-494638335.0/4294967296.0,1,-nbitq), 
to_sfixed(15035409.0/4294967296.0,1,-nbitq), 
to_sfixed(16919708.0/4294967296.0,1,-nbitq), 
to_sfixed(89339614.0/4294967296.0,1,-nbitq), 
to_sfixed(-280598048.0/4294967296.0,1,-nbitq), 
to_sfixed(185213548.0/4294967296.0,1,-nbitq), 
to_sfixed(-83118080.0/4294967296.0,1,-nbitq), 
to_sfixed(-153131159.0/4294967296.0,1,-nbitq), 
to_sfixed(-191508793.0/4294967296.0,1,-nbitq), 
to_sfixed(155433899.0/4294967296.0,1,-nbitq), 
to_sfixed(-240060798.0/4294967296.0,1,-nbitq), 
to_sfixed(-246735587.0/4294967296.0,1,-nbitq), 
to_sfixed(44679375.0/4294967296.0,1,-nbitq), 
to_sfixed(-373486588.0/4294967296.0,1,-nbitq), 
to_sfixed(5741324.0/4294967296.0,1,-nbitq), 
to_sfixed(-91938591.0/4294967296.0,1,-nbitq), 
to_sfixed(-261056527.0/4294967296.0,1,-nbitq), 
to_sfixed(294832547.0/4294967296.0,1,-nbitq), 
to_sfixed(377519789.0/4294967296.0,1,-nbitq), 
to_sfixed(-75207002.0/4294967296.0,1,-nbitq), 
to_sfixed(75771324.0/4294967296.0,1,-nbitq), 
to_sfixed(354408258.0/4294967296.0,1,-nbitq), 
to_sfixed(442865857.0/4294967296.0,1,-nbitq), 
to_sfixed(430460345.0/4294967296.0,1,-nbitq), 
to_sfixed(-266060608.0/4294967296.0,1,-nbitq), 
to_sfixed(122789402.0/4294967296.0,1,-nbitq), 
to_sfixed(-15798643.0/4294967296.0,1,-nbitq), 
to_sfixed(375587160.0/4294967296.0,1,-nbitq), 
to_sfixed(283584375.0/4294967296.0,1,-nbitq), 
to_sfixed(-50677213.0/4294967296.0,1,-nbitq), 
to_sfixed(93603081.0/4294967296.0,1,-nbitq), 
to_sfixed(345224299.0/4294967296.0,1,-nbitq), 
to_sfixed(55285040.0/4294967296.0,1,-nbitq), 
to_sfixed(309900827.0/4294967296.0,1,-nbitq), 
to_sfixed(257908069.0/4294967296.0,1,-nbitq), 
to_sfixed(-308155535.0/4294967296.0,1,-nbitq), 
to_sfixed(-246654436.0/4294967296.0,1,-nbitq), 
to_sfixed(-263822009.0/4294967296.0,1,-nbitq), 
to_sfixed(247252182.0/4294967296.0,1,-nbitq), 
to_sfixed(546155943.0/4294967296.0,1,-nbitq), 
to_sfixed(124509959.0/4294967296.0,1,-nbitq), 
to_sfixed(-174789109.0/4294967296.0,1,-nbitq), 
to_sfixed(-232073598.0/4294967296.0,1,-nbitq), 
to_sfixed(-422705143.0/4294967296.0,1,-nbitq), 
to_sfixed(-184723566.0/4294967296.0,1,-nbitq), 
to_sfixed(-111720188.0/4294967296.0,1,-nbitq), 
to_sfixed(-190694102.0/4294967296.0,1,-nbitq), 
to_sfixed(-137229834.0/4294967296.0,1,-nbitq), 
to_sfixed(-529346615.0/4294967296.0,1,-nbitq), 
to_sfixed(-52846969.0/4294967296.0,1,-nbitq), 
to_sfixed(-479959625.0/4294967296.0,1,-nbitq), 
to_sfixed(-128855814.0/4294967296.0,1,-nbitq), 
to_sfixed(283352459.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(87537418.0/4294967296.0,1,-nbitq), 
to_sfixed(-154569335.0/4294967296.0,1,-nbitq), 
to_sfixed(97921481.0/4294967296.0,1,-nbitq), 
to_sfixed(-427850174.0/4294967296.0,1,-nbitq), 
to_sfixed(485582176.0/4294967296.0,1,-nbitq), 
to_sfixed(268515551.0/4294967296.0,1,-nbitq), 
to_sfixed(-15551058.0/4294967296.0,1,-nbitq), 
to_sfixed(-232039093.0/4294967296.0,1,-nbitq), 
to_sfixed(-170242840.0/4294967296.0,1,-nbitq), 
to_sfixed(438910982.0/4294967296.0,1,-nbitq), 
to_sfixed(221391069.0/4294967296.0,1,-nbitq), 
to_sfixed(-191706602.0/4294967296.0,1,-nbitq), 
to_sfixed(-80463756.0/4294967296.0,1,-nbitq), 
to_sfixed(-207957721.0/4294967296.0,1,-nbitq), 
to_sfixed(267437922.0/4294967296.0,1,-nbitq), 
to_sfixed(199636767.0/4294967296.0,1,-nbitq), 
to_sfixed(53239286.0/4294967296.0,1,-nbitq), 
to_sfixed(381471069.0/4294967296.0,1,-nbitq), 
to_sfixed(-47538472.0/4294967296.0,1,-nbitq), 
to_sfixed(-62001655.0/4294967296.0,1,-nbitq), 
to_sfixed(-127742759.0/4294967296.0,1,-nbitq), 
to_sfixed(8963023.0/4294967296.0,1,-nbitq), 
to_sfixed(526987373.0/4294967296.0,1,-nbitq), 
to_sfixed(153889275.0/4294967296.0,1,-nbitq), 
to_sfixed(142969486.0/4294967296.0,1,-nbitq), 
to_sfixed(485187766.0/4294967296.0,1,-nbitq), 
to_sfixed(-240153019.0/4294967296.0,1,-nbitq), 
to_sfixed(-45137013.0/4294967296.0,1,-nbitq), 
to_sfixed(351680448.0/4294967296.0,1,-nbitq), 
to_sfixed(-202195457.0/4294967296.0,1,-nbitq), 
to_sfixed(-443370725.0/4294967296.0,1,-nbitq), 
to_sfixed(-32603119.0/4294967296.0,1,-nbitq), 
to_sfixed(244900225.0/4294967296.0,1,-nbitq), 
to_sfixed(17674776.0/4294967296.0,1,-nbitq), 
to_sfixed(138900434.0/4294967296.0,1,-nbitq), 
to_sfixed(-5242981.0/4294967296.0,1,-nbitq), 
to_sfixed(235769137.0/4294967296.0,1,-nbitq), 
to_sfixed(37788360.0/4294967296.0,1,-nbitq), 
to_sfixed(18942894.0/4294967296.0,1,-nbitq), 
to_sfixed(119797495.0/4294967296.0,1,-nbitq), 
to_sfixed(-371026135.0/4294967296.0,1,-nbitq), 
to_sfixed(-204867.0/4294967296.0,1,-nbitq), 
to_sfixed(-192664752.0/4294967296.0,1,-nbitq), 
to_sfixed(-217069935.0/4294967296.0,1,-nbitq), 
to_sfixed(384078153.0/4294967296.0,1,-nbitq), 
to_sfixed(399070522.0/4294967296.0,1,-nbitq), 
to_sfixed(-3746296.0/4294967296.0,1,-nbitq), 
to_sfixed(-339382271.0/4294967296.0,1,-nbitq), 
to_sfixed(-121481697.0/4294967296.0,1,-nbitq), 
to_sfixed(367452940.0/4294967296.0,1,-nbitq), 
to_sfixed(297082185.0/4294967296.0,1,-nbitq), 
to_sfixed(107177372.0/4294967296.0,1,-nbitq), 
to_sfixed(-300681397.0/4294967296.0,1,-nbitq), 
to_sfixed(-166169352.0/4294967296.0,1,-nbitq), 
to_sfixed(381686542.0/4294967296.0,1,-nbitq), 
to_sfixed(-305125834.0/4294967296.0,1,-nbitq), 
to_sfixed(306450039.0/4294967296.0,1,-nbitq), 
to_sfixed(-20894393.0/4294967296.0,1,-nbitq), 
to_sfixed(219905282.0/4294967296.0,1,-nbitq), 
to_sfixed(240655076.0/4294967296.0,1,-nbitq), 
to_sfixed(222005214.0/4294967296.0,1,-nbitq), 
to_sfixed(505384737.0/4294967296.0,1,-nbitq), 
to_sfixed(86202273.0/4294967296.0,1,-nbitq), 
to_sfixed(119730582.0/4294967296.0,1,-nbitq), 
to_sfixed(295191897.0/4294967296.0,1,-nbitq), 
to_sfixed(31175171.0/4294967296.0,1,-nbitq), 
to_sfixed(788819119.0/4294967296.0,1,-nbitq), 
to_sfixed(-241273650.0/4294967296.0,1,-nbitq), 
to_sfixed(-295254292.0/4294967296.0,1,-nbitq), 
to_sfixed(382105791.0/4294967296.0,1,-nbitq), 
to_sfixed(-30294171.0/4294967296.0,1,-nbitq), 
to_sfixed(50641957.0/4294967296.0,1,-nbitq), 
to_sfixed(138132484.0/4294967296.0,1,-nbitq), 
to_sfixed(60281797.0/4294967296.0,1,-nbitq), 
to_sfixed(489270441.0/4294967296.0,1,-nbitq), 
to_sfixed(728528.0/4294967296.0,1,-nbitq), 
to_sfixed(37675495.0/4294967296.0,1,-nbitq), 
to_sfixed(-152763661.0/4294967296.0,1,-nbitq), 
to_sfixed(-227890875.0/4294967296.0,1,-nbitq), 
to_sfixed(-2681938.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-164636443.0/4294967296.0,1,-nbitq), 
to_sfixed(201382703.0/4294967296.0,1,-nbitq), 
to_sfixed(-261855114.0/4294967296.0,1,-nbitq), 
to_sfixed(189920106.0/4294967296.0,1,-nbitq), 
to_sfixed(397293400.0/4294967296.0,1,-nbitq), 
to_sfixed(267710792.0/4294967296.0,1,-nbitq), 
to_sfixed(47523787.0/4294967296.0,1,-nbitq), 
to_sfixed(-155971076.0/4294967296.0,1,-nbitq), 
to_sfixed(200160141.0/4294967296.0,1,-nbitq), 
to_sfixed(-129564218.0/4294967296.0,1,-nbitq), 
to_sfixed(297522016.0/4294967296.0,1,-nbitq), 
to_sfixed(-140879170.0/4294967296.0,1,-nbitq), 
to_sfixed(-276286510.0/4294967296.0,1,-nbitq), 
to_sfixed(-160091670.0/4294967296.0,1,-nbitq), 
to_sfixed(-140062339.0/4294967296.0,1,-nbitq), 
to_sfixed(-407031791.0/4294967296.0,1,-nbitq), 
to_sfixed(194903023.0/4294967296.0,1,-nbitq), 
to_sfixed(139483413.0/4294967296.0,1,-nbitq), 
to_sfixed(-193900262.0/4294967296.0,1,-nbitq), 
to_sfixed(-4923166.0/4294967296.0,1,-nbitq), 
to_sfixed(-404220841.0/4294967296.0,1,-nbitq), 
to_sfixed(110054824.0/4294967296.0,1,-nbitq), 
to_sfixed(254489791.0/4294967296.0,1,-nbitq), 
to_sfixed(159572025.0/4294967296.0,1,-nbitq), 
to_sfixed(135950004.0/4294967296.0,1,-nbitq), 
to_sfixed(126866603.0/4294967296.0,1,-nbitq), 
to_sfixed(361742916.0/4294967296.0,1,-nbitq), 
to_sfixed(-73148246.0/4294967296.0,1,-nbitq), 
to_sfixed(269350542.0/4294967296.0,1,-nbitq), 
to_sfixed(62690482.0/4294967296.0,1,-nbitq), 
to_sfixed(-550747450.0/4294967296.0,1,-nbitq), 
to_sfixed(63752777.0/4294967296.0,1,-nbitq), 
to_sfixed(292577242.0/4294967296.0,1,-nbitq), 
to_sfixed(71387646.0/4294967296.0,1,-nbitq), 
to_sfixed(387885527.0/4294967296.0,1,-nbitq), 
to_sfixed(-230475104.0/4294967296.0,1,-nbitq), 
to_sfixed(-158918681.0/4294967296.0,1,-nbitq), 
to_sfixed(-101049621.0/4294967296.0,1,-nbitq), 
to_sfixed(-78793634.0/4294967296.0,1,-nbitq), 
to_sfixed(-55161983.0/4294967296.0,1,-nbitq), 
to_sfixed(87961418.0/4294967296.0,1,-nbitq), 
to_sfixed(83211950.0/4294967296.0,1,-nbitq), 
to_sfixed(173660687.0/4294967296.0,1,-nbitq), 
to_sfixed(238496151.0/4294967296.0,1,-nbitq), 
to_sfixed(22576796.0/4294967296.0,1,-nbitq), 
to_sfixed(385324510.0/4294967296.0,1,-nbitq), 
to_sfixed(310833929.0/4294967296.0,1,-nbitq), 
to_sfixed(226256631.0/4294967296.0,1,-nbitq), 
to_sfixed(-126650281.0/4294967296.0,1,-nbitq), 
to_sfixed(229264415.0/4294967296.0,1,-nbitq), 
to_sfixed(-285738957.0/4294967296.0,1,-nbitq), 
to_sfixed(274961825.0/4294967296.0,1,-nbitq), 
to_sfixed(-532300130.0/4294967296.0,1,-nbitq), 
to_sfixed(356300257.0/4294967296.0,1,-nbitq), 
to_sfixed(-104806032.0/4294967296.0,1,-nbitq), 
to_sfixed(194315239.0/4294967296.0,1,-nbitq), 
to_sfixed(358409138.0/4294967296.0,1,-nbitq), 
to_sfixed(-296157499.0/4294967296.0,1,-nbitq), 
to_sfixed(264401838.0/4294967296.0,1,-nbitq), 
to_sfixed(376098047.0/4294967296.0,1,-nbitq), 
to_sfixed(-278733928.0/4294967296.0,1,-nbitq), 
to_sfixed(409330237.0/4294967296.0,1,-nbitq), 
to_sfixed(207048638.0/4294967296.0,1,-nbitq), 
to_sfixed(152887780.0/4294967296.0,1,-nbitq), 
to_sfixed(-190424479.0/4294967296.0,1,-nbitq), 
to_sfixed(-29480392.0/4294967296.0,1,-nbitq), 
to_sfixed(520616587.0/4294967296.0,1,-nbitq), 
to_sfixed(-126653590.0/4294967296.0,1,-nbitq), 
to_sfixed(219729523.0/4294967296.0,1,-nbitq), 
to_sfixed(512554813.0/4294967296.0,1,-nbitq), 
to_sfixed(75288360.0/4294967296.0,1,-nbitq), 
to_sfixed(-83456766.0/4294967296.0,1,-nbitq), 
to_sfixed(-173967495.0/4294967296.0,1,-nbitq), 
to_sfixed(402367313.0/4294967296.0,1,-nbitq), 
to_sfixed(-178049016.0/4294967296.0,1,-nbitq), 
to_sfixed(-149586147.0/4294967296.0,1,-nbitq), 
to_sfixed(-390829251.0/4294967296.0,1,-nbitq), 
to_sfixed(-264417689.0/4294967296.0,1,-nbitq), 
to_sfixed(-94524816.0/4294967296.0,1,-nbitq), 
to_sfixed(-139522569.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(174933139.0/4294967296.0,1,-nbitq), 
to_sfixed(-209974042.0/4294967296.0,1,-nbitq), 
to_sfixed(468928074.0/4294967296.0,1,-nbitq), 
to_sfixed(-150523472.0/4294967296.0,1,-nbitq), 
to_sfixed(-85180712.0/4294967296.0,1,-nbitq), 
to_sfixed(-197041007.0/4294967296.0,1,-nbitq), 
to_sfixed(-123319031.0/4294967296.0,1,-nbitq), 
to_sfixed(197215586.0/4294967296.0,1,-nbitq), 
to_sfixed(275713861.0/4294967296.0,1,-nbitq), 
to_sfixed(25579754.0/4294967296.0,1,-nbitq), 
to_sfixed(396883382.0/4294967296.0,1,-nbitq), 
to_sfixed(452303067.0/4294967296.0,1,-nbitq), 
to_sfixed(26033717.0/4294967296.0,1,-nbitq), 
to_sfixed(337611634.0/4294967296.0,1,-nbitq), 
to_sfixed(-277891278.0/4294967296.0,1,-nbitq), 
to_sfixed(-23773714.0/4294967296.0,1,-nbitq), 
to_sfixed(-338566273.0/4294967296.0,1,-nbitq), 
to_sfixed(-341358441.0/4294967296.0,1,-nbitq), 
to_sfixed(-305176782.0/4294967296.0,1,-nbitq), 
to_sfixed(115411211.0/4294967296.0,1,-nbitq), 
to_sfixed(276329058.0/4294967296.0,1,-nbitq), 
to_sfixed(511493021.0/4294967296.0,1,-nbitq), 
to_sfixed(-85464004.0/4294967296.0,1,-nbitq), 
to_sfixed(-122419768.0/4294967296.0,1,-nbitq), 
to_sfixed(-281352570.0/4294967296.0,1,-nbitq), 
to_sfixed(119930631.0/4294967296.0,1,-nbitq), 
to_sfixed(254552367.0/4294967296.0,1,-nbitq), 
to_sfixed(-288298793.0/4294967296.0,1,-nbitq), 
to_sfixed(-175586930.0/4294967296.0,1,-nbitq), 
to_sfixed(-245717575.0/4294967296.0,1,-nbitq), 
to_sfixed(-99183268.0/4294967296.0,1,-nbitq), 
to_sfixed(-525384073.0/4294967296.0,1,-nbitq), 
to_sfixed(166606139.0/4294967296.0,1,-nbitq), 
to_sfixed(244123228.0/4294967296.0,1,-nbitq), 
to_sfixed(515283595.0/4294967296.0,1,-nbitq), 
to_sfixed(11642180.0/4294967296.0,1,-nbitq), 
to_sfixed(170775479.0/4294967296.0,1,-nbitq), 
to_sfixed(495211303.0/4294967296.0,1,-nbitq), 
to_sfixed(-174150245.0/4294967296.0,1,-nbitq), 
to_sfixed(56410533.0/4294967296.0,1,-nbitq), 
to_sfixed(-388130062.0/4294967296.0,1,-nbitq), 
to_sfixed(468911276.0/4294967296.0,1,-nbitq), 
to_sfixed(-315943411.0/4294967296.0,1,-nbitq), 
to_sfixed(240164002.0/4294967296.0,1,-nbitq), 
to_sfixed(-259410527.0/4294967296.0,1,-nbitq), 
to_sfixed(41430042.0/4294967296.0,1,-nbitq), 
to_sfixed(170860525.0/4294967296.0,1,-nbitq), 
to_sfixed(-208960897.0/4294967296.0,1,-nbitq), 
to_sfixed(-293188699.0/4294967296.0,1,-nbitq), 
to_sfixed(355042483.0/4294967296.0,1,-nbitq), 
to_sfixed(-103397255.0/4294967296.0,1,-nbitq), 
to_sfixed(-242651305.0/4294967296.0,1,-nbitq), 
to_sfixed(-556530851.0/4294967296.0,1,-nbitq), 
to_sfixed(-13728864.0/4294967296.0,1,-nbitq), 
to_sfixed(-136361336.0/4294967296.0,1,-nbitq), 
to_sfixed(-287426124.0/4294967296.0,1,-nbitq), 
to_sfixed(233595165.0/4294967296.0,1,-nbitq), 
to_sfixed(-426968534.0/4294967296.0,1,-nbitq), 
to_sfixed(387758809.0/4294967296.0,1,-nbitq), 
to_sfixed(-73065122.0/4294967296.0,1,-nbitq), 
to_sfixed(-422456468.0/4294967296.0,1,-nbitq), 
to_sfixed(524557386.0/4294967296.0,1,-nbitq), 
to_sfixed(-397785142.0/4294967296.0,1,-nbitq), 
to_sfixed(-200053348.0/4294967296.0,1,-nbitq), 
to_sfixed(29770577.0/4294967296.0,1,-nbitq), 
to_sfixed(-385735966.0/4294967296.0,1,-nbitq), 
to_sfixed(332631489.0/4294967296.0,1,-nbitq), 
to_sfixed(216244893.0/4294967296.0,1,-nbitq), 
to_sfixed(332700466.0/4294967296.0,1,-nbitq), 
to_sfixed(552693824.0/4294967296.0,1,-nbitq), 
to_sfixed(-32124639.0/4294967296.0,1,-nbitq), 
to_sfixed(-158348735.0/4294967296.0,1,-nbitq), 
to_sfixed(70310076.0/4294967296.0,1,-nbitq), 
to_sfixed(14747289.0/4294967296.0,1,-nbitq), 
to_sfixed(448530534.0/4294967296.0,1,-nbitq), 
to_sfixed(-395735976.0/4294967296.0,1,-nbitq), 
to_sfixed(321576333.0/4294967296.0,1,-nbitq), 
to_sfixed(73098598.0/4294967296.0,1,-nbitq), 
to_sfixed(-144595933.0/4294967296.0,1,-nbitq), 
to_sfixed(-270155580.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-128782811.0/4294967296.0,1,-nbitq), 
to_sfixed(-15051674.0/4294967296.0,1,-nbitq), 
to_sfixed(357697047.0/4294967296.0,1,-nbitq), 
to_sfixed(-407466703.0/4294967296.0,1,-nbitq), 
to_sfixed(348510411.0/4294967296.0,1,-nbitq), 
to_sfixed(-411171274.0/4294967296.0,1,-nbitq), 
to_sfixed(-161134304.0/4294967296.0,1,-nbitq), 
to_sfixed(-230546266.0/4294967296.0,1,-nbitq), 
to_sfixed(218164086.0/4294967296.0,1,-nbitq), 
to_sfixed(-214289340.0/4294967296.0,1,-nbitq), 
to_sfixed(-47345834.0/4294967296.0,1,-nbitq), 
to_sfixed(329069645.0/4294967296.0,1,-nbitq), 
to_sfixed(-173814221.0/4294967296.0,1,-nbitq), 
to_sfixed(-93380853.0/4294967296.0,1,-nbitq), 
to_sfixed(-200352055.0/4294967296.0,1,-nbitq), 
to_sfixed(-35627490.0/4294967296.0,1,-nbitq), 
to_sfixed(-287752115.0/4294967296.0,1,-nbitq), 
to_sfixed(197274912.0/4294967296.0,1,-nbitq), 
to_sfixed(107362659.0/4294967296.0,1,-nbitq), 
to_sfixed(216012392.0/4294967296.0,1,-nbitq), 
to_sfixed(-80079231.0/4294967296.0,1,-nbitq), 
to_sfixed(-38003908.0/4294967296.0,1,-nbitq), 
to_sfixed(102952081.0/4294967296.0,1,-nbitq), 
to_sfixed(-4719752.0/4294967296.0,1,-nbitq), 
to_sfixed(-83983099.0/4294967296.0,1,-nbitq), 
to_sfixed(289171310.0/4294967296.0,1,-nbitq), 
to_sfixed(167146153.0/4294967296.0,1,-nbitq), 
to_sfixed(-243430382.0/4294967296.0,1,-nbitq), 
to_sfixed(272361059.0/4294967296.0,1,-nbitq), 
to_sfixed(530627325.0/4294967296.0,1,-nbitq), 
to_sfixed(126618278.0/4294967296.0,1,-nbitq), 
to_sfixed(-239859537.0/4294967296.0,1,-nbitq), 
to_sfixed(-131907873.0/4294967296.0,1,-nbitq), 
to_sfixed(91708585.0/4294967296.0,1,-nbitq), 
to_sfixed(493896215.0/4294967296.0,1,-nbitq), 
to_sfixed(131543494.0/4294967296.0,1,-nbitq), 
to_sfixed(379104315.0/4294967296.0,1,-nbitq), 
to_sfixed(220794184.0/4294967296.0,1,-nbitq), 
to_sfixed(-68120497.0/4294967296.0,1,-nbitq), 
to_sfixed(-46963365.0/4294967296.0,1,-nbitq), 
to_sfixed(-323932380.0/4294967296.0,1,-nbitq), 
to_sfixed(181098807.0/4294967296.0,1,-nbitq), 
to_sfixed(86933489.0/4294967296.0,1,-nbitq), 
to_sfixed(-278241213.0/4294967296.0,1,-nbitq), 
to_sfixed(372513573.0/4294967296.0,1,-nbitq), 
to_sfixed(312099052.0/4294967296.0,1,-nbitq), 
to_sfixed(-79430979.0/4294967296.0,1,-nbitq), 
to_sfixed(-62267007.0/4294967296.0,1,-nbitq), 
to_sfixed(-140481840.0/4294967296.0,1,-nbitq), 
to_sfixed(344844362.0/4294967296.0,1,-nbitq), 
to_sfixed(107752317.0/4294967296.0,1,-nbitq), 
to_sfixed(438399107.0/4294967296.0,1,-nbitq), 
to_sfixed(-719258582.0/4294967296.0,1,-nbitq), 
to_sfixed(-32546483.0/4294967296.0,1,-nbitq), 
to_sfixed(455629599.0/4294967296.0,1,-nbitq), 
to_sfixed(74678465.0/4294967296.0,1,-nbitq), 
to_sfixed(-312200074.0/4294967296.0,1,-nbitq), 
to_sfixed(-67037396.0/4294967296.0,1,-nbitq), 
to_sfixed(220143914.0/4294967296.0,1,-nbitq), 
to_sfixed(-192793206.0/4294967296.0,1,-nbitq), 
to_sfixed(-363229021.0/4294967296.0,1,-nbitq), 
to_sfixed(398401949.0/4294967296.0,1,-nbitq), 
to_sfixed(-514394059.0/4294967296.0,1,-nbitq), 
to_sfixed(-258886033.0/4294967296.0,1,-nbitq), 
to_sfixed(251822085.0/4294967296.0,1,-nbitq), 
to_sfixed(-407124878.0/4294967296.0,1,-nbitq), 
to_sfixed(168703417.0/4294967296.0,1,-nbitq), 
to_sfixed(162397407.0/4294967296.0,1,-nbitq), 
to_sfixed(-53834503.0/4294967296.0,1,-nbitq), 
to_sfixed(25448620.0/4294967296.0,1,-nbitq), 
to_sfixed(411556022.0/4294967296.0,1,-nbitq), 
to_sfixed(12733827.0/4294967296.0,1,-nbitq), 
to_sfixed(-183485767.0/4294967296.0,1,-nbitq), 
to_sfixed(432762062.0/4294967296.0,1,-nbitq), 
to_sfixed(81900964.0/4294967296.0,1,-nbitq), 
to_sfixed(267701357.0/4294967296.0,1,-nbitq), 
to_sfixed(-258204987.0/4294967296.0,1,-nbitq), 
to_sfixed(-47636667.0/4294967296.0,1,-nbitq), 
to_sfixed(-77970979.0/4294967296.0,1,-nbitq), 
to_sfixed(235789249.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(318197733.0/4294967296.0,1,-nbitq), 
to_sfixed(-691182262.0/4294967296.0,1,-nbitq), 
to_sfixed(147140302.0/4294967296.0,1,-nbitq), 
to_sfixed(260606337.0/4294967296.0,1,-nbitq), 
to_sfixed(548176431.0/4294967296.0,1,-nbitq), 
to_sfixed(-253607756.0/4294967296.0,1,-nbitq), 
to_sfixed(465589499.0/4294967296.0,1,-nbitq), 
to_sfixed(-369653090.0/4294967296.0,1,-nbitq), 
to_sfixed(213546857.0/4294967296.0,1,-nbitq), 
to_sfixed(-337421713.0/4294967296.0,1,-nbitq), 
to_sfixed(100043014.0/4294967296.0,1,-nbitq), 
to_sfixed(201118907.0/4294967296.0,1,-nbitq), 
to_sfixed(-397240478.0/4294967296.0,1,-nbitq), 
to_sfixed(-325008707.0/4294967296.0,1,-nbitq), 
to_sfixed(-144723069.0/4294967296.0,1,-nbitq), 
to_sfixed(-280640175.0/4294967296.0,1,-nbitq), 
to_sfixed(-147501672.0/4294967296.0,1,-nbitq), 
to_sfixed(171472354.0/4294967296.0,1,-nbitq), 
to_sfixed(-447484850.0/4294967296.0,1,-nbitq), 
to_sfixed(-341711306.0/4294967296.0,1,-nbitq), 
to_sfixed(-190630655.0/4294967296.0,1,-nbitq), 
to_sfixed(442535644.0/4294967296.0,1,-nbitq), 
to_sfixed(352180792.0/4294967296.0,1,-nbitq), 
to_sfixed(-131702294.0/4294967296.0,1,-nbitq), 
to_sfixed(268528636.0/4294967296.0,1,-nbitq), 
to_sfixed(-125133704.0/4294967296.0,1,-nbitq), 
to_sfixed(153784823.0/4294967296.0,1,-nbitq), 
to_sfixed(113208954.0/4294967296.0,1,-nbitq), 
to_sfixed(107110421.0/4294967296.0,1,-nbitq), 
to_sfixed(-43353346.0/4294967296.0,1,-nbitq), 
to_sfixed(81343005.0/4294967296.0,1,-nbitq), 
to_sfixed(-224419197.0/4294967296.0,1,-nbitq), 
to_sfixed(339734507.0/4294967296.0,1,-nbitq), 
to_sfixed(-266104537.0/4294967296.0,1,-nbitq), 
to_sfixed(9995603.0/4294967296.0,1,-nbitq), 
to_sfixed(130166292.0/4294967296.0,1,-nbitq), 
to_sfixed(510149455.0/4294967296.0,1,-nbitq), 
to_sfixed(286489481.0/4294967296.0,1,-nbitq), 
to_sfixed(232721690.0/4294967296.0,1,-nbitq), 
to_sfixed(233222474.0/4294967296.0,1,-nbitq), 
to_sfixed(-119659739.0/4294967296.0,1,-nbitq), 
to_sfixed(471268655.0/4294967296.0,1,-nbitq), 
to_sfixed(403405795.0/4294967296.0,1,-nbitq), 
to_sfixed(172681995.0/4294967296.0,1,-nbitq), 
to_sfixed(-273472217.0/4294967296.0,1,-nbitq), 
to_sfixed(479292280.0/4294967296.0,1,-nbitq), 
to_sfixed(-393529198.0/4294967296.0,1,-nbitq), 
to_sfixed(-317257387.0/4294967296.0,1,-nbitq), 
to_sfixed(67050730.0/4294967296.0,1,-nbitq), 
to_sfixed(-48077725.0/4294967296.0,1,-nbitq), 
to_sfixed(259071157.0/4294967296.0,1,-nbitq), 
to_sfixed(25922512.0/4294967296.0,1,-nbitq), 
to_sfixed(-236472751.0/4294967296.0,1,-nbitq), 
to_sfixed(284804391.0/4294967296.0,1,-nbitq), 
to_sfixed(369497929.0/4294967296.0,1,-nbitq), 
to_sfixed(-9700599.0/4294967296.0,1,-nbitq), 
to_sfixed(120911797.0/4294967296.0,1,-nbitq), 
to_sfixed(127512898.0/4294967296.0,1,-nbitq), 
to_sfixed(-271535625.0/4294967296.0,1,-nbitq), 
to_sfixed(-189685410.0/4294967296.0,1,-nbitq), 
to_sfixed(-49742203.0/4294967296.0,1,-nbitq), 
to_sfixed(139796502.0/4294967296.0,1,-nbitq), 
to_sfixed(-406067452.0/4294967296.0,1,-nbitq), 
to_sfixed(409220552.0/4294967296.0,1,-nbitq), 
to_sfixed(18451857.0/4294967296.0,1,-nbitq), 
to_sfixed(262507303.0/4294967296.0,1,-nbitq), 
to_sfixed(-255221958.0/4294967296.0,1,-nbitq), 
to_sfixed(-332654738.0/4294967296.0,1,-nbitq), 
to_sfixed(44124872.0/4294967296.0,1,-nbitq), 
to_sfixed(-263028351.0/4294967296.0,1,-nbitq), 
to_sfixed(-137325558.0/4294967296.0,1,-nbitq), 
to_sfixed(-329535640.0/4294967296.0,1,-nbitq), 
to_sfixed(41633204.0/4294967296.0,1,-nbitq), 
to_sfixed(195751089.0/4294967296.0,1,-nbitq), 
to_sfixed(-77939095.0/4294967296.0,1,-nbitq), 
to_sfixed(-168403849.0/4294967296.0,1,-nbitq), 
to_sfixed(329267996.0/4294967296.0,1,-nbitq), 
to_sfixed(-169618344.0/4294967296.0,1,-nbitq), 
to_sfixed(-495837079.0/4294967296.0,1,-nbitq), 
to_sfixed(-310191835.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(39905003.0/4294967296.0,1,-nbitq), 
to_sfixed(-117813869.0/4294967296.0,1,-nbitq), 
to_sfixed(507662480.0/4294967296.0,1,-nbitq), 
to_sfixed(33147668.0/4294967296.0,1,-nbitq), 
to_sfixed(284023414.0/4294967296.0,1,-nbitq), 
to_sfixed(493253360.0/4294967296.0,1,-nbitq), 
to_sfixed(358720317.0/4294967296.0,1,-nbitq), 
to_sfixed(428057290.0/4294967296.0,1,-nbitq), 
to_sfixed(442335488.0/4294967296.0,1,-nbitq), 
to_sfixed(-275217726.0/4294967296.0,1,-nbitq), 
to_sfixed(177922208.0/4294967296.0,1,-nbitq), 
to_sfixed(671162755.0/4294967296.0,1,-nbitq), 
to_sfixed(-232730894.0/4294967296.0,1,-nbitq), 
to_sfixed(-297894499.0/4294967296.0,1,-nbitq), 
to_sfixed(-211973869.0/4294967296.0,1,-nbitq), 
to_sfixed(-224569700.0/4294967296.0,1,-nbitq), 
to_sfixed(32646496.0/4294967296.0,1,-nbitq), 
to_sfixed(-112604953.0/4294967296.0,1,-nbitq), 
to_sfixed(-292132267.0/4294967296.0,1,-nbitq), 
to_sfixed(157245934.0/4294967296.0,1,-nbitq), 
to_sfixed(-59898165.0/4294967296.0,1,-nbitq), 
to_sfixed(472494514.0/4294967296.0,1,-nbitq), 
to_sfixed(395544813.0/4294967296.0,1,-nbitq), 
to_sfixed(162649340.0/4294967296.0,1,-nbitq), 
to_sfixed(-328126608.0/4294967296.0,1,-nbitq), 
to_sfixed(-271106152.0/4294967296.0,1,-nbitq), 
to_sfixed(196521959.0/4294967296.0,1,-nbitq), 
to_sfixed(-328704639.0/4294967296.0,1,-nbitq), 
to_sfixed(-600311252.0/4294967296.0,1,-nbitq), 
to_sfixed(-116531606.0/4294967296.0,1,-nbitq), 
to_sfixed(-414964548.0/4294967296.0,1,-nbitq), 
to_sfixed(-829265399.0/4294967296.0,1,-nbitq), 
to_sfixed(-153986094.0/4294967296.0,1,-nbitq), 
to_sfixed(382374545.0/4294967296.0,1,-nbitq), 
to_sfixed(-265545062.0/4294967296.0,1,-nbitq), 
to_sfixed(-412644819.0/4294967296.0,1,-nbitq), 
to_sfixed(94072496.0/4294967296.0,1,-nbitq), 
to_sfixed(160996784.0/4294967296.0,1,-nbitq), 
to_sfixed(-207032764.0/4294967296.0,1,-nbitq), 
to_sfixed(176724867.0/4294967296.0,1,-nbitq), 
to_sfixed(-263213443.0/4294967296.0,1,-nbitq), 
to_sfixed(-35329752.0/4294967296.0,1,-nbitq), 
to_sfixed(-89783798.0/4294967296.0,1,-nbitq), 
to_sfixed(127446375.0/4294967296.0,1,-nbitq), 
to_sfixed(150488279.0/4294967296.0,1,-nbitq), 
to_sfixed(540058551.0/4294967296.0,1,-nbitq), 
to_sfixed(295854628.0/4294967296.0,1,-nbitq), 
to_sfixed(-366943934.0/4294967296.0,1,-nbitq), 
to_sfixed(101995816.0/4294967296.0,1,-nbitq), 
to_sfixed(683349589.0/4294967296.0,1,-nbitq), 
to_sfixed(-21417695.0/4294967296.0,1,-nbitq), 
to_sfixed(-130846132.0/4294967296.0,1,-nbitq), 
to_sfixed(-728581623.0/4294967296.0,1,-nbitq), 
to_sfixed(-51572063.0/4294967296.0,1,-nbitq), 
to_sfixed(114069149.0/4294967296.0,1,-nbitq), 
to_sfixed(135548726.0/4294967296.0,1,-nbitq), 
to_sfixed(136900230.0/4294967296.0,1,-nbitq), 
to_sfixed(-311996204.0/4294967296.0,1,-nbitq), 
to_sfixed(291410911.0/4294967296.0,1,-nbitq), 
to_sfixed(333813236.0/4294967296.0,1,-nbitq), 
to_sfixed(-161281538.0/4294967296.0,1,-nbitq), 
to_sfixed(-149276389.0/4294967296.0,1,-nbitq), 
to_sfixed(-626230502.0/4294967296.0,1,-nbitq), 
to_sfixed(311644663.0/4294967296.0,1,-nbitq), 
to_sfixed(-119478196.0/4294967296.0,1,-nbitq), 
to_sfixed(-449770359.0/4294967296.0,1,-nbitq), 
to_sfixed(61144935.0/4294967296.0,1,-nbitq), 
to_sfixed(-133179634.0/4294967296.0,1,-nbitq), 
to_sfixed(13115127.0/4294967296.0,1,-nbitq), 
to_sfixed(-23988142.0/4294967296.0,1,-nbitq), 
to_sfixed(510553899.0/4294967296.0,1,-nbitq), 
to_sfixed(-315366295.0/4294967296.0,1,-nbitq), 
to_sfixed(464419950.0/4294967296.0,1,-nbitq), 
to_sfixed(-212608453.0/4294967296.0,1,-nbitq), 
to_sfixed(-260904485.0/4294967296.0,1,-nbitq), 
to_sfixed(268712589.0/4294967296.0,1,-nbitq), 
to_sfixed(532680974.0/4294967296.0,1,-nbitq), 
to_sfixed(501332941.0/4294967296.0,1,-nbitq), 
to_sfixed(-586159247.0/4294967296.0,1,-nbitq), 
to_sfixed(-197490361.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(64905894.0/4294967296.0,1,-nbitq), 
to_sfixed(-588976502.0/4294967296.0,1,-nbitq), 
to_sfixed(135783019.0/4294967296.0,1,-nbitq), 
to_sfixed(-28188516.0/4294967296.0,1,-nbitq), 
to_sfixed(469029422.0/4294967296.0,1,-nbitq), 
to_sfixed(317317925.0/4294967296.0,1,-nbitq), 
to_sfixed(-328608588.0/4294967296.0,1,-nbitq), 
to_sfixed(-363382061.0/4294967296.0,1,-nbitq), 
to_sfixed(320372393.0/4294967296.0,1,-nbitq), 
to_sfixed(388244295.0/4294967296.0,1,-nbitq), 
to_sfixed(481481752.0/4294967296.0,1,-nbitq), 
to_sfixed(344644272.0/4294967296.0,1,-nbitq), 
to_sfixed(-58514739.0/4294967296.0,1,-nbitq), 
to_sfixed(-302592308.0/4294967296.0,1,-nbitq), 
to_sfixed(331101659.0/4294967296.0,1,-nbitq), 
to_sfixed(318485298.0/4294967296.0,1,-nbitq), 
to_sfixed(312790392.0/4294967296.0,1,-nbitq), 
to_sfixed(-299510189.0/4294967296.0,1,-nbitq), 
to_sfixed(-302487598.0/4294967296.0,1,-nbitq), 
to_sfixed(-20341186.0/4294967296.0,1,-nbitq), 
to_sfixed(-122815222.0/4294967296.0,1,-nbitq), 
to_sfixed(-254070948.0/4294967296.0,1,-nbitq), 
to_sfixed(411799142.0/4294967296.0,1,-nbitq), 
to_sfixed(-548987611.0/4294967296.0,1,-nbitq), 
to_sfixed(90717303.0/4294967296.0,1,-nbitq), 
to_sfixed(-583789964.0/4294967296.0,1,-nbitq), 
to_sfixed(-175694958.0/4294967296.0,1,-nbitq), 
to_sfixed(234339756.0/4294967296.0,1,-nbitq), 
to_sfixed(-182147126.0/4294967296.0,1,-nbitq), 
to_sfixed(-251262987.0/4294967296.0,1,-nbitq), 
to_sfixed(-131595215.0/4294967296.0,1,-nbitq), 
to_sfixed(-116062788.0/4294967296.0,1,-nbitq), 
to_sfixed(78643773.0/4294967296.0,1,-nbitq), 
to_sfixed(528989947.0/4294967296.0,1,-nbitq), 
to_sfixed(-423987486.0/4294967296.0,1,-nbitq), 
to_sfixed(-386762535.0/4294967296.0,1,-nbitq), 
to_sfixed(-75947149.0/4294967296.0,1,-nbitq), 
to_sfixed(-154014241.0/4294967296.0,1,-nbitq), 
to_sfixed(-318425049.0/4294967296.0,1,-nbitq), 
to_sfixed(146875650.0/4294967296.0,1,-nbitq), 
to_sfixed(296553352.0/4294967296.0,1,-nbitq), 
to_sfixed(96799259.0/4294967296.0,1,-nbitq), 
to_sfixed(-251957221.0/4294967296.0,1,-nbitq), 
to_sfixed(73481129.0/4294967296.0,1,-nbitq), 
to_sfixed(156705168.0/4294967296.0,1,-nbitq), 
to_sfixed(131646023.0/4294967296.0,1,-nbitq), 
to_sfixed(-422384040.0/4294967296.0,1,-nbitq), 
to_sfixed(430176908.0/4294967296.0,1,-nbitq), 
to_sfixed(148204259.0/4294967296.0,1,-nbitq), 
to_sfixed(-56451936.0/4294967296.0,1,-nbitq), 
to_sfixed(-104909710.0/4294967296.0,1,-nbitq), 
to_sfixed(-62466525.0/4294967296.0,1,-nbitq), 
to_sfixed(-449383696.0/4294967296.0,1,-nbitq), 
to_sfixed(-85935745.0/4294967296.0,1,-nbitq), 
to_sfixed(-525206323.0/4294967296.0,1,-nbitq), 
to_sfixed(654053021.0/4294967296.0,1,-nbitq), 
to_sfixed(149541608.0/4294967296.0,1,-nbitq), 
to_sfixed(-239412932.0/4294967296.0,1,-nbitq), 
to_sfixed(-366507382.0/4294967296.0,1,-nbitq), 
to_sfixed(67540671.0/4294967296.0,1,-nbitq), 
to_sfixed(281801919.0/4294967296.0,1,-nbitq), 
to_sfixed(-54928412.0/4294967296.0,1,-nbitq), 
to_sfixed(-453285191.0/4294967296.0,1,-nbitq), 
to_sfixed(-86670216.0/4294967296.0,1,-nbitq), 
to_sfixed(-406206530.0/4294967296.0,1,-nbitq), 
to_sfixed(122070794.0/4294967296.0,1,-nbitq), 
to_sfixed(91206694.0/4294967296.0,1,-nbitq), 
to_sfixed(-240955275.0/4294967296.0,1,-nbitq), 
to_sfixed(339787324.0/4294967296.0,1,-nbitq), 
to_sfixed(487811210.0/4294967296.0,1,-nbitq), 
to_sfixed(77461253.0/4294967296.0,1,-nbitq), 
to_sfixed(-264745241.0/4294967296.0,1,-nbitq), 
to_sfixed(177776635.0/4294967296.0,1,-nbitq), 
to_sfixed(-256743400.0/4294967296.0,1,-nbitq), 
to_sfixed(367577154.0/4294967296.0,1,-nbitq), 
to_sfixed(-289819071.0/4294967296.0,1,-nbitq), 
to_sfixed(332284308.0/4294967296.0,1,-nbitq), 
to_sfixed(219904307.0/4294967296.0,1,-nbitq), 
to_sfixed(-462859232.0/4294967296.0,1,-nbitq), 
to_sfixed(-25436373.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(326315620.0/4294967296.0,1,-nbitq), 
to_sfixed(-893632053.0/4294967296.0,1,-nbitq), 
to_sfixed(-51520234.0/4294967296.0,1,-nbitq), 
to_sfixed(-96870926.0/4294967296.0,1,-nbitq), 
to_sfixed(488757462.0/4294967296.0,1,-nbitq), 
to_sfixed(210823427.0/4294967296.0,1,-nbitq), 
to_sfixed(368091669.0/4294967296.0,1,-nbitq), 
to_sfixed(-423545330.0/4294967296.0,1,-nbitq), 
to_sfixed(629584206.0/4294967296.0,1,-nbitq), 
to_sfixed(249769121.0/4294967296.0,1,-nbitq), 
to_sfixed(264635091.0/4294967296.0,1,-nbitq), 
to_sfixed(466384496.0/4294967296.0,1,-nbitq), 
to_sfixed(-380793968.0/4294967296.0,1,-nbitq), 
to_sfixed(-183213512.0/4294967296.0,1,-nbitq), 
to_sfixed(255006485.0/4294967296.0,1,-nbitq), 
to_sfixed(-31035175.0/4294967296.0,1,-nbitq), 
to_sfixed(-281997559.0/4294967296.0,1,-nbitq), 
to_sfixed(162335678.0/4294967296.0,1,-nbitq), 
to_sfixed(-412644525.0/4294967296.0,1,-nbitq), 
to_sfixed(-271710479.0/4294967296.0,1,-nbitq), 
to_sfixed(-231716876.0/4294967296.0,1,-nbitq), 
to_sfixed(-57552575.0/4294967296.0,1,-nbitq), 
to_sfixed(404843706.0/4294967296.0,1,-nbitq), 
to_sfixed(-510524606.0/4294967296.0,1,-nbitq), 
to_sfixed(352873036.0/4294967296.0,1,-nbitq), 
to_sfixed(-208296118.0/4294967296.0,1,-nbitq), 
to_sfixed(-129278835.0/4294967296.0,1,-nbitq), 
to_sfixed(31790631.0/4294967296.0,1,-nbitq), 
to_sfixed(-11423556.0/4294967296.0,1,-nbitq), 
to_sfixed(7761103.0/4294967296.0,1,-nbitq), 
to_sfixed(-199934346.0/4294967296.0,1,-nbitq), 
to_sfixed(-526074695.0/4294967296.0,1,-nbitq), 
to_sfixed(-94209509.0/4294967296.0,1,-nbitq), 
to_sfixed(669647743.0/4294967296.0,1,-nbitq), 
to_sfixed(40654244.0/4294967296.0,1,-nbitq), 
to_sfixed(-131441795.0/4294967296.0,1,-nbitq), 
to_sfixed(21742654.0/4294967296.0,1,-nbitq), 
to_sfixed(-597839343.0/4294967296.0,1,-nbitq), 
to_sfixed(358166895.0/4294967296.0,1,-nbitq), 
to_sfixed(257207492.0/4294967296.0,1,-nbitq), 
to_sfixed(448524462.0/4294967296.0,1,-nbitq), 
to_sfixed(57773411.0/4294967296.0,1,-nbitq), 
to_sfixed(325732479.0/4294967296.0,1,-nbitq), 
to_sfixed(468521279.0/4294967296.0,1,-nbitq), 
to_sfixed(68216586.0/4294967296.0,1,-nbitq), 
to_sfixed(557259549.0/4294967296.0,1,-nbitq), 
to_sfixed(-176666299.0/4294967296.0,1,-nbitq), 
to_sfixed(415668995.0/4294967296.0,1,-nbitq), 
to_sfixed(326339061.0/4294967296.0,1,-nbitq), 
to_sfixed(152323429.0/4294967296.0,1,-nbitq), 
to_sfixed(-123807876.0/4294967296.0,1,-nbitq), 
to_sfixed(364970329.0/4294967296.0,1,-nbitq), 
to_sfixed(-650898968.0/4294967296.0,1,-nbitq), 
to_sfixed(-196882924.0/4294967296.0,1,-nbitq), 
to_sfixed(-726542081.0/4294967296.0,1,-nbitq), 
to_sfixed(725582093.0/4294967296.0,1,-nbitq), 
to_sfixed(-198804723.0/4294967296.0,1,-nbitq), 
to_sfixed(-82430434.0/4294967296.0,1,-nbitq), 
to_sfixed(-360866106.0/4294967296.0,1,-nbitq), 
to_sfixed(329435214.0/4294967296.0,1,-nbitq), 
to_sfixed(40578113.0/4294967296.0,1,-nbitq), 
to_sfixed(145098154.0/4294967296.0,1,-nbitq), 
to_sfixed(-551500706.0/4294967296.0,1,-nbitq), 
to_sfixed(528540523.0/4294967296.0,1,-nbitq), 
to_sfixed(-323397810.0/4294967296.0,1,-nbitq), 
to_sfixed(-61014595.0/4294967296.0,1,-nbitq), 
to_sfixed(-373018253.0/4294967296.0,1,-nbitq), 
to_sfixed(-324018358.0/4294967296.0,1,-nbitq), 
to_sfixed(284412950.0/4294967296.0,1,-nbitq), 
to_sfixed(283525684.0/4294967296.0,1,-nbitq), 
to_sfixed(305643219.0/4294967296.0,1,-nbitq), 
to_sfixed(131008753.0/4294967296.0,1,-nbitq), 
to_sfixed(116529311.0/4294967296.0,1,-nbitq), 
to_sfixed(420138987.0/4294967296.0,1,-nbitq), 
to_sfixed(-169467246.0/4294967296.0,1,-nbitq), 
to_sfixed(65396499.0/4294967296.0,1,-nbitq), 
to_sfixed(867619980.0/4294967296.0,1,-nbitq), 
to_sfixed(-309018279.0/4294967296.0,1,-nbitq), 
to_sfixed(-421180770.0/4294967296.0,1,-nbitq), 
to_sfixed(-174647080.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(388505582.0/4294967296.0,1,-nbitq), 
to_sfixed(-131118727.0/4294967296.0,1,-nbitq), 
to_sfixed(116657925.0/4294967296.0,1,-nbitq), 
to_sfixed(350687835.0/4294967296.0,1,-nbitq), 
to_sfixed(-139348718.0/4294967296.0,1,-nbitq), 
to_sfixed(-345429793.0/4294967296.0,1,-nbitq), 
to_sfixed(381173248.0/4294967296.0,1,-nbitq), 
to_sfixed(-48302097.0/4294967296.0,1,-nbitq), 
to_sfixed(963186679.0/4294967296.0,1,-nbitq), 
to_sfixed(-29890985.0/4294967296.0,1,-nbitq), 
to_sfixed(-147581937.0/4294967296.0,1,-nbitq), 
to_sfixed(628659127.0/4294967296.0,1,-nbitq), 
to_sfixed(-294639872.0/4294967296.0,1,-nbitq), 
to_sfixed(-684569689.0/4294967296.0,1,-nbitq), 
to_sfixed(31635739.0/4294967296.0,1,-nbitq), 
to_sfixed(67477769.0/4294967296.0,1,-nbitq), 
to_sfixed(-360965227.0/4294967296.0,1,-nbitq), 
to_sfixed(195120727.0/4294967296.0,1,-nbitq), 
to_sfixed(-837503430.0/4294967296.0,1,-nbitq), 
to_sfixed(446493676.0/4294967296.0,1,-nbitq), 
to_sfixed(-400154086.0/4294967296.0,1,-nbitq), 
to_sfixed(98950201.0/4294967296.0,1,-nbitq), 
to_sfixed(516641291.0/4294967296.0,1,-nbitq), 
to_sfixed(-531260066.0/4294967296.0,1,-nbitq), 
to_sfixed(8081987.0/4294967296.0,1,-nbitq), 
to_sfixed(-391660902.0/4294967296.0,1,-nbitq), 
to_sfixed(-72864339.0/4294967296.0,1,-nbitq), 
to_sfixed(-175132287.0/4294967296.0,1,-nbitq), 
to_sfixed(-175178173.0/4294967296.0,1,-nbitq), 
to_sfixed(-209219383.0/4294967296.0,1,-nbitq), 
to_sfixed(654371009.0/4294967296.0,1,-nbitq), 
to_sfixed(-1124783021.0/4294967296.0,1,-nbitq), 
to_sfixed(-777210135.0/4294967296.0,1,-nbitq), 
to_sfixed(543220878.0/4294967296.0,1,-nbitq), 
to_sfixed(-558031135.0/4294967296.0,1,-nbitq), 
to_sfixed(-504910524.0/4294967296.0,1,-nbitq), 
to_sfixed(458724884.0/4294967296.0,1,-nbitq), 
to_sfixed(-25114350.0/4294967296.0,1,-nbitq), 
to_sfixed(-255708744.0/4294967296.0,1,-nbitq), 
to_sfixed(243329715.0/4294967296.0,1,-nbitq), 
to_sfixed(323808287.0/4294967296.0,1,-nbitq), 
to_sfixed(-297672688.0/4294967296.0,1,-nbitq), 
to_sfixed(-144441850.0/4294967296.0,1,-nbitq), 
to_sfixed(-228291053.0/4294967296.0,1,-nbitq), 
to_sfixed(517891743.0/4294967296.0,1,-nbitq), 
to_sfixed(273241660.0/4294967296.0,1,-nbitq), 
to_sfixed(147851723.0/4294967296.0,1,-nbitq), 
to_sfixed(269543958.0/4294967296.0,1,-nbitq), 
to_sfixed(247547589.0/4294967296.0,1,-nbitq), 
to_sfixed(650051421.0/4294967296.0,1,-nbitq), 
to_sfixed(-389650916.0/4294967296.0,1,-nbitq), 
to_sfixed(323190683.0/4294967296.0,1,-nbitq), 
to_sfixed(-465948409.0/4294967296.0,1,-nbitq), 
to_sfixed(-533739618.0/4294967296.0,1,-nbitq), 
to_sfixed(-389647689.0/4294967296.0,1,-nbitq), 
to_sfixed(779875140.0/4294967296.0,1,-nbitq), 
to_sfixed(169664752.0/4294967296.0,1,-nbitq), 
to_sfixed(352885077.0/4294967296.0,1,-nbitq), 
to_sfixed(21096630.0/4294967296.0,1,-nbitq), 
to_sfixed(29661720.0/4294967296.0,1,-nbitq), 
to_sfixed(343136628.0/4294967296.0,1,-nbitq), 
to_sfixed(-575848931.0/4294967296.0,1,-nbitq), 
to_sfixed(-64881057.0/4294967296.0,1,-nbitq), 
to_sfixed(267050470.0/4294967296.0,1,-nbitq), 
to_sfixed(-149948099.0/4294967296.0,1,-nbitq), 
to_sfixed(85517714.0/4294967296.0,1,-nbitq), 
to_sfixed(-549139703.0/4294967296.0,1,-nbitq), 
to_sfixed(-503281203.0/4294967296.0,1,-nbitq), 
to_sfixed(226770427.0/4294967296.0,1,-nbitq), 
to_sfixed(649676666.0/4294967296.0,1,-nbitq), 
to_sfixed(483959955.0/4294967296.0,1,-nbitq), 
to_sfixed(-53862076.0/4294967296.0,1,-nbitq), 
to_sfixed(244425180.0/4294967296.0,1,-nbitq), 
to_sfixed(278357322.0/4294967296.0,1,-nbitq), 
to_sfixed(-7702294.0/4294967296.0,1,-nbitq), 
to_sfixed(-157911098.0/4294967296.0,1,-nbitq), 
to_sfixed(1267743381.0/4294967296.0,1,-nbitq), 
to_sfixed(-447722628.0/4294967296.0,1,-nbitq), 
to_sfixed(-689568582.0/4294967296.0,1,-nbitq), 
to_sfixed(-58727910.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-224365930.0/4294967296.0,1,-nbitq), 
to_sfixed(103675213.0/4294967296.0,1,-nbitq), 
to_sfixed(-324338223.0/4294967296.0,1,-nbitq), 
to_sfixed(510668775.0/4294967296.0,1,-nbitq), 
to_sfixed(6058589.0/4294967296.0,1,-nbitq), 
to_sfixed(-223296266.0/4294967296.0,1,-nbitq), 
to_sfixed(149489600.0/4294967296.0,1,-nbitq), 
to_sfixed(238605026.0/4294967296.0,1,-nbitq), 
to_sfixed(502653318.0/4294967296.0,1,-nbitq), 
to_sfixed(16037059.0/4294967296.0,1,-nbitq), 
to_sfixed(274729525.0/4294967296.0,1,-nbitq), 
to_sfixed(757827700.0/4294967296.0,1,-nbitq), 
to_sfixed(-150783806.0/4294967296.0,1,-nbitq), 
to_sfixed(-353103491.0/4294967296.0,1,-nbitq), 
to_sfixed(-235425333.0/4294967296.0,1,-nbitq), 
to_sfixed(-517263714.0/4294967296.0,1,-nbitq), 
to_sfixed(-7790092.0/4294967296.0,1,-nbitq), 
to_sfixed(-57720802.0/4294967296.0,1,-nbitq), 
to_sfixed(-73150878.0/4294967296.0,1,-nbitq), 
to_sfixed(499242581.0/4294967296.0,1,-nbitq), 
to_sfixed(178582158.0/4294967296.0,1,-nbitq), 
to_sfixed(-245170843.0/4294967296.0,1,-nbitq), 
to_sfixed(-56598900.0/4294967296.0,1,-nbitq), 
to_sfixed(-193528621.0/4294967296.0,1,-nbitq), 
to_sfixed(-557824.0/4294967296.0,1,-nbitq), 
to_sfixed(-107024352.0/4294967296.0,1,-nbitq), 
to_sfixed(-408452215.0/4294967296.0,1,-nbitq), 
to_sfixed(34594346.0/4294967296.0,1,-nbitq), 
to_sfixed(-126160296.0/4294967296.0,1,-nbitq), 
to_sfixed(-792437320.0/4294967296.0,1,-nbitq), 
to_sfixed(382350348.0/4294967296.0,1,-nbitq), 
to_sfixed(-1217392547.0/4294967296.0,1,-nbitq), 
to_sfixed(-137973501.0/4294967296.0,1,-nbitq), 
to_sfixed(411513351.0/4294967296.0,1,-nbitq), 
to_sfixed(-524056313.0/4294967296.0,1,-nbitq), 
to_sfixed(-730446453.0/4294967296.0,1,-nbitq), 
to_sfixed(478612711.0/4294967296.0,1,-nbitq), 
to_sfixed(-443576404.0/4294967296.0,1,-nbitq), 
to_sfixed(63193807.0/4294967296.0,1,-nbitq), 
to_sfixed(-300162597.0/4294967296.0,1,-nbitq), 
to_sfixed(111437062.0/4294967296.0,1,-nbitq), 
to_sfixed(110456431.0/4294967296.0,1,-nbitq), 
to_sfixed(380949622.0/4294967296.0,1,-nbitq), 
to_sfixed(106077776.0/4294967296.0,1,-nbitq), 
to_sfixed(220246339.0/4294967296.0,1,-nbitq), 
to_sfixed(676655496.0/4294967296.0,1,-nbitq), 
to_sfixed(-183079905.0/4294967296.0,1,-nbitq), 
to_sfixed(408259721.0/4294967296.0,1,-nbitq), 
to_sfixed(-223809367.0/4294967296.0,1,-nbitq), 
to_sfixed(19175203.0/4294967296.0,1,-nbitq), 
to_sfixed(67903975.0/4294967296.0,1,-nbitq), 
to_sfixed(340685373.0/4294967296.0,1,-nbitq), 
to_sfixed(-634196281.0/4294967296.0,1,-nbitq), 
to_sfixed(-327797417.0/4294967296.0,1,-nbitq), 
to_sfixed(-599968453.0/4294967296.0,1,-nbitq), 
to_sfixed(162180182.0/4294967296.0,1,-nbitq), 
to_sfixed(557831495.0/4294967296.0,1,-nbitq), 
to_sfixed(1047786552.0/4294967296.0,1,-nbitq), 
to_sfixed(237716884.0/4294967296.0,1,-nbitq), 
to_sfixed(291383513.0/4294967296.0,1,-nbitq), 
to_sfixed(-216685190.0/4294967296.0,1,-nbitq), 
to_sfixed(-116078083.0/4294967296.0,1,-nbitq), 
to_sfixed(-798369883.0/4294967296.0,1,-nbitq), 
to_sfixed(-60537656.0/4294967296.0,1,-nbitq), 
to_sfixed(-15866429.0/4294967296.0,1,-nbitq), 
to_sfixed(-130272892.0/4294967296.0,1,-nbitq), 
to_sfixed(-407115622.0/4294967296.0,1,-nbitq), 
to_sfixed(-178379451.0/4294967296.0,1,-nbitq), 
to_sfixed(-288645812.0/4294967296.0,1,-nbitq), 
to_sfixed(-8350133.0/4294967296.0,1,-nbitq), 
to_sfixed(200495867.0/4294967296.0,1,-nbitq), 
to_sfixed(56751565.0/4294967296.0,1,-nbitq), 
to_sfixed(135894130.0/4294967296.0,1,-nbitq), 
to_sfixed(-248615653.0/4294967296.0,1,-nbitq), 
to_sfixed(443535869.0/4294967296.0,1,-nbitq), 
to_sfixed(-311644734.0/4294967296.0,1,-nbitq), 
to_sfixed(1768600568.0/4294967296.0,1,-nbitq), 
to_sfixed(-246933501.0/4294967296.0,1,-nbitq), 
to_sfixed(-81638370.0/4294967296.0,1,-nbitq), 
to_sfixed(-290234218.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(106832838.0/4294967296.0,1,-nbitq), 
to_sfixed(526203704.0/4294967296.0,1,-nbitq), 
to_sfixed(-70793605.0/4294967296.0,1,-nbitq), 
to_sfixed(643425106.0/4294967296.0,1,-nbitq), 
to_sfixed(-262449120.0/4294967296.0,1,-nbitq), 
to_sfixed(-546896961.0/4294967296.0,1,-nbitq), 
to_sfixed(27814183.0/4294967296.0,1,-nbitq), 
to_sfixed(69673428.0/4294967296.0,1,-nbitq), 
to_sfixed(274250777.0/4294967296.0,1,-nbitq), 
to_sfixed(59942086.0/4294967296.0,1,-nbitq), 
to_sfixed(208852494.0/4294967296.0,1,-nbitq), 
to_sfixed(966716539.0/4294967296.0,1,-nbitq), 
to_sfixed(-11993083.0/4294967296.0,1,-nbitq), 
to_sfixed(-317380636.0/4294967296.0,1,-nbitq), 
to_sfixed(-189623776.0/4294967296.0,1,-nbitq), 
to_sfixed(-9368979.0/4294967296.0,1,-nbitq), 
to_sfixed(113787830.0/4294967296.0,1,-nbitq), 
to_sfixed(158777835.0/4294967296.0,1,-nbitq), 
to_sfixed(-740313232.0/4294967296.0,1,-nbitq), 
to_sfixed(-102316911.0/4294967296.0,1,-nbitq), 
to_sfixed(291637760.0/4294967296.0,1,-nbitq), 
to_sfixed(-216946247.0/4294967296.0,1,-nbitq), 
to_sfixed(199254025.0/4294967296.0,1,-nbitq), 
to_sfixed(217344561.0/4294967296.0,1,-nbitq), 
to_sfixed(243021191.0/4294967296.0,1,-nbitq), 
to_sfixed(503179248.0/4294967296.0,1,-nbitq), 
to_sfixed(-826814890.0/4294967296.0,1,-nbitq), 
to_sfixed(-21173987.0/4294967296.0,1,-nbitq), 
to_sfixed(254980729.0/4294967296.0,1,-nbitq), 
to_sfixed(-1059549039.0/4294967296.0,1,-nbitq), 
to_sfixed(196486573.0/4294967296.0,1,-nbitq), 
to_sfixed(-236543663.0/4294967296.0,1,-nbitq), 
to_sfixed(-54498886.0/4294967296.0,1,-nbitq), 
to_sfixed(14530269.0/4294967296.0,1,-nbitq), 
to_sfixed(-397237848.0/4294967296.0,1,-nbitq), 
to_sfixed(-216922809.0/4294967296.0,1,-nbitq), 
to_sfixed(226021654.0/4294967296.0,1,-nbitq), 
to_sfixed(-129246106.0/4294967296.0,1,-nbitq), 
to_sfixed(75333249.0/4294967296.0,1,-nbitq), 
to_sfixed(-321209007.0/4294967296.0,1,-nbitq), 
to_sfixed(651262821.0/4294967296.0,1,-nbitq), 
to_sfixed(364997059.0/4294967296.0,1,-nbitq), 
to_sfixed(947804485.0/4294967296.0,1,-nbitq), 
to_sfixed(725342059.0/4294967296.0,1,-nbitq), 
to_sfixed(177095367.0/4294967296.0,1,-nbitq), 
to_sfixed(940910001.0/4294967296.0,1,-nbitq), 
to_sfixed(115231175.0/4294967296.0,1,-nbitq), 
to_sfixed(94170140.0/4294967296.0,1,-nbitq), 
to_sfixed(-5073136.0/4294967296.0,1,-nbitq), 
to_sfixed(253942814.0/4294967296.0,1,-nbitq), 
to_sfixed(-21728674.0/4294967296.0,1,-nbitq), 
to_sfixed(976750412.0/4294967296.0,1,-nbitq), 
to_sfixed(-423079979.0/4294967296.0,1,-nbitq), 
to_sfixed(-99657249.0/4294967296.0,1,-nbitq), 
to_sfixed(648447106.0/4294967296.0,1,-nbitq), 
to_sfixed(465995609.0/4294967296.0,1,-nbitq), 
to_sfixed(-11974664.0/4294967296.0,1,-nbitq), 
to_sfixed(926233229.0/4294967296.0,1,-nbitq), 
to_sfixed(-204713185.0/4294967296.0,1,-nbitq), 
to_sfixed(-112679845.0/4294967296.0,1,-nbitq), 
to_sfixed(93573065.0/4294967296.0,1,-nbitq), 
to_sfixed(-204619974.0/4294967296.0,1,-nbitq), 
to_sfixed(-450703311.0/4294967296.0,1,-nbitq), 
to_sfixed(-99240767.0/4294967296.0,1,-nbitq), 
to_sfixed(-20063120.0/4294967296.0,1,-nbitq), 
to_sfixed(-68769172.0/4294967296.0,1,-nbitq), 
to_sfixed(-359646176.0/4294967296.0,1,-nbitq), 
to_sfixed(-130374050.0/4294967296.0,1,-nbitq), 
to_sfixed(52201290.0/4294967296.0,1,-nbitq), 
to_sfixed(-247313615.0/4294967296.0,1,-nbitq), 
to_sfixed(400825391.0/4294967296.0,1,-nbitq), 
to_sfixed(220658566.0/4294967296.0,1,-nbitq), 
to_sfixed(426535957.0/4294967296.0,1,-nbitq), 
to_sfixed(-655113.0/4294967296.0,1,-nbitq), 
to_sfixed(340078603.0/4294967296.0,1,-nbitq), 
to_sfixed(180328937.0/4294967296.0,1,-nbitq), 
to_sfixed(1120958127.0/4294967296.0,1,-nbitq), 
to_sfixed(-51740206.0/4294967296.0,1,-nbitq), 
to_sfixed(437535119.0/4294967296.0,1,-nbitq), 
to_sfixed(-103594719.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(404395652.0/4294967296.0,1,-nbitq), 
to_sfixed(45851325.0/4294967296.0,1,-nbitq), 
to_sfixed(-202801527.0/4294967296.0,1,-nbitq), 
to_sfixed(107767384.0/4294967296.0,1,-nbitq), 
to_sfixed(-384011945.0/4294967296.0,1,-nbitq), 
to_sfixed(-621778306.0/4294967296.0,1,-nbitq), 
to_sfixed(-181300742.0/4294967296.0,1,-nbitq), 
to_sfixed(214313697.0/4294967296.0,1,-nbitq), 
to_sfixed(851213351.0/4294967296.0,1,-nbitq), 
to_sfixed(-48921060.0/4294967296.0,1,-nbitq), 
to_sfixed(-123453034.0/4294967296.0,1,-nbitq), 
to_sfixed(673011891.0/4294967296.0,1,-nbitq), 
to_sfixed(-114818052.0/4294967296.0,1,-nbitq), 
to_sfixed(-194356257.0/4294967296.0,1,-nbitq), 
to_sfixed(235330591.0/4294967296.0,1,-nbitq), 
to_sfixed(306042691.0/4294967296.0,1,-nbitq), 
to_sfixed(-42171573.0/4294967296.0,1,-nbitq), 
to_sfixed(-147165202.0/4294967296.0,1,-nbitq), 
to_sfixed(-405105176.0/4294967296.0,1,-nbitq), 
to_sfixed(-182116005.0/4294967296.0,1,-nbitq), 
to_sfixed(-266436339.0/4294967296.0,1,-nbitq), 
to_sfixed(-3122447.0/4294967296.0,1,-nbitq), 
to_sfixed(-117776462.0/4294967296.0,1,-nbitq), 
to_sfixed(196958709.0/4294967296.0,1,-nbitq), 
to_sfixed(124246126.0/4294967296.0,1,-nbitq), 
to_sfixed(-186976809.0/4294967296.0,1,-nbitq), 
to_sfixed(-359684347.0/4294967296.0,1,-nbitq), 
to_sfixed(120668413.0/4294967296.0,1,-nbitq), 
to_sfixed(-69749820.0/4294967296.0,1,-nbitq), 
to_sfixed(-646212925.0/4294967296.0,1,-nbitq), 
to_sfixed(336453952.0/4294967296.0,1,-nbitq), 
to_sfixed(-704043442.0/4294967296.0,1,-nbitq), 
to_sfixed(318864229.0/4294967296.0,1,-nbitq), 
to_sfixed(-159994473.0/4294967296.0,1,-nbitq), 
to_sfixed(-649287362.0/4294967296.0,1,-nbitq), 
to_sfixed(-493379647.0/4294967296.0,1,-nbitq), 
to_sfixed(-110807477.0/4294967296.0,1,-nbitq), 
to_sfixed(-94128678.0/4294967296.0,1,-nbitq), 
to_sfixed(-125682864.0/4294967296.0,1,-nbitq), 
to_sfixed(47894334.0/4294967296.0,1,-nbitq), 
to_sfixed(190346900.0/4294967296.0,1,-nbitq), 
to_sfixed(3380014.0/4294967296.0,1,-nbitq), 
to_sfixed(1190606809.0/4294967296.0,1,-nbitq), 
to_sfixed(1272580194.0/4294967296.0,1,-nbitq), 
to_sfixed(93988388.0/4294967296.0,1,-nbitq), 
to_sfixed(923774045.0/4294967296.0,1,-nbitq), 
to_sfixed(117035480.0/4294967296.0,1,-nbitq), 
to_sfixed(231178958.0/4294967296.0,1,-nbitq), 
to_sfixed(-400580256.0/4294967296.0,1,-nbitq), 
to_sfixed(270932563.0/4294967296.0,1,-nbitq), 
to_sfixed(284182839.0/4294967296.0,1,-nbitq), 
to_sfixed(604608486.0/4294967296.0,1,-nbitq), 
to_sfixed(-484890623.0/4294967296.0,1,-nbitq), 
to_sfixed(59280066.0/4294967296.0,1,-nbitq), 
to_sfixed(1404803321.0/4294967296.0,1,-nbitq), 
to_sfixed(130942379.0/4294967296.0,1,-nbitq), 
to_sfixed(26071680.0/4294967296.0,1,-nbitq), 
to_sfixed(853171621.0/4294967296.0,1,-nbitq), 
to_sfixed(79050225.0/4294967296.0,1,-nbitq), 
to_sfixed(224741140.0/4294967296.0,1,-nbitq), 
to_sfixed(-5759723.0/4294967296.0,1,-nbitq), 
to_sfixed(-29765822.0/4294967296.0,1,-nbitq), 
to_sfixed(-455965121.0/4294967296.0,1,-nbitq), 
to_sfixed(116614106.0/4294967296.0,1,-nbitq), 
to_sfixed(-279739550.0/4294967296.0,1,-nbitq), 
to_sfixed(-15630964.0/4294967296.0,1,-nbitq), 
to_sfixed(-557316913.0/4294967296.0,1,-nbitq), 
to_sfixed(1042895711.0/4294967296.0,1,-nbitq), 
to_sfixed(-196829384.0/4294967296.0,1,-nbitq), 
to_sfixed(-501181721.0/4294967296.0,1,-nbitq), 
to_sfixed(336983492.0/4294967296.0,1,-nbitq), 
to_sfixed(-41818266.0/4294967296.0,1,-nbitq), 
to_sfixed(438439161.0/4294967296.0,1,-nbitq), 
to_sfixed(417515757.0/4294967296.0,1,-nbitq), 
to_sfixed(-203838263.0/4294967296.0,1,-nbitq), 
to_sfixed(-73028816.0/4294967296.0,1,-nbitq), 
to_sfixed(411568624.0/4294967296.0,1,-nbitq), 
to_sfixed(12844822.0/4294967296.0,1,-nbitq), 
to_sfixed(-6620914.0/4294967296.0,1,-nbitq), 
to_sfixed(-24895282.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(292587866.0/4294967296.0,1,-nbitq), 
to_sfixed(405636606.0/4294967296.0,1,-nbitq), 
to_sfixed(-148715615.0/4294967296.0,1,-nbitq), 
to_sfixed(569255251.0/4294967296.0,1,-nbitq), 
to_sfixed(-844861134.0/4294967296.0,1,-nbitq), 
to_sfixed(-536470417.0/4294967296.0,1,-nbitq), 
to_sfixed(531897246.0/4294967296.0,1,-nbitq), 
to_sfixed(-285789356.0/4294967296.0,1,-nbitq), 
to_sfixed(-426341396.0/4294967296.0,1,-nbitq), 
to_sfixed(204776226.0/4294967296.0,1,-nbitq), 
to_sfixed(647516532.0/4294967296.0,1,-nbitq), 
to_sfixed(36800566.0/4294967296.0,1,-nbitq), 
to_sfixed(-242012464.0/4294967296.0,1,-nbitq), 
to_sfixed(549490558.0/4294967296.0,1,-nbitq), 
to_sfixed(112571642.0/4294967296.0,1,-nbitq), 
to_sfixed(269790265.0/4294967296.0,1,-nbitq), 
to_sfixed(292000565.0/4294967296.0,1,-nbitq), 
to_sfixed(209181840.0/4294967296.0,1,-nbitq), 
to_sfixed(-367161338.0/4294967296.0,1,-nbitq), 
to_sfixed(-56253349.0/4294967296.0,1,-nbitq), 
to_sfixed(316330489.0/4294967296.0,1,-nbitq), 
to_sfixed(-187024594.0/4294967296.0,1,-nbitq), 
to_sfixed(674406199.0/4294967296.0,1,-nbitq), 
to_sfixed(34652831.0/4294967296.0,1,-nbitq), 
to_sfixed(-270202689.0/4294967296.0,1,-nbitq), 
to_sfixed(314070301.0/4294967296.0,1,-nbitq), 
to_sfixed(20722823.0/4294967296.0,1,-nbitq), 
to_sfixed(-494048641.0/4294967296.0,1,-nbitq), 
to_sfixed(-109615721.0/4294967296.0,1,-nbitq), 
to_sfixed(-185106112.0/4294967296.0,1,-nbitq), 
to_sfixed(805315710.0/4294967296.0,1,-nbitq), 
to_sfixed(-154582348.0/4294967296.0,1,-nbitq), 
to_sfixed(179463145.0/4294967296.0,1,-nbitq), 
to_sfixed(385421811.0/4294967296.0,1,-nbitq), 
to_sfixed(-337090851.0/4294967296.0,1,-nbitq), 
to_sfixed(-620572453.0/4294967296.0,1,-nbitq), 
to_sfixed(26542852.0/4294967296.0,1,-nbitq), 
to_sfixed(-12327453.0/4294967296.0,1,-nbitq), 
to_sfixed(60356270.0/4294967296.0,1,-nbitq), 
to_sfixed(-326426917.0/4294967296.0,1,-nbitq), 
to_sfixed(101989995.0/4294967296.0,1,-nbitq), 
to_sfixed(-403006630.0/4294967296.0,1,-nbitq), 
to_sfixed(894889054.0/4294967296.0,1,-nbitq), 
to_sfixed(861149774.0/4294967296.0,1,-nbitq), 
to_sfixed(-156714968.0/4294967296.0,1,-nbitq), 
to_sfixed(737206487.0/4294967296.0,1,-nbitq), 
to_sfixed(-165656084.0/4294967296.0,1,-nbitq), 
to_sfixed(424375982.0/4294967296.0,1,-nbitq), 
to_sfixed(-584133220.0/4294967296.0,1,-nbitq), 
to_sfixed(-197976024.0/4294967296.0,1,-nbitq), 
to_sfixed(399160434.0/4294967296.0,1,-nbitq), 
to_sfixed(451598264.0/4294967296.0,1,-nbitq), 
to_sfixed(6147226.0/4294967296.0,1,-nbitq), 
to_sfixed(331527101.0/4294967296.0,1,-nbitq), 
to_sfixed(622257301.0/4294967296.0,1,-nbitq), 
to_sfixed(-292554472.0/4294967296.0,1,-nbitq), 
to_sfixed(593046543.0/4294967296.0,1,-nbitq), 
to_sfixed(630489034.0/4294967296.0,1,-nbitq), 
to_sfixed(-179080286.0/4294967296.0,1,-nbitq), 
to_sfixed(321835846.0/4294967296.0,1,-nbitq), 
to_sfixed(356681741.0/4294967296.0,1,-nbitq), 
to_sfixed(-110410789.0/4294967296.0,1,-nbitq), 
to_sfixed(-195639874.0/4294967296.0,1,-nbitq), 
to_sfixed(376746160.0/4294967296.0,1,-nbitq), 
to_sfixed(-367670171.0/4294967296.0,1,-nbitq), 
to_sfixed(-89484817.0/4294967296.0,1,-nbitq), 
to_sfixed(-286289322.0/4294967296.0,1,-nbitq), 
to_sfixed(562159646.0/4294967296.0,1,-nbitq), 
to_sfixed(426879899.0/4294967296.0,1,-nbitq), 
to_sfixed(-899319090.0/4294967296.0,1,-nbitq), 
to_sfixed(-499706988.0/4294967296.0,1,-nbitq), 
to_sfixed(-419284173.0/4294967296.0,1,-nbitq), 
to_sfixed(541597620.0/4294967296.0,1,-nbitq), 
to_sfixed(-55155895.0/4294967296.0,1,-nbitq), 
to_sfixed(34930072.0/4294967296.0,1,-nbitq), 
to_sfixed(-266310480.0/4294967296.0,1,-nbitq), 
to_sfixed(229745421.0/4294967296.0,1,-nbitq), 
to_sfixed(-32915889.0/4294967296.0,1,-nbitq), 
to_sfixed(580642941.0/4294967296.0,1,-nbitq), 
to_sfixed(-430649716.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(689393197.0/4294967296.0,1,-nbitq), 
to_sfixed(417186169.0/4294967296.0,1,-nbitq), 
to_sfixed(-827952038.0/4294967296.0,1,-nbitq), 
to_sfixed(165562345.0/4294967296.0,1,-nbitq), 
to_sfixed(-1315065989.0/4294967296.0,1,-nbitq), 
to_sfixed(-339217620.0/4294967296.0,1,-nbitq), 
to_sfixed(135949220.0/4294967296.0,1,-nbitq), 
to_sfixed(-270279433.0/4294967296.0,1,-nbitq), 
to_sfixed(279164113.0/4294967296.0,1,-nbitq), 
to_sfixed(14835158.0/4294967296.0,1,-nbitq), 
to_sfixed(442969292.0/4294967296.0,1,-nbitq), 
to_sfixed(219072821.0/4294967296.0,1,-nbitq), 
to_sfixed(-17950090.0/4294967296.0,1,-nbitq), 
to_sfixed(1309724724.0/4294967296.0,1,-nbitq), 
to_sfixed(360595411.0/4294967296.0,1,-nbitq), 
to_sfixed(-136533464.0/4294967296.0,1,-nbitq), 
to_sfixed(338637154.0/4294967296.0,1,-nbitq), 
to_sfixed(-251598394.0/4294967296.0,1,-nbitq), 
to_sfixed(-32902275.0/4294967296.0,1,-nbitq), 
to_sfixed(-513825645.0/4294967296.0,1,-nbitq), 
to_sfixed(-419355483.0/4294967296.0,1,-nbitq), 
to_sfixed(-219505451.0/4294967296.0,1,-nbitq), 
to_sfixed(701689373.0/4294967296.0,1,-nbitq), 
to_sfixed(554128150.0/4294967296.0,1,-nbitq), 
to_sfixed(273271288.0/4294967296.0,1,-nbitq), 
to_sfixed(656353842.0/4294967296.0,1,-nbitq), 
to_sfixed(-404141940.0/4294967296.0,1,-nbitq), 
to_sfixed(-38624139.0/4294967296.0,1,-nbitq), 
to_sfixed(-362263496.0/4294967296.0,1,-nbitq), 
to_sfixed(231601662.0/4294967296.0,1,-nbitq), 
to_sfixed(14654279.0/4294967296.0,1,-nbitq), 
to_sfixed(-688671713.0/4294967296.0,1,-nbitq), 
to_sfixed(-523396583.0/4294967296.0,1,-nbitq), 
to_sfixed(-161291653.0/4294967296.0,1,-nbitq), 
to_sfixed(107233915.0/4294967296.0,1,-nbitq), 
to_sfixed(-484631886.0/4294967296.0,1,-nbitq), 
to_sfixed(-200622525.0/4294967296.0,1,-nbitq), 
to_sfixed(189347465.0/4294967296.0,1,-nbitq), 
to_sfixed(306722727.0/4294967296.0,1,-nbitq), 
to_sfixed(-11901059.0/4294967296.0,1,-nbitq), 
to_sfixed(320685911.0/4294967296.0,1,-nbitq), 
to_sfixed(-517162760.0/4294967296.0,1,-nbitq), 
to_sfixed(1346560097.0/4294967296.0,1,-nbitq), 
to_sfixed(1045940914.0/4294967296.0,1,-nbitq), 
to_sfixed(452233006.0/4294967296.0,1,-nbitq), 
to_sfixed(196576555.0/4294967296.0,1,-nbitq), 
to_sfixed(225431607.0/4294967296.0,1,-nbitq), 
to_sfixed(549673317.0/4294967296.0,1,-nbitq), 
to_sfixed(-447714030.0/4294967296.0,1,-nbitq), 
to_sfixed(67056564.0/4294967296.0,1,-nbitq), 
to_sfixed(363652678.0/4294967296.0,1,-nbitq), 
to_sfixed(463810832.0/4294967296.0,1,-nbitq), 
to_sfixed(-695886542.0/4294967296.0,1,-nbitq), 
to_sfixed(855129469.0/4294967296.0,1,-nbitq), 
to_sfixed(426866041.0/4294967296.0,1,-nbitq), 
to_sfixed(-754026439.0/4294967296.0,1,-nbitq), 
to_sfixed(518500115.0/4294967296.0,1,-nbitq), 
to_sfixed(-15249024.0/4294967296.0,1,-nbitq), 
to_sfixed(-253587460.0/4294967296.0,1,-nbitq), 
to_sfixed(218433034.0/4294967296.0,1,-nbitq), 
to_sfixed(98254233.0/4294967296.0,1,-nbitq), 
to_sfixed(82774700.0/4294967296.0,1,-nbitq), 
to_sfixed(-609918102.0/4294967296.0,1,-nbitq), 
to_sfixed(122084453.0/4294967296.0,1,-nbitq), 
to_sfixed(111439951.0/4294967296.0,1,-nbitq), 
to_sfixed(158726150.0/4294967296.0,1,-nbitq), 
to_sfixed(93554867.0/4294967296.0,1,-nbitq), 
to_sfixed(379149512.0/4294967296.0,1,-nbitq), 
to_sfixed(-42754399.0/4294967296.0,1,-nbitq), 
to_sfixed(-1313610089.0/4294967296.0,1,-nbitq), 
to_sfixed(-69173953.0/4294967296.0,1,-nbitq), 
to_sfixed(118991311.0/4294967296.0,1,-nbitq), 
to_sfixed(707744954.0/4294967296.0,1,-nbitq), 
to_sfixed(-226231778.0/4294967296.0,1,-nbitq), 
to_sfixed(-451420494.0/4294967296.0,1,-nbitq), 
to_sfixed(-451991935.0/4294967296.0,1,-nbitq), 
to_sfixed(-303590498.0/4294967296.0,1,-nbitq), 
to_sfixed(139024395.0/4294967296.0,1,-nbitq), 
to_sfixed(-75818090.0/4294967296.0,1,-nbitq), 
to_sfixed(-154554983.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(784907104.0/4294967296.0,1,-nbitq), 
to_sfixed(1463330819.0/4294967296.0,1,-nbitq), 
to_sfixed(-802904931.0/4294967296.0,1,-nbitq), 
to_sfixed(428178660.0/4294967296.0,1,-nbitq), 
to_sfixed(-1108608394.0/4294967296.0,1,-nbitq), 
to_sfixed(-580119176.0/4294967296.0,1,-nbitq), 
to_sfixed(43341220.0/4294967296.0,1,-nbitq), 
to_sfixed(-28528788.0/4294967296.0,1,-nbitq), 
to_sfixed(-243739023.0/4294967296.0,1,-nbitq), 
to_sfixed(-1117913.0/4294967296.0,1,-nbitq), 
to_sfixed(767888701.0/4294967296.0,1,-nbitq), 
to_sfixed(-29856485.0/4294967296.0,1,-nbitq), 
to_sfixed(-373709572.0/4294967296.0,1,-nbitq), 
to_sfixed(876754135.0/4294967296.0,1,-nbitq), 
to_sfixed(-57336349.0/4294967296.0,1,-nbitq), 
to_sfixed(-207089371.0/4294967296.0,1,-nbitq), 
to_sfixed(288725776.0/4294967296.0,1,-nbitq), 
to_sfixed(-159869438.0/4294967296.0,1,-nbitq), 
to_sfixed(-363582680.0/4294967296.0,1,-nbitq), 
to_sfixed(34055786.0/4294967296.0,1,-nbitq), 
to_sfixed(228689403.0/4294967296.0,1,-nbitq), 
to_sfixed(-894615603.0/4294967296.0,1,-nbitq), 
to_sfixed(-97276074.0/4294967296.0,1,-nbitq), 
to_sfixed(213940207.0/4294967296.0,1,-nbitq), 
to_sfixed(289158921.0/4294967296.0,1,-nbitq), 
to_sfixed(991989261.0/4294967296.0,1,-nbitq), 
to_sfixed(-34601899.0/4294967296.0,1,-nbitq), 
to_sfixed(-289328365.0/4294967296.0,1,-nbitq), 
to_sfixed(63340342.0/4294967296.0,1,-nbitq), 
to_sfixed(408351802.0/4294967296.0,1,-nbitq), 
to_sfixed(293237958.0/4294967296.0,1,-nbitq), 
to_sfixed(-517216464.0/4294967296.0,1,-nbitq), 
to_sfixed(-102693600.0/4294967296.0,1,-nbitq), 
to_sfixed(-291138521.0/4294967296.0,1,-nbitq), 
to_sfixed(-142567247.0/4294967296.0,1,-nbitq), 
to_sfixed(-61992045.0/4294967296.0,1,-nbitq), 
to_sfixed(-412696697.0/4294967296.0,1,-nbitq), 
to_sfixed(-62670368.0/4294967296.0,1,-nbitq), 
to_sfixed(327218534.0/4294967296.0,1,-nbitq), 
to_sfixed(-493971772.0/4294967296.0,1,-nbitq), 
to_sfixed(-150542995.0/4294967296.0,1,-nbitq), 
to_sfixed(-355294159.0/4294967296.0,1,-nbitq), 
to_sfixed(1317959573.0/4294967296.0,1,-nbitq), 
to_sfixed(1218736405.0/4294967296.0,1,-nbitq), 
to_sfixed(507689110.0/4294967296.0,1,-nbitq), 
to_sfixed(-171170238.0/4294967296.0,1,-nbitq), 
to_sfixed(177686635.0/4294967296.0,1,-nbitq), 
to_sfixed(651856129.0/4294967296.0,1,-nbitq), 
to_sfixed(-7862910.0/4294967296.0,1,-nbitq), 
to_sfixed(544051285.0/4294967296.0,1,-nbitq), 
to_sfixed(421616288.0/4294967296.0,1,-nbitq), 
to_sfixed(125867125.0/4294967296.0,1,-nbitq), 
to_sfixed(-271077412.0/4294967296.0,1,-nbitq), 
to_sfixed(228496086.0/4294967296.0,1,-nbitq), 
to_sfixed(1148329438.0/4294967296.0,1,-nbitq), 
to_sfixed(-477413650.0/4294967296.0,1,-nbitq), 
to_sfixed(99585430.0/4294967296.0,1,-nbitq), 
to_sfixed(431074468.0/4294967296.0,1,-nbitq), 
to_sfixed(-60921105.0/4294967296.0,1,-nbitq), 
to_sfixed(-320917523.0/4294967296.0,1,-nbitq), 
to_sfixed(-59952051.0/4294967296.0,1,-nbitq), 
to_sfixed(-541847881.0/4294967296.0,1,-nbitq), 
to_sfixed(-292487653.0/4294967296.0,1,-nbitq), 
to_sfixed(8723785.0/4294967296.0,1,-nbitq), 
to_sfixed(-78725280.0/4294967296.0,1,-nbitq), 
to_sfixed(328541819.0/4294967296.0,1,-nbitq), 
to_sfixed(-649364009.0/4294967296.0,1,-nbitq), 
to_sfixed(1151415129.0/4294967296.0,1,-nbitq), 
to_sfixed(83550467.0/4294967296.0,1,-nbitq), 
to_sfixed(-385255059.0/4294967296.0,1,-nbitq), 
to_sfixed(284850784.0/4294967296.0,1,-nbitq), 
to_sfixed(-446257903.0/4294967296.0,1,-nbitq), 
to_sfixed(482569162.0/4294967296.0,1,-nbitq), 
to_sfixed(64641946.0/4294967296.0,1,-nbitq), 
to_sfixed(-76315349.0/4294967296.0,1,-nbitq), 
to_sfixed(-263574464.0/4294967296.0,1,-nbitq), 
to_sfixed(-302617252.0/4294967296.0,1,-nbitq), 
to_sfixed(138959330.0/4294967296.0,1,-nbitq), 
to_sfixed(217616293.0/4294967296.0,1,-nbitq), 
to_sfixed(199560089.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(314561069.0/4294967296.0,1,-nbitq), 
to_sfixed(1242432709.0/4294967296.0,1,-nbitq), 
to_sfixed(-618543424.0/4294967296.0,1,-nbitq), 
to_sfixed(367354611.0/4294967296.0,1,-nbitq), 
to_sfixed(-821019116.0/4294967296.0,1,-nbitq), 
to_sfixed(-566887435.0/4294967296.0,1,-nbitq), 
to_sfixed(-479863712.0/4294967296.0,1,-nbitq), 
to_sfixed(-2080122.0/4294967296.0,1,-nbitq), 
to_sfixed(23499773.0/4294967296.0,1,-nbitq), 
to_sfixed(400630151.0/4294967296.0,1,-nbitq), 
to_sfixed(715173705.0/4294967296.0,1,-nbitq), 
to_sfixed(-83907386.0/4294967296.0,1,-nbitq), 
to_sfixed(-46229943.0/4294967296.0,1,-nbitq), 
to_sfixed(463475101.0/4294967296.0,1,-nbitq), 
to_sfixed(-239479430.0/4294967296.0,1,-nbitq), 
to_sfixed(-320269966.0/4294967296.0,1,-nbitq), 
to_sfixed(115987208.0/4294967296.0,1,-nbitq), 
to_sfixed(177523176.0/4294967296.0,1,-nbitq), 
to_sfixed(-134242566.0/4294967296.0,1,-nbitq), 
to_sfixed(-71032684.0/4294967296.0,1,-nbitq), 
to_sfixed(20426797.0/4294967296.0,1,-nbitq), 
to_sfixed(-628192197.0/4294967296.0,1,-nbitq), 
to_sfixed(286614873.0/4294967296.0,1,-nbitq), 
to_sfixed(273208334.0/4294967296.0,1,-nbitq), 
to_sfixed(160467265.0/4294967296.0,1,-nbitq), 
to_sfixed(299861824.0/4294967296.0,1,-nbitq), 
to_sfixed(504908450.0/4294967296.0,1,-nbitq), 
to_sfixed(551442435.0/4294967296.0,1,-nbitq), 
to_sfixed(7199776.0/4294967296.0,1,-nbitq), 
to_sfixed(551844905.0/4294967296.0,1,-nbitq), 
to_sfixed(283178279.0/4294967296.0,1,-nbitq), 
to_sfixed(251628784.0/4294967296.0,1,-nbitq), 
to_sfixed(362218079.0/4294967296.0,1,-nbitq), 
to_sfixed(-175760672.0/4294967296.0,1,-nbitq), 
to_sfixed(14175847.0/4294967296.0,1,-nbitq), 
to_sfixed(127646442.0/4294967296.0,1,-nbitq), 
to_sfixed(-376874840.0/4294967296.0,1,-nbitq), 
to_sfixed(55633239.0/4294967296.0,1,-nbitq), 
to_sfixed(-357327223.0/4294967296.0,1,-nbitq), 
to_sfixed(-330459849.0/4294967296.0,1,-nbitq), 
to_sfixed(261047118.0/4294967296.0,1,-nbitq), 
to_sfixed(-104149233.0/4294967296.0,1,-nbitq), 
to_sfixed(688442561.0/4294967296.0,1,-nbitq), 
to_sfixed(1050534064.0/4294967296.0,1,-nbitq), 
to_sfixed(790395536.0/4294967296.0,1,-nbitq), 
to_sfixed(487230304.0/4294967296.0,1,-nbitq), 
to_sfixed(145154944.0/4294967296.0,1,-nbitq), 
to_sfixed(430378523.0/4294967296.0,1,-nbitq), 
to_sfixed(-287697095.0/4294967296.0,1,-nbitq), 
to_sfixed(811857929.0/4294967296.0,1,-nbitq), 
to_sfixed(449414975.0/4294967296.0,1,-nbitq), 
to_sfixed(-543182031.0/4294967296.0,1,-nbitq), 
to_sfixed(-351699242.0/4294967296.0,1,-nbitq), 
to_sfixed(134424635.0/4294967296.0,1,-nbitq), 
to_sfixed(1097414248.0/4294967296.0,1,-nbitq), 
to_sfixed(-763747757.0/4294967296.0,1,-nbitq), 
to_sfixed(461094477.0/4294967296.0,1,-nbitq), 
to_sfixed(134543879.0/4294967296.0,1,-nbitq), 
to_sfixed(389994614.0/4294967296.0,1,-nbitq), 
to_sfixed(-97325461.0/4294967296.0,1,-nbitq), 
to_sfixed(-55706062.0/4294967296.0,1,-nbitq), 
to_sfixed(-540865621.0/4294967296.0,1,-nbitq), 
to_sfixed(-96834325.0/4294967296.0,1,-nbitq), 
to_sfixed(-657109733.0/4294967296.0,1,-nbitq), 
to_sfixed(-128569605.0/4294967296.0,1,-nbitq), 
to_sfixed(165077913.0/4294967296.0,1,-nbitq), 
to_sfixed(-123336281.0/4294967296.0,1,-nbitq), 
to_sfixed(1559068896.0/4294967296.0,1,-nbitq), 
to_sfixed(-162966006.0/4294967296.0,1,-nbitq), 
to_sfixed(14821256.0/4294967296.0,1,-nbitq), 
to_sfixed(1068424314.0/4294967296.0,1,-nbitq), 
to_sfixed(-367625809.0/4294967296.0,1,-nbitq), 
to_sfixed(1142948495.0/4294967296.0,1,-nbitq), 
to_sfixed(-159414596.0/4294967296.0,1,-nbitq), 
to_sfixed(53925600.0/4294967296.0,1,-nbitq), 
to_sfixed(293084386.0/4294967296.0,1,-nbitq), 
to_sfixed(-885967424.0/4294967296.0,1,-nbitq), 
to_sfixed(127597891.0/4294967296.0,1,-nbitq), 
to_sfixed(430899242.0/4294967296.0,1,-nbitq), 
to_sfixed(280853742.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(168589985.0/4294967296.0,1,-nbitq), 
to_sfixed(436046814.0/4294967296.0,1,-nbitq), 
to_sfixed(-46430240.0/4294967296.0,1,-nbitq), 
to_sfixed(274817535.0/4294967296.0,1,-nbitq), 
to_sfixed(-163764244.0/4294967296.0,1,-nbitq), 
to_sfixed(-256878430.0/4294967296.0,1,-nbitq), 
to_sfixed(-69919145.0/4294967296.0,1,-nbitq), 
to_sfixed(-306065977.0/4294967296.0,1,-nbitq), 
to_sfixed(295911451.0/4294967296.0,1,-nbitq), 
to_sfixed(57949732.0/4294967296.0,1,-nbitq), 
to_sfixed(1161327863.0/4294967296.0,1,-nbitq), 
to_sfixed(392567049.0/4294967296.0,1,-nbitq), 
to_sfixed(-212168605.0/4294967296.0,1,-nbitq), 
to_sfixed(1054928701.0/4294967296.0,1,-nbitq), 
to_sfixed(-53301767.0/4294967296.0,1,-nbitq), 
to_sfixed(252307595.0/4294967296.0,1,-nbitq), 
to_sfixed(-33697395.0/4294967296.0,1,-nbitq), 
to_sfixed(-112324141.0/4294967296.0,1,-nbitq), 
to_sfixed(427272048.0/4294967296.0,1,-nbitq), 
to_sfixed(34092939.0/4294967296.0,1,-nbitq), 
to_sfixed(93370453.0/4294967296.0,1,-nbitq), 
to_sfixed(-886484601.0/4294967296.0,1,-nbitq), 
to_sfixed(476942902.0/4294967296.0,1,-nbitq), 
to_sfixed(314447359.0/4294967296.0,1,-nbitq), 
to_sfixed(146400548.0/4294967296.0,1,-nbitq), 
to_sfixed(314390072.0/4294967296.0,1,-nbitq), 
to_sfixed(-92730638.0/4294967296.0,1,-nbitq), 
to_sfixed(554904232.0/4294967296.0,1,-nbitq), 
to_sfixed(205890746.0/4294967296.0,1,-nbitq), 
to_sfixed(648089554.0/4294967296.0,1,-nbitq), 
to_sfixed(-414598707.0/4294967296.0,1,-nbitq), 
to_sfixed(-168346262.0/4294967296.0,1,-nbitq), 
to_sfixed(-355253511.0/4294967296.0,1,-nbitq), 
to_sfixed(-462823913.0/4294967296.0,1,-nbitq), 
to_sfixed(-155364681.0/4294967296.0,1,-nbitq), 
to_sfixed(-222491270.0/4294967296.0,1,-nbitq), 
to_sfixed(254297034.0/4294967296.0,1,-nbitq), 
to_sfixed(466396900.0/4294967296.0,1,-nbitq), 
to_sfixed(-215120561.0/4294967296.0,1,-nbitq), 
to_sfixed(12327345.0/4294967296.0,1,-nbitq), 
to_sfixed(-152062567.0/4294967296.0,1,-nbitq), 
to_sfixed(9162334.0/4294967296.0,1,-nbitq), 
to_sfixed(478904455.0/4294967296.0,1,-nbitq), 
to_sfixed(1336386110.0/4294967296.0,1,-nbitq), 
to_sfixed(782030130.0/4294967296.0,1,-nbitq), 
to_sfixed(463725710.0/4294967296.0,1,-nbitq), 
to_sfixed(-207087447.0/4294967296.0,1,-nbitq), 
to_sfixed(1119489317.0/4294967296.0,1,-nbitq), 
to_sfixed(213790894.0/4294967296.0,1,-nbitq), 
to_sfixed(485811923.0/4294967296.0,1,-nbitq), 
to_sfixed(246574030.0/4294967296.0,1,-nbitq), 
to_sfixed(-442362977.0/4294967296.0,1,-nbitq), 
to_sfixed(150880923.0/4294967296.0,1,-nbitq), 
to_sfixed(559884184.0/4294967296.0,1,-nbitq), 
to_sfixed(832953084.0/4294967296.0,1,-nbitq), 
to_sfixed(-406085842.0/4294967296.0,1,-nbitq), 
to_sfixed(353819678.0/4294967296.0,1,-nbitq), 
to_sfixed(-172243874.0/4294967296.0,1,-nbitq), 
to_sfixed(66555832.0/4294967296.0,1,-nbitq), 
to_sfixed(174090907.0/4294967296.0,1,-nbitq), 
to_sfixed(213249545.0/4294967296.0,1,-nbitq), 
to_sfixed(-326707288.0/4294967296.0,1,-nbitq), 
to_sfixed(32548699.0/4294967296.0,1,-nbitq), 
to_sfixed(-50094894.0/4294967296.0,1,-nbitq), 
to_sfixed(-28094452.0/4294967296.0,1,-nbitq), 
to_sfixed(71912361.0/4294967296.0,1,-nbitq), 
to_sfixed(-340308854.0/4294967296.0,1,-nbitq), 
to_sfixed(1878104400.0/4294967296.0,1,-nbitq), 
to_sfixed(169251959.0/4294967296.0,1,-nbitq), 
to_sfixed(-89598808.0/4294967296.0,1,-nbitq), 
to_sfixed(662167698.0/4294967296.0,1,-nbitq), 
to_sfixed(-248360396.0/4294967296.0,1,-nbitq), 
to_sfixed(401121977.0/4294967296.0,1,-nbitq), 
to_sfixed(376357482.0/4294967296.0,1,-nbitq), 
to_sfixed(131312702.0/4294967296.0,1,-nbitq), 
to_sfixed(816812020.0/4294967296.0,1,-nbitq), 
to_sfixed(-602024329.0/4294967296.0,1,-nbitq), 
to_sfixed(214392250.0/4294967296.0,1,-nbitq), 
to_sfixed(584694669.0/4294967296.0,1,-nbitq), 
to_sfixed(-392944038.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-207349245.0/4294967296.0,1,-nbitq), 
to_sfixed(585837790.0/4294967296.0,1,-nbitq), 
to_sfixed(-484403485.0/4294967296.0,1,-nbitq), 
to_sfixed(989781729.0/4294967296.0,1,-nbitq), 
to_sfixed(-473688585.0/4294967296.0,1,-nbitq), 
to_sfixed(-217526199.0/4294967296.0,1,-nbitq), 
to_sfixed(-345787548.0/4294967296.0,1,-nbitq), 
to_sfixed(246360615.0/4294967296.0,1,-nbitq), 
to_sfixed(634169887.0/4294967296.0,1,-nbitq), 
to_sfixed(443629613.0/4294967296.0,1,-nbitq), 
to_sfixed(839055356.0/4294967296.0,1,-nbitq), 
to_sfixed(295953392.0/4294967296.0,1,-nbitq), 
to_sfixed(250574474.0/4294967296.0,1,-nbitq), 
to_sfixed(-141609823.0/4294967296.0,1,-nbitq), 
to_sfixed(-219963821.0/4294967296.0,1,-nbitq), 
to_sfixed(301899398.0/4294967296.0,1,-nbitq), 
to_sfixed(-239079727.0/4294967296.0,1,-nbitq), 
to_sfixed(77134061.0/4294967296.0,1,-nbitq), 
to_sfixed(-245047605.0/4294967296.0,1,-nbitq), 
to_sfixed(380906809.0/4294967296.0,1,-nbitq), 
to_sfixed(-21878267.0/4294967296.0,1,-nbitq), 
to_sfixed(5007007.0/4294967296.0,1,-nbitq), 
to_sfixed(381488929.0/4294967296.0,1,-nbitq), 
to_sfixed(72497452.0/4294967296.0,1,-nbitq), 
to_sfixed(-92810601.0/4294967296.0,1,-nbitq), 
to_sfixed(-197679065.0/4294967296.0,1,-nbitq), 
to_sfixed(-238753495.0/4294967296.0,1,-nbitq), 
to_sfixed(90566878.0/4294967296.0,1,-nbitq), 
to_sfixed(-520211715.0/4294967296.0,1,-nbitq), 
to_sfixed(258557918.0/4294967296.0,1,-nbitq), 
to_sfixed(56619109.0/4294967296.0,1,-nbitq), 
to_sfixed(-308738944.0/4294967296.0,1,-nbitq), 
to_sfixed(492804893.0/4294967296.0,1,-nbitq), 
to_sfixed(-557383273.0/4294967296.0,1,-nbitq), 
to_sfixed(199921117.0/4294967296.0,1,-nbitq), 
to_sfixed(296706947.0/4294967296.0,1,-nbitq), 
to_sfixed(276798434.0/4294967296.0,1,-nbitq), 
to_sfixed(239610399.0/4294967296.0,1,-nbitq), 
to_sfixed(-165385044.0/4294967296.0,1,-nbitq), 
to_sfixed(336915584.0/4294967296.0,1,-nbitq), 
to_sfixed(-380296043.0/4294967296.0,1,-nbitq), 
to_sfixed(188258182.0/4294967296.0,1,-nbitq), 
to_sfixed(554459845.0/4294967296.0,1,-nbitq), 
to_sfixed(638958564.0/4294967296.0,1,-nbitq), 
to_sfixed(578403078.0/4294967296.0,1,-nbitq), 
to_sfixed(1050195510.0/4294967296.0,1,-nbitq), 
to_sfixed(250308777.0/4294967296.0,1,-nbitq), 
to_sfixed(499464069.0/4294967296.0,1,-nbitq), 
to_sfixed(81157704.0/4294967296.0,1,-nbitq), 
to_sfixed(308377414.0/4294967296.0,1,-nbitq), 
to_sfixed(-45979464.0/4294967296.0,1,-nbitq), 
to_sfixed(-36901942.0/4294967296.0,1,-nbitq), 
to_sfixed(-22603573.0/4294967296.0,1,-nbitq), 
to_sfixed(149411095.0/4294967296.0,1,-nbitq), 
to_sfixed(902206503.0/4294967296.0,1,-nbitq), 
to_sfixed(-230247947.0/4294967296.0,1,-nbitq), 
to_sfixed(-207208723.0/4294967296.0,1,-nbitq), 
to_sfixed(68139144.0/4294967296.0,1,-nbitq), 
to_sfixed(284367105.0/4294967296.0,1,-nbitq), 
to_sfixed(270047307.0/4294967296.0,1,-nbitq), 
to_sfixed(-206698754.0/4294967296.0,1,-nbitq), 
to_sfixed(41808344.0/4294967296.0,1,-nbitq), 
to_sfixed(304472871.0/4294967296.0,1,-nbitq), 
to_sfixed(-460519967.0/4294967296.0,1,-nbitq), 
to_sfixed(375075784.0/4294967296.0,1,-nbitq), 
to_sfixed(-84604528.0/4294967296.0,1,-nbitq), 
to_sfixed(-786679799.0/4294967296.0,1,-nbitq), 
to_sfixed(1763069131.0/4294967296.0,1,-nbitq), 
to_sfixed(390579943.0/4294967296.0,1,-nbitq), 
to_sfixed(-104047528.0/4294967296.0,1,-nbitq), 
to_sfixed(490997729.0/4294967296.0,1,-nbitq), 
to_sfixed(-65547728.0/4294967296.0,1,-nbitq), 
to_sfixed(326923952.0/4294967296.0,1,-nbitq), 
to_sfixed(274622300.0/4294967296.0,1,-nbitq), 
to_sfixed(-17820685.0/4294967296.0,1,-nbitq), 
to_sfixed(532222375.0/4294967296.0,1,-nbitq), 
to_sfixed(-652090354.0/4294967296.0,1,-nbitq), 
to_sfixed(444260930.0/4294967296.0,1,-nbitq), 
to_sfixed(35911306.0/4294967296.0,1,-nbitq), 
to_sfixed(198655648.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(170461242.0/4294967296.0,1,-nbitq), 
to_sfixed(278542816.0/4294967296.0,1,-nbitq), 
to_sfixed(449261974.0/4294967296.0,1,-nbitq), 
to_sfixed(817700488.0/4294967296.0,1,-nbitq), 
to_sfixed(-573663581.0/4294967296.0,1,-nbitq), 
to_sfixed(881303214.0/4294967296.0,1,-nbitq), 
to_sfixed(100632108.0/4294967296.0,1,-nbitq), 
to_sfixed(223944200.0/4294967296.0,1,-nbitq), 
to_sfixed(285139998.0/4294967296.0,1,-nbitq), 
to_sfixed(-146192500.0/4294967296.0,1,-nbitq), 
to_sfixed(36394273.0/4294967296.0,1,-nbitq), 
to_sfixed(584744655.0/4294967296.0,1,-nbitq), 
to_sfixed(88400783.0/4294967296.0,1,-nbitq), 
to_sfixed(-167334434.0/4294967296.0,1,-nbitq), 
to_sfixed(-84456723.0/4294967296.0,1,-nbitq), 
to_sfixed(-91470511.0/4294967296.0,1,-nbitq), 
to_sfixed(70228975.0/4294967296.0,1,-nbitq), 
to_sfixed(-314579707.0/4294967296.0,1,-nbitq), 
to_sfixed(761048304.0/4294967296.0,1,-nbitq), 
to_sfixed(-197006454.0/4294967296.0,1,-nbitq), 
to_sfixed(-75927786.0/4294967296.0,1,-nbitq), 
to_sfixed(-124909438.0/4294967296.0,1,-nbitq), 
to_sfixed(601934953.0/4294967296.0,1,-nbitq), 
to_sfixed(38881618.0/4294967296.0,1,-nbitq), 
to_sfixed(369340337.0/4294967296.0,1,-nbitq), 
to_sfixed(293255919.0/4294967296.0,1,-nbitq), 
to_sfixed(-90223417.0/4294967296.0,1,-nbitq), 
to_sfixed(738941947.0/4294967296.0,1,-nbitq), 
to_sfixed(-521967438.0/4294967296.0,1,-nbitq), 
to_sfixed(-216832240.0/4294967296.0,1,-nbitq), 
to_sfixed(-167854143.0/4294967296.0,1,-nbitq), 
to_sfixed(-95237671.0/4294967296.0,1,-nbitq), 
to_sfixed(-229144641.0/4294967296.0,1,-nbitq), 
to_sfixed(-531754260.0/4294967296.0,1,-nbitq), 
to_sfixed(507626179.0/4294967296.0,1,-nbitq), 
to_sfixed(498724913.0/4294967296.0,1,-nbitq), 
to_sfixed(483986215.0/4294967296.0,1,-nbitq), 
to_sfixed(-110183487.0/4294967296.0,1,-nbitq), 
to_sfixed(-383017920.0/4294967296.0,1,-nbitq), 
to_sfixed(245274917.0/4294967296.0,1,-nbitq), 
to_sfixed(78528444.0/4294967296.0,1,-nbitq), 
to_sfixed(764375619.0/4294967296.0,1,-nbitq), 
to_sfixed(817352992.0/4294967296.0,1,-nbitq), 
to_sfixed(1131250887.0/4294967296.0,1,-nbitq), 
to_sfixed(634755531.0/4294967296.0,1,-nbitq), 
to_sfixed(538829200.0/4294967296.0,1,-nbitq), 
to_sfixed(-188892133.0/4294967296.0,1,-nbitq), 
to_sfixed(171031953.0/4294967296.0,1,-nbitq), 
to_sfixed(-142093904.0/4294967296.0,1,-nbitq), 
to_sfixed(315510534.0/4294967296.0,1,-nbitq), 
to_sfixed(372045952.0/4294967296.0,1,-nbitq), 
to_sfixed(78296068.0/4294967296.0,1,-nbitq), 
to_sfixed(-573856122.0/4294967296.0,1,-nbitq), 
to_sfixed(160126616.0/4294967296.0,1,-nbitq), 
to_sfixed(61699724.0/4294967296.0,1,-nbitq), 
to_sfixed(96955776.0/4294967296.0,1,-nbitq), 
to_sfixed(-946968955.0/4294967296.0,1,-nbitq), 
to_sfixed(250460975.0/4294967296.0,1,-nbitq), 
to_sfixed(291576988.0/4294967296.0,1,-nbitq), 
to_sfixed(141159997.0/4294967296.0,1,-nbitq), 
to_sfixed(284705199.0/4294967296.0,1,-nbitq), 
to_sfixed(-287693123.0/4294967296.0,1,-nbitq), 
to_sfixed(326200834.0/4294967296.0,1,-nbitq), 
to_sfixed(-391445076.0/4294967296.0,1,-nbitq), 
to_sfixed(206547471.0/4294967296.0,1,-nbitq), 
to_sfixed(178437158.0/4294967296.0,1,-nbitq), 
to_sfixed(-231893437.0/4294967296.0,1,-nbitq), 
to_sfixed(1182988694.0/4294967296.0,1,-nbitq), 
to_sfixed(312014257.0/4294967296.0,1,-nbitq), 
to_sfixed(-177254732.0/4294967296.0,1,-nbitq), 
to_sfixed(227577237.0/4294967296.0,1,-nbitq), 
to_sfixed(174484307.0/4294967296.0,1,-nbitq), 
to_sfixed(-592291675.0/4294967296.0,1,-nbitq), 
to_sfixed(-137463574.0/4294967296.0,1,-nbitq), 
to_sfixed(157587518.0/4294967296.0,1,-nbitq), 
to_sfixed(170423893.0/4294967296.0,1,-nbitq), 
to_sfixed(-327200202.0/4294967296.0,1,-nbitq), 
to_sfixed(146870488.0/4294967296.0,1,-nbitq), 
to_sfixed(72257225.0/4294967296.0,1,-nbitq), 
to_sfixed(188909640.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-346191140.0/4294967296.0,1,-nbitq), 
to_sfixed(231793905.0/4294967296.0,1,-nbitq), 
to_sfixed(-31266556.0/4294967296.0,1,-nbitq), 
to_sfixed(629217959.0/4294967296.0,1,-nbitq), 
to_sfixed(-597285157.0/4294967296.0,1,-nbitq), 
to_sfixed(547008890.0/4294967296.0,1,-nbitq), 
to_sfixed(138540093.0/4294967296.0,1,-nbitq), 
to_sfixed(-46228053.0/4294967296.0,1,-nbitq), 
to_sfixed(-395940857.0/4294967296.0,1,-nbitq), 
to_sfixed(204553738.0/4294967296.0,1,-nbitq), 
to_sfixed(257492338.0/4294967296.0,1,-nbitq), 
to_sfixed(183185573.0/4294967296.0,1,-nbitq), 
to_sfixed(-212969337.0/4294967296.0,1,-nbitq), 
to_sfixed(18457319.0/4294967296.0,1,-nbitq), 
to_sfixed(-187389795.0/4294967296.0,1,-nbitq), 
to_sfixed(68234689.0/4294967296.0,1,-nbitq), 
to_sfixed(55751089.0/4294967296.0,1,-nbitq), 
to_sfixed(94149153.0/4294967296.0,1,-nbitq), 
to_sfixed(983173061.0/4294967296.0,1,-nbitq), 
to_sfixed(267173606.0/4294967296.0,1,-nbitq), 
to_sfixed(131827989.0/4294967296.0,1,-nbitq), 
to_sfixed(726819677.0/4294967296.0,1,-nbitq), 
to_sfixed(293793732.0/4294967296.0,1,-nbitq), 
to_sfixed(-140176188.0/4294967296.0,1,-nbitq), 
to_sfixed(421614856.0/4294967296.0,1,-nbitq), 
to_sfixed(351810453.0/4294967296.0,1,-nbitq), 
to_sfixed(-515859957.0/4294967296.0,1,-nbitq), 
to_sfixed(227972283.0/4294967296.0,1,-nbitq), 
to_sfixed(-318398808.0/4294967296.0,1,-nbitq), 
to_sfixed(-85880032.0/4294967296.0,1,-nbitq), 
to_sfixed(257566734.0/4294967296.0,1,-nbitq), 
to_sfixed(-612098728.0/4294967296.0,1,-nbitq), 
to_sfixed(-150055353.0/4294967296.0,1,-nbitq), 
to_sfixed(-653479179.0/4294967296.0,1,-nbitq), 
to_sfixed(321006499.0/4294967296.0,1,-nbitq), 
to_sfixed(325377234.0/4294967296.0,1,-nbitq), 
to_sfixed(186480113.0/4294967296.0,1,-nbitq), 
to_sfixed(113697557.0/4294967296.0,1,-nbitq), 
to_sfixed(291263220.0/4294967296.0,1,-nbitq), 
to_sfixed(-273992804.0/4294967296.0,1,-nbitq), 
to_sfixed(-381516312.0/4294967296.0,1,-nbitq), 
to_sfixed(722049344.0/4294967296.0,1,-nbitq), 
to_sfixed(274148775.0/4294967296.0,1,-nbitq), 
to_sfixed(691487767.0/4294967296.0,1,-nbitq), 
to_sfixed(93418454.0/4294967296.0,1,-nbitq), 
to_sfixed(421519953.0/4294967296.0,1,-nbitq), 
to_sfixed(189097558.0/4294967296.0,1,-nbitq), 
to_sfixed(-271820873.0/4294967296.0,1,-nbitq), 
to_sfixed(9475796.0/4294967296.0,1,-nbitq), 
to_sfixed(-216301208.0/4294967296.0,1,-nbitq), 
to_sfixed(70030138.0/4294967296.0,1,-nbitq), 
to_sfixed(-169858882.0/4294967296.0,1,-nbitq), 
to_sfixed(-331403089.0/4294967296.0,1,-nbitq), 
to_sfixed(539997340.0/4294967296.0,1,-nbitq), 
to_sfixed(-349502655.0/4294967296.0,1,-nbitq), 
to_sfixed(332176630.0/4294967296.0,1,-nbitq), 
to_sfixed(-221287287.0/4294967296.0,1,-nbitq), 
to_sfixed(-222227012.0/4294967296.0,1,-nbitq), 
to_sfixed(-266155547.0/4294967296.0,1,-nbitq), 
to_sfixed(376548429.0/4294967296.0,1,-nbitq), 
to_sfixed(74684415.0/4294967296.0,1,-nbitq), 
to_sfixed(286422560.0/4294967296.0,1,-nbitq), 
to_sfixed(-299019903.0/4294967296.0,1,-nbitq), 
to_sfixed(336408826.0/4294967296.0,1,-nbitq), 
to_sfixed(107241717.0/4294967296.0,1,-nbitq), 
to_sfixed(-218797228.0/4294967296.0,1,-nbitq), 
to_sfixed(-689868454.0/4294967296.0,1,-nbitq), 
to_sfixed(415602560.0/4294967296.0,1,-nbitq), 
to_sfixed(79756972.0/4294967296.0,1,-nbitq), 
to_sfixed(-98443616.0/4294967296.0,1,-nbitq), 
to_sfixed(-51271932.0/4294967296.0,1,-nbitq), 
to_sfixed(-62238506.0/4294967296.0,1,-nbitq), 
to_sfixed(-892251411.0/4294967296.0,1,-nbitq), 
to_sfixed(-277361415.0/4294967296.0,1,-nbitq), 
to_sfixed(104259016.0/4294967296.0,1,-nbitq), 
to_sfixed(-23307053.0/4294967296.0,1,-nbitq), 
to_sfixed(-83288097.0/4294967296.0,1,-nbitq), 
to_sfixed(-42348537.0/4294967296.0,1,-nbitq), 
to_sfixed(218672432.0/4294967296.0,1,-nbitq), 
to_sfixed(-262725325.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-52509964.0/4294967296.0,1,-nbitq), 
to_sfixed(-47943233.0/4294967296.0,1,-nbitq), 
to_sfixed(248611915.0/4294967296.0,1,-nbitq), 
to_sfixed(-193475121.0/4294967296.0,1,-nbitq), 
to_sfixed(60265632.0/4294967296.0,1,-nbitq), 
to_sfixed(240115382.0/4294967296.0,1,-nbitq), 
to_sfixed(208619721.0/4294967296.0,1,-nbitq), 
to_sfixed(-101731005.0/4294967296.0,1,-nbitq), 
to_sfixed(-211548582.0/4294967296.0,1,-nbitq), 
to_sfixed(-325923750.0/4294967296.0,1,-nbitq), 
to_sfixed(-211107311.0/4294967296.0,1,-nbitq), 
to_sfixed(199467934.0/4294967296.0,1,-nbitq), 
to_sfixed(-519550792.0/4294967296.0,1,-nbitq), 
to_sfixed(269948117.0/4294967296.0,1,-nbitq), 
to_sfixed(-112782147.0/4294967296.0,1,-nbitq), 
to_sfixed(-78338828.0/4294967296.0,1,-nbitq), 
to_sfixed(-39179625.0/4294967296.0,1,-nbitq), 
to_sfixed(-104637520.0/4294967296.0,1,-nbitq), 
to_sfixed(526449295.0/4294967296.0,1,-nbitq), 
to_sfixed(-333446746.0/4294967296.0,1,-nbitq), 
to_sfixed(373290303.0/4294967296.0,1,-nbitq), 
to_sfixed(623613904.0/4294967296.0,1,-nbitq), 
to_sfixed(702231525.0/4294967296.0,1,-nbitq), 
to_sfixed(201675530.0/4294967296.0,1,-nbitq), 
to_sfixed(-240186213.0/4294967296.0,1,-nbitq), 
to_sfixed(471430611.0/4294967296.0,1,-nbitq), 
to_sfixed(62969608.0/4294967296.0,1,-nbitq), 
to_sfixed(381848222.0/4294967296.0,1,-nbitq), 
to_sfixed(-297055133.0/4294967296.0,1,-nbitq), 
to_sfixed(-169586701.0/4294967296.0,1,-nbitq), 
to_sfixed(26857781.0/4294967296.0,1,-nbitq), 
to_sfixed(-378424411.0/4294967296.0,1,-nbitq), 
to_sfixed(564854278.0/4294967296.0,1,-nbitq), 
to_sfixed(-153199593.0/4294967296.0,1,-nbitq), 
to_sfixed(72761176.0/4294967296.0,1,-nbitq), 
to_sfixed(291542625.0/4294967296.0,1,-nbitq), 
to_sfixed(-67497884.0/4294967296.0,1,-nbitq), 
to_sfixed(-500510907.0/4294967296.0,1,-nbitq), 
to_sfixed(12682314.0/4294967296.0,1,-nbitq), 
to_sfixed(110633293.0/4294967296.0,1,-nbitq), 
to_sfixed(-428406741.0/4294967296.0,1,-nbitq), 
to_sfixed(-43355136.0/4294967296.0,1,-nbitq), 
to_sfixed(515575327.0/4294967296.0,1,-nbitq), 
to_sfixed(-165085619.0/4294967296.0,1,-nbitq), 
to_sfixed(253771642.0/4294967296.0,1,-nbitq), 
to_sfixed(253812701.0/4294967296.0,1,-nbitq), 
to_sfixed(-4335950.0/4294967296.0,1,-nbitq), 
to_sfixed(-33768660.0/4294967296.0,1,-nbitq), 
to_sfixed(-12654517.0/4294967296.0,1,-nbitq), 
to_sfixed(241612681.0/4294967296.0,1,-nbitq), 
to_sfixed(466415703.0/4294967296.0,1,-nbitq), 
to_sfixed(258579234.0/4294967296.0,1,-nbitq), 
to_sfixed(148495323.0/4294967296.0,1,-nbitq), 
to_sfixed(558474456.0/4294967296.0,1,-nbitq), 
to_sfixed(-212746931.0/4294967296.0,1,-nbitq), 
to_sfixed(419362986.0/4294967296.0,1,-nbitq), 
to_sfixed(-309699350.0/4294967296.0,1,-nbitq), 
to_sfixed(-171093023.0/4294967296.0,1,-nbitq), 
to_sfixed(373437785.0/4294967296.0,1,-nbitq), 
to_sfixed(156823204.0/4294967296.0,1,-nbitq), 
to_sfixed(387050497.0/4294967296.0,1,-nbitq), 
to_sfixed(160118495.0/4294967296.0,1,-nbitq), 
to_sfixed(-19133369.0/4294967296.0,1,-nbitq), 
to_sfixed(32476636.0/4294967296.0,1,-nbitq), 
to_sfixed(334819388.0/4294967296.0,1,-nbitq), 
to_sfixed(329234959.0/4294967296.0,1,-nbitq), 
to_sfixed(41547277.0/4294967296.0,1,-nbitq), 
to_sfixed(351683769.0/4294967296.0,1,-nbitq), 
to_sfixed(-97166541.0/4294967296.0,1,-nbitq), 
to_sfixed(-389355713.0/4294967296.0,1,-nbitq), 
to_sfixed(58033419.0/4294967296.0,1,-nbitq), 
to_sfixed(459044515.0/4294967296.0,1,-nbitq), 
to_sfixed(-211716484.0/4294967296.0,1,-nbitq), 
to_sfixed(-259958659.0/4294967296.0,1,-nbitq), 
to_sfixed(165404469.0/4294967296.0,1,-nbitq), 
to_sfixed(155673419.0/4294967296.0,1,-nbitq), 
to_sfixed(-43412608.0/4294967296.0,1,-nbitq), 
to_sfixed(270682209.0/4294967296.0,1,-nbitq), 
to_sfixed(215673193.0/4294967296.0,1,-nbitq), 
to_sfixed(-207709542.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-64766151.0/4294967296.0,1,-nbitq), 
to_sfixed(-270626941.0/4294967296.0,1,-nbitq), 
to_sfixed(612582648.0/4294967296.0,1,-nbitq), 
to_sfixed(149996648.0/4294967296.0,1,-nbitq), 
to_sfixed(-176643344.0/4294967296.0,1,-nbitq), 
to_sfixed(671858308.0/4294967296.0,1,-nbitq), 
to_sfixed(-229248282.0/4294967296.0,1,-nbitq), 
to_sfixed(-200447909.0/4294967296.0,1,-nbitq), 
to_sfixed(-509694730.0/4294967296.0,1,-nbitq), 
to_sfixed(302634039.0/4294967296.0,1,-nbitq), 
to_sfixed(-224072619.0/4294967296.0,1,-nbitq), 
to_sfixed(390760016.0/4294967296.0,1,-nbitq), 
to_sfixed(152679131.0/4294967296.0,1,-nbitq), 
to_sfixed(470754911.0/4294967296.0,1,-nbitq), 
to_sfixed(103505245.0/4294967296.0,1,-nbitq), 
to_sfixed(298844553.0/4294967296.0,1,-nbitq), 
to_sfixed(-109804487.0/4294967296.0,1,-nbitq), 
to_sfixed(-218331923.0/4294967296.0,1,-nbitq), 
to_sfixed(392957221.0/4294967296.0,1,-nbitq), 
to_sfixed(-229879238.0/4294967296.0,1,-nbitq), 
to_sfixed(-30486084.0/4294967296.0,1,-nbitq), 
to_sfixed(7021274.0/4294967296.0,1,-nbitq), 
to_sfixed(169487280.0/4294967296.0,1,-nbitq), 
to_sfixed(-355918696.0/4294967296.0,1,-nbitq), 
to_sfixed(-266639569.0/4294967296.0,1,-nbitq), 
to_sfixed(-1329434.0/4294967296.0,1,-nbitq), 
to_sfixed(342931358.0/4294967296.0,1,-nbitq), 
to_sfixed(-28936583.0/4294967296.0,1,-nbitq), 
to_sfixed(-153979563.0/4294967296.0,1,-nbitq), 
to_sfixed(32312221.0/4294967296.0,1,-nbitq), 
to_sfixed(-97561144.0/4294967296.0,1,-nbitq), 
to_sfixed(171399248.0/4294967296.0,1,-nbitq), 
to_sfixed(559198212.0/4294967296.0,1,-nbitq), 
to_sfixed(198343247.0/4294967296.0,1,-nbitq), 
to_sfixed(120248865.0/4294967296.0,1,-nbitq), 
to_sfixed(244652026.0/4294967296.0,1,-nbitq), 
to_sfixed(47379793.0/4294967296.0,1,-nbitq), 
to_sfixed(-290096492.0/4294967296.0,1,-nbitq), 
to_sfixed(-378985806.0/4294967296.0,1,-nbitq), 
to_sfixed(365447957.0/4294967296.0,1,-nbitq), 
to_sfixed(-346620928.0/4294967296.0,1,-nbitq), 
to_sfixed(235487420.0/4294967296.0,1,-nbitq), 
to_sfixed(502097699.0/4294967296.0,1,-nbitq), 
to_sfixed(155628071.0/4294967296.0,1,-nbitq), 
to_sfixed(331765438.0/4294967296.0,1,-nbitq), 
to_sfixed(-381497604.0/4294967296.0,1,-nbitq), 
to_sfixed(-380206607.0/4294967296.0,1,-nbitq), 
to_sfixed(-376803602.0/4294967296.0,1,-nbitq), 
to_sfixed(5026419.0/4294967296.0,1,-nbitq), 
to_sfixed(-58910619.0/4294967296.0,1,-nbitq), 
to_sfixed(-258787257.0/4294967296.0,1,-nbitq), 
to_sfixed(-16530226.0/4294967296.0,1,-nbitq), 
to_sfixed(-148166026.0/4294967296.0,1,-nbitq), 
to_sfixed(85399113.0/4294967296.0,1,-nbitq), 
to_sfixed(63677347.0/4294967296.0,1,-nbitq), 
to_sfixed(-60609764.0/4294967296.0,1,-nbitq), 
to_sfixed(-93382616.0/4294967296.0,1,-nbitq), 
to_sfixed(9115352.0/4294967296.0,1,-nbitq), 
to_sfixed(-188687048.0/4294967296.0,1,-nbitq), 
to_sfixed(-124380418.0/4294967296.0,1,-nbitq), 
to_sfixed(-52383905.0/4294967296.0,1,-nbitq), 
to_sfixed(64855660.0/4294967296.0,1,-nbitq), 
to_sfixed(-76436680.0/4294967296.0,1,-nbitq), 
to_sfixed(-52724111.0/4294967296.0,1,-nbitq), 
to_sfixed(139234790.0/4294967296.0,1,-nbitq), 
to_sfixed(18022393.0/4294967296.0,1,-nbitq), 
to_sfixed(442321894.0/4294967296.0,1,-nbitq), 
to_sfixed(-486086083.0/4294967296.0,1,-nbitq), 
to_sfixed(-328909342.0/4294967296.0,1,-nbitq), 
to_sfixed(513592359.0/4294967296.0,1,-nbitq), 
to_sfixed(174640576.0/4294967296.0,1,-nbitq), 
to_sfixed(-257985950.0/4294967296.0,1,-nbitq), 
to_sfixed(-749330522.0/4294967296.0,1,-nbitq), 
to_sfixed(395100989.0/4294967296.0,1,-nbitq), 
to_sfixed(-259442736.0/4294967296.0,1,-nbitq), 
to_sfixed(-311242812.0/4294967296.0,1,-nbitq), 
to_sfixed(-238332925.0/4294967296.0,1,-nbitq), 
to_sfixed(-58549195.0/4294967296.0,1,-nbitq), 
to_sfixed(-211889661.0/4294967296.0,1,-nbitq), 
to_sfixed(-30403948.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-382278827.0/4294967296.0,1,-nbitq), 
to_sfixed(-324799736.0/4294967296.0,1,-nbitq), 
to_sfixed(-107608303.0/4294967296.0,1,-nbitq), 
to_sfixed(78387703.0/4294967296.0,1,-nbitq), 
to_sfixed(-254112770.0/4294967296.0,1,-nbitq), 
to_sfixed(176239601.0/4294967296.0,1,-nbitq), 
to_sfixed(194902935.0/4294967296.0,1,-nbitq), 
to_sfixed(260236092.0/4294967296.0,1,-nbitq), 
to_sfixed(-29090253.0/4294967296.0,1,-nbitq), 
to_sfixed(60448419.0/4294967296.0,1,-nbitq), 
to_sfixed(349206980.0/4294967296.0,1,-nbitq), 
to_sfixed(-154163052.0/4294967296.0,1,-nbitq), 
to_sfixed(57037161.0/4294967296.0,1,-nbitq), 
to_sfixed(38608782.0/4294967296.0,1,-nbitq), 
to_sfixed(-320727103.0/4294967296.0,1,-nbitq), 
to_sfixed(454424722.0/4294967296.0,1,-nbitq), 
to_sfixed(-169633314.0/4294967296.0,1,-nbitq), 
to_sfixed(243481316.0/4294967296.0,1,-nbitq), 
to_sfixed(85738962.0/4294967296.0,1,-nbitq), 
to_sfixed(-69236412.0/4294967296.0,1,-nbitq), 
to_sfixed(-332816763.0/4294967296.0,1,-nbitq), 
to_sfixed(541696510.0/4294967296.0,1,-nbitq), 
to_sfixed(338354639.0/4294967296.0,1,-nbitq), 
to_sfixed(-80259971.0/4294967296.0,1,-nbitq), 
to_sfixed(-93466758.0/4294967296.0,1,-nbitq), 
to_sfixed(191835927.0/4294967296.0,1,-nbitq), 
to_sfixed(-380574839.0/4294967296.0,1,-nbitq), 
to_sfixed(-107180557.0/4294967296.0,1,-nbitq), 
to_sfixed(154273917.0/4294967296.0,1,-nbitq), 
to_sfixed(-54479384.0/4294967296.0,1,-nbitq), 
to_sfixed(-25458689.0/4294967296.0,1,-nbitq), 
to_sfixed(-92489467.0/4294967296.0,1,-nbitq), 
to_sfixed(274579520.0/4294967296.0,1,-nbitq), 
to_sfixed(152426733.0/4294967296.0,1,-nbitq), 
to_sfixed(288739948.0/4294967296.0,1,-nbitq), 
to_sfixed(383323384.0/4294967296.0,1,-nbitq), 
to_sfixed(-266077669.0/4294967296.0,1,-nbitq), 
to_sfixed(-292241415.0/4294967296.0,1,-nbitq), 
to_sfixed(195280756.0/4294967296.0,1,-nbitq), 
to_sfixed(137620137.0/4294967296.0,1,-nbitq), 
to_sfixed(-397510794.0/4294967296.0,1,-nbitq), 
to_sfixed(73690174.0/4294967296.0,1,-nbitq), 
to_sfixed(-2284887.0/4294967296.0,1,-nbitq), 
to_sfixed(45688517.0/4294967296.0,1,-nbitq), 
to_sfixed(-31823174.0/4294967296.0,1,-nbitq), 
to_sfixed(331942510.0/4294967296.0,1,-nbitq), 
to_sfixed(158535484.0/4294967296.0,1,-nbitq), 
to_sfixed(155824713.0/4294967296.0,1,-nbitq), 
to_sfixed(-82840309.0/4294967296.0,1,-nbitq), 
to_sfixed(-300312257.0/4294967296.0,1,-nbitq), 
to_sfixed(429154009.0/4294967296.0,1,-nbitq), 
to_sfixed(-216005953.0/4294967296.0,1,-nbitq), 
to_sfixed(-616666453.0/4294967296.0,1,-nbitq), 
to_sfixed(3976491.0/4294967296.0,1,-nbitq), 
to_sfixed(-55346036.0/4294967296.0,1,-nbitq), 
to_sfixed(12533555.0/4294967296.0,1,-nbitq), 
to_sfixed(-199947593.0/4294967296.0,1,-nbitq), 
to_sfixed(-28641687.0/4294967296.0,1,-nbitq), 
to_sfixed(295940034.0/4294967296.0,1,-nbitq), 
to_sfixed(145915543.0/4294967296.0,1,-nbitq), 
to_sfixed(19802880.0/4294967296.0,1,-nbitq), 
to_sfixed(179276669.0/4294967296.0,1,-nbitq), 
to_sfixed(-448932795.0/4294967296.0,1,-nbitq), 
to_sfixed(-202322992.0/4294967296.0,1,-nbitq), 
to_sfixed(-64321816.0/4294967296.0,1,-nbitq), 
to_sfixed(85717880.0/4294967296.0,1,-nbitq), 
to_sfixed(203975077.0/4294967296.0,1,-nbitq), 
to_sfixed(-282891464.0/4294967296.0,1,-nbitq), 
to_sfixed(-3223321.0/4294967296.0,1,-nbitq), 
to_sfixed(327768193.0/4294967296.0,1,-nbitq), 
to_sfixed(290553516.0/4294967296.0,1,-nbitq), 
to_sfixed(407620049.0/4294967296.0,1,-nbitq), 
to_sfixed(-313773371.0/4294967296.0,1,-nbitq), 
to_sfixed(293868516.0/4294967296.0,1,-nbitq), 
to_sfixed(88440986.0/4294967296.0,1,-nbitq), 
to_sfixed(-376310393.0/4294967296.0,1,-nbitq), 
to_sfixed(152355558.0/4294967296.0,1,-nbitq), 
to_sfixed(-167635180.0/4294967296.0,1,-nbitq), 
to_sfixed(236093466.0/4294967296.0,1,-nbitq), 
to_sfixed(-245036412.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-44608319.0/4294967296.0,1,-nbitq), 
to_sfixed(-156550840.0/4294967296.0,1,-nbitq), 
to_sfixed(302568602.0/4294967296.0,1,-nbitq), 
to_sfixed(-355948731.0/4294967296.0,1,-nbitq), 
to_sfixed(-126208252.0/4294967296.0,1,-nbitq), 
to_sfixed(-21386310.0/4294967296.0,1,-nbitq), 
to_sfixed(-44077125.0/4294967296.0,1,-nbitq), 
to_sfixed(35357152.0/4294967296.0,1,-nbitq), 
to_sfixed(196490747.0/4294967296.0,1,-nbitq), 
to_sfixed(209326487.0/4294967296.0,1,-nbitq), 
to_sfixed(171148514.0/4294967296.0,1,-nbitq), 
to_sfixed(351665712.0/4294967296.0,1,-nbitq), 
to_sfixed(48829487.0/4294967296.0,1,-nbitq), 
to_sfixed(294590824.0/4294967296.0,1,-nbitq), 
to_sfixed(241488085.0/4294967296.0,1,-nbitq), 
to_sfixed(-154807083.0/4294967296.0,1,-nbitq), 
to_sfixed(-44160900.0/4294967296.0,1,-nbitq), 
to_sfixed(-162579945.0/4294967296.0,1,-nbitq), 
to_sfixed(-69748748.0/4294967296.0,1,-nbitq), 
to_sfixed(57483825.0/4294967296.0,1,-nbitq), 
to_sfixed(-279883262.0/4294967296.0,1,-nbitq), 
to_sfixed(434963316.0/4294967296.0,1,-nbitq), 
to_sfixed(250594086.0/4294967296.0,1,-nbitq), 
to_sfixed(-118595148.0/4294967296.0,1,-nbitq), 
to_sfixed(-11026806.0/4294967296.0,1,-nbitq), 
to_sfixed(549878160.0/4294967296.0,1,-nbitq), 
to_sfixed(274406894.0/4294967296.0,1,-nbitq), 
to_sfixed(-284320795.0/4294967296.0,1,-nbitq), 
to_sfixed(60415537.0/4294967296.0,1,-nbitq), 
to_sfixed(93146289.0/4294967296.0,1,-nbitq), 
to_sfixed(-599902489.0/4294967296.0,1,-nbitq), 
to_sfixed(-154835013.0/4294967296.0,1,-nbitq), 
to_sfixed(-284981400.0/4294967296.0,1,-nbitq), 
to_sfixed(-345624739.0/4294967296.0,1,-nbitq), 
to_sfixed(-109401683.0/4294967296.0,1,-nbitq), 
to_sfixed(246301006.0/4294967296.0,1,-nbitq), 
to_sfixed(365710522.0/4294967296.0,1,-nbitq), 
to_sfixed(18394656.0/4294967296.0,1,-nbitq), 
to_sfixed(-125217724.0/4294967296.0,1,-nbitq), 
to_sfixed(336204188.0/4294967296.0,1,-nbitq), 
to_sfixed(-458144692.0/4294967296.0,1,-nbitq), 
to_sfixed(28055389.0/4294967296.0,1,-nbitq), 
to_sfixed(-70152040.0/4294967296.0,1,-nbitq), 
to_sfixed(329899060.0/4294967296.0,1,-nbitq), 
to_sfixed(215341617.0/4294967296.0,1,-nbitq), 
to_sfixed(364105589.0/4294967296.0,1,-nbitq), 
to_sfixed(153437060.0/4294967296.0,1,-nbitq), 
to_sfixed(-394640872.0/4294967296.0,1,-nbitq), 
to_sfixed(16142128.0/4294967296.0,1,-nbitq), 
to_sfixed(317341803.0/4294967296.0,1,-nbitq), 
to_sfixed(-89432104.0/4294967296.0,1,-nbitq), 
to_sfixed(-306104912.0/4294967296.0,1,-nbitq), 
to_sfixed(-3081509.0/4294967296.0,1,-nbitq), 
to_sfixed(450954410.0/4294967296.0,1,-nbitq), 
to_sfixed(349758719.0/4294967296.0,1,-nbitq), 
to_sfixed(-247250618.0/4294967296.0,1,-nbitq), 
to_sfixed(-321056325.0/4294967296.0,1,-nbitq), 
to_sfixed(-135965704.0/4294967296.0,1,-nbitq), 
to_sfixed(-188981067.0/4294967296.0,1,-nbitq), 
to_sfixed(120322421.0/4294967296.0,1,-nbitq), 
to_sfixed(-234258594.0/4294967296.0,1,-nbitq), 
to_sfixed(-248546608.0/4294967296.0,1,-nbitq), 
to_sfixed(-454092803.0/4294967296.0,1,-nbitq), 
to_sfixed(241210245.0/4294967296.0,1,-nbitq), 
to_sfixed(168975585.0/4294967296.0,1,-nbitq), 
to_sfixed(292057103.0/4294967296.0,1,-nbitq), 
to_sfixed(583197095.0/4294967296.0,1,-nbitq), 
to_sfixed(-123011028.0/4294967296.0,1,-nbitq), 
to_sfixed(-327062363.0/4294967296.0,1,-nbitq), 
to_sfixed(569353798.0/4294967296.0,1,-nbitq), 
to_sfixed(-434805559.0/4294967296.0,1,-nbitq), 
to_sfixed(186690875.0/4294967296.0,1,-nbitq), 
to_sfixed(-531890163.0/4294967296.0,1,-nbitq), 
to_sfixed(122440418.0/4294967296.0,1,-nbitq), 
to_sfixed(264356093.0/4294967296.0,1,-nbitq), 
to_sfixed(-53871546.0/4294967296.0,1,-nbitq), 
to_sfixed(105803201.0/4294967296.0,1,-nbitq), 
to_sfixed(112544149.0/4294967296.0,1,-nbitq), 
to_sfixed(-438679464.0/4294967296.0,1,-nbitq), 
to_sfixed(-280420689.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(202137801.0/4294967296.0,1,-nbitq), 
to_sfixed(-8183375.0/4294967296.0,1,-nbitq), 
to_sfixed(-329041496.0/4294967296.0,1,-nbitq), 
to_sfixed(-331114772.0/4294967296.0,1,-nbitq), 
to_sfixed(496129534.0/4294967296.0,1,-nbitq), 
to_sfixed(-321932764.0/4294967296.0,1,-nbitq), 
to_sfixed(-117422541.0/4294967296.0,1,-nbitq), 
to_sfixed(-256494666.0/4294967296.0,1,-nbitq), 
to_sfixed(-15207230.0/4294967296.0,1,-nbitq), 
to_sfixed(-312308122.0/4294967296.0,1,-nbitq), 
to_sfixed(236790314.0/4294967296.0,1,-nbitq), 
to_sfixed(-165805822.0/4294967296.0,1,-nbitq), 
to_sfixed(-145526938.0/4294967296.0,1,-nbitq), 
to_sfixed(-200792918.0/4294967296.0,1,-nbitq), 
to_sfixed(-260630797.0/4294967296.0,1,-nbitq), 
to_sfixed(-373899763.0/4294967296.0,1,-nbitq), 
to_sfixed(215034757.0/4294967296.0,1,-nbitq), 
to_sfixed(-354272878.0/4294967296.0,1,-nbitq), 
to_sfixed(57155404.0/4294967296.0,1,-nbitq), 
to_sfixed(-418218496.0/4294967296.0,1,-nbitq), 
to_sfixed(-120590509.0/4294967296.0,1,-nbitq), 
to_sfixed(-26161665.0/4294967296.0,1,-nbitq), 
to_sfixed(463141082.0/4294967296.0,1,-nbitq), 
to_sfixed(-322960155.0/4294967296.0,1,-nbitq), 
to_sfixed(325861688.0/4294967296.0,1,-nbitq), 
to_sfixed(521986349.0/4294967296.0,1,-nbitq), 
to_sfixed(-108690910.0/4294967296.0,1,-nbitq), 
to_sfixed(-345957559.0/4294967296.0,1,-nbitq), 
to_sfixed(-47955922.0/4294967296.0,1,-nbitq), 
to_sfixed(-230552226.0/4294967296.0,1,-nbitq), 
to_sfixed(-119877779.0/4294967296.0,1,-nbitq), 
to_sfixed(-21090005.0/4294967296.0,1,-nbitq), 
to_sfixed(176352995.0/4294967296.0,1,-nbitq), 
to_sfixed(-250486950.0/4294967296.0,1,-nbitq), 
to_sfixed(-168420278.0/4294967296.0,1,-nbitq), 
to_sfixed(-20372646.0/4294967296.0,1,-nbitq), 
to_sfixed(58519914.0/4294967296.0,1,-nbitq), 
to_sfixed(3731827.0/4294967296.0,1,-nbitq), 
to_sfixed(-371333238.0/4294967296.0,1,-nbitq), 
to_sfixed(260329738.0/4294967296.0,1,-nbitq), 
to_sfixed(233501045.0/4294967296.0,1,-nbitq), 
to_sfixed(147248020.0/4294967296.0,1,-nbitq), 
to_sfixed(-163311309.0/4294967296.0,1,-nbitq), 
to_sfixed(99276898.0/4294967296.0,1,-nbitq), 
to_sfixed(234721850.0/4294967296.0,1,-nbitq), 
to_sfixed(-235936080.0/4294967296.0,1,-nbitq), 
to_sfixed(15233460.0/4294967296.0,1,-nbitq), 
to_sfixed(-202021573.0/4294967296.0,1,-nbitq), 
to_sfixed(127514165.0/4294967296.0,1,-nbitq), 
to_sfixed(52680600.0/4294967296.0,1,-nbitq), 
to_sfixed(75047232.0/4294967296.0,1,-nbitq), 
to_sfixed(9644640.0/4294967296.0,1,-nbitq), 
to_sfixed(-79402930.0/4294967296.0,1,-nbitq), 
to_sfixed(212081673.0/4294967296.0,1,-nbitq), 
to_sfixed(-76243856.0/4294967296.0,1,-nbitq), 
to_sfixed(-81606093.0/4294967296.0,1,-nbitq), 
to_sfixed(-305233306.0/4294967296.0,1,-nbitq), 
to_sfixed(111246606.0/4294967296.0,1,-nbitq), 
to_sfixed(105758533.0/4294967296.0,1,-nbitq), 
to_sfixed(280287130.0/4294967296.0,1,-nbitq), 
to_sfixed(-264173672.0/4294967296.0,1,-nbitq), 
to_sfixed(458868810.0/4294967296.0,1,-nbitq), 
to_sfixed(242340095.0/4294967296.0,1,-nbitq), 
to_sfixed(-267668010.0/4294967296.0,1,-nbitq), 
to_sfixed(437756881.0/4294967296.0,1,-nbitq), 
to_sfixed(-94030405.0/4294967296.0,1,-nbitq), 
to_sfixed(326465647.0/4294967296.0,1,-nbitq), 
to_sfixed(-344314232.0/4294967296.0,1,-nbitq), 
to_sfixed(-262043454.0/4294967296.0,1,-nbitq), 
to_sfixed(-27306244.0/4294967296.0,1,-nbitq), 
to_sfixed(142007807.0/4294967296.0,1,-nbitq), 
to_sfixed(-104462890.0/4294967296.0,1,-nbitq), 
to_sfixed(-329999589.0/4294967296.0,1,-nbitq), 
to_sfixed(64845631.0/4294967296.0,1,-nbitq), 
to_sfixed(-198690743.0/4294967296.0,1,-nbitq), 
to_sfixed(92345731.0/4294967296.0,1,-nbitq), 
to_sfixed(149177277.0/4294967296.0,1,-nbitq), 
to_sfixed(-374123785.0/4294967296.0,1,-nbitq), 
to_sfixed(-7593044.0/4294967296.0,1,-nbitq), 
to_sfixed(381426623.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-240900154.0/4294967296.0,1,-nbitq), 
to_sfixed(-220055907.0/4294967296.0,1,-nbitq), 
to_sfixed(309397630.0/4294967296.0,1,-nbitq), 
to_sfixed(233613977.0/4294967296.0,1,-nbitq), 
to_sfixed(339838587.0/4294967296.0,1,-nbitq), 
to_sfixed(-338734781.0/4294967296.0,1,-nbitq), 
to_sfixed(369211715.0/4294967296.0,1,-nbitq), 
to_sfixed(-290200525.0/4294967296.0,1,-nbitq), 
to_sfixed(-317025964.0/4294967296.0,1,-nbitq), 
to_sfixed(-241935488.0/4294967296.0,1,-nbitq), 
to_sfixed(-263674062.0/4294967296.0,1,-nbitq), 
to_sfixed(514028317.0/4294967296.0,1,-nbitq), 
to_sfixed(-82599124.0/4294967296.0,1,-nbitq), 
to_sfixed(183181329.0/4294967296.0,1,-nbitq), 
to_sfixed(125638925.0/4294967296.0,1,-nbitq), 
to_sfixed(44557123.0/4294967296.0,1,-nbitq), 
to_sfixed(-213430839.0/4294967296.0,1,-nbitq), 
to_sfixed(341021967.0/4294967296.0,1,-nbitq), 
to_sfixed(-146302570.0/4294967296.0,1,-nbitq), 
to_sfixed(-420405252.0/4294967296.0,1,-nbitq), 
to_sfixed(-199819790.0/4294967296.0,1,-nbitq), 
to_sfixed(464368663.0/4294967296.0,1,-nbitq), 
to_sfixed(147471108.0/4294967296.0,1,-nbitq), 
to_sfixed(-334014565.0/4294967296.0,1,-nbitq), 
to_sfixed(-157887656.0/4294967296.0,1,-nbitq), 
to_sfixed(5649014.0/4294967296.0,1,-nbitq), 
to_sfixed(-67113209.0/4294967296.0,1,-nbitq), 
to_sfixed(-381302048.0/4294967296.0,1,-nbitq), 
to_sfixed(-252770438.0/4294967296.0,1,-nbitq), 
to_sfixed(-20429574.0/4294967296.0,1,-nbitq), 
to_sfixed(-489098595.0/4294967296.0,1,-nbitq), 
to_sfixed(-501681232.0/4294967296.0,1,-nbitq), 
to_sfixed(140087019.0/4294967296.0,1,-nbitq), 
to_sfixed(-488642685.0/4294967296.0,1,-nbitq), 
to_sfixed(462893522.0/4294967296.0,1,-nbitq), 
to_sfixed(329017365.0/4294967296.0,1,-nbitq), 
to_sfixed(7527470.0/4294967296.0,1,-nbitq), 
to_sfixed(-207590900.0/4294967296.0,1,-nbitq), 
to_sfixed(93333600.0/4294967296.0,1,-nbitq), 
to_sfixed(484873237.0/4294967296.0,1,-nbitq), 
to_sfixed(51733298.0/4294967296.0,1,-nbitq), 
to_sfixed(515416991.0/4294967296.0,1,-nbitq), 
to_sfixed(148807120.0/4294967296.0,1,-nbitq), 
to_sfixed(289668530.0/4294967296.0,1,-nbitq), 
to_sfixed(-314948412.0/4294967296.0,1,-nbitq), 
to_sfixed(263887403.0/4294967296.0,1,-nbitq), 
to_sfixed(-153719054.0/4294967296.0,1,-nbitq), 
to_sfixed(-28923006.0/4294967296.0,1,-nbitq), 
to_sfixed(-128164961.0/4294967296.0,1,-nbitq), 
to_sfixed(384456263.0/4294967296.0,1,-nbitq), 
to_sfixed(-253429344.0/4294967296.0,1,-nbitq), 
to_sfixed(25116131.0/4294967296.0,1,-nbitq), 
to_sfixed(-307224069.0/4294967296.0,1,-nbitq), 
to_sfixed(283255930.0/4294967296.0,1,-nbitq), 
to_sfixed(-203911900.0/4294967296.0,1,-nbitq), 
to_sfixed(175552812.0/4294967296.0,1,-nbitq), 
to_sfixed(-322860231.0/4294967296.0,1,-nbitq), 
to_sfixed(13060006.0/4294967296.0,1,-nbitq), 
to_sfixed(-46995411.0/4294967296.0,1,-nbitq), 
to_sfixed(-162137745.0/4294967296.0,1,-nbitq), 
to_sfixed(-267607019.0/4294967296.0,1,-nbitq), 
to_sfixed(389958030.0/4294967296.0,1,-nbitq), 
to_sfixed(-123992647.0/4294967296.0,1,-nbitq), 
to_sfixed(-33366554.0/4294967296.0,1,-nbitq), 
to_sfixed(-145738843.0/4294967296.0,1,-nbitq), 
to_sfixed(-115158838.0/4294967296.0,1,-nbitq), 
to_sfixed(721702965.0/4294967296.0,1,-nbitq), 
to_sfixed(-66169416.0/4294967296.0,1,-nbitq), 
to_sfixed(31924046.0/4294967296.0,1,-nbitq), 
to_sfixed(-131535265.0/4294967296.0,1,-nbitq), 
to_sfixed(44368619.0/4294967296.0,1,-nbitq), 
to_sfixed(-59829210.0/4294967296.0,1,-nbitq), 
to_sfixed(-355503598.0/4294967296.0,1,-nbitq), 
to_sfixed(-155047974.0/4294967296.0,1,-nbitq), 
to_sfixed(-21651318.0/4294967296.0,1,-nbitq), 
to_sfixed(-128844893.0/4294967296.0,1,-nbitq), 
to_sfixed(155707633.0/4294967296.0,1,-nbitq), 
to_sfixed(334884422.0/4294967296.0,1,-nbitq), 
to_sfixed(-591761727.0/4294967296.0,1,-nbitq), 
to_sfixed(204366164.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(190535618.0/4294967296.0,1,-nbitq), 
to_sfixed(-90019855.0/4294967296.0,1,-nbitq), 
to_sfixed(237150784.0/4294967296.0,1,-nbitq), 
to_sfixed(-26722979.0/4294967296.0,1,-nbitq), 
to_sfixed(-84502605.0/4294967296.0,1,-nbitq), 
to_sfixed(-116270334.0/4294967296.0,1,-nbitq), 
to_sfixed(495881503.0/4294967296.0,1,-nbitq), 
to_sfixed(17785331.0/4294967296.0,1,-nbitq), 
to_sfixed(180439310.0/4294967296.0,1,-nbitq), 
to_sfixed(384235143.0/4294967296.0,1,-nbitq), 
to_sfixed(315695460.0/4294967296.0,1,-nbitq), 
to_sfixed(460477883.0/4294967296.0,1,-nbitq), 
to_sfixed(-229383552.0/4294967296.0,1,-nbitq), 
to_sfixed(-129669417.0/4294967296.0,1,-nbitq), 
to_sfixed(-299395958.0/4294967296.0,1,-nbitq), 
to_sfixed(244600898.0/4294967296.0,1,-nbitq), 
to_sfixed(108283388.0/4294967296.0,1,-nbitq), 
to_sfixed(-119296642.0/4294967296.0,1,-nbitq), 
to_sfixed(-240278053.0/4294967296.0,1,-nbitq), 
to_sfixed(-314443786.0/4294967296.0,1,-nbitq), 
to_sfixed(6659550.0/4294967296.0,1,-nbitq), 
to_sfixed(150613727.0/4294967296.0,1,-nbitq), 
to_sfixed(-81196586.0/4294967296.0,1,-nbitq), 
to_sfixed(-194764323.0/4294967296.0,1,-nbitq), 
to_sfixed(-37696336.0/4294967296.0,1,-nbitq), 
to_sfixed(-370950901.0/4294967296.0,1,-nbitq), 
to_sfixed(-170856557.0/4294967296.0,1,-nbitq), 
to_sfixed(-328531249.0/4294967296.0,1,-nbitq), 
to_sfixed(336108308.0/4294967296.0,1,-nbitq), 
to_sfixed(310948924.0/4294967296.0,1,-nbitq), 
to_sfixed(-469923787.0/4294967296.0,1,-nbitq), 
to_sfixed(-274250476.0/4294967296.0,1,-nbitq), 
to_sfixed(35317877.0/4294967296.0,1,-nbitq), 
to_sfixed(-8445949.0/4294967296.0,1,-nbitq), 
to_sfixed(259178508.0/4294967296.0,1,-nbitq), 
to_sfixed(-91667446.0/4294967296.0,1,-nbitq), 
to_sfixed(501651939.0/4294967296.0,1,-nbitq), 
to_sfixed(1306878.0/4294967296.0,1,-nbitq), 
to_sfixed(-415897144.0/4294967296.0,1,-nbitq), 
to_sfixed(-109021152.0/4294967296.0,1,-nbitq), 
to_sfixed(-275265224.0/4294967296.0,1,-nbitq), 
to_sfixed(33668682.0/4294967296.0,1,-nbitq), 
to_sfixed(108004058.0/4294967296.0,1,-nbitq), 
to_sfixed(-178096908.0/4294967296.0,1,-nbitq), 
to_sfixed(4063902.0/4294967296.0,1,-nbitq), 
to_sfixed(155992205.0/4294967296.0,1,-nbitq), 
to_sfixed(-323970796.0/4294967296.0,1,-nbitq), 
to_sfixed(-164456321.0/4294967296.0,1,-nbitq), 
to_sfixed(-5243382.0/4294967296.0,1,-nbitq), 
to_sfixed(-47484743.0/4294967296.0,1,-nbitq), 
to_sfixed(346927488.0/4294967296.0,1,-nbitq), 
to_sfixed(358794129.0/4294967296.0,1,-nbitq), 
to_sfixed(-164152241.0/4294967296.0,1,-nbitq), 
to_sfixed(-1714145.0/4294967296.0,1,-nbitq), 
to_sfixed(313887018.0/4294967296.0,1,-nbitq), 
to_sfixed(-8504312.0/4294967296.0,1,-nbitq), 
to_sfixed(-62167004.0/4294967296.0,1,-nbitq), 
to_sfixed(-561441215.0/4294967296.0,1,-nbitq), 
to_sfixed(385708980.0/4294967296.0,1,-nbitq), 
to_sfixed(429279773.0/4294967296.0,1,-nbitq), 
to_sfixed(-81023774.0/4294967296.0,1,-nbitq), 
to_sfixed(-12852716.0/4294967296.0,1,-nbitq), 
to_sfixed(-560237937.0/4294967296.0,1,-nbitq), 
to_sfixed(365455784.0/4294967296.0,1,-nbitq), 
to_sfixed(-371753458.0/4294967296.0,1,-nbitq), 
to_sfixed(-381925177.0/4294967296.0,1,-nbitq), 
to_sfixed(57805032.0/4294967296.0,1,-nbitq), 
to_sfixed(42909647.0/4294967296.0,1,-nbitq), 
to_sfixed(337909087.0/4294967296.0,1,-nbitq), 
to_sfixed(143428846.0/4294967296.0,1,-nbitq), 
to_sfixed(165404826.0/4294967296.0,1,-nbitq), 
to_sfixed(264620355.0/4294967296.0,1,-nbitq), 
to_sfixed(-336005180.0/4294967296.0,1,-nbitq), 
to_sfixed(247871086.0/4294967296.0,1,-nbitq), 
to_sfixed(39692478.0/4294967296.0,1,-nbitq), 
to_sfixed(213329591.0/4294967296.0,1,-nbitq), 
to_sfixed(155388127.0/4294967296.0,1,-nbitq), 
to_sfixed(119045665.0/4294967296.0,1,-nbitq), 
to_sfixed(-530639032.0/4294967296.0,1,-nbitq), 
to_sfixed(89476060.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-213148446.0/4294967296.0,1,-nbitq), 
to_sfixed(-647251896.0/4294967296.0,1,-nbitq), 
to_sfixed(405107889.0/4294967296.0,1,-nbitq), 
to_sfixed(-309033823.0/4294967296.0,1,-nbitq), 
to_sfixed(221596470.0/4294967296.0,1,-nbitq), 
to_sfixed(89243418.0/4294967296.0,1,-nbitq), 
to_sfixed(164522387.0/4294967296.0,1,-nbitq), 
to_sfixed(-125054033.0/4294967296.0,1,-nbitq), 
to_sfixed(347205130.0/4294967296.0,1,-nbitq), 
to_sfixed(160940048.0/4294967296.0,1,-nbitq), 
to_sfixed(239847655.0/4294967296.0,1,-nbitq), 
to_sfixed(190577375.0/4294967296.0,1,-nbitq), 
to_sfixed(-367509668.0/4294967296.0,1,-nbitq), 
to_sfixed(-659077600.0/4294967296.0,1,-nbitq), 
to_sfixed(251633948.0/4294967296.0,1,-nbitq), 
to_sfixed(176527599.0/4294967296.0,1,-nbitq), 
to_sfixed(270933270.0/4294967296.0,1,-nbitq), 
to_sfixed(-128964788.0/4294967296.0,1,-nbitq), 
to_sfixed(-197428671.0/4294967296.0,1,-nbitq), 
to_sfixed(199840359.0/4294967296.0,1,-nbitq), 
to_sfixed(268500221.0/4294967296.0,1,-nbitq), 
to_sfixed(409048682.0/4294967296.0,1,-nbitq), 
to_sfixed(275818889.0/4294967296.0,1,-nbitq), 
to_sfixed(-564947163.0/4294967296.0,1,-nbitq), 
to_sfixed(165669921.0/4294967296.0,1,-nbitq), 
to_sfixed(405679062.0/4294967296.0,1,-nbitq), 
to_sfixed(132586883.0/4294967296.0,1,-nbitq), 
to_sfixed(-456337831.0/4294967296.0,1,-nbitq), 
to_sfixed(83698838.0/4294967296.0,1,-nbitq), 
to_sfixed(150793542.0/4294967296.0,1,-nbitq), 
to_sfixed(-179688403.0/4294967296.0,1,-nbitq), 
to_sfixed(-210229753.0/4294967296.0,1,-nbitq), 
to_sfixed(-98013443.0/4294967296.0,1,-nbitq), 
to_sfixed(-67303993.0/4294967296.0,1,-nbitq), 
to_sfixed(106735217.0/4294967296.0,1,-nbitq), 
to_sfixed(89677891.0/4294967296.0,1,-nbitq), 
to_sfixed(484251116.0/4294967296.0,1,-nbitq), 
to_sfixed(-224465631.0/4294967296.0,1,-nbitq), 
to_sfixed(-282368718.0/4294967296.0,1,-nbitq), 
to_sfixed(29261599.0/4294967296.0,1,-nbitq), 
to_sfixed(-132073700.0/4294967296.0,1,-nbitq), 
to_sfixed(-240452567.0/4294967296.0,1,-nbitq), 
to_sfixed(119021625.0/4294967296.0,1,-nbitq), 
to_sfixed(-76043851.0/4294967296.0,1,-nbitq), 
to_sfixed(-280691154.0/4294967296.0,1,-nbitq), 
to_sfixed(405553704.0/4294967296.0,1,-nbitq), 
to_sfixed(186019404.0/4294967296.0,1,-nbitq), 
to_sfixed(-174408489.0/4294967296.0,1,-nbitq), 
to_sfixed(-267258719.0/4294967296.0,1,-nbitq), 
to_sfixed(700149583.0/4294967296.0,1,-nbitq), 
to_sfixed(350940189.0/4294967296.0,1,-nbitq), 
to_sfixed(340693033.0/4294967296.0,1,-nbitq), 
to_sfixed(-15055977.0/4294967296.0,1,-nbitq), 
to_sfixed(179168256.0/4294967296.0,1,-nbitq), 
to_sfixed(429923047.0/4294967296.0,1,-nbitq), 
to_sfixed(1814956.0/4294967296.0,1,-nbitq), 
to_sfixed(-233825882.0/4294967296.0,1,-nbitq), 
to_sfixed(181634598.0/4294967296.0,1,-nbitq), 
to_sfixed(72876085.0/4294967296.0,1,-nbitq), 
to_sfixed(-253071523.0/4294967296.0,1,-nbitq), 
to_sfixed(-81071600.0/4294967296.0,1,-nbitq), 
to_sfixed(-250276665.0/4294967296.0,1,-nbitq), 
to_sfixed(-206210023.0/4294967296.0,1,-nbitq), 
to_sfixed(129859182.0/4294967296.0,1,-nbitq), 
to_sfixed(-254591488.0/4294967296.0,1,-nbitq), 
to_sfixed(-238860138.0/4294967296.0,1,-nbitq), 
to_sfixed(-59412474.0/4294967296.0,1,-nbitq), 
to_sfixed(-437248767.0/4294967296.0,1,-nbitq), 
to_sfixed(-193913123.0/4294967296.0,1,-nbitq), 
to_sfixed(-136316836.0/4294967296.0,1,-nbitq), 
to_sfixed(182012018.0/4294967296.0,1,-nbitq), 
to_sfixed(-19057356.0/4294967296.0,1,-nbitq), 
to_sfixed(-230838282.0/4294967296.0,1,-nbitq), 
to_sfixed(221042808.0/4294967296.0,1,-nbitq), 
to_sfixed(80219047.0/4294967296.0,1,-nbitq), 
to_sfixed(-400628413.0/4294967296.0,1,-nbitq), 
to_sfixed(332181868.0/4294967296.0,1,-nbitq), 
to_sfixed(25017893.0/4294967296.0,1,-nbitq), 
to_sfixed(-96570492.0/4294967296.0,1,-nbitq), 
to_sfixed(307723649.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-96501308.0/4294967296.0,1,-nbitq), 
to_sfixed(-138383361.0/4294967296.0,1,-nbitq), 
to_sfixed(337780833.0/4294967296.0,1,-nbitq), 
to_sfixed(-79730026.0/4294967296.0,1,-nbitq), 
to_sfixed(338616038.0/4294967296.0,1,-nbitq), 
to_sfixed(359196394.0/4294967296.0,1,-nbitq), 
to_sfixed(235932535.0/4294967296.0,1,-nbitq), 
to_sfixed(274300666.0/4294967296.0,1,-nbitq), 
to_sfixed(118406683.0/4294967296.0,1,-nbitq), 
to_sfixed(-111845565.0/4294967296.0,1,-nbitq), 
to_sfixed(144590597.0/4294967296.0,1,-nbitq), 
to_sfixed(649192798.0/4294967296.0,1,-nbitq), 
to_sfixed(-71316680.0/4294967296.0,1,-nbitq), 
to_sfixed(4819079.0/4294967296.0,1,-nbitq), 
to_sfixed(294141643.0/4294967296.0,1,-nbitq), 
to_sfixed(-93832301.0/4294967296.0,1,-nbitq), 
to_sfixed(-183284617.0/4294967296.0,1,-nbitq), 
to_sfixed(80110636.0/4294967296.0,1,-nbitq), 
to_sfixed(-570650637.0/4294967296.0,1,-nbitq), 
to_sfixed(356815281.0/4294967296.0,1,-nbitq), 
to_sfixed(-214479656.0/4294967296.0,1,-nbitq), 
to_sfixed(-226514685.0/4294967296.0,1,-nbitq), 
to_sfixed(447616364.0/4294967296.0,1,-nbitq), 
to_sfixed(-155981387.0/4294967296.0,1,-nbitq), 
to_sfixed(182971189.0/4294967296.0,1,-nbitq), 
to_sfixed(-158714126.0/4294967296.0,1,-nbitq), 
to_sfixed(-392535328.0/4294967296.0,1,-nbitq), 
to_sfixed(-130268717.0/4294967296.0,1,-nbitq), 
to_sfixed(-774340684.0/4294967296.0,1,-nbitq), 
to_sfixed(100044219.0/4294967296.0,1,-nbitq), 
to_sfixed(-167050610.0/4294967296.0,1,-nbitq), 
to_sfixed(-798587625.0/4294967296.0,1,-nbitq), 
to_sfixed(-28984040.0/4294967296.0,1,-nbitq), 
to_sfixed(-15251935.0/4294967296.0,1,-nbitq), 
to_sfixed(-211099926.0/4294967296.0,1,-nbitq), 
to_sfixed(-37534560.0/4294967296.0,1,-nbitq), 
to_sfixed(505651987.0/4294967296.0,1,-nbitq), 
to_sfixed(-260552635.0/4294967296.0,1,-nbitq), 
to_sfixed(-140420564.0/4294967296.0,1,-nbitq), 
to_sfixed(-61482660.0/4294967296.0,1,-nbitq), 
to_sfixed(-52775190.0/4294967296.0,1,-nbitq), 
to_sfixed(192458061.0/4294967296.0,1,-nbitq), 
to_sfixed(197933644.0/4294967296.0,1,-nbitq), 
to_sfixed(-306762150.0/4294967296.0,1,-nbitq), 
to_sfixed(-154166963.0/4294967296.0,1,-nbitq), 
to_sfixed(233585760.0/4294967296.0,1,-nbitq), 
to_sfixed(252532458.0/4294967296.0,1,-nbitq), 
to_sfixed(-306584028.0/4294967296.0,1,-nbitq), 
to_sfixed(142577978.0/4294967296.0,1,-nbitq), 
to_sfixed(-15068691.0/4294967296.0,1,-nbitq), 
to_sfixed(-114810430.0/4294967296.0,1,-nbitq), 
to_sfixed(-91535801.0/4294967296.0,1,-nbitq), 
to_sfixed(-45105229.0/4294967296.0,1,-nbitq), 
to_sfixed(259611877.0/4294967296.0,1,-nbitq), 
to_sfixed(133943599.0/4294967296.0,1,-nbitq), 
to_sfixed(512607615.0/4294967296.0,1,-nbitq), 
to_sfixed(22619699.0/4294967296.0,1,-nbitq), 
to_sfixed(-285924460.0/4294967296.0,1,-nbitq), 
to_sfixed(-1942819.0/4294967296.0,1,-nbitq), 
to_sfixed(-157535530.0/4294967296.0,1,-nbitq), 
to_sfixed(181756599.0/4294967296.0,1,-nbitq), 
to_sfixed(-149960082.0/4294967296.0,1,-nbitq), 
to_sfixed(-556696440.0/4294967296.0,1,-nbitq), 
to_sfixed(-278456531.0/4294967296.0,1,-nbitq), 
to_sfixed(141621058.0/4294967296.0,1,-nbitq), 
to_sfixed(84595897.0/4294967296.0,1,-nbitq), 
to_sfixed(-557958339.0/4294967296.0,1,-nbitq), 
to_sfixed(-86469633.0/4294967296.0,1,-nbitq), 
to_sfixed(402747432.0/4294967296.0,1,-nbitq), 
to_sfixed(403046285.0/4294967296.0,1,-nbitq), 
to_sfixed(207108877.0/4294967296.0,1,-nbitq), 
to_sfixed(42534891.0/4294967296.0,1,-nbitq), 
to_sfixed(314574048.0/4294967296.0,1,-nbitq), 
to_sfixed(291856281.0/4294967296.0,1,-nbitq), 
to_sfixed(-49214121.0/4294967296.0,1,-nbitq), 
to_sfixed(145269686.0/4294967296.0,1,-nbitq), 
to_sfixed(151326259.0/4294967296.0,1,-nbitq), 
to_sfixed(434536498.0/4294967296.0,1,-nbitq), 
to_sfixed(-520628755.0/4294967296.0,1,-nbitq), 
to_sfixed(-276635443.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(220544189.0/4294967296.0,1,-nbitq), 
to_sfixed(-522345312.0/4294967296.0,1,-nbitq), 
to_sfixed(519176928.0/4294967296.0,1,-nbitq), 
to_sfixed(-56594876.0/4294967296.0,1,-nbitq), 
to_sfixed(-43371268.0/4294967296.0,1,-nbitq), 
to_sfixed(258870356.0/4294967296.0,1,-nbitq), 
to_sfixed(360665953.0/4294967296.0,1,-nbitq), 
to_sfixed(-191289498.0/4294967296.0,1,-nbitq), 
to_sfixed(774174229.0/4294967296.0,1,-nbitq), 
to_sfixed(34364603.0/4294967296.0,1,-nbitq), 
to_sfixed(9940881.0/4294967296.0,1,-nbitq), 
to_sfixed(266002506.0/4294967296.0,1,-nbitq), 
to_sfixed(-77646305.0/4294967296.0,1,-nbitq), 
to_sfixed(-559275002.0/4294967296.0,1,-nbitq), 
to_sfixed(-417653130.0/4294967296.0,1,-nbitq), 
to_sfixed(-37786187.0/4294967296.0,1,-nbitq), 
to_sfixed(120225638.0/4294967296.0,1,-nbitq), 
to_sfixed(77423921.0/4294967296.0,1,-nbitq), 
to_sfixed(-386216666.0/4294967296.0,1,-nbitq), 
to_sfixed(417729240.0/4294967296.0,1,-nbitq), 
to_sfixed(73685081.0/4294967296.0,1,-nbitq), 
to_sfixed(563300257.0/4294967296.0,1,-nbitq), 
to_sfixed(593202837.0/4294967296.0,1,-nbitq), 
to_sfixed(-553239367.0/4294967296.0,1,-nbitq), 
to_sfixed(110864188.0/4294967296.0,1,-nbitq), 
to_sfixed(-539868439.0/4294967296.0,1,-nbitq), 
to_sfixed(139910018.0/4294967296.0,1,-nbitq), 
to_sfixed(459643287.0/4294967296.0,1,-nbitq), 
to_sfixed(83597696.0/4294967296.0,1,-nbitq), 
to_sfixed(31511098.0/4294967296.0,1,-nbitq), 
to_sfixed(19342495.0/4294967296.0,1,-nbitq), 
to_sfixed(-886723581.0/4294967296.0,1,-nbitq), 
to_sfixed(124327782.0/4294967296.0,1,-nbitq), 
to_sfixed(575224009.0/4294967296.0,1,-nbitq), 
to_sfixed(-73613924.0/4294967296.0,1,-nbitq), 
to_sfixed(-113111810.0/4294967296.0,1,-nbitq), 
to_sfixed(419589511.0/4294967296.0,1,-nbitq), 
to_sfixed(-677933550.0/4294967296.0,1,-nbitq), 
to_sfixed(-159644825.0/4294967296.0,1,-nbitq), 
to_sfixed(212631012.0/4294967296.0,1,-nbitq), 
to_sfixed(-36261708.0/4294967296.0,1,-nbitq), 
to_sfixed(-244163439.0/4294967296.0,1,-nbitq), 
to_sfixed(-138607676.0/4294967296.0,1,-nbitq), 
to_sfixed(-428463336.0/4294967296.0,1,-nbitq), 
to_sfixed(613318240.0/4294967296.0,1,-nbitq), 
to_sfixed(462672766.0/4294967296.0,1,-nbitq), 
to_sfixed(-16923334.0/4294967296.0,1,-nbitq), 
to_sfixed(238389279.0/4294967296.0,1,-nbitq), 
to_sfixed(-25938925.0/4294967296.0,1,-nbitq), 
to_sfixed(550670206.0/4294967296.0,1,-nbitq), 
to_sfixed(-155623830.0/4294967296.0,1,-nbitq), 
to_sfixed(665048398.0/4294967296.0,1,-nbitq), 
to_sfixed(-139557644.0/4294967296.0,1,-nbitq), 
to_sfixed(84684103.0/4294967296.0,1,-nbitq), 
to_sfixed(-798114909.0/4294967296.0,1,-nbitq), 
to_sfixed(830962540.0/4294967296.0,1,-nbitq), 
to_sfixed(419322551.0/4294967296.0,1,-nbitq), 
to_sfixed(83132054.0/4294967296.0,1,-nbitq), 
to_sfixed(255203858.0/4294967296.0,1,-nbitq), 
to_sfixed(45768030.0/4294967296.0,1,-nbitq), 
to_sfixed(-408917938.0/4294967296.0,1,-nbitq), 
to_sfixed(2214633.0/4294967296.0,1,-nbitq), 
to_sfixed(-396818501.0/4294967296.0,1,-nbitq), 
to_sfixed(36710591.0/4294967296.0,1,-nbitq), 
to_sfixed(-47512325.0/4294967296.0,1,-nbitq), 
to_sfixed(-339238818.0/4294967296.0,1,-nbitq), 
to_sfixed(-994621510.0/4294967296.0,1,-nbitq), 
to_sfixed(-121452504.0/4294967296.0,1,-nbitq), 
to_sfixed(-96413852.0/4294967296.0,1,-nbitq), 
to_sfixed(234801215.0/4294967296.0,1,-nbitq), 
to_sfixed(206608787.0/4294967296.0,1,-nbitq), 
to_sfixed(-472534847.0/4294967296.0,1,-nbitq), 
to_sfixed(406370299.0/4294967296.0,1,-nbitq), 
to_sfixed(200260805.0/4294967296.0,1,-nbitq), 
to_sfixed(494724157.0/4294967296.0,1,-nbitq), 
to_sfixed(103733271.0/4294967296.0,1,-nbitq), 
to_sfixed(620623725.0/4294967296.0,1,-nbitq), 
to_sfixed(-45317858.0/4294967296.0,1,-nbitq), 
to_sfixed(-506546019.0/4294967296.0,1,-nbitq), 
to_sfixed(-141185888.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-63993779.0/4294967296.0,1,-nbitq), 
to_sfixed(-583094897.0/4294967296.0,1,-nbitq), 
to_sfixed(-170063852.0/4294967296.0,1,-nbitq), 
to_sfixed(311336061.0/4294967296.0,1,-nbitq), 
to_sfixed(302587989.0/4294967296.0,1,-nbitq), 
to_sfixed(-429167208.0/4294967296.0,1,-nbitq), 
to_sfixed(-24772543.0/4294967296.0,1,-nbitq), 
to_sfixed(65255653.0/4294967296.0,1,-nbitq), 
to_sfixed(931462592.0/4294967296.0,1,-nbitq), 
to_sfixed(159956287.0/4294967296.0,1,-nbitq), 
to_sfixed(-188976541.0/4294967296.0,1,-nbitq), 
to_sfixed(634300718.0/4294967296.0,1,-nbitq), 
to_sfixed(-202236152.0/4294967296.0,1,-nbitq), 
to_sfixed(-703724118.0/4294967296.0,1,-nbitq), 
to_sfixed(4187693.0/4294967296.0,1,-nbitq), 
to_sfixed(418293557.0/4294967296.0,1,-nbitq), 
to_sfixed(-378800604.0/4294967296.0,1,-nbitq), 
to_sfixed(317166769.0/4294967296.0,1,-nbitq), 
to_sfixed(-540963233.0/4294967296.0,1,-nbitq), 
to_sfixed(277118397.0/4294967296.0,1,-nbitq), 
to_sfixed(314746342.0/4294967296.0,1,-nbitq), 
to_sfixed(581162445.0/4294967296.0,1,-nbitq), 
to_sfixed(202965175.0/4294967296.0,1,-nbitq), 
to_sfixed(-433127441.0/4294967296.0,1,-nbitq), 
to_sfixed(-111111824.0/4294967296.0,1,-nbitq), 
to_sfixed(-783037564.0/4294967296.0,1,-nbitq), 
to_sfixed(-121516244.0/4294967296.0,1,-nbitq), 
to_sfixed(-12482010.0/4294967296.0,1,-nbitq), 
to_sfixed(-53102833.0/4294967296.0,1,-nbitq), 
to_sfixed(-179814605.0/4294967296.0,1,-nbitq), 
to_sfixed(8610115.0/4294967296.0,1,-nbitq), 
to_sfixed(-1111803125.0/4294967296.0,1,-nbitq), 
to_sfixed(-578804466.0/4294967296.0,1,-nbitq), 
to_sfixed(615833650.0/4294967296.0,1,-nbitq), 
to_sfixed(-662013437.0/4294967296.0,1,-nbitq), 
to_sfixed(-318539036.0/4294967296.0,1,-nbitq), 
to_sfixed(256523015.0/4294967296.0,1,-nbitq), 
to_sfixed(-412284746.0/4294967296.0,1,-nbitq), 
to_sfixed(105847767.0/4294967296.0,1,-nbitq), 
to_sfixed(304344939.0/4294967296.0,1,-nbitq), 
to_sfixed(394267096.0/4294967296.0,1,-nbitq), 
to_sfixed(81733324.0/4294967296.0,1,-nbitq), 
to_sfixed(-20369540.0/4294967296.0,1,-nbitq), 
to_sfixed(74271637.0/4294967296.0,1,-nbitq), 
to_sfixed(238493194.0/4294967296.0,1,-nbitq), 
to_sfixed(271912569.0/4294967296.0,1,-nbitq), 
to_sfixed(266575678.0/4294967296.0,1,-nbitq), 
to_sfixed(246600001.0/4294967296.0,1,-nbitq), 
to_sfixed(113412297.0/4294967296.0,1,-nbitq), 
to_sfixed(59211452.0/4294967296.0,1,-nbitq), 
to_sfixed(40030576.0/4294967296.0,1,-nbitq), 
to_sfixed(690551733.0/4294967296.0,1,-nbitq), 
to_sfixed(-300932357.0/4294967296.0,1,-nbitq), 
to_sfixed(-138295396.0/4294967296.0,1,-nbitq), 
to_sfixed(-815411175.0/4294967296.0,1,-nbitq), 
to_sfixed(1056573810.0/4294967296.0,1,-nbitq), 
to_sfixed(382654862.0/4294967296.0,1,-nbitq), 
to_sfixed(428912234.0/4294967296.0,1,-nbitq), 
to_sfixed(-105695966.0/4294967296.0,1,-nbitq), 
to_sfixed(18318001.0/4294967296.0,1,-nbitq), 
to_sfixed(-131982491.0/4294967296.0,1,-nbitq), 
to_sfixed(173793217.0/4294967296.0,1,-nbitq), 
to_sfixed(-152069471.0/4294967296.0,1,-nbitq), 
to_sfixed(331856671.0/4294967296.0,1,-nbitq), 
to_sfixed(-143268269.0/4294967296.0,1,-nbitq), 
to_sfixed(-233414653.0/4294967296.0,1,-nbitq), 
to_sfixed(-394566610.0/4294967296.0,1,-nbitq), 
to_sfixed(-694652241.0/4294967296.0,1,-nbitq), 
to_sfixed(-270251983.0/4294967296.0,1,-nbitq), 
to_sfixed(794948738.0/4294967296.0,1,-nbitq), 
to_sfixed(156680675.0/4294967296.0,1,-nbitq), 
to_sfixed(-222559116.0/4294967296.0,1,-nbitq), 
to_sfixed(579549007.0/4294967296.0,1,-nbitq), 
to_sfixed(195368568.0/4294967296.0,1,-nbitq), 
to_sfixed(290808654.0/4294967296.0,1,-nbitq), 
to_sfixed(491912483.0/4294967296.0,1,-nbitq), 
to_sfixed(5348631.0/4294967296.0,1,-nbitq), 
to_sfixed(323336954.0/4294967296.0,1,-nbitq), 
to_sfixed(-166887338.0/4294967296.0,1,-nbitq), 
to_sfixed(315387506.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(470072181.0/4294967296.0,1,-nbitq), 
to_sfixed(104389444.0/4294967296.0,1,-nbitq), 
to_sfixed(40952036.0/4294967296.0,1,-nbitq), 
to_sfixed(524396616.0/4294967296.0,1,-nbitq), 
to_sfixed(428077148.0/4294967296.0,1,-nbitq), 
to_sfixed(-810627936.0/4294967296.0,1,-nbitq), 
to_sfixed(-113589192.0/4294967296.0,1,-nbitq), 
to_sfixed(42538362.0/4294967296.0,1,-nbitq), 
to_sfixed(1367532668.0/4294967296.0,1,-nbitq), 
to_sfixed(23502552.0/4294967296.0,1,-nbitq), 
to_sfixed(-54605658.0/4294967296.0,1,-nbitq), 
to_sfixed(280322978.0/4294967296.0,1,-nbitq), 
to_sfixed(-167972758.0/4294967296.0,1,-nbitq), 
to_sfixed(-751938296.0/4294967296.0,1,-nbitq), 
to_sfixed(-245587186.0/4294967296.0,1,-nbitq), 
to_sfixed(-307056500.0/4294967296.0,1,-nbitq), 
to_sfixed(216030486.0/4294967296.0,1,-nbitq), 
to_sfixed(89571829.0/4294967296.0,1,-nbitq), 
to_sfixed(-223909709.0/4294967296.0,1,-nbitq), 
to_sfixed(386134783.0/4294967296.0,1,-nbitq), 
to_sfixed(-233101738.0/4294967296.0,1,-nbitq), 
to_sfixed(419440959.0/4294967296.0,1,-nbitq), 
to_sfixed(-540057960.0/4294967296.0,1,-nbitq), 
to_sfixed(-564601097.0/4294967296.0,1,-nbitq), 
to_sfixed(-72623261.0/4294967296.0,1,-nbitq), 
to_sfixed(-873572885.0/4294967296.0,1,-nbitq), 
to_sfixed(-359335256.0/4294967296.0,1,-nbitq), 
to_sfixed(-352840700.0/4294967296.0,1,-nbitq), 
to_sfixed(-174389685.0/4294967296.0,1,-nbitq), 
to_sfixed(-554651078.0/4294967296.0,1,-nbitq), 
to_sfixed(522462920.0/4294967296.0,1,-nbitq), 
to_sfixed(-575696491.0/4294967296.0,1,-nbitq), 
to_sfixed(209130146.0/4294967296.0,1,-nbitq), 
to_sfixed(636759392.0/4294967296.0,1,-nbitq), 
to_sfixed(-756335928.0/4294967296.0,1,-nbitq), 
to_sfixed(-290280870.0/4294967296.0,1,-nbitq), 
to_sfixed(112739707.0/4294967296.0,1,-nbitq), 
to_sfixed(-751266105.0/4294967296.0,1,-nbitq), 
to_sfixed(31728853.0/4294967296.0,1,-nbitq), 
to_sfixed(203071854.0/4294967296.0,1,-nbitq), 
to_sfixed(603428473.0/4294967296.0,1,-nbitq), 
to_sfixed(-564803154.0/4294967296.0,1,-nbitq), 
to_sfixed(-904560056.0/4294967296.0,1,-nbitq), 
to_sfixed(426532799.0/4294967296.0,1,-nbitq), 
to_sfixed(-387972029.0/4294967296.0,1,-nbitq), 
to_sfixed(367446983.0/4294967296.0,1,-nbitq), 
to_sfixed(295528280.0/4294967296.0,1,-nbitq), 
to_sfixed(505565847.0/4294967296.0,1,-nbitq), 
to_sfixed(-455601819.0/4294967296.0,1,-nbitq), 
to_sfixed(-280872465.0/4294967296.0,1,-nbitq), 
to_sfixed(-347076716.0/4294967296.0,1,-nbitq), 
to_sfixed(849228220.0/4294967296.0,1,-nbitq), 
to_sfixed(-106893686.0/4294967296.0,1,-nbitq), 
to_sfixed(-259377199.0/4294967296.0,1,-nbitq), 
to_sfixed(-331636421.0/4294967296.0,1,-nbitq), 
to_sfixed(681297487.0/4294967296.0,1,-nbitq), 
to_sfixed(-254025895.0/4294967296.0,1,-nbitq), 
to_sfixed(960962784.0/4294967296.0,1,-nbitq), 
to_sfixed(-354205966.0/4294967296.0,1,-nbitq), 
to_sfixed(181518790.0/4294967296.0,1,-nbitq), 
to_sfixed(-116297056.0/4294967296.0,1,-nbitq), 
to_sfixed(462707098.0/4294967296.0,1,-nbitq), 
to_sfixed(-221726254.0/4294967296.0,1,-nbitq), 
to_sfixed(-434908466.0/4294967296.0,1,-nbitq), 
to_sfixed(132913507.0/4294967296.0,1,-nbitq), 
to_sfixed(-75409108.0/4294967296.0,1,-nbitq), 
to_sfixed(-456992111.0/4294967296.0,1,-nbitq), 
to_sfixed(47274483.0/4294967296.0,1,-nbitq), 
to_sfixed(114504131.0/4294967296.0,1,-nbitq), 
to_sfixed(896847214.0/4294967296.0,1,-nbitq), 
to_sfixed(180037277.0/4294967296.0,1,-nbitq), 
to_sfixed(340210899.0/4294967296.0,1,-nbitq), 
to_sfixed(137920331.0/4294967296.0,1,-nbitq), 
to_sfixed(317158725.0/4294967296.0,1,-nbitq), 
to_sfixed(-173248857.0/4294967296.0,1,-nbitq), 
to_sfixed(1104461697.0/4294967296.0,1,-nbitq), 
to_sfixed(1256207686.0/4294967296.0,1,-nbitq), 
to_sfixed(-185031826.0/4294967296.0,1,-nbitq), 
to_sfixed(-82538391.0/4294967296.0,1,-nbitq), 
to_sfixed(76576599.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(566217419.0/4294967296.0,1,-nbitq), 
to_sfixed(-253412473.0/4294967296.0,1,-nbitq), 
to_sfixed(-288193624.0/4294967296.0,1,-nbitq), 
to_sfixed(508144026.0/4294967296.0,1,-nbitq), 
to_sfixed(524631011.0/4294967296.0,1,-nbitq), 
to_sfixed(-494746962.0/4294967296.0,1,-nbitq), 
to_sfixed(325449179.0/4294967296.0,1,-nbitq), 
to_sfixed(-17031008.0/4294967296.0,1,-nbitq), 
to_sfixed(1339880250.0/4294967296.0,1,-nbitq), 
to_sfixed(166289899.0/4294967296.0,1,-nbitq), 
to_sfixed(-61891970.0/4294967296.0,1,-nbitq), 
to_sfixed(417664026.0/4294967296.0,1,-nbitq), 
to_sfixed(-211413824.0/4294967296.0,1,-nbitq), 
to_sfixed(-1136389954.0/4294967296.0,1,-nbitq), 
to_sfixed(-477663186.0/4294967296.0,1,-nbitq), 
to_sfixed(-94288417.0/4294967296.0,1,-nbitq), 
to_sfixed(-439939788.0/4294967296.0,1,-nbitq), 
to_sfixed(222046007.0/4294967296.0,1,-nbitq), 
to_sfixed(-19422289.0/4294967296.0,1,-nbitq), 
to_sfixed(357336436.0/4294967296.0,1,-nbitq), 
to_sfixed(-12886541.0/4294967296.0,1,-nbitq), 
to_sfixed(224895555.0/4294967296.0,1,-nbitq), 
to_sfixed(122868291.0/4294967296.0,1,-nbitq), 
to_sfixed(-312753280.0/4294967296.0,1,-nbitq), 
to_sfixed(-106817201.0/4294967296.0,1,-nbitq), 
to_sfixed(-255901916.0/4294967296.0,1,-nbitq), 
to_sfixed(-236284627.0/4294967296.0,1,-nbitq), 
to_sfixed(-365805178.0/4294967296.0,1,-nbitq), 
to_sfixed(177209369.0/4294967296.0,1,-nbitq), 
to_sfixed(-1497496627.0/4294967296.0,1,-nbitq), 
to_sfixed(343556877.0/4294967296.0,1,-nbitq), 
to_sfixed(-765945629.0/4294967296.0,1,-nbitq), 
to_sfixed(113410874.0/4294967296.0,1,-nbitq), 
to_sfixed(269857939.0/4294967296.0,1,-nbitq), 
to_sfixed(-611152414.0/4294967296.0,1,-nbitq), 
to_sfixed(-667320127.0/4294967296.0,1,-nbitq), 
to_sfixed(107732849.0/4294967296.0,1,-nbitq), 
to_sfixed(-481082926.0/4294967296.0,1,-nbitq), 
to_sfixed(124931604.0/4294967296.0,1,-nbitq), 
to_sfixed(-346200130.0/4294967296.0,1,-nbitq), 
to_sfixed(400171256.0/4294967296.0,1,-nbitq), 
to_sfixed(-315123301.0/4294967296.0,1,-nbitq), 
to_sfixed(-1278719.0/4294967296.0,1,-nbitq), 
to_sfixed(810702800.0/4294967296.0,1,-nbitq), 
to_sfixed(-52605909.0/4294967296.0,1,-nbitq), 
to_sfixed(1401142558.0/4294967296.0,1,-nbitq), 
to_sfixed(55483783.0/4294967296.0,1,-nbitq), 
to_sfixed(73250335.0/4294967296.0,1,-nbitq), 
to_sfixed(-245807351.0/4294967296.0,1,-nbitq), 
to_sfixed(-466215600.0/4294967296.0,1,-nbitq), 
to_sfixed(-189378760.0/4294967296.0,1,-nbitq), 
to_sfixed(927731496.0/4294967296.0,1,-nbitq), 
to_sfixed(-187102652.0/4294967296.0,1,-nbitq), 
to_sfixed(101598080.0/4294967296.0,1,-nbitq), 
to_sfixed(475659404.0/4294967296.0,1,-nbitq), 
to_sfixed(1034017166.0/4294967296.0,1,-nbitq), 
to_sfixed(-143570820.0/4294967296.0,1,-nbitq), 
to_sfixed(292473087.0/4294967296.0,1,-nbitq), 
to_sfixed(301906179.0/4294967296.0,1,-nbitq), 
to_sfixed(-213470316.0/4294967296.0,1,-nbitq), 
to_sfixed(-235631611.0/4294967296.0,1,-nbitq), 
to_sfixed(-97245229.0/4294967296.0,1,-nbitq), 
to_sfixed(-314701096.0/4294967296.0,1,-nbitq), 
to_sfixed(-67768941.0/4294967296.0,1,-nbitq), 
to_sfixed(239824830.0/4294967296.0,1,-nbitq), 
to_sfixed(240052640.0/4294967296.0,1,-nbitq), 
to_sfixed(-270275886.0/4294967296.0,1,-nbitq), 
to_sfixed(360084729.0/4294967296.0,1,-nbitq), 
to_sfixed(-256622921.0/4294967296.0,1,-nbitq), 
to_sfixed(11476473.0/4294967296.0,1,-nbitq), 
to_sfixed(187345989.0/4294967296.0,1,-nbitq), 
to_sfixed(342431660.0/4294967296.0,1,-nbitq), 
to_sfixed(951053081.0/4294967296.0,1,-nbitq), 
to_sfixed(106888462.0/4294967296.0,1,-nbitq), 
to_sfixed(-132816213.0/4294967296.0,1,-nbitq), 
to_sfixed(478367888.0/4294967296.0,1,-nbitq), 
to_sfixed(1345783528.0/4294967296.0,1,-nbitq), 
to_sfixed(-406931718.0/4294967296.0,1,-nbitq), 
to_sfixed(28102886.0/4294967296.0,1,-nbitq), 
to_sfixed(-204303634.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(642766239.0/4294967296.0,1,-nbitq), 
to_sfixed(-663086000.0/4294967296.0,1,-nbitq), 
to_sfixed(-283520620.0/4294967296.0,1,-nbitq), 
to_sfixed(953502194.0/4294967296.0,1,-nbitq), 
to_sfixed(181442131.0/4294967296.0,1,-nbitq), 
to_sfixed(-882031652.0/4294967296.0,1,-nbitq), 
to_sfixed(227615018.0/4294967296.0,1,-nbitq), 
to_sfixed(-163994524.0/4294967296.0,1,-nbitq), 
to_sfixed(685400102.0/4294967296.0,1,-nbitq), 
to_sfixed(169015310.0/4294967296.0,1,-nbitq), 
to_sfixed(-202424274.0/4294967296.0,1,-nbitq), 
to_sfixed(900913204.0/4294967296.0,1,-nbitq), 
to_sfixed(-368894942.0/4294967296.0,1,-nbitq), 
to_sfixed(-677639740.0/4294967296.0,1,-nbitq), 
to_sfixed(-112681865.0/4294967296.0,1,-nbitq), 
to_sfixed(209887919.0/4294967296.0,1,-nbitq), 
to_sfixed(-275782389.0/4294967296.0,1,-nbitq), 
to_sfixed(148559810.0/4294967296.0,1,-nbitq), 
to_sfixed(-155309447.0/4294967296.0,1,-nbitq), 
to_sfixed(-178151443.0/4294967296.0,1,-nbitq), 
to_sfixed(145376039.0/4294967296.0,1,-nbitq), 
to_sfixed(-40448850.0/4294967296.0,1,-nbitq), 
to_sfixed(21132726.0/4294967296.0,1,-nbitq), 
to_sfixed(-120518712.0/4294967296.0,1,-nbitq), 
to_sfixed(142915704.0/4294967296.0,1,-nbitq), 
to_sfixed(-461000103.0/4294967296.0,1,-nbitq), 
to_sfixed(-128129127.0/4294967296.0,1,-nbitq), 
to_sfixed(149222971.0/4294967296.0,1,-nbitq), 
to_sfixed(76268586.0/4294967296.0,1,-nbitq), 
to_sfixed(-576179524.0/4294967296.0,1,-nbitq), 
to_sfixed(1038456193.0/4294967296.0,1,-nbitq), 
to_sfixed(-170917031.0/4294967296.0,1,-nbitq), 
to_sfixed(-369321416.0/4294967296.0,1,-nbitq), 
to_sfixed(105864760.0/4294967296.0,1,-nbitq), 
to_sfixed(-710474362.0/4294967296.0,1,-nbitq), 
to_sfixed(-809989108.0/4294967296.0,1,-nbitq), 
to_sfixed(-47464.0/4294967296.0,1,-nbitq), 
to_sfixed(-502632646.0/4294967296.0,1,-nbitq), 
to_sfixed(-217440846.0/4294967296.0,1,-nbitq), 
to_sfixed(192961892.0/4294967296.0,1,-nbitq), 
to_sfixed(414500101.0/4294967296.0,1,-nbitq), 
to_sfixed(23715319.0/4294967296.0,1,-nbitq), 
to_sfixed(236704503.0/4294967296.0,1,-nbitq), 
to_sfixed(890752206.0/4294967296.0,1,-nbitq), 
to_sfixed(-227019373.0/4294967296.0,1,-nbitq), 
to_sfixed(1563288141.0/4294967296.0,1,-nbitq), 
to_sfixed(-9258439.0/4294967296.0,1,-nbitq), 
to_sfixed(503260482.0/4294967296.0,1,-nbitq), 
to_sfixed(-619087145.0/4294967296.0,1,-nbitq), 
to_sfixed(-81411742.0/4294967296.0,1,-nbitq), 
to_sfixed(-101073368.0/4294967296.0,1,-nbitq), 
to_sfixed(1279912003.0/4294967296.0,1,-nbitq), 
to_sfixed(-21732802.0/4294967296.0,1,-nbitq), 
to_sfixed(60790559.0/4294967296.0,1,-nbitq), 
to_sfixed(744929362.0/4294967296.0,1,-nbitq), 
to_sfixed(578508012.0/4294967296.0,1,-nbitq), 
to_sfixed(303614815.0/4294967296.0,1,-nbitq), 
to_sfixed(519981582.0/4294967296.0,1,-nbitq), 
to_sfixed(-385504518.0/4294967296.0,1,-nbitq), 
to_sfixed(221305208.0/4294967296.0,1,-nbitq), 
to_sfixed(31286156.0/4294967296.0,1,-nbitq), 
to_sfixed(655192174.0/4294967296.0,1,-nbitq), 
to_sfixed(-345011720.0/4294967296.0,1,-nbitq), 
to_sfixed(-235680523.0/4294967296.0,1,-nbitq), 
to_sfixed(-208368249.0/4294967296.0,1,-nbitq), 
to_sfixed(-144100272.0/4294967296.0,1,-nbitq), 
to_sfixed(-196019616.0/4294967296.0,1,-nbitq), 
to_sfixed(614386486.0/4294967296.0,1,-nbitq), 
to_sfixed(-305374584.0/4294967296.0,1,-nbitq), 
to_sfixed(59631049.0/4294967296.0,1,-nbitq), 
to_sfixed(-707692111.0/4294967296.0,1,-nbitq), 
to_sfixed(315378998.0/4294967296.0,1,-nbitq), 
to_sfixed(849059664.0/4294967296.0,1,-nbitq), 
to_sfixed(327931247.0/4294967296.0,1,-nbitq), 
to_sfixed(-274007073.0/4294967296.0,1,-nbitq), 
to_sfixed(58456976.0/4294967296.0,1,-nbitq), 
to_sfixed(636292901.0/4294967296.0,1,-nbitq), 
to_sfixed(26765878.0/4294967296.0,1,-nbitq), 
to_sfixed(-374852836.0/4294967296.0,1,-nbitq), 
to_sfixed(72798572.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(55406888.0/4294967296.0,1,-nbitq), 
to_sfixed(-637238103.0/4294967296.0,1,-nbitq), 
to_sfixed(-730121626.0/4294967296.0,1,-nbitq), 
to_sfixed(700425938.0/4294967296.0,1,-nbitq), 
to_sfixed(-170511371.0/4294967296.0,1,-nbitq), 
to_sfixed(-840405173.0/4294967296.0,1,-nbitq), 
to_sfixed(144541968.0/4294967296.0,1,-nbitq), 
to_sfixed(-106808417.0/4294967296.0,1,-nbitq), 
to_sfixed(-62628919.0/4294967296.0,1,-nbitq), 
to_sfixed(26408673.0/4294967296.0,1,-nbitq), 
to_sfixed(123842813.0/4294967296.0,1,-nbitq), 
to_sfixed(910060628.0/4294967296.0,1,-nbitq), 
to_sfixed(-37028281.0/4294967296.0,1,-nbitq), 
to_sfixed(-164793112.0/4294967296.0,1,-nbitq), 
to_sfixed(-32249009.0/4294967296.0,1,-nbitq), 
to_sfixed(402591089.0/4294967296.0,1,-nbitq), 
to_sfixed(-124737193.0/4294967296.0,1,-nbitq), 
to_sfixed(139782514.0/4294967296.0,1,-nbitq), 
to_sfixed(5667767.0/4294967296.0,1,-nbitq), 
to_sfixed(-354429641.0/4294967296.0,1,-nbitq), 
to_sfixed(-412121802.0/4294967296.0,1,-nbitq), 
to_sfixed(-213504762.0/4294967296.0,1,-nbitq), 
to_sfixed(451615379.0/4294967296.0,1,-nbitq), 
to_sfixed(-233364321.0/4294967296.0,1,-nbitq), 
to_sfixed(-140517958.0/4294967296.0,1,-nbitq), 
to_sfixed(-621342599.0/4294967296.0,1,-nbitq), 
to_sfixed(-247300299.0/4294967296.0,1,-nbitq), 
to_sfixed(-348468017.0/4294967296.0,1,-nbitq), 
to_sfixed(-288225473.0/4294967296.0,1,-nbitq), 
to_sfixed(-957833648.0/4294967296.0,1,-nbitq), 
to_sfixed(791528817.0/4294967296.0,1,-nbitq), 
to_sfixed(-265639820.0/4294967296.0,1,-nbitq), 
to_sfixed(23942629.0/4294967296.0,1,-nbitq), 
to_sfixed(-381380812.0/4294967296.0,1,-nbitq), 
to_sfixed(-255451674.0/4294967296.0,1,-nbitq), 
to_sfixed(-511656370.0/4294967296.0,1,-nbitq), 
to_sfixed(444740673.0/4294967296.0,1,-nbitq), 
to_sfixed(-721626662.0/4294967296.0,1,-nbitq), 
to_sfixed(58542685.0/4294967296.0,1,-nbitq), 
to_sfixed(95154679.0/4294967296.0,1,-nbitq), 
to_sfixed(325610253.0/4294967296.0,1,-nbitq), 
to_sfixed(-272007601.0/4294967296.0,1,-nbitq), 
to_sfixed(576225874.0/4294967296.0,1,-nbitq), 
to_sfixed(1093728930.0/4294967296.0,1,-nbitq), 
to_sfixed(35397974.0/4294967296.0,1,-nbitq), 
to_sfixed(206477722.0/4294967296.0,1,-nbitq), 
to_sfixed(97713674.0/4294967296.0,1,-nbitq), 
to_sfixed(228729476.0/4294967296.0,1,-nbitq), 
to_sfixed(-717624223.0/4294967296.0,1,-nbitq), 
to_sfixed(310673868.0/4294967296.0,1,-nbitq), 
to_sfixed(337032025.0/4294967296.0,1,-nbitq), 
to_sfixed(1244016176.0/4294967296.0,1,-nbitq), 
to_sfixed(-42211413.0/4294967296.0,1,-nbitq), 
to_sfixed(-316886546.0/4294967296.0,1,-nbitq), 
to_sfixed(-151535879.0/4294967296.0,1,-nbitq), 
to_sfixed(42168986.0/4294967296.0,1,-nbitq), 
to_sfixed(-101362866.0/4294967296.0,1,-nbitq), 
to_sfixed(946929794.0/4294967296.0,1,-nbitq), 
to_sfixed(181104407.0/4294967296.0,1,-nbitq), 
to_sfixed(3796854.0/4294967296.0,1,-nbitq), 
to_sfixed(-348773693.0/4294967296.0,1,-nbitq), 
to_sfixed(595622721.0/4294967296.0,1,-nbitq), 
to_sfixed(-110872184.0/4294967296.0,1,-nbitq), 
to_sfixed(-254982304.0/4294967296.0,1,-nbitq), 
to_sfixed(-320357680.0/4294967296.0,1,-nbitq), 
to_sfixed(378009257.0/4294967296.0,1,-nbitq), 
to_sfixed(43055836.0/4294967296.0,1,-nbitq), 
to_sfixed(359949249.0/4294967296.0,1,-nbitq), 
to_sfixed(-344814520.0/4294967296.0,1,-nbitq), 
to_sfixed(-10850816.0/4294967296.0,1,-nbitq), 
to_sfixed(-537341401.0/4294967296.0,1,-nbitq), 
to_sfixed(-373739291.0/4294967296.0,1,-nbitq), 
to_sfixed(1037191019.0/4294967296.0,1,-nbitq), 
to_sfixed(-235162043.0/4294967296.0,1,-nbitq), 
to_sfixed(-296016323.0/4294967296.0,1,-nbitq), 
to_sfixed(-403971004.0/4294967296.0,1,-nbitq), 
to_sfixed(-191553996.0/4294967296.0,1,-nbitq), 
to_sfixed(314293996.0/4294967296.0,1,-nbitq), 
to_sfixed(-132960994.0/4294967296.0,1,-nbitq), 
to_sfixed(239869096.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(519754253.0/4294967296.0,1,-nbitq), 
to_sfixed(-892049452.0/4294967296.0,1,-nbitq), 
to_sfixed(246851661.0/4294967296.0,1,-nbitq), 
to_sfixed(957159634.0/4294967296.0,1,-nbitq), 
to_sfixed(-421662556.0/4294967296.0,1,-nbitq), 
to_sfixed(-605469399.0/4294967296.0,1,-nbitq), 
to_sfixed(-18163251.0/4294967296.0,1,-nbitq), 
to_sfixed(-188241550.0/4294967296.0,1,-nbitq), 
to_sfixed(-368574385.0/4294967296.0,1,-nbitq), 
to_sfixed(-101481788.0/4294967296.0,1,-nbitq), 
to_sfixed(794988086.0/4294967296.0,1,-nbitq), 
to_sfixed(48885814.0/4294967296.0,1,-nbitq), 
to_sfixed(14908353.0/4294967296.0,1,-nbitq), 
to_sfixed(642132930.0/4294967296.0,1,-nbitq), 
to_sfixed(304482980.0/4294967296.0,1,-nbitq), 
to_sfixed(159452428.0/4294967296.0,1,-nbitq), 
to_sfixed(-74806123.0/4294967296.0,1,-nbitq), 
to_sfixed(180561255.0/4294967296.0,1,-nbitq), 
to_sfixed(232928510.0/4294967296.0,1,-nbitq), 
to_sfixed(-147705104.0/4294967296.0,1,-nbitq), 
to_sfixed(101364322.0/4294967296.0,1,-nbitq), 
to_sfixed(200211234.0/4294967296.0,1,-nbitq), 
to_sfixed(749468979.0/4294967296.0,1,-nbitq), 
to_sfixed(-267109478.0/4294967296.0,1,-nbitq), 
to_sfixed(-286960911.0/4294967296.0,1,-nbitq), 
to_sfixed(-435615322.0/4294967296.0,1,-nbitq), 
to_sfixed(-144985570.0/4294967296.0,1,-nbitq), 
to_sfixed(-154512324.0/4294967296.0,1,-nbitq), 
to_sfixed(-243827299.0/4294967296.0,1,-nbitq), 
to_sfixed(-349136966.0/4294967296.0,1,-nbitq), 
to_sfixed(722622389.0/4294967296.0,1,-nbitq), 
to_sfixed(407105915.0/4294967296.0,1,-nbitq), 
to_sfixed(58673208.0/4294967296.0,1,-nbitq), 
to_sfixed(-178364925.0/4294967296.0,1,-nbitq), 
to_sfixed(126803009.0/4294967296.0,1,-nbitq), 
to_sfixed(27346384.0/4294967296.0,1,-nbitq), 
to_sfixed(40232564.0/4294967296.0,1,-nbitq), 
to_sfixed(155551366.0/4294967296.0,1,-nbitq), 
to_sfixed(346872693.0/4294967296.0,1,-nbitq), 
to_sfixed(-224748802.0/4294967296.0,1,-nbitq), 
to_sfixed(-183590099.0/4294967296.0,1,-nbitq), 
to_sfixed(-459150916.0/4294967296.0,1,-nbitq), 
to_sfixed(778545689.0/4294967296.0,1,-nbitq), 
to_sfixed(1099776434.0/4294967296.0,1,-nbitq), 
to_sfixed(494591128.0/4294967296.0,1,-nbitq), 
to_sfixed(-42134870.0/4294967296.0,1,-nbitq), 
to_sfixed(202946544.0/4294967296.0,1,-nbitq), 
to_sfixed(228872871.0/4294967296.0,1,-nbitq), 
to_sfixed(-518692820.0/4294967296.0,1,-nbitq), 
to_sfixed(460125109.0/4294967296.0,1,-nbitq), 
to_sfixed(124706866.0/4294967296.0,1,-nbitq), 
to_sfixed(136569589.0/4294967296.0,1,-nbitq), 
to_sfixed(12419337.0/4294967296.0,1,-nbitq), 
to_sfixed(372986136.0/4294967296.0,1,-nbitq), 
to_sfixed(590316292.0/4294967296.0,1,-nbitq), 
to_sfixed(-28259595.0/4294967296.0,1,-nbitq), 
to_sfixed(-159239422.0/4294967296.0,1,-nbitq), 
to_sfixed(521076427.0/4294967296.0,1,-nbitq), 
to_sfixed(-123290701.0/4294967296.0,1,-nbitq), 
to_sfixed(361664361.0/4294967296.0,1,-nbitq), 
to_sfixed(-362615078.0/4294967296.0,1,-nbitq), 
to_sfixed(397828131.0/4294967296.0,1,-nbitq), 
to_sfixed(-277294669.0/4294967296.0,1,-nbitq), 
to_sfixed(-748568535.0/4294967296.0,1,-nbitq), 
to_sfixed(279049719.0/4294967296.0,1,-nbitq), 
to_sfixed(328883007.0/4294967296.0,1,-nbitq), 
to_sfixed(468508578.0/4294967296.0,1,-nbitq), 
to_sfixed(134605560.0/4294967296.0,1,-nbitq), 
to_sfixed(367122219.0/4294967296.0,1,-nbitq), 
to_sfixed(105262931.0/4294967296.0,1,-nbitq), 
to_sfixed(-646676301.0/4294967296.0,1,-nbitq), 
to_sfixed(240808740.0/4294967296.0,1,-nbitq), 
to_sfixed(416809680.0/4294967296.0,1,-nbitq), 
to_sfixed(314166050.0/4294967296.0,1,-nbitq), 
to_sfixed(246303100.0/4294967296.0,1,-nbitq), 
to_sfixed(-643613961.0/4294967296.0,1,-nbitq), 
to_sfixed(470638643.0/4294967296.0,1,-nbitq), 
to_sfixed(154453125.0/4294967296.0,1,-nbitq), 
to_sfixed(114598794.0/4294967296.0,1,-nbitq), 
to_sfixed(316168494.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(346411241.0/4294967296.0,1,-nbitq), 
to_sfixed(695789189.0/4294967296.0,1,-nbitq), 
to_sfixed(-130797142.0/4294967296.0,1,-nbitq), 
to_sfixed(703926753.0/4294967296.0,1,-nbitq), 
to_sfixed(-801833961.0/4294967296.0,1,-nbitq), 
to_sfixed(-130043367.0/4294967296.0,1,-nbitq), 
to_sfixed(218751249.0/4294967296.0,1,-nbitq), 
to_sfixed(-465293848.0/4294967296.0,1,-nbitq), 
to_sfixed(70115485.0/4294967296.0,1,-nbitq), 
to_sfixed(272381464.0/4294967296.0,1,-nbitq), 
to_sfixed(1159692686.0/4294967296.0,1,-nbitq), 
to_sfixed(348672658.0/4294967296.0,1,-nbitq), 
to_sfixed(481112933.0/4294967296.0,1,-nbitq), 
to_sfixed(1180130607.0/4294967296.0,1,-nbitq), 
to_sfixed(148382376.0/4294967296.0,1,-nbitq), 
to_sfixed(192172257.0/4294967296.0,1,-nbitq), 
to_sfixed(170031964.0/4294967296.0,1,-nbitq), 
to_sfixed(350336591.0/4294967296.0,1,-nbitq), 
to_sfixed(402499997.0/4294967296.0,1,-nbitq), 
to_sfixed(-613608468.0/4294967296.0,1,-nbitq), 
to_sfixed(350837315.0/4294967296.0,1,-nbitq), 
to_sfixed(-103492843.0/4294967296.0,1,-nbitq), 
to_sfixed(168478949.0/4294967296.0,1,-nbitq), 
to_sfixed(414375737.0/4294967296.0,1,-nbitq), 
to_sfixed(-334486452.0/4294967296.0,1,-nbitq), 
to_sfixed(-225140059.0/4294967296.0,1,-nbitq), 
to_sfixed(-560716794.0/4294967296.0,1,-nbitq), 
to_sfixed(-450779994.0/4294967296.0,1,-nbitq), 
to_sfixed(-1034466217.0/4294967296.0,1,-nbitq), 
to_sfixed(395497283.0/4294967296.0,1,-nbitq), 
to_sfixed(205027685.0/4294967296.0,1,-nbitq), 
to_sfixed(-261224911.0/4294967296.0,1,-nbitq), 
to_sfixed(1011906276.0/4294967296.0,1,-nbitq), 
to_sfixed(-164760186.0/4294967296.0,1,-nbitq), 
to_sfixed(-256508397.0/4294967296.0,1,-nbitq), 
to_sfixed(-24184970.0/4294967296.0,1,-nbitq), 
to_sfixed(62692849.0/4294967296.0,1,-nbitq), 
to_sfixed(408290084.0/4294967296.0,1,-nbitq), 
to_sfixed(-262729049.0/4294967296.0,1,-nbitq), 
to_sfixed(-240021070.0/4294967296.0,1,-nbitq), 
to_sfixed(32414655.0/4294967296.0,1,-nbitq), 
to_sfixed(-301437269.0/4294967296.0,1,-nbitq), 
to_sfixed(1630809048.0/4294967296.0,1,-nbitq), 
to_sfixed(1001696011.0/4294967296.0,1,-nbitq), 
to_sfixed(106364743.0/4294967296.0,1,-nbitq), 
to_sfixed(-440912633.0/4294967296.0,1,-nbitq), 
to_sfixed(-437443298.0/4294967296.0,1,-nbitq), 
to_sfixed(348767874.0/4294967296.0,1,-nbitq), 
to_sfixed(-782514085.0/4294967296.0,1,-nbitq), 
to_sfixed(1002828622.0/4294967296.0,1,-nbitq), 
to_sfixed(240711682.0/4294967296.0,1,-nbitq), 
to_sfixed(-6878738.0/4294967296.0,1,-nbitq), 
to_sfixed(626799426.0/4294967296.0,1,-nbitq), 
to_sfixed(568413187.0/4294967296.0,1,-nbitq), 
to_sfixed(1463752794.0/4294967296.0,1,-nbitq), 
to_sfixed(410343081.0/4294967296.0,1,-nbitq), 
to_sfixed(-87224340.0/4294967296.0,1,-nbitq), 
to_sfixed(-412671931.0/4294967296.0,1,-nbitq), 
to_sfixed(-197073324.0/4294967296.0,1,-nbitq), 
to_sfixed(-147620871.0/4294967296.0,1,-nbitq), 
to_sfixed(150162440.0/4294967296.0,1,-nbitq), 
to_sfixed(735573028.0/4294967296.0,1,-nbitq), 
to_sfixed(-416260601.0/4294967296.0,1,-nbitq), 
to_sfixed(-487121623.0/4294967296.0,1,-nbitq), 
to_sfixed(-126774083.0/4294967296.0,1,-nbitq), 
to_sfixed(214486389.0/4294967296.0,1,-nbitq), 
to_sfixed(-233737117.0/4294967296.0,1,-nbitq), 
to_sfixed(1116936694.0/4294967296.0,1,-nbitq), 
to_sfixed(13960339.0/4294967296.0,1,-nbitq), 
to_sfixed(-198927674.0/4294967296.0,1,-nbitq), 
to_sfixed(-160667148.0/4294967296.0,1,-nbitq), 
to_sfixed(17444348.0/4294967296.0,1,-nbitq), 
to_sfixed(331331820.0/4294967296.0,1,-nbitq), 
to_sfixed(149409700.0/4294967296.0,1,-nbitq), 
to_sfixed(147468193.0/4294967296.0,1,-nbitq), 
to_sfixed(-248382605.0/4294967296.0,1,-nbitq), 
to_sfixed(76785318.0/4294967296.0,1,-nbitq), 
to_sfixed(372201473.0/4294967296.0,1,-nbitq), 
to_sfixed(-93199873.0/4294967296.0,1,-nbitq), 
to_sfixed(-373924095.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(90427738.0/4294967296.0,1,-nbitq), 
to_sfixed(896594586.0/4294967296.0,1,-nbitq), 
to_sfixed(82167182.0/4294967296.0,1,-nbitq), 
to_sfixed(799887413.0/4294967296.0,1,-nbitq), 
to_sfixed(-499731356.0/4294967296.0,1,-nbitq), 
to_sfixed(-221685255.0/4294967296.0,1,-nbitq), 
to_sfixed(442394110.0/4294967296.0,1,-nbitq), 
to_sfixed(-270504882.0/4294967296.0,1,-nbitq), 
to_sfixed(383682804.0/4294967296.0,1,-nbitq), 
to_sfixed(311693132.0/4294967296.0,1,-nbitq), 
to_sfixed(1290422429.0/4294967296.0,1,-nbitq), 
to_sfixed(187123074.0/4294967296.0,1,-nbitq), 
to_sfixed(-335767874.0/4294967296.0,1,-nbitq), 
to_sfixed(363482332.0/4294967296.0,1,-nbitq), 
to_sfixed(41097922.0/4294967296.0,1,-nbitq), 
to_sfixed(-392869039.0/4294967296.0,1,-nbitq), 
to_sfixed(51211958.0/4294967296.0,1,-nbitq), 
to_sfixed(-132313756.0/4294967296.0,1,-nbitq), 
to_sfixed(246313967.0/4294967296.0,1,-nbitq), 
to_sfixed(-500759242.0/4294967296.0,1,-nbitq), 
to_sfixed(162618010.0/4294967296.0,1,-nbitq), 
to_sfixed(-478166529.0/4294967296.0,1,-nbitq), 
to_sfixed(416222286.0/4294967296.0,1,-nbitq), 
to_sfixed(834451504.0/4294967296.0,1,-nbitq), 
to_sfixed(100193602.0/4294967296.0,1,-nbitq), 
to_sfixed(298932956.0/4294967296.0,1,-nbitq), 
to_sfixed(-478070258.0/4294967296.0,1,-nbitq), 
to_sfixed(-117677877.0/4294967296.0,1,-nbitq), 
to_sfixed(-338430942.0/4294967296.0,1,-nbitq), 
to_sfixed(364914958.0/4294967296.0,1,-nbitq), 
to_sfixed(-178292795.0/4294967296.0,1,-nbitq), 
to_sfixed(28397394.0/4294967296.0,1,-nbitq), 
to_sfixed(892744914.0/4294967296.0,1,-nbitq), 
to_sfixed(51813170.0/4294967296.0,1,-nbitq), 
to_sfixed(468915012.0/4294967296.0,1,-nbitq), 
to_sfixed(477861553.0/4294967296.0,1,-nbitq), 
to_sfixed(-40237318.0/4294967296.0,1,-nbitq), 
to_sfixed(846367280.0/4294967296.0,1,-nbitq), 
to_sfixed(-454347440.0/4294967296.0,1,-nbitq), 
to_sfixed(191103386.0/4294967296.0,1,-nbitq), 
to_sfixed(-49272971.0/4294967296.0,1,-nbitq), 
to_sfixed(-261953464.0/4294967296.0,1,-nbitq), 
to_sfixed(1344379759.0/4294967296.0,1,-nbitq), 
to_sfixed(938943510.0/4294967296.0,1,-nbitq), 
to_sfixed(174618206.0/4294967296.0,1,-nbitq), 
to_sfixed(-50346227.0/4294967296.0,1,-nbitq), 
to_sfixed(-141569331.0/4294967296.0,1,-nbitq), 
to_sfixed(250446689.0/4294967296.0,1,-nbitq), 
to_sfixed(-412261923.0/4294967296.0,1,-nbitq), 
to_sfixed(84425404.0/4294967296.0,1,-nbitq), 
to_sfixed(-68569444.0/4294967296.0,1,-nbitq), 
to_sfixed(-17396379.0/4294967296.0,1,-nbitq), 
to_sfixed(-177183558.0/4294967296.0,1,-nbitq), 
to_sfixed(504714264.0/4294967296.0,1,-nbitq), 
to_sfixed(1213406401.0/4294967296.0,1,-nbitq), 
to_sfixed(-457429902.0/4294967296.0,1,-nbitq), 
to_sfixed(9144838.0/4294967296.0,1,-nbitq), 
to_sfixed(-438004470.0/4294967296.0,1,-nbitq), 
to_sfixed(-19722903.0/4294967296.0,1,-nbitq), 
to_sfixed(155959808.0/4294967296.0,1,-nbitq), 
to_sfixed(-211025256.0/4294967296.0,1,-nbitq), 
to_sfixed(394774798.0/4294967296.0,1,-nbitq), 
to_sfixed(-540394119.0/4294967296.0,1,-nbitq), 
to_sfixed(-139924991.0/4294967296.0,1,-nbitq), 
to_sfixed(-299496996.0/4294967296.0,1,-nbitq), 
to_sfixed(-159027855.0/4294967296.0,1,-nbitq), 
to_sfixed(-60008398.0/4294967296.0,1,-nbitq), 
to_sfixed(1213423036.0/4294967296.0,1,-nbitq), 
to_sfixed(279174471.0/4294967296.0,1,-nbitq), 
to_sfixed(-541515030.0/4294967296.0,1,-nbitq), 
to_sfixed(917381291.0/4294967296.0,1,-nbitq), 
to_sfixed(144490038.0/4294967296.0,1,-nbitq), 
to_sfixed(635670685.0/4294967296.0,1,-nbitq), 
to_sfixed(-4662568.0/4294967296.0,1,-nbitq), 
to_sfixed(-157085148.0/4294967296.0,1,-nbitq), 
to_sfixed(-574863528.0/4294967296.0,1,-nbitq), 
to_sfixed(116984568.0/4294967296.0,1,-nbitq), 
to_sfixed(71532887.0/4294967296.0,1,-nbitq), 
to_sfixed(354982499.0/4294967296.0,1,-nbitq), 
to_sfixed(43753774.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(844448777.0/4294967296.0,1,-nbitq), 
to_sfixed(303614192.0/4294967296.0,1,-nbitq), 
to_sfixed(937461732.0/4294967296.0,1,-nbitq), 
to_sfixed(-74011873.0/4294967296.0,1,-nbitq), 
to_sfixed(-679256170.0/4294967296.0,1,-nbitq), 
to_sfixed(-661750766.0/4294967296.0,1,-nbitq), 
to_sfixed(258172614.0/4294967296.0,1,-nbitq), 
to_sfixed(-390803100.0/4294967296.0,1,-nbitq), 
to_sfixed(1257610203.0/4294967296.0,1,-nbitq), 
to_sfixed(315780042.0/4294967296.0,1,-nbitq), 
to_sfixed(589314057.0/4294967296.0,1,-nbitq), 
to_sfixed(-101284154.0/4294967296.0,1,-nbitq), 
to_sfixed(-830004706.0/4294967296.0,1,-nbitq), 
to_sfixed(1030783640.0/4294967296.0,1,-nbitq), 
to_sfixed(-380837377.0/4294967296.0,1,-nbitq), 
to_sfixed(-327175633.0/4294967296.0,1,-nbitq), 
to_sfixed(-429722181.0/4294967296.0,1,-nbitq), 
to_sfixed(-186753221.0/4294967296.0,1,-nbitq), 
to_sfixed(892753113.0/4294967296.0,1,-nbitq), 
to_sfixed(-3798083.0/4294967296.0,1,-nbitq), 
to_sfixed(85254805.0/4294967296.0,1,-nbitq), 
to_sfixed(-425912801.0/4294967296.0,1,-nbitq), 
to_sfixed(-390805949.0/4294967296.0,1,-nbitq), 
to_sfixed(333027064.0/4294967296.0,1,-nbitq), 
to_sfixed(302239722.0/4294967296.0,1,-nbitq), 
to_sfixed(367975062.0/4294967296.0,1,-nbitq), 
to_sfixed(-104398413.0/4294967296.0,1,-nbitq), 
to_sfixed(-99668735.0/4294967296.0,1,-nbitq), 
to_sfixed(-107276333.0/4294967296.0,1,-nbitq), 
to_sfixed(-714653727.0/4294967296.0,1,-nbitq), 
to_sfixed(91055287.0/4294967296.0,1,-nbitq), 
to_sfixed(-890813092.0/4294967296.0,1,-nbitq), 
to_sfixed(944928239.0/4294967296.0,1,-nbitq), 
to_sfixed(-191594280.0/4294967296.0,1,-nbitq), 
to_sfixed(432106162.0/4294967296.0,1,-nbitq), 
to_sfixed(402500681.0/4294967296.0,1,-nbitq), 
to_sfixed(-68736313.0/4294967296.0,1,-nbitq), 
to_sfixed(538575362.0/4294967296.0,1,-nbitq), 
to_sfixed(-136349179.0/4294967296.0,1,-nbitq), 
to_sfixed(-211835200.0/4294967296.0,1,-nbitq), 
to_sfixed(-132028404.0/4294967296.0,1,-nbitq), 
to_sfixed(-735615334.0/4294967296.0,1,-nbitq), 
to_sfixed(1050354000.0/4294967296.0,1,-nbitq), 
to_sfixed(1414646444.0/4294967296.0,1,-nbitq), 
to_sfixed(585707290.0/4294967296.0,1,-nbitq), 
to_sfixed(613411706.0/4294967296.0,1,-nbitq), 
to_sfixed(-37137896.0/4294967296.0,1,-nbitq), 
to_sfixed(765393398.0/4294967296.0,1,-nbitq), 
to_sfixed(-341915167.0/4294967296.0,1,-nbitq), 
to_sfixed(-30807926.0/4294967296.0,1,-nbitq), 
to_sfixed(23838473.0/4294967296.0,1,-nbitq), 
to_sfixed(229488691.0/4294967296.0,1,-nbitq), 
to_sfixed(-938983022.0/4294967296.0,1,-nbitq), 
to_sfixed(717962909.0/4294967296.0,1,-nbitq), 
to_sfixed(1223926095.0/4294967296.0,1,-nbitq), 
to_sfixed(-757576633.0/4294967296.0,1,-nbitq), 
to_sfixed(-301718851.0/4294967296.0,1,-nbitq), 
to_sfixed(111789044.0/4294967296.0,1,-nbitq), 
to_sfixed(218500929.0/4294967296.0,1,-nbitq), 
to_sfixed(276049855.0/4294967296.0,1,-nbitq), 
to_sfixed(-330811116.0/4294967296.0,1,-nbitq), 
to_sfixed(653773844.0/4294967296.0,1,-nbitq), 
to_sfixed(-1221511020.0/4294967296.0,1,-nbitq), 
to_sfixed(-457658928.0/4294967296.0,1,-nbitq), 
to_sfixed(164555411.0/4294967296.0,1,-nbitq), 
to_sfixed(-34707766.0/4294967296.0,1,-nbitq), 
to_sfixed(-744516837.0/4294967296.0,1,-nbitq), 
to_sfixed(1053740068.0/4294967296.0,1,-nbitq), 
to_sfixed(-318483307.0/4294967296.0,1,-nbitq), 
to_sfixed(-657251922.0/4294967296.0,1,-nbitq), 
to_sfixed(132471760.0/4294967296.0,1,-nbitq), 
to_sfixed(-199033614.0/4294967296.0,1,-nbitq), 
to_sfixed(682745909.0/4294967296.0,1,-nbitq), 
to_sfixed(288791350.0/4294967296.0,1,-nbitq), 
to_sfixed(-174536529.0/4294967296.0,1,-nbitq), 
to_sfixed(-245153489.0/4294967296.0,1,-nbitq), 
to_sfixed(216605325.0/4294967296.0,1,-nbitq), 
to_sfixed(-135621669.0/4294967296.0,1,-nbitq), 
to_sfixed(48057697.0/4294967296.0,1,-nbitq), 
to_sfixed(-46076649.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(614567023.0/4294967296.0,1,-nbitq), 
to_sfixed(669216696.0/4294967296.0,1,-nbitq), 
to_sfixed(488399963.0/4294967296.0,1,-nbitq), 
to_sfixed(-140333630.0/4294967296.0,1,-nbitq), 
to_sfixed(-1009460724.0/4294967296.0,1,-nbitq), 
to_sfixed(-612847220.0/4294967296.0,1,-nbitq), 
to_sfixed(-289060727.0/4294967296.0,1,-nbitq), 
to_sfixed(132014382.0/4294967296.0,1,-nbitq), 
to_sfixed(945882673.0/4294967296.0,1,-nbitq), 
to_sfixed(90156655.0/4294967296.0,1,-nbitq), 
to_sfixed(947734105.0/4294967296.0,1,-nbitq), 
to_sfixed(-207215020.0/4294967296.0,1,-nbitq), 
to_sfixed(-816382961.0/4294967296.0,1,-nbitq), 
to_sfixed(1204603632.0/4294967296.0,1,-nbitq), 
to_sfixed(49920162.0/4294967296.0,1,-nbitq), 
to_sfixed(-225109235.0/4294967296.0,1,-nbitq), 
to_sfixed(193035784.0/4294967296.0,1,-nbitq), 
to_sfixed(-159449050.0/4294967296.0,1,-nbitq), 
to_sfixed(875819960.0/4294967296.0,1,-nbitq), 
to_sfixed(65611675.0/4294967296.0,1,-nbitq), 
to_sfixed(-228515482.0/4294967296.0,1,-nbitq), 
to_sfixed(-583955655.0/4294967296.0,1,-nbitq), 
to_sfixed(-56718129.0/4294967296.0,1,-nbitq), 
to_sfixed(353297531.0/4294967296.0,1,-nbitq), 
to_sfixed(363152358.0/4294967296.0,1,-nbitq), 
to_sfixed(-355242619.0/4294967296.0,1,-nbitq), 
to_sfixed(233003052.0/4294967296.0,1,-nbitq), 
to_sfixed(152728045.0/4294967296.0,1,-nbitq), 
to_sfixed(39158312.0/4294967296.0,1,-nbitq), 
to_sfixed(-258078652.0/4294967296.0,1,-nbitq), 
to_sfixed(-90041659.0/4294967296.0,1,-nbitq), 
to_sfixed(47725422.0/4294967296.0,1,-nbitq), 
to_sfixed(169542532.0/4294967296.0,1,-nbitq), 
to_sfixed(-427702642.0/4294967296.0,1,-nbitq), 
to_sfixed(90321021.0/4294967296.0,1,-nbitq), 
to_sfixed(440584150.0/4294967296.0,1,-nbitq), 
to_sfixed(-477393460.0/4294967296.0,1,-nbitq), 
to_sfixed(742207581.0/4294967296.0,1,-nbitq), 
to_sfixed(-433495476.0/4294967296.0,1,-nbitq), 
to_sfixed(-57784822.0/4294967296.0,1,-nbitq), 
to_sfixed(306500366.0/4294967296.0,1,-nbitq), 
to_sfixed(-758899744.0/4294967296.0,1,-nbitq), 
to_sfixed(1102698834.0/4294967296.0,1,-nbitq), 
to_sfixed(1509323169.0/4294967296.0,1,-nbitq), 
to_sfixed(62189308.0/4294967296.0,1,-nbitq), 
to_sfixed(279924119.0/4294967296.0,1,-nbitq), 
to_sfixed(-336863212.0/4294967296.0,1,-nbitq), 
to_sfixed(566796326.0/4294967296.0,1,-nbitq), 
to_sfixed(-437411096.0/4294967296.0,1,-nbitq), 
to_sfixed(249183296.0/4294967296.0,1,-nbitq), 
to_sfixed(356608901.0/4294967296.0,1,-nbitq), 
to_sfixed(443638991.0/4294967296.0,1,-nbitq), 
to_sfixed(-212276696.0/4294967296.0,1,-nbitq), 
to_sfixed(418806738.0/4294967296.0,1,-nbitq), 
to_sfixed(1140053348.0/4294967296.0,1,-nbitq), 
to_sfixed(-565544858.0/4294967296.0,1,-nbitq), 
to_sfixed(191244628.0/4294967296.0,1,-nbitq), 
to_sfixed(-552125173.0/4294967296.0,1,-nbitq), 
to_sfixed(391303536.0/4294967296.0,1,-nbitq), 
to_sfixed(42614476.0/4294967296.0,1,-nbitq), 
to_sfixed(305870511.0/4294967296.0,1,-nbitq), 
to_sfixed(430998736.0/4294967296.0,1,-nbitq), 
to_sfixed(-560671805.0/4294967296.0,1,-nbitq), 
to_sfixed(-477869715.0/4294967296.0,1,-nbitq), 
to_sfixed(-219411820.0/4294967296.0,1,-nbitq), 
to_sfixed(-138083580.0/4294967296.0,1,-nbitq), 
to_sfixed(-68191031.0/4294967296.0,1,-nbitq), 
to_sfixed(1847697517.0/4294967296.0,1,-nbitq), 
to_sfixed(-901919.0/4294967296.0,1,-nbitq), 
to_sfixed(-386414490.0/4294967296.0,1,-nbitq), 
to_sfixed(574457877.0/4294967296.0,1,-nbitq), 
to_sfixed(157386465.0/4294967296.0,1,-nbitq), 
to_sfixed(535078719.0/4294967296.0,1,-nbitq), 
to_sfixed(-8506096.0/4294967296.0,1,-nbitq), 
to_sfixed(333395991.0/4294967296.0,1,-nbitq), 
to_sfixed(89013607.0/4294967296.0,1,-nbitq), 
to_sfixed(-19817320.0/4294967296.0,1,-nbitq), 
to_sfixed(52040382.0/4294967296.0,1,-nbitq), 
to_sfixed(697139951.0/4294967296.0,1,-nbitq), 
to_sfixed(-67011983.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-82994290.0/4294967296.0,1,-nbitq), 
to_sfixed(905147035.0/4294967296.0,1,-nbitq), 
to_sfixed(346070323.0/4294967296.0,1,-nbitq), 
to_sfixed(122956796.0/4294967296.0,1,-nbitq), 
to_sfixed(-296707983.0/4294967296.0,1,-nbitq), 
to_sfixed(-242426693.0/4294967296.0,1,-nbitq), 
to_sfixed(128747772.0/4294967296.0,1,-nbitq), 
to_sfixed(-68827382.0/4294967296.0,1,-nbitq), 
to_sfixed(680833511.0/4294967296.0,1,-nbitq), 
to_sfixed(240045168.0/4294967296.0,1,-nbitq), 
to_sfixed(826205588.0/4294967296.0,1,-nbitq), 
to_sfixed(282389555.0/4294967296.0,1,-nbitq), 
to_sfixed(-14978606.0/4294967296.0,1,-nbitq), 
to_sfixed(1275500364.0/4294967296.0,1,-nbitq), 
to_sfixed(-458823307.0/4294967296.0,1,-nbitq), 
to_sfixed(-315755930.0/4294967296.0,1,-nbitq), 
to_sfixed(285880644.0/4294967296.0,1,-nbitq), 
to_sfixed(-298669314.0/4294967296.0,1,-nbitq), 
to_sfixed(1370901002.0/4294967296.0,1,-nbitq), 
to_sfixed(-323211964.0/4294967296.0,1,-nbitq), 
to_sfixed(170079001.0/4294967296.0,1,-nbitq), 
to_sfixed(-602760628.0/4294967296.0,1,-nbitq), 
to_sfixed(583122470.0/4294967296.0,1,-nbitq), 
to_sfixed(807923547.0/4294967296.0,1,-nbitq), 
to_sfixed(9026815.0/4294967296.0,1,-nbitq), 
to_sfixed(-657598679.0/4294967296.0,1,-nbitq), 
to_sfixed(88409851.0/4294967296.0,1,-nbitq), 
to_sfixed(686779560.0/4294967296.0,1,-nbitq), 
to_sfixed(-307201264.0/4294967296.0,1,-nbitq), 
to_sfixed(-696204390.0/4294967296.0,1,-nbitq), 
to_sfixed(-706636714.0/4294967296.0,1,-nbitq), 
to_sfixed(174480724.0/4294967296.0,1,-nbitq), 
to_sfixed(-152067893.0/4294967296.0,1,-nbitq), 
to_sfixed(-659810897.0/4294967296.0,1,-nbitq), 
to_sfixed(-590515549.0/4294967296.0,1,-nbitq), 
to_sfixed(259812245.0/4294967296.0,1,-nbitq), 
to_sfixed(-177043165.0/4294967296.0,1,-nbitq), 
to_sfixed(-131093713.0/4294967296.0,1,-nbitq), 
to_sfixed(88054760.0/4294967296.0,1,-nbitq), 
to_sfixed(201380722.0/4294967296.0,1,-nbitq), 
to_sfixed(549412753.0/4294967296.0,1,-nbitq), 
to_sfixed(37599879.0/4294967296.0,1,-nbitq), 
to_sfixed(201774626.0/4294967296.0,1,-nbitq), 
to_sfixed(1079969094.0/4294967296.0,1,-nbitq), 
to_sfixed(546752450.0/4294967296.0,1,-nbitq), 
to_sfixed(340232609.0/4294967296.0,1,-nbitq), 
to_sfixed(50646702.0/4294967296.0,1,-nbitq), 
to_sfixed(950635494.0/4294967296.0,1,-nbitq), 
to_sfixed(76020010.0/4294967296.0,1,-nbitq), 
to_sfixed(59230837.0/4294967296.0,1,-nbitq), 
to_sfixed(312595965.0/4294967296.0,1,-nbitq), 
to_sfixed(197235986.0/4294967296.0,1,-nbitq), 
to_sfixed(-713518750.0/4294967296.0,1,-nbitq), 
to_sfixed(92699756.0/4294967296.0,1,-nbitq), 
to_sfixed(402113350.0/4294967296.0,1,-nbitq), 
to_sfixed(-165945605.0/4294967296.0,1,-nbitq), 
to_sfixed(174744696.0/4294967296.0,1,-nbitq), 
to_sfixed(-433543326.0/4294967296.0,1,-nbitq), 
to_sfixed(-3400079.0/4294967296.0,1,-nbitq), 
to_sfixed(-68586657.0/4294967296.0,1,-nbitq), 
to_sfixed(163601547.0/4294967296.0,1,-nbitq), 
to_sfixed(388701778.0/4294967296.0,1,-nbitq), 
to_sfixed(186852285.0/4294967296.0,1,-nbitq), 
to_sfixed(-516235675.0/4294967296.0,1,-nbitq), 
to_sfixed(88076769.0/4294967296.0,1,-nbitq), 
to_sfixed(186605036.0/4294967296.0,1,-nbitq), 
to_sfixed(-384849712.0/4294967296.0,1,-nbitq), 
to_sfixed(1654457244.0/4294967296.0,1,-nbitq), 
to_sfixed(-167430228.0/4294967296.0,1,-nbitq), 
to_sfixed(-387713709.0/4294967296.0,1,-nbitq), 
to_sfixed(-453600823.0/4294967296.0,1,-nbitq), 
to_sfixed(323984656.0/4294967296.0,1,-nbitq), 
to_sfixed(150679050.0/4294967296.0,1,-nbitq), 
to_sfixed(184626963.0/4294967296.0,1,-nbitq), 
to_sfixed(-445233868.0/4294967296.0,1,-nbitq), 
to_sfixed(941881511.0/4294967296.0,1,-nbitq), 
to_sfixed(-909438691.0/4294967296.0,1,-nbitq), 
to_sfixed(127068166.0/4294967296.0,1,-nbitq), 
to_sfixed(280178759.0/4294967296.0,1,-nbitq), 
to_sfixed(236550037.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(84157247.0/4294967296.0,1,-nbitq), 
to_sfixed(521478369.0/4294967296.0,1,-nbitq), 
to_sfixed(-914085668.0/4294967296.0,1,-nbitq), 
to_sfixed(545859262.0/4294967296.0,1,-nbitq), 
to_sfixed(-778040102.0/4294967296.0,1,-nbitq), 
to_sfixed(277327581.0/4294967296.0,1,-nbitq), 
to_sfixed(66426665.0/4294967296.0,1,-nbitq), 
to_sfixed(-371463587.0/4294967296.0,1,-nbitq), 
to_sfixed(409771005.0/4294967296.0,1,-nbitq), 
to_sfixed(168562212.0/4294967296.0,1,-nbitq), 
to_sfixed(588420998.0/4294967296.0,1,-nbitq), 
to_sfixed(-196752333.0/4294967296.0,1,-nbitq), 
to_sfixed(-70754212.0/4294967296.0,1,-nbitq), 
to_sfixed(736845867.0/4294967296.0,1,-nbitq), 
to_sfixed(112613664.0/4294967296.0,1,-nbitq), 
to_sfixed(6812219.0/4294967296.0,1,-nbitq), 
to_sfixed(-101136861.0/4294967296.0,1,-nbitq), 
to_sfixed(-279257312.0/4294967296.0,1,-nbitq), 
to_sfixed(619646466.0/4294967296.0,1,-nbitq), 
to_sfixed(-136555149.0/4294967296.0,1,-nbitq), 
to_sfixed(40883697.0/4294967296.0,1,-nbitq), 
to_sfixed(-628921085.0/4294967296.0,1,-nbitq), 
to_sfixed(641301150.0/4294967296.0,1,-nbitq), 
to_sfixed(-72365298.0/4294967296.0,1,-nbitq), 
to_sfixed(-59786402.0/4294967296.0,1,-nbitq), 
to_sfixed(17410220.0/4294967296.0,1,-nbitq), 
to_sfixed(-630366601.0/4294967296.0,1,-nbitq), 
to_sfixed(523884136.0/4294967296.0,1,-nbitq), 
to_sfixed(-310593182.0/4294967296.0,1,-nbitq), 
to_sfixed(-158244228.0/4294967296.0,1,-nbitq), 
to_sfixed(-495934219.0/4294967296.0,1,-nbitq), 
to_sfixed(-392123969.0/4294967296.0,1,-nbitq), 
to_sfixed(-95374432.0/4294967296.0,1,-nbitq), 
to_sfixed(-448811816.0/4294967296.0,1,-nbitq), 
to_sfixed(553193494.0/4294967296.0,1,-nbitq), 
to_sfixed(-342313301.0/4294967296.0,1,-nbitq), 
to_sfixed(-253846121.0/4294967296.0,1,-nbitq), 
to_sfixed(556914571.0/4294967296.0,1,-nbitq), 
to_sfixed(130421700.0/4294967296.0,1,-nbitq), 
to_sfixed(-158342825.0/4294967296.0,1,-nbitq), 
to_sfixed(272736126.0/4294967296.0,1,-nbitq), 
to_sfixed(60254223.0/4294967296.0,1,-nbitq), 
to_sfixed(-12682829.0/4294967296.0,1,-nbitq), 
to_sfixed(1276927353.0/4294967296.0,1,-nbitq), 
to_sfixed(517707319.0/4294967296.0,1,-nbitq), 
to_sfixed(-146987258.0/4294967296.0,1,-nbitq), 
to_sfixed(-226040586.0/4294967296.0,1,-nbitq), 
to_sfixed(684361149.0/4294967296.0,1,-nbitq), 
to_sfixed(302717444.0/4294967296.0,1,-nbitq), 
to_sfixed(441308747.0/4294967296.0,1,-nbitq), 
to_sfixed(542771485.0/4294967296.0,1,-nbitq), 
to_sfixed(215641990.0/4294967296.0,1,-nbitq), 
to_sfixed(-398775195.0/4294967296.0,1,-nbitq), 
to_sfixed(269734833.0/4294967296.0,1,-nbitq), 
to_sfixed(65423954.0/4294967296.0,1,-nbitq), 
to_sfixed(416009182.0/4294967296.0,1,-nbitq), 
to_sfixed(-81260431.0/4294967296.0,1,-nbitq), 
to_sfixed(-343630498.0/4294967296.0,1,-nbitq), 
to_sfixed(259469278.0/4294967296.0,1,-nbitq), 
to_sfixed(-9449812.0/4294967296.0,1,-nbitq), 
to_sfixed(334584137.0/4294967296.0,1,-nbitq), 
to_sfixed(89528035.0/4294967296.0,1,-nbitq), 
to_sfixed(-2161460.0/4294967296.0,1,-nbitq), 
to_sfixed(-465276074.0/4294967296.0,1,-nbitq), 
to_sfixed(197573094.0/4294967296.0,1,-nbitq), 
to_sfixed(105083734.0/4294967296.0,1,-nbitq), 
to_sfixed(166497716.0/4294967296.0,1,-nbitq), 
to_sfixed(1211996704.0/4294967296.0,1,-nbitq), 
to_sfixed(260053458.0/4294967296.0,1,-nbitq), 
to_sfixed(-252427180.0/4294967296.0,1,-nbitq), 
to_sfixed(-739912116.0/4294967296.0,1,-nbitq), 
to_sfixed(-125154127.0/4294967296.0,1,-nbitq), 
to_sfixed(-232191699.0/4294967296.0,1,-nbitq), 
to_sfixed(-250803535.0/4294967296.0,1,-nbitq), 
to_sfixed(-525430145.0/4294967296.0,1,-nbitq), 
to_sfixed(576780742.0/4294967296.0,1,-nbitq), 
to_sfixed(-1430430866.0/4294967296.0,1,-nbitq), 
to_sfixed(260588666.0/4294967296.0,1,-nbitq), 
to_sfixed(159044930.0/4294967296.0,1,-nbitq), 
to_sfixed(-322002131.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-428869053.0/4294967296.0,1,-nbitq), 
to_sfixed(11238514.0/4294967296.0,1,-nbitq), 
to_sfixed(648775951.0/4294967296.0,1,-nbitq), 
to_sfixed(409209466.0/4294967296.0,1,-nbitq), 
to_sfixed(-653878759.0/4294967296.0,1,-nbitq), 
to_sfixed(629555379.0/4294967296.0,1,-nbitq), 
to_sfixed(-360868977.0/4294967296.0,1,-nbitq), 
to_sfixed(-484632465.0/4294967296.0,1,-nbitq), 
to_sfixed(184835707.0/4294967296.0,1,-nbitq), 
to_sfixed(398121268.0/4294967296.0,1,-nbitq), 
to_sfixed(106270278.0/4294967296.0,1,-nbitq), 
to_sfixed(689505182.0/4294967296.0,1,-nbitq), 
to_sfixed(-173740676.0/4294967296.0,1,-nbitq), 
to_sfixed(717993674.0/4294967296.0,1,-nbitq), 
to_sfixed(-332080666.0/4294967296.0,1,-nbitq), 
to_sfixed(-269138211.0/4294967296.0,1,-nbitq), 
to_sfixed(152917645.0/4294967296.0,1,-nbitq), 
to_sfixed(-2065189.0/4294967296.0,1,-nbitq), 
to_sfixed(827697071.0/4294967296.0,1,-nbitq), 
to_sfixed(-86747752.0/4294967296.0,1,-nbitq), 
to_sfixed(132406068.0/4294967296.0,1,-nbitq), 
to_sfixed(141540706.0/4294967296.0,1,-nbitq), 
to_sfixed(318457272.0/4294967296.0,1,-nbitq), 
to_sfixed(342729865.0/4294967296.0,1,-nbitq), 
to_sfixed(203271178.0/4294967296.0,1,-nbitq), 
to_sfixed(-147768547.0/4294967296.0,1,-nbitq), 
to_sfixed(-355337865.0/4294967296.0,1,-nbitq), 
to_sfixed(754788347.0/4294967296.0,1,-nbitq), 
to_sfixed(-136459199.0/4294967296.0,1,-nbitq), 
to_sfixed(139598244.0/4294967296.0,1,-nbitq), 
to_sfixed(102787085.0/4294967296.0,1,-nbitq), 
to_sfixed(-83436420.0/4294967296.0,1,-nbitq), 
to_sfixed(-154402444.0/4294967296.0,1,-nbitq), 
to_sfixed(-803858430.0/4294967296.0,1,-nbitq), 
to_sfixed(245958427.0/4294967296.0,1,-nbitq), 
to_sfixed(-268316924.0/4294967296.0,1,-nbitq), 
to_sfixed(-180886089.0/4294967296.0,1,-nbitq), 
to_sfixed(-306139362.0/4294967296.0,1,-nbitq), 
to_sfixed(240749071.0/4294967296.0,1,-nbitq), 
to_sfixed(-263139531.0/4294967296.0,1,-nbitq), 
to_sfixed(-92846254.0/4294967296.0,1,-nbitq), 
to_sfixed(219250935.0/4294967296.0,1,-nbitq), 
to_sfixed(358550192.0/4294967296.0,1,-nbitq), 
to_sfixed(540779633.0/4294967296.0,1,-nbitq), 
to_sfixed(824752791.0/4294967296.0,1,-nbitq), 
to_sfixed(186985824.0/4294967296.0,1,-nbitq), 
to_sfixed(-62845567.0/4294967296.0,1,-nbitq), 
to_sfixed(207383447.0/4294967296.0,1,-nbitq), 
to_sfixed(358201990.0/4294967296.0,1,-nbitq), 
to_sfixed(656238138.0/4294967296.0,1,-nbitq), 
to_sfixed(514083858.0/4294967296.0,1,-nbitq), 
to_sfixed(84097359.0/4294967296.0,1,-nbitq), 
to_sfixed(72522035.0/4294967296.0,1,-nbitq), 
to_sfixed(544970239.0/4294967296.0,1,-nbitq), 
to_sfixed(-296973022.0/4294967296.0,1,-nbitq), 
to_sfixed(759702311.0/4294967296.0,1,-nbitq), 
to_sfixed(-58786361.0/4294967296.0,1,-nbitq), 
to_sfixed(-1126517002.0/4294967296.0,1,-nbitq), 
to_sfixed(340318371.0/4294967296.0,1,-nbitq), 
to_sfixed(168667319.0/4294967296.0,1,-nbitq), 
to_sfixed(-71101527.0/4294967296.0,1,-nbitq), 
to_sfixed(-58024576.0/4294967296.0,1,-nbitq), 
to_sfixed(-98009865.0/4294967296.0,1,-nbitq), 
to_sfixed(-623566479.0/4294967296.0,1,-nbitq), 
to_sfixed(431214360.0/4294967296.0,1,-nbitq), 
to_sfixed(207015295.0/4294967296.0,1,-nbitq), 
to_sfixed(-104276685.0/4294967296.0,1,-nbitq), 
to_sfixed(492162170.0/4294967296.0,1,-nbitq), 
to_sfixed(282691168.0/4294967296.0,1,-nbitq), 
to_sfixed(289018461.0/4294967296.0,1,-nbitq), 
to_sfixed(-356907612.0/4294967296.0,1,-nbitq), 
to_sfixed(-4617715.0/4294967296.0,1,-nbitq), 
to_sfixed(-826310896.0/4294967296.0,1,-nbitq), 
to_sfixed(-2778781.0/4294967296.0,1,-nbitq), 
to_sfixed(28568123.0/4294967296.0,1,-nbitq), 
to_sfixed(369300718.0/4294967296.0,1,-nbitq), 
to_sfixed(-419653469.0/4294967296.0,1,-nbitq), 
to_sfixed(30179687.0/4294967296.0,1,-nbitq), 
to_sfixed(-58227962.0/4294967296.0,1,-nbitq), 
to_sfixed(294287020.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(282683222.0/4294967296.0,1,-nbitq), 
to_sfixed(165673433.0/4294967296.0,1,-nbitq), 
to_sfixed(606352900.0/4294967296.0,1,-nbitq), 
to_sfixed(500345263.0/4294967296.0,1,-nbitq), 
to_sfixed(-18474635.0/4294967296.0,1,-nbitq), 
to_sfixed(1149701369.0/4294967296.0,1,-nbitq), 
to_sfixed(398967250.0/4294967296.0,1,-nbitq), 
to_sfixed(150959593.0/4294967296.0,1,-nbitq), 
to_sfixed(-225898454.0/4294967296.0,1,-nbitq), 
to_sfixed(-149271162.0/4294967296.0,1,-nbitq), 
to_sfixed(-331501375.0/4294967296.0,1,-nbitq), 
to_sfixed(597417487.0/4294967296.0,1,-nbitq), 
to_sfixed(9217907.0/4294967296.0,1,-nbitq), 
to_sfixed(504249537.0/4294967296.0,1,-nbitq), 
to_sfixed(-309259543.0/4294967296.0,1,-nbitq), 
to_sfixed(254320247.0/4294967296.0,1,-nbitq), 
to_sfixed(-181013086.0/4294967296.0,1,-nbitq), 
to_sfixed(60702421.0/4294967296.0,1,-nbitq), 
to_sfixed(14973850.0/4294967296.0,1,-nbitq), 
to_sfixed(-321992514.0/4294967296.0,1,-nbitq), 
to_sfixed(349546478.0/4294967296.0,1,-nbitq), 
to_sfixed(263575453.0/4294967296.0,1,-nbitq), 
to_sfixed(10266953.0/4294967296.0,1,-nbitq), 
to_sfixed(34634266.0/4294967296.0,1,-nbitq), 
to_sfixed(-145302651.0/4294967296.0,1,-nbitq), 
to_sfixed(-41964133.0/4294967296.0,1,-nbitq), 
to_sfixed(-527199560.0/4294967296.0,1,-nbitq), 
to_sfixed(150042841.0/4294967296.0,1,-nbitq), 
to_sfixed(98703205.0/4294967296.0,1,-nbitq), 
to_sfixed(465083967.0/4294967296.0,1,-nbitq), 
to_sfixed(-51387453.0/4294967296.0,1,-nbitq), 
to_sfixed(-435931825.0/4294967296.0,1,-nbitq), 
to_sfixed(61811194.0/4294967296.0,1,-nbitq), 
to_sfixed(-638227299.0/4294967296.0,1,-nbitq), 
to_sfixed(75860391.0/4294967296.0,1,-nbitq), 
to_sfixed(-188878299.0/4294967296.0,1,-nbitq), 
to_sfixed(51088951.0/4294967296.0,1,-nbitq), 
to_sfixed(-431496533.0/4294967296.0,1,-nbitq), 
to_sfixed(369944456.0/4294967296.0,1,-nbitq), 
to_sfixed(174196406.0/4294967296.0,1,-nbitq), 
to_sfixed(170843337.0/4294967296.0,1,-nbitq), 
to_sfixed(746150982.0/4294967296.0,1,-nbitq), 
to_sfixed(17312265.0/4294967296.0,1,-nbitq), 
to_sfixed(384789043.0/4294967296.0,1,-nbitq), 
to_sfixed(-28287940.0/4294967296.0,1,-nbitq), 
to_sfixed(-88020673.0/4294967296.0,1,-nbitq), 
to_sfixed(224194141.0/4294967296.0,1,-nbitq), 
to_sfixed(-297282846.0/4294967296.0,1,-nbitq), 
to_sfixed(68975055.0/4294967296.0,1,-nbitq), 
to_sfixed(164877430.0/4294967296.0,1,-nbitq), 
to_sfixed(454201175.0/4294967296.0,1,-nbitq), 
to_sfixed(-121321399.0/4294967296.0,1,-nbitq), 
to_sfixed(-344262397.0/4294967296.0,1,-nbitq), 
to_sfixed(650773663.0/4294967296.0,1,-nbitq), 
to_sfixed(85278212.0/4294967296.0,1,-nbitq), 
to_sfixed(506913628.0/4294967296.0,1,-nbitq), 
to_sfixed(229085232.0/4294967296.0,1,-nbitq), 
to_sfixed(-822290826.0/4294967296.0,1,-nbitq), 
to_sfixed(-85268554.0/4294967296.0,1,-nbitq), 
to_sfixed(-1363953.0/4294967296.0,1,-nbitq), 
to_sfixed(-73811141.0/4294967296.0,1,-nbitq), 
to_sfixed(166854505.0/4294967296.0,1,-nbitq), 
to_sfixed(-223552033.0/4294967296.0,1,-nbitq), 
to_sfixed(-57601317.0/4294967296.0,1,-nbitq), 
to_sfixed(423226382.0/4294967296.0,1,-nbitq), 
to_sfixed(-214369912.0/4294967296.0,1,-nbitq), 
to_sfixed(-470839913.0/4294967296.0,1,-nbitq), 
to_sfixed(285884665.0/4294967296.0,1,-nbitq), 
to_sfixed(-62829291.0/4294967296.0,1,-nbitq), 
to_sfixed(265128411.0/4294967296.0,1,-nbitq), 
to_sfixed(-382657048.0/4294967296.0,1,-nbitq), 
to_sfixed(456527020.0/4294967296.0,1,-nbitq), 
to_sfixed(-352137428.0/4294967296.0,1,-nbitq), 
to_sfixed(137100502.0/4294967296.0,1,-nbitq), 
to_sfixed(168789100.0/4294967296.0,1,-nbitq), 
to_sfixed(161127757.0/4294967296.0,1,-nbitq), 
to_sfixed(-194111153.0/4294967296.0,1,-nbitq), 
to_sfixed(66882059.0/4294967296.0,1,-nbitq), 
to_sfixed(-338902236.0/4294967296.0,1,-nbitq), 
to_sfixed(63284635.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-170642506.0/4294967296.0,1,-nbitq), 
to_sfixed(200703583.0/4294967296.0,1,-nbitq), 
to_sfixed(727085265.0/4294967296.0,1,-nbitq), 
to_sfixed(213367757.0/4294967296.0,1,-nbitq), 
to_sfixed(163977993.0/4294967296.0,1,-nbitq), 
to_sfixed(170973205.0/4294967296.0,1,-nbitq), 
to_sfixed(5725136.0/4294967296.0,1,-nbitq), 
to_sfixed(138418663.0/4294967296.0,1,-nbitq), 
to_sfixed(17641506.0/4294967296.0,1,-nbitq), 
to_sfixed(7779998.0/4294967296.0,1,-nbitq), 
to_sfixed(73666070.0/4294967296.0,1,-nbitq), 
to_sfixed(155336910.0/4294967296.0,1,-nbitq), 
to_sfixed(-383166685.0/4294967296.0,1,-nbitq), 
to_sfixed(282302995.0/4294967296.0,1,-nbitq), 
to_sfixed(354171036.0/4294967296.0,1,-nbitq), 
to_sfixed(102783928.0/4294967296.0,1,-nbitq), 
to_sfixed(59860978.0/4294967296.0,1,-nbitq), 
to_sfixed(82661543.0/4294967296.0,1,-nbitq), 
to_sfixed(444620239.0/4294967296.0,1,-nbitq), 
to_sfixed(-154834677.0/4294967296.0,1,-nbitq), 
to_sfixed(-361250934.0/4294967296.0,1,-nbitq), 
to_sfixed(333134999.0/4294967296.0,1,-nbitq), 
to_sfixed(-76659442.0/4294967296.0,1,-nbitq), 
to_sfixed(372451955.0/4294967296.0,1,-nbitq), 
to_sfixed(135005221.0/4294967296.0,1,-nbitq), 
to_sfixed(-299403841.0/4294967296.0,1,-nbitq), 
to_sfixed(60303618.0/4294967296.0,1,-nbitq), 
to_sfixed(89546764.0/4294967296.0,1,-nbitq), 
to_sfixed(-41099254.0/4294967296.0,1,-nbitq), 
to_sfixed(569033580.0/4294967296.0,1,-nbitq), 
to_sfixed(148088319.0/4294967296.0,1,-nbitq), 
to_sfixed(-367411354.0/4294967296.0,1,-nbitq), 
to_sfixed(484434638.0/4294967296.0,1,-nbitq), 
to_sfixed(335328730.0/4294967296.0,1,-nbitq), 
to_sfixed(244743537.0/4294967296.0,1,-nbitq), 
to_sfixed(-448952592.0/4294967296.0,1,-nbitq), 
to_sfixed(-219505046.0/4294967296.0,1,-nbitq), 
to_sfixed(-30230502.0/4294967296.0,1,-nbitq), 
to_sfixed(266961838.0/4294967296.0,1,-nbitq), 
to_sfixed(-135017609.0/4294967296.0,1,-nbitq), 
to_sfixed(-22286108.0/4294967296.0,1,-nbitq), 
to_sfixed(4072862.0/4294967296.0,1,-nbitq), 
to_sfixed(491840685.0/4294967296.0,1,-nbitq), 
to_sfixed(-285770780.0/4294967296.0,1,-nbitq), 
to_sfixed(-76138581.0/4294967296.0,1,-nbitq), 
to_sfixed(-52322378.0/4294967296.0,1,-nbitq), 
to_sfixed(-184896320.0/4294967296.0,1,-nbitq), 
to_sfixed(70105853.0/4294967296.0,1,-nbitq), 
to_sfixed(27141337.0/4294967296.0,1,-nbitq), 
to_sfixed(-264210162.0/4294967296.0,1,-nbitq), 
to_sfixed(105066791.0/4294967296.0,1,-nbitq), 
to_sfixed(208250475.0/4294967296.0,1,-nbitq), 
to_sfixed(85474486.0/4294967296.0,1,-nbitq), 
to_sfixed(466541218.0/4294967296.0,1,-nbitq), 
to_sfixed(-112071244.0/4294967296.0,1,-nbitq), 
to_sfixed(-144254348.0/4294967296.0,1,-nbitq), 
to_sfixed(285194564.0/4294967296.0,1,-nbitq), 
to_sfixed(-752202061.0/4294967296.0,1,-nbitq), 
to_sfixed(122636489.0/4294967296.0,1,-nbitq), 
to_sfixed(-198553896.0/4294967296.0,1,-nbitq), 
to_sfixed(367657235.0/4294967296.0,1,-nbitq), 
to_sfixed(408992050.0/4294967296.0,1,-nbitq), 
to_sfixed(97511929.0/4294967296.0,1,-nbitq), 
to_sfixed(85009543.0/4294967296.0,1,-nbitq), 
to_sfixed(233702424.0/4294967296.0,1,-nbitq), 
to_sfixed(-327712579.0/4294967296.0,1,-nbitq), 
to_sfixed(-342776221.0/4294967296.0,1,-nbitq), 
to_sfixed(-22062341.0/4294967296.0,1,-nbitq), 
to_sfixed(183675005.0/4294967296.0,1,-nbitq), 
to_sfixed(134757172.0/4294967296.0,1,-nbitq), 
to_sfixed(-152136481.0/4294967296.0,1,-nbitq), 
to_sfixed(-167210473.0/4294967296.0,1,-nbitq), 
to_sfixed(-419244975.0/4294967296.0,1,-nbitq), 
to_sfixed(325285589.0/4294967296.0,1,-nbitq), 
to_sfixed(-2324176.0/4294967296.0,1,-nbitq), 
to_sfixed(-37849237.0/4294967296.0,1,-nbitq), 
to_sfixed(176457629.0/4294967296.0,1,-nbitq), 
to_sfixed(279454673.0/4294967296.0,1,-nbitq), 
to_sfixed(239742582.0/4294967296.0,1,-nbitq), 
to_sfixed(203417102.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(65291120.0/4294967296.0,1,-nbitq), 
to_sfixed(-247075668.0/4294967296.0,1,-nbitq), 
to_sfixed(667587434.0/4294967296.0,1,-nbitq), 
to_sfixed(-256004990.0/4294967296.0,1,-nbitq), 
to_sfixed(22549530.0/4294967296.0,1,-nbitq), 
to_sfixed(-544823477.0/4294967296.0,1,-nbitq), 
to_sfixed(-16356700.0/4294967296.0,1,-nbitq), 
to_sfixed(154329331.0/4294967296.0,1,-nbitq), 
to_sfixed(-316575789.0/4294967296.0,1,-nbitq), 
to_sfixed(34793089.0/4294967296.0,1,-nbitq), 
to_sfixed(237151214.0/4294967296.0,1,-nbitq), 
to_sfixed(55190871.0/4294967296.0,1,-nbitq), 
to_sfixed(76538416.0/4294967296.0,1,-nbitq), 
to_sfixed(190543513.0/4294967296.0,1,-nbitq), 
to_sfixed(114089425.0/4294967296.0,1,-nbitq), 
to_sfixed(203983067.0/4294967296.0,1,-nbitq), 
to_sfixed(197699764.0/4294967296.0,1,-nbitq), 
to_sfixed(-314029705.0/4294967296.0,1,-nbitq), 
to_sfixed(260430881.0/4294967296.0,1,-nbitq), 
to_sfixed(157240537.0/4294967296.0,1,-nbitq), 
to_sfixed(-393983345.0/4294967296.0,1,-nbitq), 
to_sfixed(2691925.0/4294967296.0,1,-nbitq), 
to_sfixed(413612950.0/4294967296.0,1,-nbitq), 
to_sfixed(-26776973.0/4294967296.0,1,-nbitq), 
to_sfixed(27481712.0/4294967296.0,1,-nbitq), 
to_sfixed(-3213395.0/4294967296.0,1,-nbitq), 
to_sfixed(37407649.0/4294967296.0,1,-nbitq), 
to_sfixed(-98916160.0/4294967296.0,1,-nbitq), 
to_sfixed(162421111.0/4294967296.0,1,-nbitq), 
to_sfixed(404685834.0/4294967296.0,1,-nbitq), 
to_sfixed(-160310160.0/4294967296.0,1,-nbitq), 
to_sfixed(-163596891.0/4294967296.0,1,-nbitq), 
to_sfixed(385770995.0/4294967296.0,1,-nbitq), 
to_sfixed(-240472969.0/4294967296.0,1,-nbitq), 
to_sfixed(443860988.0/4294967296.0,1,-nbitq), 
to_sfixed(-312577859.0/4294967296.0,1,-nbitq), 
to_sfixed(50365241.0/4294967296.0,1,-nbitq), 
to_sfixed(-340520158.0/4294967296.0,1,-nbitq), 
to_sfixed(-105461859.0/4294967296.0,1,-nbitq), 
to_sfixed(298314218.0/4294967296.0,1,-nbitq), 
to_sfixed(-183312836.0/4294967296.0,1,-nbitq), 
to_sfixed(238014844.0/4294967296.0,1,-nbitq), 
to_sfixed(238811395.0/4294967296.0,1,-nbitq), 
to_sfixed(284652657.0/4294967296.0,1,-nbitq), 
to_sfixed(399146542.0/4294967296.0,1,-nbitq), 
to_sfixed(155478449.0/4294967296.0,1,-nbitq), 
to_sfixed(-340829410.0/4294967296.0,1,-nbitq), 
to_sfixed(249098910.0/4294967296.0,1,-nbitq), 
to_sfixed(28896290.0/4294967296.0,1,-nbitq), 
to_sfixed(-153129413.0/4294967296.0,1,-nbitq), 
to_sfixed(432937528.0/4294967296.0,1,-nbitq), 
to_sfixed(340155102.0/4294967296.0,1,-nbitq), 
to_sfixed(-110863555.0/4294967296.0,1,-nbitq), 
to_sfixed(-244748954.0/4294967296.0,1,-nbitq), 
to_sfixed(-45233600.0/4294967296.0,1,-nbitq), 
to_sfixed(69085146.0/4294967296.0,1,-nbitq), 
to_sfixed(265373026.0/4294967296.0,1,-nbitq), 
to_sfixed(-386716992.0/4294967296.0,1,-nbitq), 
to_sfixed(-302009989.0/4294967296.0,1,-nbitq), 
to_sfixed(68125717.0/4294967296.0,1,-nbitq), 
to_sfixed(-170621658.0/4294967296.0,1,-nbitq), 
to_sfixed(-130694282.0/4294967296.0,1,-nbitq), 
to_sfixed(-110629114.0/4294967296.0,1,-nbitq), 
to_sfixed(-110891153.0/4294967296.0,1,-nbitq), 
to_sfixed(-243791228.0/4294967296.0,1,-nbitq), 
to_sfixed(140814477.0/4294967296.0,1,-nbitq), 
to_sfixed(-42769370.0/4294967296.0,1,-nbitq), 
to_sfixed(-312415511.0/4294967296.0,1,-nbitq), 
to_sfixed(-182947830.0/4294967296.0,1,-nbitq), 
to_sfixed(21858421.0/4294967296.0,1,-nbitq), 
to_sfixed(89011857.0/4294967296.0,1,-nbitq), 
to_sfixed(149481302.0/4294967296.0,1,-nbitq), 
to_sfixed(-168116241.0/4294967296.0,1,-nbitq), 
to_sfixed(315336018.0/4294967296.0,1,-nbitq), 
to_sfixed(-44586246.0/4294967296.0,1,-nbitq), 
to_sfixed(-241409056.0/4294967296.0,1,-nbitq), 
to_sfixed(157637411.0/4294967296.0,1,-nbitq), 
to_sfixed(157935351.0/4294967296.0,1,-nbitq), 
to_sfixed(16955195.0/4294967296.0,1,-nbitq), 
to_sfixed(316242689.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-227539995.0/4294967296.0,1,-nbitq), 
to_sfixed(-458779129.0/4294967296.0,1,-nbitq), 
to_sfixed(119912141.0/4294967296.0,1,-nbitq), 
to_sfixed(-168858703.0/4294967296.0,1,-nbitq), 
to_sfixed(316592559.0/4294967296.0,1,-nbitq), 
to_sfixed(180852753.0/4294967296.0,1,-nbitq), 
to_sfixed(12481817.0/4294967296.0,1,-nbitq), 
to_sfixed(-207008291.0/4294967296.0,1,-nbitq), 
to_sfixed(-87811600.0/4294967296.0,1,-nbitq), 
to_sfixed(204015085.0/4294967296.0,1,-nbitq), 
to_sfixed(-262790581.0/4294967296.0,1,-nbitq), 
to_sfixed(449619057.0/4294967296.0,1,-nbitq), 
to_sfixed(-603106286.0/4294967296.0,1,-nbitq), 
to_sfixed(-67997888.0/4294967296.0,1,-nbitq), 
to_sfixed(-193650826.0/4294967296.0,1,-nbitq), 
to_sfixed(-142300852.0/4294967296.0,1,-nbitq), 
to_sfixed(-227687552.0/4294967296.0,1,-nbitq), 
to_sfixed(39183066.0/4294967296.0,1,-nbitq), 
to_sfixed(-357597540.0/4294967296.0,1,-nbitq), 
to_sfixed(-44342422.0/4294967296.0,1,-nbitq), 
to_sfixed(-215547396.0/4294967296.0,1,-nbitq), 
to_sfixed(546214208.0/4294967296.0,1,-nbitq), 
to_sfixed(473560751.0/4294967296.0,1,-nbitq), 
to_sfixed(390080007.0/4294967296.0,1,-nbitq), 
to_sfixed(370642226.0/4294967296.0,1,-nbitq), 
to_sfixed(-157321556.0/4294967296.0,1,-nbitq), 
to_sfixed(-266617812.0/4294967296.0,1,-nbitq), 
to_sfixed(-277452583.0/4294967296.0,1,-nbitq), 
to_sfixed(-223101810.0/4294967296.0,1,-nbitq), 
to_sfixed(86918862.0/4294967296.0,1,-nbitq), 
to_sfixed(115422959.0/4294967296.0,1,-nbitq), 
to_sfixed(-520847025.0/4294967296.0,1,-nbitq), 
to_sfixed(311457011.0/4294967296.0,1,-nbitq), 
to_sfixed(-478130248.0/4294967296.0,1,-nbitq), 
to_sfixed(193622630.0/4294967296.0,1,-nbitq), 
to_sfixed(-135476955.0/4294967296.0,1,-nbitq), 
to_sfixed(155162116.0/4294967296.0,1,-nbitq), 
to_sfixed(51255605.0/4294967296.0,1,-nbitq), 
to_sfixed(-68619542.0/4294967296.0,1,-nbitq), 
to_sfixed(474390507.0/4294967296.0,1,-nbitq), 
to_sfixed(138805546.0/4294967296.0,1,-nbitq), 
to_sfixed(171545769.0/4294967296.0,1,-nbitq), 
to_sfixed(432999207.0/4294967296.0,1,-nbitq), 
to_sfixed(-97467999.0/4294967296.0,1,-nbitq), 
to_sfixed(477129.0/4294967296.0,1,-nbitq), 
to_sfixed(-2730047.0/4294967296.0,1,-nbitq), 
to_sfixed(-194040003.0/4294967296.0,1,-nbitq), 
to_sfixed(102378228.0/4294967296.0,1,-nbitq), 
to_sfixed(-159185421.0/4294967296.0,1,-nbitq), 
to_sfixed(87183330.0/4294967296.0,1,-nbitq), 
to_sfixed(-263486998.0/4294967296.0,1,-nbitq), 
to_sfixed(45477436.0/4294967296.0,1,-nbitq), 
to_sfixed(-468787188.0/4294967296.0,1,-nbitq), 
to_sfixed(328653580.0/4294967296.0,1,-nbitq), 
to_sfixed(-190956613.0/4294967296.0,1,-nbitq), 
to_sfixed(192671013.0/4294967296.0,1,-nbitq), 
to_sfixed(-130005009.0/4294967296.0,1,-nbitq), 
to_sfixed(62435129.0/4294967296.0,1,-nbitq), 
to_sfixed(183130186.0/4294967296.0,1,-nbitq), 
to_sfixed(-273876230.0/4294967296.0,1,-nbitq), 
to_sfixed(383745816.0/4294967296.0,1,-nbitq), 
to_sfixed(9353634.0/4294967296.0,1,-nbitq), 
to_sfixed(-384185329.0/4294967296.0,1,-nbitq), 
to_sfixed(-26031293.0/4294967296.0,1,-nbitq), 
to_sfixed(-265553604.0/4294967296.0,1,-nbitq), 
to_sfixed(46919166.0/4294967296.0,1,-nbitq), 
to_sfixed(6400859.0/4294967296.0,1,-nbitq), 
to_sfixed(-53450099.0/4294967296.0,1,-nbitq), 
to_sfixed(310237173.0/4294967296.0,1,-nbitq), 
to_sfixed(50382562.0/4294967296.0,1,-nbitq), 
to_sfixed(-134075339.0/4294967296.0,1,-nbitq), 
to_sfixed(-145367559.0/4294967296.0,1,-nbitq), 
to_sfixed(-645357982.0/4294967296.0,1,-nbitq), 
to_sfixed(400423000.0/4294967296.0,1,-nbitq), 
to_sfixed(329226885.0/4294967296.0,1,-nbitq), 
to_sfixed(-557250523.0/4294967296.0,1,-nbitq), 
to_sfixed(-94291276.0/4294967296.0,1,-nbitq), 
to_sfixed(222240938.0/4294967296.0,1,-nbitq), 
to_sfixed(-509066405.0/4294967296.0,1,-nbitq), 
to_sfixed(-130901694.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(10980949.0/4294967296.0,1,-nbitq), 
to_sfixed(148681416.0/4294967296.0,1,-nbitq), 
to_sfixed(197509062.0/4294967296.0,1,-nbitq), 
to_sfixed(-23767544.0/4294967296.0,1,-nbitq), 
to_sfixed(68436049.0/4294967296.0,1,-nbitq), 
to_sfixed(-234523443.0/4294967296.0,1,-nbitq), 
to_sfixed(231573009.0/4294967296.0,1,-nbitq), 
to_sfixed(-18287458.0/4294967296.0,1,-nbitq), 
to_sfixed(-28981410.0/4294967296.0,1,-nbitq), 
to_sfixed(-72732819.0/4294967296.0,1,-nbitq), 
to_sfixed(128942039.0/4294967296.0,1,-nbitq), 
to_sfixed(579719016.0/4294967296.0,1,-nbitq), 
to_sfixed(145787333.0/4294967296.0,1,-nbitq), 
to_sfixed(-138076811.0/4294967296.0,1,-nbitq), 
to_sfixed(303240432.0/4294967296.0,1,-nbitq), 
to_sfixed(278750059.0/4294967296.0,1,-nbitq), 
to_sfixed(-255581199.0/4294967296.0,1,-nbitq), 
to_sfixed(-153906148.0/4294967296.0,1,-nbitq), 
to_sfixed(-171895509.0/4294967296.0,1,-nbitq), 
to_sfixed(363716971.0/4294967296.0,1,-nbitq), 
to_sfixed(-407052460.0/4294967296.0,1,-nbitq), 
to_sfixed(248337871.0/4294967296.0,1,-nbitq), 
to_sfixed(-137832730.0/4294967296.0,1,-nbitq), 
to_sfixed(-297844962.0/4294967296.0,1,-nbitq), 
to_sfixed(-238556078.0/4294967296.0,1,-nbitq), 
to_sfixed(275727528.0/4294967296.0,1,-nbitq), 
to_sfixed(-53730071.0/4294967296.0,1,-nbitq), 
to_sfixed(-400812206.0/4294967296.0,1,-nbitq), 
to_sfixed(-101422566.0/4294967296.0,1,-nbitq), 
to_sfixed(161825327.0/4294967296.0,1,-nbitq), 
to_sfixed(-186953937.0/4294967296.0,1,-nbitq), 
to_sfixed(-454723846.0/4294967296.0,1,-nbitq), 
to_sfixed(366639419.0/4294967296.0,1,-nbitq), 
to_sfixed(159790953.0/4294967296.0,1,-nbitq), 
to_sfixed(191728027.0/4294967296.0,1,-nbitq), 
to_sfixed(363555496.0/4294967296.0,1,-nbitq), 
to_sfixed(172012809.0/4294967296.0,1,-nbitq), 
to_sfixed(78302227.0/4294967296.0,1,-nbitq), 
to_sfixed(-231183448.0/4294967296.0,1,-nbitq), 
to_sfixed(76076054.0/4294967296.0,1,-nbitq), 
to_sfixed(104431319.0/4294967296.0,1,-nbitq), 
to_sfixed(384739722.0/4294967296.0,1,-nbitq), 
to_sfixed(49131388.0/4294967296.0,1,-nbitq), 
to_sfixed(29873181.0/4294967296.0,1,-nbitq), 
to_sfixed(73459824.0/4294967296.0,1,-nbitq), 
to_sfixed(-239378492.0/4294967296.0,1,-nbitq), 
to_sfixed(49652729.0/4294967296.0,1,-nbitq), 
to_sfixed(120822708.0/4294967296.0,1,-nbitq), 
to_sfixed(-369669632.0/4294967296.0,1,-nbitq), 
to_sfixed(218532895.0/4294967296.0,1,-nbitq), 
to_sfixed(349576933.0/4294967296.0,1,-nbitq), 
to_sfixed(368373835.0/4294967296.0,1,-nbitq), 
to_sfixed(42706197.0/4294967296.0,1,-nbitq), 
to_sfixed(-127442504.0/4294967296.0,1,-nbitq), 
to_sfixed(470949744.0/4294967296.0,1,-nbitq), 
to_sfixed(299609666.0/4294967296.0,1,-nbitq), 
to_sfixed(129023380.0/4294967296.0,1,-nbitq), 
to_sfixed(-133074317.0/4294967296.0,1,-nbitq), 
to_sfixed(194578902.0/4294967296.0,1,-nbitq), 
to_sfixed(-144632816.0/4294967296.0,1,-nbitq), 
to_sfixed(-261925797.0/4294967296.0,1,-nbitq), 
to_sfixed(-119471466.0/4294967296.0,1,-nbitq), 
to_sfixed(-220198100.0/4294967296.0,1,-nbitq), 
to_sfixed(332872120.0/4294967296.0,1,-nbitq), 
to_sfixed(93977133.0/4294967296.0,1,-nbitq), 
to_sfixed(-127081686.0/4294967296.0,1,-nbitq), 
to_sfixed(647635732.0/4294967296.0,1,-nbitq), 
to_sfixed(117124395.0/4294967296.0,1,-nbitq), 
to_sfixed(234780519.0/4294967296.0,1,-nbitq), 
to_sfixed(453229863.0/4294967296.0,1,-nbitq), 
to_sfixed(256482544.0/4294967296.0,1,-nbitq), 
to_sfixed(-175629262.0/4294967296.0,1,-nbitq), 
to_sfixed(-324952972.0/4294967296.0,1,-nbitq), 
to_sfixed(-285790509.0/4294967296.0,1,-nbitq), 
to_sfixed(-257328661.0/4294967296.0,1,-nbitq), 
to_sfixed(-127108576.0/4294967296.0,1,-nbitq), 
to_sfixed(-185249997.0/4294967296.0,1,-nbitq), 
to_sfixed(-102389134.0/4294967296.0,1,-nbitq), 
to_sfixed(-274555895.0/4294967296.0,1,-nbitq), 
to_sfixed(12279564.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-153241480.0/4294967296.0,1,-nbitq), 
to_sfixed(-1465804.0/4294967296.0,1,-nbitq), 
to_sfixed(-125056801.0/4294967296.0,1,-nbitq), 
to_sfixed(-196551760.0/4294967296.0,1,-nbitq), 
to_sfixed(-191763203.0/4294967296.0,1,-nbitq), 
to_sfixed(-440873514.0/4294967296.0,1,-nbitq), 
to_sfixed(-259051240.0/4294967296.0,1,-nbitq), 
to_sfixed(-401731555.0/4294967296.0,1,-nbitq), 
to_sfixed(-292240797.0/4294967296.0,1,-nbitq), 
to_sfixed(-188154578.0/4294967296.0,1,-nbitq), 
to_sfixed(222973899.0/4294967296.0,1,-nbitq), 
to_sfixed(-40995155.0/4294967296.0,1,-nbitq), 
to_sfixed(-54116432.0/4294967296.0,1,-nbitq), 
to_sfixed(181506929.0/4294967296.0,1,-nbitq), 
to_sfixed(145317427.0/4294967296.0,1,-nbitq), 
to_sfixed(-401357615.0/4294967296.0,1,-nbitq), 
to_sfixed(-385280173.0/4294967296.0,1,-nbitq), 
to_sfixed(250712540.0/4294967296.0,1,-nbitq), 
to_sfixed(-41436744.0/4294967296.0,1,-nbitq), 
to_sfixed(265619127.0/4294967296.0,1,-nbitq), 
to_sfixed(-245397437.0/4294967296.0,1,-nbitq), 
to_sfixed(-74752458.0/4294967296.0,1,-nbitq), 
to_sfixed(130698886.0/4294967296.0,1,-nbitq), 
to_sfixed(-186174909.0/4294967296.0,1,-nbitq), 
to_sfixed(350992733.0/4294967296.0,1,-nbitq), 
to_sfixed(-45971027.0/4294967296.0,1,-nbitq), 
to_sfixed(-251010831.0/4294967296.0,1,-nbitq), 
to_sfixed(-643169323.0/4294967296.0,1,-nbitq), 
to_sfixed(-9585242.0/4294967296.0,1,-nbitq), 
to_sfixed(-234664349.0/4294967296.0,1,-nbitq), 
to_sfixed(-29642773.0/4294967296.0,1,-nbitq), 
to_sfixed(-198655573.0/4294967296.0,1,-nbitq), 
to_sfixed(79935628.0/4294967296.0,1,-nbitq), 
to_sfixed(54476386.0/4294967296.0,1,-nbitq), 
to_sfixed(562251891.0/4294967296.0,1,-nbitq), 
to_sfixed(286697583.0/4294967296.0,1,-nbitq), 
to_sfixed(38898538.0/4294967296.0,1,-nbitq), 
to_sfixed(375639307.0/4294967296.0,1,-nbitq), 
to_sfixed(-322975066.0/4294967296.0,1,-nbitq), 
to_sfixed(324612469.0/4294967296.0,1,-nbitq), 
to_sfixed(211816022.0/4294967296.0,1,-nbitq), 
to_sfixed(67714064.0/4294967296.0,1,-nbitq), 
to_sfixed(-23201290.0/4294967296.0,1,-nbitq), 
to_sfixed(-12739429.0/4294967296.0,1,-nbitq), 
to_sfixed(367798233.0/4294967296.0,1,-nbitq), 
to_sfixed(-22677061.0/4294967296.0,1,-nbitq), 
to_sfixed(-39279639.0/4294967296.0,1,-nbitq), 
to_sfixed(-472970324.0/4294967296.0,1,-nbitq), 
to_sfixed(-33306880.0/4294967296.0,1,-nbitq), 
to_sfixed(47489156.0/4294967296.0,1,-nbitq), 
to_sfixed(101163999.0/4294967296.0,1,-nbitq), 
to_sfixed(-195955268.0/4294967296.0,1,-nbitq), 
to_sfixed(-152943775.0/4294967296.0,1,-nbitq), 
to_sfixed(242492698.0/4294967296.0,1,-nbitq), 
to_sfixed(449841100.0/4294967296.0,1,-nbitq), 
to_sfixed(-144593885.0/4294967296.0,1,-nbitq), 
to_sfixed(184854033.0/4294967296.0,1,-nbitq), 
to_sfixed(-146992351.0/4294967296.0,1,-nbitq), 
to_sfixed(3910143.0/4294967296.0,1,-nbitq), 
to_sfixed(410931335.0/4294967296.0,1,-nbitq), 
to_sfixed(-82424971.0/4294967296.0,1,-nbitq), 
to_sfixed(299308749.0/4294967296.0,1,-nbitq), 
to_sfixed(-176509328.0/4294967296.0,1,-nbitq), 
to_sfixed(-72236553.0/4294967296.0,1,-nbitq), 
to_sfixed(-216636080.0/4294967296.0,1,-nbitq), 
to_sfixed(-169256651.0/4294967296.0,1,-nbitq), 
to_sfixed(442446335.0/4294967296.0,1,-nbitq), 
to_sfixed(-233055245.0/4294967296.0,1,-nbitq), 
to_sfixed(271831856.0/4294967296.0,1,-nbitq), 
to_sfixed(67300591.0/4294967296.0,1,-nbitq), 
to_sfixed(171527117.0/4294967296.0,1,-nbitq), 
to_sfixed(373648333.0/4294967296.0,1,-nbitq), 
to_sfixed(-295571802.0/4294967296.0,1,-nbitq), 
to_sfixed(214317038.0/4294967296.0,1,-nbitq), 
to_sfixed(-148742030.0/4294967296.0,1,-nbitq), 
to_sfixed(105513667.0/4294967296.0,1,-nbitq), 
to_sfixed(98151175.0/4294967296.0,1,-nbitq), 
to_sfixed(-4085772.0/4294967296.0,1,-nbitq), 
to_sfixed(-443194260.0/4294967296.0,1,-nbitq), 
to_sfixed(-33851161.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(45087273.0/4294967296.0,1,-nbitq), 
to_sfixed(40043042.0/4294967296.0,1,-nbitq), 
to_sfixed(218886910.0/4294967296.0,1,-nbitq), 
to_sfixed(-284291483.0/4294967296.0,1,-nbitq), 
to_sfixed(-143261647.0/4294967296.0,1,-nbitq), 
to_sfixed(-427246961.0/4294967296.0,1,-nbitq), 
to_sfixed(-24878919.0/4294967296.0,1,-nbitq), 
to_sfixed(-150996011.0/4294967296.0,1,-nbitq), 
to_sfixed(145436768.0/4294967296.0,1,-nbitq), 
to_sfixed(48643087.0/4294967296.0,1,-nbitq), 
to_sfixed(-111054645.0/4294967296.0,1,-nbitq), 
to_sfixed(-89218302.0/4294967296.0,1,-nbitq), 
to_sfixed(224014846.0/4294967296.0,1,-nbitq), 
to_sfixed(-197707810.0/4294967296.0,1,-nbitq), 
to_sfixed(324617347.0/4294967296.0,1,-nbitq), 
to_sfixed(-303416920.0/4294967296.0,1,-nbitq), 
to_sfixed(83723681.0/4294967296.0,1,-nbitq), 
to_sfixed(2565304.0/4294967296.0,1,-nbitq), 
to_sfixed(333305572.0/4294967296.0,1,-nbitq), 
to_sfixed(-108616322.0/4294967296.0,1,-nbitq), 
to_sfixed(112900214.0/4294967296.0,1,-nbitq), 
to_sfixed(-89451535.0/4294967296.0,1,-nbitq), 
to_sfixed(472573245.0/4294967296.0,1,-nbitq), 
to_sfixed(204958127.0/4294967296.0,1,-nbitq), 
to_sfixed(-117083649.0/4294967296.0,1,-nbitq), 
to_sfixed(85203088.0/4294967296.0,1,-nbitq), 
to_sfixed(357094343.0/4294967296.0,1,-nbitq), 
to_sfixed(81973246.0/4294967296.0,1,-nbitq), 
to_sfixed(376296255.0/4294967296.0,1,-nbitq), 
to_sfixed(-163385786.0/4294967296.0,1,-nbitq), 
to_sfixed(-244659267.0/4294967296.0,1,-nbitq), 
to_sfixed(-149378991.0/4294967296.0,1,-nbitq), 
to_sfixed(146618932.0/4294967296.0,1,-nbitq), 
to_sfixed(-104485036.0/4294967296.0,1,-nbitq), 
to_sfixed(-72122531.0/4294967296.0,1,-nbitq), 
to_sfixed(-115341407.0/4294967296.0,1,-nbitq), 
to_sfixed(-21569678.0/4294967296.0,1,-nbitq), 
to_sfixed(376143785.0/4294967296.0,1,-nbitq), 
to_sfixed(362260369.0/4294967296.0,1,-nbitq), 
to_sfixed(157425715.0/4294967296.0,1,-nbitq), 
to_sfixed(-465230476.0/4294967296.0,1,-nbitq), 
to_sfixed(13675081.0/4294967296.0,1,-nbitq), 
to_sfixed(-57922470.0/4294967296.0,1,-nbitq), 
to_sfixed(-179754987.0/4294967296.0,1,-nbitq), 
to_sfixed(222114473.0/4294967296.0,1,-nbitq), 
to_sfixed(58637998.0/4294967296.0,1,-nbitq), 
to_sfixed(-298671465.0/4294967296.0,1,-nbitq), 
to_sfixed(84215308.0/4294967296.0,1,-nbitq), 
to_sfixed(55234209.0/4294967296.0,1,-nbitq), 
to_sfixed(333833970.0/4294967296.0,1,-nbitq), 
to_sfixed(-133936133.0/4294967296.0,1,-nbitq), 
to_sfixed(-152271487.0/4294967296.0,1,-nbitq), 
to_sfixed(-586726565.0/4294967296.0,1,-nbitq), 
to_sfixed(-123518042.0/4294967296.0,1,-nbitq), 
to_sfixed(-93533007.0/4294967296.0,1,-nbitq), 
to_sfixed(264018938.0/4294967296.0,1,-nbitq), 
to_sfixed(-93506913.0/4294967296.0,1,-nbitq), 
to_sfixed(218184144.0/4294967296.0,1,-nbitq), 
to_sfixed(181901435.0/4294967296.0,1,-nbitq), 
to_sfixed(-133490051.0/4294967296.0,1,-nbitq), 
to_sfixed(-196737759.0/4294967296.0,1,-nbitq), 
to_sfixed(383703571.0/4294967296.0,1,-nbitq), 
to_sfixed(272866145.0/4294967296.0,1,-nbitq), 
to_sfixed(62527336.0/4294967296.0,1,-nbitq), 
to_sfixed(209905245.0/4294967296.0,1,-nbitq), 
to_sfixed(-51366546.0/4294967296.0,1,-nbitq), 
to_sfixed(316621390.0/4294967296.0,1,-nbitq), 
to_sfixed(-429667651.0/4294967296.0,1,-nbitq), 
to_sfixed(73179332.0/4294967296.0,1,-nbitq), 
to_sfixed(22720460.0/4294967296.0,1,-nbitq), 
to_sfixed(-338366609.0/4294967296.0,1,-nbitq), 
to_sfixed(-116009820.0/4294967296.0,1,-nbitq), 
to_sfixed(-244374704.0/4294967296.0,1,-nbitq), 
to_sfixed(27278984.0/4294967296.0,1,-nbitq), 
to_sfixed(397951084.0/4294967296.0,1,-nbitq), 
to_sfixed(-146561605.0/4294967296.0,1,-nbitq), 
to_sfixed(-31188201.0/4294967296.0,1,-nbitq), 
to_sfixed(-332747939.0/4294967296.0,1,-nbitq), 
to_sfixed(108263602.0/4294967296.0,1,-nbitq), 
to_sfixed(-20784994.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-61558876.0/4294967296.0,1,-nbitq), 
to_sfixed(-108237295.0/4294967296.0,1,-nbitq), 
to_sfixed(-130830922.0/4294967296.0,1,-nbitq), 
to_sfixed(-283966076.0/4294967296.0,1,-nbitq), 
to_sfixed(43669268.0/4294967296.0,1,-nbitq), 
to_sfixed(-166624024.0/4294967296.0,1,-nbitq), 
to_sfixed(3091382.0/4294967296.0,1,-nbitq), 
to_sfixed(203919985.0/4294967296.0,1,-nbitq), 
to_sfixed(346862545.0/4294967296.0,1,-nbitq), 
to_sfixed(262309940.0/4294967296.0,1,-nbitq), 
to_sfixed(-62263787.0/4294967296.0,1,-nbitq), 
to_sfixed(91463780.0/4294967296.0,1,-nbitq), 
to_sfixed(-257151861.0/4294967296.0,1,-nbitq), 
to_sfixed(-195219015.0/4294967296.0,1,-nbitq), 
to_sfixed(19233700.0/4294967296.0,1,-nbitq), 
to_sfixed(-54389388.0/4294967296.0,1,-nbitq), 
to_sfixed(-100230399.0/4294967296.0,1,-nbitq), 
to_sfixed(358366341.0/4294967296.0,1,-nbitq), 
to_sfixed(289897656.0/4294967296.0,1,-nbitq), 
to_sfixed(100636089.0/4294967296.0,1,-nbitq), 
to_sfixed(-188790260.0/4294967296.0,1,-nbitq), 
to_sfixed(327353290.0/4294967296.0,1,-nbitq), 
to_sfixed(204062030.0/4294967296.0,1,-nbitq), 
to_sfixed(289654646.0/4294967296.0,1,-nbitq), 
to_sfixed(139017384.0/4294967296.0,1,-nbitq), 
to_sfixed(506639499.0/4294967296.0,1,-nbitq), 
to_sfixed(213255902.0/4294967296.0,1,-nbitq), 
to_sfixed(-437185754.0/4294967296.0,1,-nbitq), 
to_sfixed(-110746295.0/4294967296.0,1,-nbitq), 
to_sfixed(25764349.0/4294967296.0,1,-nbitq), 
to_sfixed(-235684398.0/4294967296.0,1,-nbitq), 
to_sfixed(196992644.0/4294967296.0,1,-nbitq), 
to_sfixed(333712629.0/4294967296.0,1,-nbitq), 
to_sfixed(-166573506.0/4294967296.0,1,-nbitq), 
to_sfixed(299815814.0/4294967296.0,1,-nbitq), 
to_sfixed(143203673.0/4294967296.0,1,-nbitq), 
to_sfixed(-315309292.0/4294967296.0,1,-nbitq), 
to_sfixed(33542647.0/4294967296.0,1,-nbitq), 
to_sfixed(-293604814.0/4294967296.0,1,-nbitq), 
to_sfixed(395696560.0/4294967296.0,1,-nbitq), 
to_sfixed(-228059796.0/4294967296.0,1,-nbitq), 
to_sfixed(260467054.0/4294967296.0,1,-nbitq), 
to_sfixed(-339675746.0/4294967296.0,1,-nbitq), 
to_sfixed(327774506.0/4294967296.0,1,-nbitq), 
to_sfixed(-352615414.0/4294967296.0,1,-nbitq), 
to_sfixed(283278648.0/4294967296.0,1,-nbitq), 
to_sfixed(190794127.0/4294967296.0,1,-nbitq), 
to_sfixed(-451925862.0/4294967296.0,1,-nbitq), 
to_sfixed(-111411656.0/4294967296.0,1,-nbitq), 
to_sfixed(402850600.0/4294967296.0,1,-nbitq), 
to_sfixed(99188261.0/4294967296.0,1,-nbitq), 
to_sfixed(-110684973.0/4294967296.0,1,-nbitq), 
to_sfixed(-177838253.0/4294967296.0,1,-nbitq), 
to_sfixed(183051918.0/4294967296.0,1,-nbitq), 
to_sfixed(-147908879.0/4294967296.0,1,-nbitq), 
to_sfixed(244468270.0/4294967296.0,1,-nbitq), 
to_sfixed(-34540908.0/4294967296.0,1,-nbitq), 
to_sfixed(-36128597.0/4294967296.0,1,-nbitq), 
to_sfixed(91164873.0/4294967296.0,1,-nbitq), 
to_sfixed(-126239392.0/4294967296.0,1,-nbitq), 
to_sfixed(-289118686.0/4294967296.0,1,-nbitq), 
to_sfixed(-127060297.0/4294967296.0,1,-nbitq), 
to_sfixed(-339175469.0/4294967296.0,1,-nbitq), 
to_sfixed(363208128.0/4294967296.0,1,-nbitq), 
to_sfixed(405943516.0/4294967296.0,1,-nbitq), 
to_sfixed(168332529.0/4294967296.0,1,-nbitq), 
to_sfixed(634657445.0/4294967296.0,1,-nbitq), 
to_sfixed(226128044.0/4294967296.0,1,-nbitq), 
to_sfixed(132470766.0/4294967296.0,1,-nbitq), 
to_sfixed(-256336212.0/4294967296.0,1,-nbitq), 
to_sfixed(-79955153.0/4294967296.0,1,-nbitq), 
to_sfixed(-6282641.0/4294967296.0,1,-nbitq), 
to_sfixed(-299848224.0/4294967296.0,1,-nbitq), 
to_sfixed(425275202.0/4294967296.0,1,-nbitq), 
to_sfixed(113510872.0/4294967296.0,1,-nbitq), 
to_sfixed(170556439.0/4294967296.0,1,-nbitq), 
to_sfixed(236069408.0/4294967296.0,1,-nbitq), 
to_sfixed(-275399460.0/4294967296.0,1,-nbitq), 
to_sfixed(-268414391.0/4294967296.0,1,-nbitq), 
to_sfixed(-234210154.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(310372397.0/4294967296.0,1,-nbitq), 
to_sfixed(-645102565.0/4294967296.0,1,-nbitq), 
to_sfixed(-327400917.0/4294967296.0,1,-nbitq), 
to_sfixed(571058136.0/4294967296.0,1,-nbitq), 
to_sfixed(386514941.0/4294967296.0,1,-nbitq), 
to_sfixed(307613004.0/4294967296.0,1,-nbitq), 
to_sfixed(-194427466.0/4294967296.0,1,-nbitq), 
to_sfixed(-319847559.0/4294967296.0,1,-nbitq), 
to_sfixed(226397630.0/4294967296.0,1,-nbitq), 
to_sfixed(-352859377.0/4294967296.0,1,-nbitq), 
to_sfixed(-325032825.0/4294967296.0,1,-nbitq), 
to_sfixed(146950848.0/4294967296.0,1,-nbitq), 
to_sfixed(-244377990.0/4294967296.0,1,-nbitq), 
to_sfixed(213303672.0/4294967296.0,1,-nbitq), 
to_sfixed(-268132575.0/4294967296.0,1,-nbitq), 
to_sfixed(-322828090.0/4294967296.0,1,-nbitq), 
to_sfixed(139056239.0/4294967296.0,1,-nbitq), 
to_sfixed(-358670004.0/4294967296.0,1,-nbitq), 
to_sfixed(-424084616.0/4294967296.0,1,-nbitq), 
to_sfixed(14357164.0/4294967296.0,1,-nbitq), 
to_sfixed(319198716.0/4294967296.0,1,-nbitq), 
to_sfixed(56242033.0/4294967296.0,1,-nbitq), 
to_sfixed(355507438.0/4294967296.0,1,-nbitq), 
to_sfixed(362959675.0/4294967296.0,1,-nbitq), 
to_sfixed(-335657899.0/4294967296.0,1,-nbitq), 
to_sfixed(145586062.0/4294967296.0,1,-nbitq), 
to_sfixed(-109750825.0/4294967296.0,1,-nbitq), 
to_sfixed(-331744373.0/4294967296.0,1,-nbitq), 
to_sfixed(-365437634.0/4294967296.0,1,-nbitq), 
to_sfixed(-294838597.0/4294967296.0,1,-nbitq), 
to_sfixed(-514795273.0/4294967296.0,1,-nbitq), 
to_sfixed(-558117872.0/4294967296.0,1,-nbitq), 
to_sfixed(13078833.0/4294967296.0,1,-nbitq), 
to_sfixed(-135847545.0/4294967296.0,1,-nbitq), 
to_sfixed(-39130956.0/4294967296.0,1,-nbitq), 
to_sfixed(153024936.0/4294967296.0,1,-nbitq), 
to_sfixed(254892066.0/4294967296.0,1,-nbitq), 
to_sfixed(133575230.0/4294967296.0,1,-nbitq), 
to_sfixed(-329578731.0/4294967296.0,1,-nbitq), 
to_sfixed(479593535.0/4294967296.0,1,-nbitq), 
to_sfixed(-476434363.0/4294967296.0,1,-nbitq), 
to_sfixed(-135232200.0/4294967296.0,1,-nbitq), 
to_sfixed(56154118.0/4294967296.0,1,-nbitq), 
to_sfixed(408504704.0/4294967296.0,1,-nbitq), 
to_sfixed(-189774764.0/4294967296.0,1,-nbitq), 
to_sfixed(-336388495.0/4294967296.0,1,-nbitq), 
to_sfixed(-40059678.0/4294967296.0,1,-nbitq), 
to_sfixed(63647969.0/4294967296.0,1,-nbitq), 
to_sfixed(11241503.0/4294967296.0,1,-nbitq), 
to_sfixed(-57415552.0/4294967296.0,1,-nbitq), 
to_sfixed(-212039906.0/4294967296.0,1,-nbitq), 
to_sfixed(-57544824.0/4294967296.0,1,-nbitq), 
to_sfixed(-759209651.0/4294967296.0,1,-nbitq), 
to_sfixed(42932629.0/4294967296.0,1,-nbitq), 
to_sfixed(102511610.0/4294967296.0,1,-nbitq), 
to_sfixed(163945479.0/4294967296.0,1,-nbitq), 
to_sfixed(228609313.0/4294967296.0,1,-nbitq), 
to_sfixed(-243652727.0/4294967296.0,1,-nbitq), 
to_sfixed(185014916.0/4294967296.0,1,-nbitq), 
to_sfixed(-124434602.0/4294967296.0,1,-nbitq), 
to_sfixed(22049167.0/4294967296.0,1,-nbitq), 
to_sfixed(194537400.0/4294967296.0,1,-nbitq), 
to_sfixed(27232650.0/4294967296.0,1,-nbitq), 
to_sfixed(342371374.0/4294967296.0,1,-nbitq), 
to_sfixed(-293663165.0/4294967296.0,1,-nbitq), 
to_sfixed(222340230.0/4294967296.0,1,-nbitq), 
to_sfixed(526972533.0/4294967296.0,1,-nbitq), 
to_sfixed(-139829484.0/4294967296.0,1,-nbitq), 
to_sfixed(313128847.0/4294967296.0,1,-nbitq), 
to_sfixed(-39554080.0/4294967296.0,1,-nbitq), 
to_sfixed(-135989638.0/4294967296.0,1,-nbitq), 
to_sfixed(302245549.0/4294967296.0,1,-nbitq), 
to_sfixed(222661728.0/4294967296.0,1,-nbitq), 
to_sfixed(215004243.0/4294967296.0,1,-nbitq), 
to_sfixed(53880567.0/4294967296.0,1,-nbitq), 
to_sfixed(-337463914.0/4294967296.0,1,-nbitq), 
to_sfixed(169068741.0/4294967296.0,1,-nbitq), 
to_sfixed(225630911.0/4294967296.0,1,-nbitq), 
to_sfixed(-562946136.0/4294967296.0,1,-nbitq), 
to_sfixed(-217764400.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-387089605.0/4294967296.0,1,-nbitq), 
to_sfixed(-703125950.0/4294967296.0,1,-nbitq), 
to_sfixed(-574114210.0/4294967296.0,1,-nbitq), 
to_sfixed(-297230045.0/4294967296.0,1,-nbitq), 
to_sfixed(399817878.0/4294967296.0,1,-nbitq), 
to_sfixed(101021901.0/4294967296.0,1,-nbitq), 
to_sfixed(85721233.0/4294967296.0,1,-nbitq), 
to_sfixed(276376256.0/4294967296.0,1,-nbitq), 
to_sfixed(316671614.0/4294967296.0,1,-nbitq), 
to_sfixed(55825225.0/4294967296.0,1,-nbitq), 
to_sfixed(273012221.0/4294967296.0,1,-nbitq), 
to_sfixed(700321546.0/4294967296.0,1,-nbitq), 
to_sfixed(-553098761.0/4294967296.0,1,-nbitq), 
to_sfixed(34568830.0/4294967296.0,1,-nbitq), 
to_sfixed(-212005910.0/4294967296.0,1,-nbitq), 
to_sfixed(82493268.0/4294967296.0,1,-nbitq), 
to_sfixed(212581954.0/4294967296.0,1,-nbitq), 
to_sfixed(-325786800.0/4294967296.0,1,-nbitq), 
to_sfixed(-395147844.0/4294967296.0,1,-nbitq), 
to_sfixed(55523177.0/4294967296.0,1,-nbitq), 
to_sfixed(-103538198.0/4294967296.0,1,-nbitq), 
to_sfixed(-85917231.0/4294967296.0,1,-nbitq), 
to_sfixed(213602120.0/4294967296.0,1,-nbitq), 
to_sfixed(-258220256.0/4294967296.0,1,-nbitq), 
to_sfixed(316654947.0/4294967296.0,1,-nbitq), 
to_sfixed(-188275690.0/4294967296.0,1,-nbitq), 
to_sfixed(-250575194.0/4294967296.0,1,-nbitq), 
to_sfixed(-75907779.0/4294967296.0,1,-nbitq), 
to_sfixed(-295226694.0/4294967296.0,1,-nbitq), 
to_sfixed(-465273275.0/4294967296.0,1,-nbitq), 
to_sfixed(61408159.0/4294967296.0,1,-nbitq), 
to_sfixed(35995112.0/4294967296.0,1,-nbitq), 
to_sfixed(282659976.0/4294967296.0,1,-nbitq), 
to_sfixed(-435610757.0/4294967296.0,1,-nbitq), 
to_sfixed(359505086.0/4294967296.0,1,-nbitq), 
to_sfixed(365527845.0/4294967296.0,1,-nbitq), 
to_sfixed(542348920.0/4294967296.0,1,-nbitq), 
to_sfixed(395246392.0/4294967296.0,1,-nbitq), 
to_sfixed(138737260.0/4294967296.0,1,-nbitq), 
to_sfixed(296401091.0/4294967296.0,1,-nbitq), 
to_sfixed(-496499757.0/4294967296.0,1,-nbitq), 
to_sfixed(-73521707.0/4294967296.0,1,-nbitq), 
to_sfixed(159606805.0/4294967296.0,1,-nbitq), 
to_sfixed(116216135.0/4294967296.0,1,-nbitq), 
to_sfixed(-204681842.0/4294967296.0,1,-nbitq), 
to_sfixed(-42177487.0/4294967296.0,1,-nbitq), 
to_sfixed(30639170.0/4294967296.0,1,-nbitq), 
to_sfixed(241518380.0/4294967296.0,1,-nbitq), 
to_sfixed(-229416508.0/4294967296.0,1,-nbitq), 
to_sfixed(321673253.0/4294967296.0,1,-nbitq), 
to_sfixed(-279748426.0/4294967296.0,1,-nbitq), 
to_sfixed(440260301.0/4294967296.0,1,-nbitq), 
to_sfixed(40592090.0/4294967296.0,1,-nbitq), 
to_sfixed(284557236.0/4294967296.0,1,-nbitq), 
to_sfixed(186134416.0/4294967296.0,1,-nbitq), 
to_sfixed(245572139.0/4294967296.0,1,-nbitq), 
to_sfixed(-236594566.0/4294967296.0,1,-nbitq), 
to_sfixed(-173692536.0/4294967296.0,1,-nbitq), 
to_sfixed(-146322235.0/4294967296.0,1,-nbitq), 
to_sfixed(-44511968.0/4294967296.0,1,-nbitq), 
to_sfixed(-11842906.0/4294967296.0,1,-nbitq), 
to_sfixed(-279172598.0/4294967296.0,1,-nbitq), 
to_sfixed(-204826906.0/4294967296.0,1,-nbitq), 
to_sfixed(-342809002.0/4294967296.0,1,-nbitq), 
to_sfixed(-86464133.0/4294967296.0,1,-nbitq), 
to_sfixed(-86974039.0/4294967296.0,1,-nbitq), 
to_sfixed(-168518469.0/4294967296.0,1,-nbitq), 
to_sfixed(-35706708.0/4294967296.0,1,-nbitq), 
to_sfixed(272788978.0/4294967296.0,1,-nbitq), 
to_sfixed(-257969915.0/4294967296.0,1,-nbitq), 
to_sfixed(223476995.0/4294967296.0,1,-nbitq), 
to_sfixed(42989767.0/4294967296.0,1,-nbitq), 
to_sfixed(-380576911.0/4294967296.0,1,-nbitq), 
to_sfixed(384875563.0/4294967296.0,1,-nbitq), 
to_sfixed(407664359.0/4294967296.0,1,-nbitq), 
to_sfixed(164145723.0/4294967296.0,1,-nbitq), 
to_sfixed(331946512.0/4294967296.0,1,-nbitq), 
to_sfixed(-165699428.0/4294967296.0,1,-nbitq), 
to_sfixed(-558571819.0/4294967296.0,1,-nbitq), 
to_sfixed(165831386.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-163163246.0/4294967296.0,1,-nbitq), 
to_sfixed(-370852330.0/4294967296.0,1,-nbitq), 
to_sfixed(-48178838.0/4294967296.0,1,-nbitq), 
to_sfixed(-442058154.0/4294967296.0,1,-nbitq), 
to_sfixed(232035197.0/4294967296.0,1,-nbitq), 
to_sfixed(530837958.0/4294967296.0,1,-nbitq), 
to_sfixed(248574527.0/4294967296.0,1,-nbitq), 
to_sfixed(-124064474.0/4294967296.0,1,-nbitq), 
to_sfixed(97546141.0/4294967296.0,1,-nbitq), 
to_sfixed(-298249047.0/4294967296.0,1,-nbitq), 
to_sfixed(305203169.0/4294967296.0,1,-nbitq), 
to_sfixed(265179353.0/4294967296.0,1,-nbitq), 
to_sfixed(-564717657.0/4294967296.0,1,-nbitq), 
to_sfixed(-381193723.0/4294967296.0,1,-nbitq), 
to_sfixed(385372717.0/4294967296.0,1,-nbitq), 
to_sfixed(378543859.0/4294967296.0,1,-nbitq), 
to_sfixed(-266443573.0/4294967296.0,1,-nbitq), 
to_sfixed(320354165.0/4294967296.0,1,-nbitq), 
to_sfixed(-365625873.0/4294967296.0,1,-nbitq), 
to_sfixed(41295642.0/4294967296.0,1,-nbitq), 
to_sfixed(15755400.0/4294967296.0,1,-nbitq), 
to_sfixed(-89875748.0/4294967296.0,1,-nbitq), 
to_sfixed(362045417.0/4294967296.0,1,-nbitq), 
to_sfixed(96601269.0/4294967296.0,1,-nbitq), 
to_sfixed(272247620.0/4294967296.0,1,-nbitq), 
to_sfixed(-302263650.0/4294967296.0,1,-nbitq), 
to_sfixed(47594955.0/4294967296.0,1,-nbitq), 
to_sfixed(-92587682.0/4294967296.0,1,-nbitq), 
to_sfixed(-111706219.0/4294967296.0,1,-nbitq), 
to_sfixed(-743277872.0/4294967296.0,1,-nbitq), 
to_sfixed(241299982.0/4294967296.0,1,-nbitq), 
to_sfixed(-307505203.0/4294967296.0,1,-nbitq), 
to_sfixed(125504006.0/4294967296.0,1,-nbitq), 
to_sfixed(-145059448.0/4294967296.0,1,-nbitq), 
to_sfixed(67781745.0/4294967296.0,1,-nbitq), 
to_sfixed(30320078.0/4294967296.0,1,-nbitq), 
to_sfixed(-131606175.0/4294967296.0,1,-nbitq), 
to_sfixed(35360634.0/4294967296.0,1,-nbitq), 
to_sfixed(-163809081.0/4294967296.0,1,-nbitq), 
to_sfixed(62252643.0/4294967296.0,1,-nbitq), 
to_sfixed(-261324893.0/4294967296.0,1,-nbitq), 
to_sfixed(-508838839.0/4294967296.0,1,-nbitq), 
to_sfixed(966076.0/4294967296.0,1,-nbitq), 
to_sfixed(-143791693.0/4294967296.0,1,-nbitq), 
to_sfixed(359612700.0/4294967296.0,1,-nbitq), 
to_sfixed(418033738.0/4294967296.0,1,-nbitq), 
to_sfixed(-414104176.0/4294967296.0,1,-nbitq), 
to_sfixed(-49804479.0/4294967296.0,1,-nbitq), 
to_sfixed(230732538.0/4294967296.0,1,-nbitq), 
to_sfixed(-239818603.0/4294967296.0,1,-nbitq), 
to_sfixed(-49451729.0/4294967296.0,1,-nbitq), 
to_sfixed(611464069.0/4294967296.0,1,-nbitq), 
to_sfixed(264614039.0/4294967296.0,1,-nbitq), 
to_sfixed(484406399.0/4294967296.0,1,-nbitq), 
to_sfixed(-201396584.0/4294967296.0,1,-nbitq), 
to_sfixed(78520692.0/4294967296.0,1,-nbitq), 
to_sfixed(278652446.0/4294967296.0,1,-nbitq), 
to_sfixed(-683011364.0/4294967296.0,1,-nbitq), 
to_sfixed(-108432955.0/4294967296.0,1,-nbitq), 
to_sfixed(-131361953.0/4294967296.0,1,-nbitq), 
to_sfixed(-487158006.0/4294967296.0,1,-nbitq), 
to_sfixed(162644974.0/4294967296.0,1,-nbitq), 
to_sfixed(273248620.0/4294967296.0,1,-nbitq), 
to_sfixed(-52187413.0/4294967296.0,1,-nbitq), 
to_sfixed(383354477.0/4294967296.0,1,-nbitq), 
to_sfixed(-281530243.0/4294967296.0,1,-nbitq), 
to_sfixed(-388597531.0/4294967296.0,1,-nbitq), 
to_sfixed(-618582765.0/4294967296.0,1,-nbitq), 
to_sfixed(380362214.0/4294967296.0,1,-nbitq), 
to_sfixed(-371452715.0/4294967296.0,1,-nbitq), 
to_sfixed(112613471.0/4294967296.0,1,-nbitq), 
to_sfixed(-318355926.0/4294967296.0,1,-nbitq), 
to_sfixed(-284304720.0/4294967296.0,1,-nbitq), 
to_sfixed(331513422.0/4294967296.0,1,-nbitq), 
to_sfixed(-217050614.0/4294967296.0,1,-nbitq), 
to_sfixed(392425390.0/4294967296.0,1,-nbitq), 
to_sfixed(550099417.0/4294967296.0,1,-nbitq), 
to_sfixed(133207566.0/4294967296.0,1,-nbitq), 
to_sfixed(-536700196.0/4294967296.0,1,-nbitq), 
to_sfixed(-270265415.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(300714277.0/4294967296.0,1,-nbitq), 
to_sfixed(-381425790.0/4294967296.0,1,-nbitq), 
to_sfixed(94818558.0/4294967296.0,1,-nbitq), 
to_sfixed(100003131.0/4294967296.0,1,-nbitq), 
to_sfixed(167582786.0/4294967296.0,1,-nbitq), 
to_sfixed(273183933.0/4294967296.0,1,-nbitq), 
to_sfixed(358218075.0/4294967296.0,1,-nbitq), 
to_sfixed(623011090.0/4294967296.0,1,-nbitq), 
to_sfixed(131029141.0/4294967296.0,1,-nbitq), 
to_sfixed(213846485.0/4294967296.0,1,-nbitq), 
to_sfixed(-8077976.0/4294967296.0,1,-nbitq), 
to_sfixed(390167461.0/4294967296.0,1,-nbitq), 
to_sfixed(-459928163.0/4294967296.0,1,-nbitq), 
to_sfixed(-645449039.0/4294967296.0,1,-nbitq), 
to_sfixed(-220361530.0/4294967296.0,1,-nbitq), 
to_sfixed(339532442.0/4294967296.0,1,-nbitq), 
to_sfixed(125886168.0/4294967296.0,1,-nbitq), 
to_sfixed(84553951.0/4294967296.0,1,-nbitq), 
to_sfixed(-113988601.0/4294967296.0,1,-nbitq), 
to_sfixed(487835914.0/4294967296.0,1,-nbitq), 
to_sfixed(193968727.0/4294967296.0,1,-nbitq), 
to_sfixed(-122628334.0/4294967296.0,1,-nbitq), 
to_sfixed(44514820.0/4294967296.0,1,-nbitq), 
to_sfixed(-377399579.0/4294967296.0,1,-nbitq), 
to_sfixed(-224125499.0/4294967296.0,1,-nbitq), 
to_sfixed(-537815461.0/4294967296.0,1,-nbitq), 
to_sfixed(397416677.0/4294967296.0,1,-nbitq), 
to_sfixed(129565021.0/4294967296.0,1,-nbitq), 
to_sfixed(-150726143.0/4294967296.0,1,-nbitq), 
to_sfixed(-491147408.0/4294967296.0,1,-nbitq), 
to_sfixed(213330472.0/4294967296.0,1,-nbitq), 
to_sfixed(-465199510.0/4294967296.0,1,-nbitq), 
to_sfixed(-82023680.0/4294967296.0,1,-nbitq), 
to_sfixed(298206117.0/4294967296.0,1,-nbitq), 
to_sfixed(54346517.0/4294967296.0,1,-nbitq), 
to_sfixed(-806200611.0/4294967296.0,1,-nbitq), 
to_sfixed(369641908.0/4294967296.0,1,-nbitq), 
to_sfixed(80548241.0/4294967296.0,1,-nbitq), 
to_sfixed(304846055.0/4294967296.0,1,-nbitq), 
to_sfixed(70084394.0/4294967296.0,1,-nbitq), 
to_sfixed(694708142.0/4294967296.0,1,-nbitq), 
to_sfixed(-687150931.0/4294967296.0,1,-nbitq), 
to_sfixed(511829918.0/4294967296.0,1,-nbitq), 
to_sfixed(-314583672.0/4294967296.0,1,-nbitq), 
to_sfixed(139501494.0/4294967296.0,1,-nbitq), 
to_sfixed(-17049907.0/4294967296.0,1,-nbitq), 
to_sfixed(95343020.0/4294967296.0,1,-nbitq), 
to_sfixed(-38187505.0/4294967296.0,1,-nbitq), 
to_sfixed(173589765.0/4294967296.0,1,-nbitq), 
to_sfixed(-132415390.0/4294967296.0,1,-nbitq), 
to_sfixed(-319723919.0/4294967296.0,1,-nbitq), 
to_sfixed(904362219.0/4294967296.0,1,-nbitq), 
to_sfixed(-265226626.0/4294967296.0,1,-nbitq), 
to_sfixed(228956334.0/4294967296.0,1,-nbitq), 
to_sfixed(-791146042.0/4294967296.0,1,-nbitq), 
to_sfixed(1026014046.0/4294967296.0,1,-nbitq), 
to_sfixed(119666310.0/4294967296.0,1,-nbitq), 
to_sfixed(84007634.0/4294967296.0,1,-nbitq), 
to_sfixed(-90490434.0/4294967296.0,1,-nbitq), 
to_sfixed(256090898.0/4294967296.0,1,-nbitq), 
to_sfixed(20089551.0/4294967296.0,1,-nbitq), 
to_sfixed(-107041439.0/4294967296.0,1,-nbitq), 
to_sfixed(-279128586.0/4294967296.0,1,-nbitq), 
to_sfixed(-279378964.0/4294967296.0,1,-nbitq), 
to_sfixed(-271353664.0/4294967296.0,1,-nbitq), 
to_sfixed(240169149.0/4294967296.0,1,-nbitq), 
to_sfixed(-762800980.0/4294967296.0,1,-nbitq), 
to_sfixed(-560524888.0/4294967296.0,1,-nbitq), 
to_sfixed(212158795.0/4294967296.0,1,-nbitq), 
to_sfixed(461761897.0/4294967296.0,1,-nbitq), 
to_sfixed(-293510933.0/4294967296.0,1,-nbitq), 
to_sfixed(-220215508.0/4294967296.0,1,-nbitq), 
to_sfixed(225315069.0/4294967296.0,1,-nbitq), 
to_sfixed(-75491675.0/4294967296.0,1,-nbitq), 
to_sfixed(408074830.0/4294967296.0,1,-nbitq), 
to_sfixed(477358878.0/4294967296.0,1,-nbitq), 
to_sfixed(-265901771.0/4294967296.0,1,-nbitq), 
to_sfixed(-499819116.0/4294967296.0,1,-nbitq), 
to_sfixed(-911177316.0/4294967296.0,1,-nbitq), 
to_sfixed(177753795.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(235170443.0/4294967296.0,1,-nbitq), 
to_sfixed(-399796514.0/4294967296.0,1,-nbitq), 
to_sfixed(-786914335.0/4294967296.0,1,-nbitq), 
to_sfixed(941879545.0/4294967296.0,1,-nbitq), 
to_sfixed(366677720.0/4294967296.0,1,-nbitq), 
to_sfixed(-46677534.0/4294967296.0,1,-nbitq), 
to_sfixed(42599536.0/4294967296.0,1,-nbitq), 
to_sfixed(97125014.0/4294967296.0,1,-nbitq), 
to_sfixed(991570976.0/4294967296.0,1,-nbitq), 
to_sfixed(-255503416.0/4294967296.0,1,-nbitq), 
to_sfixed(-457423273.0/4294967296.0,1,-nbitq), 
to_sfixed(207707033.0/4294967296.0,1,-nbitq), 
to_sfixed(-35571568.0/4294967296.0,1,-nbitq), 
to_sfixed(-1164280171.0/4294967296.0,1,-nbitq), 
to_sfixed(312775340.0/4294967296.0,1,-nbitq), 
to_sfixed(567928668.0/4294967296.0,1,-nbitq), 
to_sfixed(-272837105.0/4294967296.0,1,-nbitq), 
to_sfixed(-104835012.0/4294967296.0,1,-nbitq), 
to_sfixed(284353666.0/4294967296.0,1,-nbitq), 
to_sfixed(223540265.0/4294967296.0,1,-nbitq), 
to_sfixed(-331270182.0/4294967296.0,1,-nbitq), 
to_sfixed(544312637.0/4294967296.0,1,-nbitq), 
to_sfixed(17508119.0/4294967296.0,1,-nbitq), 
to_sfixed(-286394651.0/4294967296.0,1,-nbitq), 
to_sfixed(-305331347.0/4294967296.0,1,-nbitq), 
to_sfixed(-376856945.0/4294967296.0,1,-nbitq), 
to_sfixed(-103712495.0/4294967296.0,1,-nbitq), 
to_sfixed(39511843.0/4294967296.0,1,-nbitq), 
to_sfixed(567148591.0/4294967296.0,1,-nbitq), 
to_sfixed(-963556819.0/4294967296.0,1,-nbitq), 
to_sfixed(612296919.0/4294967296.0,1,-nbitq), 
to_sfixed(-404228135.0/4294967296.0,1,-nbitq), 
to_sfixed(336669825.0/4294967296.0,1,-nbitq), 
to_sfixed(-70491643.0/4294967296.0,1,-nbitq), 
to_sfixed(-651875330.0/4294967296.0,1,-nbitq), 
to_sfixed(-383627328.0/4294967296.0,1,-nbitq), 
to_sfixed(-79939252.0/4294967296.0,1,-nbitq), 
to_sfixed(-504443870.0/4294967296.0,1,-nbitq), 
to_sfixed(-249333755.0/4294967296.0,1,-nbitq), 
to_sfixed(45636357.0/4294967296.0,1,-nbitq), 
to_sfixed(483754476.0/4294967296.0,1,-nbitq), 
to_sfixed(-629883736.0/4294967296.0,1,-nbitq), 
to_sfixed(-113288616.0/4294967296.0,1,-nbitq), 
to_sfixed(311851075.0/4294967296.0,1,-nbitq), 
to_sfixed(367594441.0/4294967296.0,1,-nbitq), 
to_sfixed(296764535.0/4294967296.0,1,-nbitq), 
to_sfixed(-23667971.0/4294967296.0,1,-nbitq), 
to_sfixed(516610437.0/4294967296.0,1,-nbitq), 
to_sfixed(272468590.0/4294967296.0,1,-nbitq), 
to_sfixed(-92638368.0/4294967296.0,1,-nbitq), 
to_sfixed(-699229279.0/4294967296.0,1,-nbitq), 
to_sfixed(767731790.0/4294967296.0,1,-nbitq), 
to_sfixed(259246220.0/4294967296.0,1,-nbitq), 
to_sfixed(-234963727.0/4294967296.0,1,-nbitq), 
to_sfixed(-363062839.0/4294967296.0,1,-nbitq), 
to_sfixed(1145122734.0/4294967296.0,1,-nbitq), 
to_sfixed(-44814210.0/4294967296.0,1,-nbitq), 
to_sfixed(241014304.0/4294967296.0,1,-nbitq), 
to_sfixed(311332312.0/4294967296.0,1,-nbitq), 
to_sfixed(-106096344.0/4294967296.0,1,-nbitq), 
to_sfixed(26709448.0/4294967296.0,1,-nbitq), 
to_sfixed(124931058.0/4294967296.0,1,-nbitq), 
to_sfixed(-579438417.0/4294967296.0,1,-nbitq), 
to_sfixed(152250603.0/4294967296.0,1,-nbitq), 
to_sfixed(-237959811.0/4294967296.0,1,-nbitq), 
to_sfixed(-30170800.0/4294967296.0,1,-nbitq), 
to_sfixed(-665579483.0/4294967296.0,1,-nbitq), 
to_sfixed(-770337246.0/4294967296.0,1,-nbitq), 
to_sfixed(-231822397.0/4294967296.0,1,-nbitq), 
to_sfixed(423755422.0/4294967296.0,1,-nbitq), 
to_sfixed(77643694.0/4294967296.0,1,-nbitq), 
to_sfixed(-315516086.0/4294967296.0,1,-nbitq), 
to_sfixed(300922088.0/4294967296.0,1,-nbitq), 
to_sfixed(235705272.0/4294967296.0,1,-nbitq), 
to_sfixed(-259099114.0/4294967296.0,1,-nbitq), 
to_sfixed(570154335.0/4294967296.0,1,-nbitq), 
to_sfixed(358915300.0/4294967296.0,1,-nbitq), 
to_sfixed(70251250.0/4294967296.0,1,-nbitq), 
to_sfixed(-592280957.0/4294967296.0,1,-nbitq), 
to_sfixed(34852141.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(502023138.0/4294967296.0,1,-nbitq), 
to_sfixed(-68280641.0/4294967296.0,1,-nbitq), 
to_sfixed(-584895356.0/4294967296.0,1,-nbitq), 
to_sfixed(505764619.0/4294967296.0,1,-nbitq), 
to_sfixed(758411300.0/4294967296.0,1,-nbitq), 
to_sfixed(-649836790.0/4294967296.0,1,-nbitq), 
to_sfixed(-262553266.0/4294967296.0,1,-nbitq), 
to_sfixed(481360576.0/4294967296.0,1,-nbitq), 
to_sfixed(519418846.0/4294967296.0,1,-nbitq), 
to_sfixed(121079970.0/4294967296.0,1,-nbitq), 
to_sfixed(140841330.0/4294967296.0,1,-nbitq), 
to_sfixed(401430760.0/4294967296.0,1,-nbitq), 
to_sfixed(-554332899.0/4294967296.0,1,-nbitq), 
to_sfixed(-1006484158.0/4294967296.0,1,-nbitq), 
to_sfixed(337817034.0/4294967296.0,1,-nbitq), 
to_sfixed(99031982.0/4294967296.0,1,-nbitq), 
to_sfixed(3625093.0/4294967296.0,1,-nbitq), 
to_sfixed(-108132507.0/4294967296.0,1,-nbitq), 
to_sfixed(264965.0/4294967296.0,1,-nbitq), 
to_sfixed(318895765.0/4294967296.0,1,-nbitq), 
to_sfixed(-204219315.0/4294967296.0,1,-nbitq), 
to_sfixed(172026542.0/4294967296.0,1,-nbitq), 
to_sfixed(-8661956.0/4294967296.0,1,-nbitq), 
to_sfixed(-27370063.0/4294967296.0,1,-nbitq), 
to_sfixed(-79958028.0/4294967296.0,1,-nbitq), 
to_sfixed(-352768540.0/4294967296.0,1,-nbitq), 
to_sfixed(-741792920.0/4294967296.0,1,-nbitq), 
to_sfixed(481572597.0/4294967296.0,1,-nbitq), 
to_sfixed(221705295.0/4294967296.0,1,-nbitq), 
to_sfixed(-907600554.0/4294967296.0,1,-nbitq), 
to_sfixed(691221993.0/4294967296.0,1,-nbitq), 
to_sfixed(88614130.0/4294967296.0,1,-nbitq), 
to_sfixed(410878182.0/4294967296.0,1,-nbitq), 
to_sfixed(20902269.0/4294967296.0,1,-nbitq), 
to_sfixed(-1140218630.0/4294967296.0,1,-nbitq), 
to_sfixed(-316241082.0/4294967296.0,1,-nbitq), 
to_sfixed(207586090.0/4294967296.0,1,-nbitq), 
to_sfixed(-459344236.0/4294967296.0,1,-nbitq), 
to_sfixed(-182328305.0/4294967296.0,1,-nbitq), 
to_sfixed(-45819823.0/4294967296.0,1,-nbitq), 
to_sfixed(185608576.0/4294967296.0,1,-nbitq), 
to_sfixed(-498747918.0/4294967296.0,1,-nbitq), 
to_sfixed(99715722.0/4294967296.0,1,-nbitq), 
to_sfixed(307029309.0/4294967296.0,1,-nbitq), 
to_sfixed(-14056594.0/4294967296.0,1,-nbitq), 
to_sfixed(497057923.0/4294967296.0,1,-nbitq), 
to_sfixed(-195271182.0/4294967296.0,1,-nbitq), 
to_sfixed(467237457.0/4294967296.0,1,-nbitq), 
to_sfixed(-126510419.0/4294967296.0,1,-nbitq), 
to_sfixed(-894846295.0/4294967296.0,1,-nbitq), 
to_sfixed(-268111455.0/4294967296.0,1,-nbitq), 
to_sfixed(962445688.0/4294967296.0,1,-nbitq), 
to_sfixed(-474675770.0/4294967296.0,1,-nbitq), 
to_sfixed(71607515.0/4294967296.0,1,-nbitq), 
to_sfixed(26234191.0/4294967296.0,1,-nbitq), 
to_sfixed(668829746.0/4294967296.0,1,-nbitq), 
to_sfixed(146561968.0/4294967296.0,1,-nbitq), 
to_sfixed(271958963.0/4294967296.0,1,-nbitq), 
to_sfixed(320552102.0/4294967296.0,1,-nbitq), 
to_sfixed(333458846.0/4294967296.0,1,-nbitq), 
to_sfixed(238157887.0/4294967296.0,1,-nbitq), 
to_sfixed(-298054672.0/4294967296.0,1,-nbitq), 
to_sfixed(-718557549.0/4294967296.0,1,-nbitq), 
to_sfixed(-679431207.0/4294967296.0,1,-nbitq), 
to_sfixed(-187292627.0/4294967296.0,1,-nbitq), 
to_sfixed(-203381981.0/4294967296.0,1,-nbitq), 
to_sfixed(-723258358.0/4294967296.0,1,-nbitq), 
to_sfixed(-684962879.0/4294967296.0,1,-nbitq), 
to_sfixed(71712113.0/4294967296.0,1,-nbitq), 
to_sfixed(287473471.0/4294967296.0,1,-nbitq), 
to_sfixed(413723694.0/4294967296.0,1,-nbitq), 
to_sfixed(-31804958.0/4294967296.0,1,-nbitq), 
to_sfixed(457497327.0/4294967296.0,1,-nbitq), 
to_sfixed(-264314863.0/4294967296.0,1,-nbitq), 
to_sfixed(-224357315.0/4294967296.0,1,-nbitq), 
to_sfixed(-23817510.0/4294967296.0,1,-nbitq), 
to_sfixed(859580505.0/4294967296.0,1,-nbitq), 
to_sfixed(-253624626.0/4294967296.0,1,-nbitq), 
to_sfixed(508253295.0/4294967296.0,1,-nbitq), 
to_sfixed(-150669734.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(526363007.0/4294967296.0,1,-nbitq), 
to_sfixed(-265350981.0/4294967296.0,1,-nbitq), 
to_sfixed(-621658869.0/4294967296.0,1,-nbitq), 
to_sfixed(572190411.0/4294967296.0,1,-nbitq), 
to_sfixed(97136409.0/4294967296.0,1,-nbitq), 
to_sfixed(-717731731.0/4294967296.0,1,-nbitq), 
to_sfixed(22652134.0/4294967296.0,1,-nbitq), 
to_sfixed(742657256.0/4294967296.0,1,-nbitq), 
to_sfixed(1249590206.0/4294967296.0,1,-nbitq), 
to_sfixed(11364579.0/4294967296.0,1,-nbitq), 
to_sfixed(-279828583.0/4294967296.0,1,-nbitq), 
to_sfixed(524071147.0/4294967296.0,1,-nbitq), 
to_sfixed(214172271.0/4294967296.0,1,-nbitq), 
to_sfixed(-1400046182.0/4294967296.0,1,-nbitq), 
to_sfixed(-318536881.0/4294967296.0,1,-nbitq), 
to_sfixed(72338025.0/4294967296.0,1,-nbitq), 
to_sfixed(123773735.0/4294967296.0,1,-nbitq), 
to_sfixed(268384224.0/4294967296.0,1,-nbitq), 
to_sfixed(-51722471.0/4294967296.0,1,-nbitq), 
to_sfixed(-28327909.0/4294967296.0,1,-nbitq), 
to_sfixed(-221179084.0/4294967296.0,1,-nbitq), 
to_sfixed(172279731.0/4294967296.0,1,-nbitq), 
to_sfixed(400014049.0/4294967296.0,1,-nbitq), 
to_sfixed(-861435735.0/4294967296.0,1,-nbitq), 
to_sfixed(-298791795.0/4294967296.0,1,-nbitq), 
to_sfixed(-463403587.0/4294967296.0,1,-nbitq), 
to_sfixed(-125193816.0/4294967296.0,1,-nbitq), 
to_sfixed(320021822.0/4294967296.0,1,-nbitq), 
to_sfixed(123827248.0/4294967296.0,1,-nbitq), 
to_sfixed(-724034338.0/4294967296.0,1,-nbitq), 
to_sfixed(889308327.0/4294967296.0,1,-nbitq), 
to_sfixed(310716424.0/4294967296.0,1,-nbitq), 
to_sfixed(-83157351.0/4294967296.0,1,-nbitq), 
to_sfixed(-421399158.0/4294967296.0,1,-nbitq), 
to_sfixed(-1397993484.0/4294967296.0,1,-nbitq), 
to_sfixed(-903887119.0/4294967296.0,1,-nbitq), 
to_sfixed(168570636.0/4294967296.0,1,-nbitq), 
to_sfixed(-824723078.0/4294967296.0,1,-nbitq), 
to_sfixed(475094388.0/4294967296.0,1,-nbitq), 
to_sfixed(-42298973.0/4294967296.0,1,-nbitq), 
to_sfixed(343275351.0/4294967296.0,1,-nbitq), 
to_sfixed(-458388807.0/4294967296.0,1,-nbitq), 
to_sfixed(137881145.0/4294967296.0,1,-nbitq), 
to_sfixed(318743447.0/4294967296.0,1,-nbitq), 
to_sfixed(-569692490.0/4294967296.0,1,-nbitq), 
to_sfixed(468252884.0/4294967296.0,1,-nbitq), 
to_sfixed(308227184.0/4294967296.0,1,-nbitq), 
to_sfixed(14552869.0/4294967296.0,1,-nbitq), 
to_sfixed(-153324920.0/4294967296.0,1,-nbitq), 
to_sfixed(-1151827104.0/4294967296.0,1,-nbitq), 
to_sfixed(147608651.0/4294967296.0,1,-nbitq), 
to_sfixed(942609344.0/4294967296.0,1,-nbitq), 
to_sfixed(136388126.0/4294967296.0,1,-nbitq), 
to_sfixed(575519928.0/4294967296.0,1,-nbitq), 
to_sfixed(418783710.0/4294967296.0,1,-nbitq), 
to_sfixed(1654731233.0/4294967296.0,1,-nbitq), 
to_sfixed(-38918888.0/4294967296.0,1,-nbitq), 
to_sfixed(140357755.0/4294967296.0,1,-nbitq), 
to_sfixed(249790296.0/4294967296.0,1,-nbitq), 
to_sfixed(-396796424.0/4294967296.0,1,-nbitq), 
to_sfixed(-287812774.0/4294967296.0,1,-nbitq), 
to_sfixed(-579355381.0/4294967296.0,1,-nbitq), 
to_sfixed(-761247831.0/4294967296.0,1,-nbitq), 
to_sfixed(-638931485.0/4294967296.0,1,-nbitq), 
to_sfixed(77458749.0/4294967296.0,1,-nbitq), 
to_sfixed(57194019.0/4294967296.0,1,-nbitq), 
to_sfixed(-246330343.0/4294967296.0,1,-nbitq), 
to_sfixed(24966690.0/4294967296.0,1,-nbitq), 
to_sfixed(-54186798.0/4294967296.0,1,-nbitq), 
to_sfixed(367323872.0/4294967296.0,1,-nbitq), 
to_sfixed(-779318242.0/4294967296.0,1,-nbitq), 
to_sfixed(-322091331.0/4294967296.0,1,-nbitq), 
to_sfixed(873651120.0/4294967296.0,1,-nbitq), 
to_sfixed(-228537265.0/4294967296.0,1,-nbitq), 
to_sfixed(434099042.0/4294967296.0,1,-nbitq), 
to_sfixed(-638664623.0/4294967296.0,1,-nbitq), 
to_sfixed(620321882.0/4294967296.0,1,-nbitq), 
to_sfixed(-920057221.0/4294967296.0,1,-nbitq), 
to_sfixed(308437980.0/4294967296.0,1,-nbitq), 
to_sfixed(-422068339.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(658690668.0/4294967296.0,1,-nbitq), 
to_sfixed(-1323346022.0/4294967296.0,1,-nbitq), 
to_sfixed(-793277344.0/4294967296.0,1,-nbitq), 
to_sfixed(915042304.0/4294967296.0,1,-nbitq), 
to_sfixed(-182172585.0/4294967296.0,1,-nbitq), 
to_sfixed(-14294108.0/4294967296.0,1,-nbitq), 
to_sfixed(159884605.0/4294967296.0,1,-nbitq), 
to_sfixed(298958460.0/4294967296.0,1,-nbitq), 
to_sfixed(211572099.0/4294967296.0,1,-nbitq), 
to_sfixed(-182608053.0/4294967296.0,1,-nbitq), 
to_sfixed(152386033.0/4294967296.0,1,-nbitq), 
to_sfixed(741480803.0/4294967296.0,1,-nbitq), 
to_sfixed(-204657055.0/4294967296.0,1,-nbitq), 
to_sfixed(-386801517.0/4294967296.0,1,-nbitq), 
to_sfixed(373105913.0/4294967296.0,1,-nbitq), 
to_sfixed(131788145.0/4294967296.0,1,-nbitq), 
to_sfixed(-234823408.0/4294967296.0,1,-nbitq), 
to_sfixed(165478715.0/4294967296.0,1,-nbitq), 
to_sfixed(-455936894.0/4294967296.0,1,-nbitq), 
to_sfixed(-338190692.0/4294967296.0,1,-nbitq), 
to_sfixed(-297699795.0/4294967296.0,1,-nbitq), 
to_sfixed(-200149308.0/4294967296.0,1,-nbitq), 
to_sfixed(568456261.0/4294967296.0,1,-nbitq), 
to_sfixed(-475579926.0/4294967296.0,1,-nbitq), 
to_sfixed(219223654.0/4294967296.0,1,-nbitq), 
to_sfixed(-1189744308.0/4294967296.0,1,-nbitq), 
to_sfixed(6832129.0/4294967296.0,1,-nbitq), 
to_sfixed(-226956555.0/4294967296.0,1,-nbitq), 
to_sfixed(119211633.0/4294967296.0,1,-nbitq), 
to_sfixed(-247474104.0/4294967296.0,1,-nbitq), 
to_sfixed(738484637.0/4294967296.0,1,-nbitq), 
to_sfixed(620643355.0/4294967296.0,1,-nbitq), 
to_sfixed(62436162.0/4294967296.0,1,-nbitq), 
to_sfixed(-838345444.0/4294967296.0,1,-nbitq), 
to_sfixed(-758267959.0/4294967296.0,1,-nbitq), 
to_sfixed(-1582099310.0/4294967296.0,1,-nbitq), 
to_sfixed(127724805.0/4294967296.0,1,-nbitq), 
to_sfixed(-1155025717.0/4294967296.0,1,-nbitq), 
to_sfixed(-35761542.0/4294967296.0,1,-nbitq), 
to_sfixed(150753618.0/4294967296.0,1,-nbitq), 
to_sfixed(288885299.0/4294967296.0,1,-nbitq), 
to_sfixed(-851092696.0/4294967296.0,1,-nbitq), 
to_sfixed(843846799.0/4294967296.0,1,-nbitq), 
to_sfixed(152444649.0/4294967296.0,1,-nbitq), 
to_sfixed(-159918824.0/4294967296.0,1,-nbitq), 
to_sfixed(74067164.0/4294967296.0,1,-nbitq), 
to_sfixed(-342919515.0/4294967296.0,1,-nbitq), 
to_sfixed(-9439474.0/4294967296.0,1,-nbitq), 
to_sfixed(-340161998.0/4294967296.0,1,-nbitq), 
to_sfixed(-788001329.0/4294967296.0,1,-nbitq), 
to_sfixed(138760267.0/4294967296.0,1,-nbitq), 
to_sfixed(1431918921.0/4294967296.0,1,-nbitq), 
to_sfixed(-175455202.0/4294967296.0,1,-nbitq), 
to_sfixed(330057272.0/4294967296.0,1,-nbitq), 
to_sfixed(-1015884240.0/4294967296.0,1,-nbitq), 
to_sfixed(731838684.0/4294967296.0,1,-nbitq), 
to_sfixed(-44844597.0/4294967296.0,1,-nbitq), 
to_sfixed(-550999050.0/4294967296.0,1,-nbitq), 
to_sfixed(49285338.0/4294967296.0,1,-nbitq), 
to_sfixed(349317383.0/4294967296.0,1,-nbitq), 
to_sfixed(-158758875.0/4294967296.0,1,-nbitq), 
to_sfixed(-1835733.0/4294967296.0,1,-nbitq), 
to_sfixed(-1006971778.0/4294967296.0,1,-nbitq), 
to_sfixed(-325228816.0/4294967296.0,1,-nbitq), 
to_sfixed(21002826.0/4294967296.0,1,-nbitq), 
to_sfixed(-99450409.0/4294967296.0,1,-nbitq), 
to_sfixed(416486567.0/4294967296.0,1,-nbitq), 
to_sfixed(-183669821.0/4294967296.0,1,-nbitq), 
to_sfixed(-333904161.0/4294967296.0,1,-nbitq), 
to_sfixed(303702204.0/4294967296.0,1,-nbitq), 
to_sfixed(-1156912681.0/4294967296.0,1,-nbitq), 
to_sfixed(222712358.0/4294967296.0,1,-nbitq), 
to_sfixed(1168419741.0/4294967296.0,1,-nbitq), 
to_sfixed(-267851577.0/4294967296.0,1,-nbitq), 
to_sfixed(-53611704.0/4294967296.0,1,-nbitq), 
to_sfixed(-628121283.0/4294967296.0,1,-nbitq), 
to_sfixed(-430413140.0/4294967296.0,1,-nbitq), 
to_sfixed(-469066084.0/4294967296.0,1,-nbitq), 
to_sfixed(-80715222.0/4294967296.0,1,-nbitq), 
to_sfixed(207774773.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(727552624.0/4294967296.0,1,-nbitq), 
to_sfixed(-1713131785.0/4294967296.0,1,-nbitq), 
to_sfixed(92293116.0/4294967296.0,1,-nbitq), 
to_sfixed(1340463285.0/4294967296.0,1,-nbitq), 
to_sfixed(-574665043.0/4294967296.0,1,-nbitq), 
to_sfixed(-460726915.0/4294967296.0,1,-nbitq), 
to_sfixed(-215996074.0/4294967296.0,1,-nbitq), 
to_sfixed(-406967988.0/4294967296.0,1,-nbitq), 
to_sfixed(-1933232.0/4294967296.0,1,-nbitq), 
to_sfixed(266733046.0/4294967296.0,1,-nbitq), 
to_sfixed(-228955556.0/4294967296.0,1,-nbitq), 
to_sfixed(596008748.0/4294967296.0,1,-nbitq), 
to_sfixed(-482582531.0/4294967296.0,1,-nbitq), 
to_sfixed(28550305.0/4294967296.0,1,-nbitq), 
to_sfixed(427852656.0/4294967296.0,1,-nbitq), 
to_sfixed(419995589.0/4294967296.0,1,-nbitq), 
to_sfixed(155129928.0/4294967296.0,1,-nbitq), 
to_sfixed(-363135728.0/4294967296.0,1,-nbitq), 
to_sfixed(237576510.0/4294967296.0,1,-nbitq), 
to_sfixed(-738839552.0/4294967296.0,1,-nbitq), 
to_sfixed(-345552193.0/4294967296.0,1,-nbitq), 
to_sfixed(113452270.0/4294967296.0,1,-nbitq), 
to_sfixed(812576702.0/4294967296.0,1,-nbitq), 
to_sfixed(-47362221.0/4294967296.0,1,-nbitq), 
to_sfixed(210762688.0/4294967296.0,1,-nbitq), 
to_sfixed(-863129170.0/4294967296.0,1,-nbitq), 
to_sfixed(-146064240.0/4294967296.0,1,-nbitq), 
to_sfixed(209698987.0/4294967296.0,1,-nbitq), 
to_sfixed(-160998432.0/4294967296.0,1,-nbitq), 
to_sfixed(-401425207.0/4294967296.0,1,-nbitq), 
to_sfixed(735702043.0/4294967296.0,1,-nbitq), 
to_sfixed(-277344227.0/4294967296.0,1,-nbitq), 
to_sfixed(505365519.0/4294967296.0,1,-nbitq), 
to_sfixed(-925819900.0/4294967296.0,1,-nbitq), 
to_sfixed(-112015848.0/4294967296.0,1,-nbitq), 
to_sfixed(-200626275.0/4294967296.0,1,-nbitq), 
to_sfixed(287728819.0/4294967296.0,1,-nbitq), 
to_sfixed(-996321736.0/4294967296.0,1,-nbitq), 
to_sfixed(44093602.0/4294967296.0,1,-nbitq), 
to_sfixed(-73318582.0/4294967296.0,1,-nbitq), 
to_sfixed(-55375102.0/4294967296.0,1,-nbitq), 
to_sfixed(-293270763.0/4294967296.0,1,-nbitq), 
to_sfixed(1474609987.0/4294967296.0,1,-nbitq), 
to_sfixed(872009650.0/4294967296.0,1,-nbitq), 
to_sfixed(332453760.0/4294967296.0,1,-nbitq), 
to_sfixed(-383180852.0/4294967296.0,1,-nbitq), 
to_sfixed(-241919149.0/4294967296.0,1,-nbitq), 
to_sfixed(18440892.0/4294967296.0,1,-nbitq), 
to_sfixed(-464944885.0/4294967296.0,1,-nbitq), 
to_sfixed(-530409397.0/4294967296.0,1,-nbitq), 
to_sfixed(-394447809.0/4294967296.0,1,-nbitq), 
to_sfixed(386596240.0/4294967296.0,1,-nbitq), 
to_sfixed(-390877098.0/4294967296.0,1,-nbitq), 
to_sfixed(-249250654.0/4294967296.0,1,-nbitq), 
to_sfixed(-360558789.0/4294967296.0,1,-nbitq), 
to_sfixed(-35134585.0/4294967296.0,1,-nbitq), 
to_sfixed(-59650023.0/4294967296.0,1,-nbitq), 
to_sfixed(97134374.0/4294967296.0,1,-nbitq), 
to_sfixed(243934022.0/4294967296.0,1,-nbitq), 
to_sfixed(76668196.0/4294967296.0,1,-nbitq), 
to_sfixed(-42385072.0/4294967296.0,1,-nbitq), 
to_sfixed(-134515835.0/4294967296.0,1,-nbitq), 
to_sfixed(-800520095.0/4294967296.0,1,-nbitq), 
to_sfixed(-657220868.0/4294967296.0,1,-nbitq), 
to_sfixed(78534807.0/4294967296.0,1,-nbitq), 
to_sfixed(181013129.0/4294967296.0,1,-nbitq), 
to_sfixed(1007731953.0/4294967296.0,1,-nbitq), 
to_sfixed(495823812.0/4294967296.0,1,-nbitq), 
to_sfixed(103963608.0/4294967296.0,1,-nbitq), 
to_sfixed(234973688.0/4294967296.0,1,-nbitq), 
to_sfixed(-1960892411.0/4294967296.0,1,-nbitq), 
to_sfixed(277172078.0/4294967296.0,1,-nbitq), 
to_sfixed(496317696.0/4294967296.0,1,-nbitq), 
to_sfixed(-70778759.0/4294967296.0,1,-nbitq), 
to_sfixed(-473935586.0/4294967296.0,1,-nbitq), 
to_sfixed(19288879.0/4294967296.0,1,-nbitq), 
to_sfixed(-51658841.0/4294967296.0,1,-nbitq), 
to_sfixed(138055614.0/4294967296.0,1,-nbitq), 
to_sfixed(-113221973.0/4294967296.0,1,-nbitq), 
to_sfixed(-6330844.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(689188744.0/4294967296.0,1,-nbitq), 
to_sfixed(-1091874331.0/4294967296.0,1,-nbitq), 
to_sfixed(-11964185.0/4294967296.0,1,-nbitq), 
to_sfixed(729144743.0/4294967296.0,1,-nbitq), 
to_sfixed(-1292028674.0/4294967296.0,1,-nbitq), 
to_sfixed(-877289189.0/4294967296.0,1,-nbitq), 
to_sfixed(12672581.0/4294967296.0,1,-nbitq), 
to_sfixed(-811217426.0/4294967296.0,1,-nbitq), 
to_sfixed(-830389268.0/4294967296.0,1,-nbitq), 
to_sfixed(-265239859.0/4294967296.0,1,-nbitq), 
to_sfixed(-500535456.0/4294967296.0,1,-nbitq), 
to_sfixed(853269656.0/4294967296.0,1,-nbitq), 
to_sfixed(-708617906.0/4294967296.0,1,-nbitq), 
to_sfixed(-190758235.0/4294967296.0,1,-nbitq), 
to_sfixed(-175661018.0/4294967296.0,1,-nbitq), 
to_sfixed(81897301.0/4294967296.0,1,-nbitq), 
to_sfixed(167749522.0/4294967296.0,1,-nbitq), 
to_sfixed(-39277560.0/4294967296.0,1,-nbitq), 
to_sfixed(715263170.0/4294967296.0,1,-nbitq), 
to_sfixed(-844153833.0/4294967296.0,1,-nbitq), 
to_sfixed(5994054.0/4294967296.0,1,-nbitq), 
to_sfixed(499989309.0/4294967296.0,1,-nbitq), 
to_sfixed(516309002.0/4294967296.0,1,-nbitq), 
to_sfixed(-136576539.0/4294967296.0,1,-nbitq), 
to_sfixed(150202607.0/4294967296.0,1,-nbitq), 
to_sfixed(-898655176.0/4294967296.0,1,-nbitq), 
to_sfixed(-108560013.0/4294967296.0,1,-nbitq), 
to_sfixed(-780125370.0/4294967296.0,1,-nbitq), 
to_sfixed(-406579817.0/4294967296.0,1,-nbitq), 
to_sfixed(307813867.0/4294967296.0,1,-nbitq), 
to_sfixed(560274397.0/4294967296.0,1,-nbitq), 
to_sfixed(-244263074.0/4294967296.0,1,-nbitq), 
to_sfixed(704668530.0/4294967296.0,1,-nbitq), 
to_sfixed(-254717049.0/4294967296.0,1,-nbitq), 
to_sfixed(239070334.0/4294967296.0,1,-nbitq), 
to_sfixed(993146331.0/4294967296.0,1,-nbitq), 
to_sfixed(175161786.0/4294967296.0,1,-nbitq), 
to_sfixed(-294776305.0/4294967296.0,1,-nbitq), 
to_sfixed(189333356.0/4294967296.0,1,-nbitq), 
to_sfixed(99513147.0/4294967296.0,1,-nbitq), 
to_sfixed(-375460404.0/4294967296.0,1,-nbitq), 
to_sfixed(-291544032.0/4294967296.0,1,-nbitq), 
to_sfixed(1082207488.0/4294967296.0,1,-nbitq), 
to_sfixed(616217585.0/4294967296.0,1,-nbitq), 
to_sfixed(165337252.0/4294967296.0,1,-nbitq), 
to_sfixed(-242021892.0/4294967296.0,1,-nbitq), 
to_sfixed(-238088086.0/4294967296.0,1,-nbitq), 
to_sfixed(463193130.0/4294967296.0,1,-nbitq), 
to_sfixed(-478253435.0/4294967296.0,1,-nbitq), 
to_sfixed(1007356905.0/4294967296.0,1,-nbitq), 
to_sfixed(225254855.0/4294967296.0,1,-nbitq), 
to_sfixed(820390695.0/4294967296.0,1,-nbitq), 
to_sfixed(521035092.0/4294967296.0,1,-nbitq), 
to_sfixed(131277608.0/4294967296.0,1,-nbitq), 
to_sfixed(65139529.0/4294967296.0,1,-nbitq), 
to_sfixed(220332186.0/4294967296.0,1,-nbitq), 
to_sfixed(-268695634.0/4294967296.0,1,-nbitq), 
to_sfixed(34091002.0/4294967296.0,1,-nbitq), 
to_sfixed(211108590.0/4294967296.0,1,-nbitq), 
to_sfixed(167836318.0/4294967296.0,1,-nbitq), 
to_sfixed(213656995.0/4294967296.0,1,-nbitq), 
to_sfixed(725481363.0/4294967296.0,1,-nbitq), 
to_sfixed(-236386191.0/4294967296.0,1,-nbitq), 
to_sfixed(-232408314.0/4294967296.0,1,-nbitq), 
to_sfixed(146898269.0/4294967296.0,1,-nbitq), 
to_sfixed(398500760.0/4294967296.0,1,-nbitq), 
to_sfixed(-52874364.0/4294967296.0,1,-nbitq), 
to_sfixed(1066756146.0/4294967296.0,1,-nbitq), 
to_sfixed(94813141.0/4294967296.0,1,-nbitq), 
to_sfixed(354762266.0/4294967296.0,1,-nbitq), 
to_sfixed(-1141630596.0/4294967296.0,1,-nbitq), 
to_sfixed(27557636.0/4294967296.0,1,-nbitq), 
to_sfixed(-313646332.0/4294967296.0,1,-nbitq), 
to_sfixed(-58751511.0/4294967296.0,1,-nbitq), 
to_sfixed(245590415.0/4294967296.0,1,-nbitq), 
to_sfixed(1077054790.0/4294967296.0,1,-nbitq), 
to_sfixed(484544503.0/4294967296.0,1,-nbitq), 
to_sfixed(72588524.0/4294967296.0,1,-nbitq), 
to_sfixed(-36062235.0/4294967296.0,1,-nbitq), 
to_sfixed(-251466491.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(274510123.0/4294967296.0,1,-nbitq), 
to_sfixed(531307984.0/4294967296.0,1,-nbitq), 
to_sfixed(-1305201867.0/4294967296.0,1,-nbitq), 
to_sfixed(566531988.0/4294967296.0,1,-nbitq), 
to_sfixed(-638256663.0/4294967296.0,1,-nbitq), 
to_sfixed(-785883622.0/4294967296.0,1,-nbitq), 
to_sfixed(388216735.0/4294967296.0,1,-nbitq), 
to_sfixed(-99876297.0/4294967296.0,1,-nbitq), 
to_sfixed(-536633622.0/4294967296.0,1,-nbitq), 
to_sfixed(-203916283.0/4294967296.0,1,-nbitq), 
to_sfixed(319848710.0/4294967296.0,1,-nbitq), 
to_sfixed(371667101.0/4294967296.0,1,-nbitq), 
to_sfixed(-175033815.0/4294967296.0,1,-nbitq), 
to_sfixed(684726274.0/4294967296.0,1,-nbitq), 
to_sfixed(-272759853.0/4294967296.0,1,-nbitq), 
to_sfixed(48518933.0/4294967296.0,1,-nbitq), 
to_sfixed(-65714842.0/4294967296.0,1,-nbitq), 
to_sfixed(-203597292.0/4294967296.0,1,-nbitq), 
to_sfixed(1143743716.0/4294967296.0,1,-nbitq), 
to_sfixed(-600913195.0/4294967296.0,1,-nbitq), 
to_sfixed(-63532163.0/4294967296.0,1,-nbitq), 
to_sfixed(-419991651.0/4294967296.0,1,-nbitq), 
to_sfixed(349118324.0/4294967296.0,1,-nbitq), 
to_sfixed(302100220.0/4294967296.0,1,-nbitq), 
to_sfixed(-57203684.0/4294967296.0,1,-nbitq), 
to_sfixed(-289190020.0/4294967296.0,1,-nbitq), 
to_sfixed(-460027410.0/4294967296.0,1,-nbitq), 
to_sfixed(-586266021.0/4294967296.0,1,-nbitq), 
to_sfixed(-291991502.0/4294967296.0,1,-nbitq), 
to_sfixed(667436468.0/4294967296.0,1,-nbitq), 
to_sfixed(-541529677.0/4294967296.0,1,-nbitq), 
to_sfixed(-237151597.0/4294967296.0,1,-nbitq), 
to_sfixed(679546621.0/4294967296.0,1,-nbitq), 
to_sfixed(235376582.0/4294967296.0,1,-nbitq), 
to_sfixed(535659017.0/4294967296.0,1,-nbitq), 
to_sfixed(1237553932.0/4294967296.0,1,-nbitq), 
to_sfixed(66368753.0/4294967296.0,1,-nbitq), 
to_sfixed(-2002191.0/4294967296.0,1,-nbitq), 
to_sfixed(-11789251.0/4294967296.0,1,-nbitq), 
to_sfixed(16405834.0/4294967296.0,1,-nbitq), 
to_sfixed(285902726.0/4294967296.0,1,-nbitq), 
to_sfixed(-527301102.0/4294967296.0,1,-nbitq), 
to_sfixed(893369992.0/4294967296.0,1,-nbitq), 
to_sfixed(801859023.0/4294967296.0,1,-nbitq), 
to_sfixed(465869096.0/4294967296.0,1,-nbitq), 
to_sfixed(-975335047.0/4294967296.0,1,-nbitq), 
to_sfixed(330533431.0/4294967296.0,1,-nbitq), 
to_sfixed(292060850.0/4294967296.0,1,-nbitq), 
to_sfixed(-522008303.0/4294967296.0,1,-nbitq), 
to_sfixed(1118991662.0/4294967296.0,1,-nbitq), 
to_sfixed(138725689.0/4294967296.0,1,-nbitq), 
to_sfixed(20636576.0/4294967296.0,1,-nbitq), 
to_sfixed(1017533184.0/4294967296.0,1,-nbitq), 
to_sfixed(382999329.0/4294967296.0,1,-nbitq), 
to_sfixed(387270920.0/4294967296.0,1,-nbitq), 
to_sfixed(658000151.0/4294967296.0,1,-nbitq), 
to_sfixed(-568626751.0/4294967296.0,1,-nbitq), 
to_sfixed(-59841096.0/4294967296.0,1,-nbitq), 
to_sfixed(-129937562.0/4294967296.0,1,-nbitq), 
to_sfixed(267565521.0/4294967296.0,1,-nbitq), 
to_sfixed(88620502.0/4294967296.0,1,-nbitq), 
to_sfixed(582975572.0/4294967296.0,1,-nbitq), 
to_sfixed(327448609.0/4294967296.0,1,-nbitq), 
to_sfixed(-221492570.0/4294967296.0,1,-nbitq), 
to_sfixed(-459213519.0/4294967296.0,1,-nbitq), 
to_sfixed(-267314241.0/4294967296.0,1,-nbitq), 
to_sfixed(368852437.0/4294967296.0,1,-nbitq), 
to_sfixed(998297642.0/4294967296.0,1,-nbitq), 
to_sfixed(-172523840.0/4294967296.0,1,-nbitq), 
to_sfixed(98439061.0/4294967296.0,1,-nbitq), 
to_sfixed(-261797544.0/4294967296.0,1,-nbitq), 
to_sfixed(-392487978.0/4294967296.0,1,-nbitq), 
to_sfixed(288778559.0/4294967296.0,1,-nbitq), 
to_sfixed(274090729.0/4294967296.0,1,-nbitq), 
to_sfixed(-408505523.0/4294967296.0,1,-nbitq), 
to_sfixed(437068331.0/4294967296.0,1,-nbitq), 
to_sfixed(-440386462.0/4294967296.0,1,-nbitq), 
to_sfixed(-147244764.0/4294967296.0,1,-nbitq), 
to_sfixed(100676268.0/4294967296.0,1,-nbitq), 
to_sfixed(-393056785.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(25272749.0/4294967296.0,1,-nbitq), 
to_sfixed(170112490.0/4294967296.0,1,-nbitq), 
to_sfixed(-206735392.0/4294967296.0,1,-nbitq), 
to_sfixed(666025061.0/4294967296.0,1,-nbitq), 
to_sfixed(-329810617.0/4294967296.0,1,-nbitq), 
to_sfixed(-632776523.0/4294967296.0,1,-nbitq), 
to_sfixed(117564511.0/4294967296.0,1,-nbitq), 
to_sfixed(-404867133.0/4294967296.0,1,-nbitq), 
to_sfixed(630476920.0/4294967296.0,1,-nbitq), 
to_sfixed(122307379.0/4294967296.0,1,-nbitq), 
to_sfixed(599112989.0/4294967296.0,1,-nbitq), 
to_sfixed(366418773.0/4294967296.0,1,-nbitq), 
to_sfixed(-508759491.0/4294967296.0,1,-nbitq), 
to_sfixed(1276218145.0/4294967296.0,1,-nbitq), 
to_sfixed(312301743.0/4294967296.0,1,-nbitq), 
to_sfixed(-212782274.0/4294967296.0,1,-nbitq), 
to_sfixed(313895221.0/4294967296.0,1,-nbitq), 
to_sfixed(-331837310.0/4294967296.0,1,-nbitq), 
to_sfixed(934190655.0/4294967296.0,1,-nbitq), 
to_sfixed(-213445558.0/4294967296.0,1,-nbitq), 
to_sfixed(32593024.0/4294967296.0,1,-nbitq), 
to_sfixed(-474470735.0/4294967296.0,1,-nbitq), 
to_sfixed(504398886.0/4294967296.0,1,-nbitq), 
to_sfixed(301389562.0/4294967296.0,1,-nbitq), 
to_sfixed(-121985131.0/4294967296.0,1,-nbitq), 
to_sfixed(-191884880.0/4294967296.0,1,-nbitq), 
to_sfixed(-316454678.0/4294967296.0,1,-nbitq), 
to_sfixed(-884925813.0/4294967296.0,1,-nbitq), 
to_sfixed(-498521401.0/4294967296.0,1,-nbitq), 
to_sfixed(-579494538.0/4294967296.0,1,-nbitq), 
to_sfixed(-696379966.0/4294967296.0,1,-nbitq), 
to_sfixed(-107204126.0/4294967296.0,1,-nbitq), 
to_sfixed(529154514.0/4294967296.0,1,-nbitq), 
to_sfixed(285919610.0/4294967296.0,1,-nbitq), 
to_sfixed(684833994.0/4294967296.0,1,-nbitq), 
to_sfixed(901848157.0/4294967296.0,1,-nbitq), 
to_sfixed(1096708671.0/4294967296.0,1,-nbitq), 
to_sfixed(-121534104.0/4294967296.0,1,-nbitq), 
to_sfixed(-347389898.0/4294967296.0,1,-nbitq), 
to_sfixed(-16096769.0/4294967296.0,1,-nbitq), 
to_sfixed(-272136994.0/4294967296.0,1,-nbitq), 
to_sfixed(-206869887.0/4294967296.0,1,-nbitq), 
to_sfixed(1290468033.0/4294967296.0,1,-nbitq), 
to_sfixed(941635981.0/4294967296.0,1,-nbitq), 
to_sfixed(92927851.0/4294967296.0,1,-nbitq), 
to_sfixed(109406751.0/4294967296.0,1,-nbitq), 
to_sfixed(-148566988.0/4294967296.0,1,-nbitq), 
to_sfixed(695921337.0/4294967296.0,1,-nbitq), 
to_sfixed(-119116028.0/4294967296.0,1,-nbitq), 
to_sfixed(652131758.0/4294967296.0,1,-nbitq), 
to_sfixed(-503997148.0/4294967296.0,1,-nbitq), 
to_sfixed(103496396.0/4294967296.0,1,-nbitq), 
to_sfixed(-667938771.0/4294967296.0,1,-nbitq), 
to_sfixed(950240852.0/4294967296.0,1,-nbitq), 
to_sfixed(1050970473.0/4294967296.0,1,-nbitq), 
to_sfixed(748968828.0/4294967296.0,1,-nbitq), 
to_sfixed(-260341076.0/4294967296.0,1,-nbitq), 
to_sfixed(-761048298.0/4294967296.0,1,-nbitq), 
to_sfixed(310266946.0/4294967296.0,1,-nbitq), 
to_sfixed(2551450.0/4294967296.0,1,-nbitq), 
to_sfixed(138201568.0/4294967296.0,1,-nbitq), 
to_sfixed(504924342.0/4294967296.0,1,-nbitq), 
to_sfixed(19861553.0/4294967296.0,1,-nbitq), 
to_sfixed(-126973346.0/4294967296.0,1,-nbitq), 
to_sfixed(-540449252.0/4294967296.0,1,-nbitq), 
to_sfixed(154489554.0/4294967296.0,1,-nbitq), 
to_sfixed(-328131868.0/4294967296.0,1,-nbitq), 
to_sfixed(739610015.0/4294967296.0,1,-nbitq), 
to_sfixed(20881033.0/4294967296.0,1,-nbitq), 
to_sfixed(-967542469.0/4294967296.0,1,-nbitq), 
to_sfixed(-717962827.0/4294967296.0,1,-nbitq), 
to_sfixed(-180320179.0/4294967296.0,1,-nbitq), 
to_sfixed(-344655062.0/4294967296.0,1,-nbitq), 
to_sfixed(182008378.0/4294967296.0,1,-nbitq), 
to_sfixed(-83459476.0/4294967296.0,1,-nbitq), 
to_sfixed(497326918.0/4294967296.0,1,-nbitq), 
to_sfixed(195340281.0/4294967296.0,1,-nbitq), 
to_sfixed(285415747.0/4294967296.0,1,-nbitq), 
to_sfixed(234537026.0/4294967296.0,1,-nbitq), 
to_sfixed(201611504.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(15632145.0/4294967296.0,1,-nbitq), 
to_sfixed(216611204.0/4294967296.0,1,-nbitq), 
to_sfixed(-8346952.0/4294967296.0,1,-nbitq), 
to_sfixed(-56145882.0/4294967296.0,1,-nbitq), 
to_sfixed(-753627832.0/4294967296.0,1,-nbitq), 
to_sfixed(-313635226.0/4294967296.0,1,-nbitq), 
to_sfixed(132925948.0/4294967296.0,1,-nbitq), 
to_sfixed(-534953435.0/4294967296.0,1,-nbitq), 
to_sfixed(245116937.0/4294967296.0,1,-nbitq), 
to_sfixed(-389363728.0/4294967296.0,1,-nbitq), 
to_sfixed(760478959.0/4294967296.0,1,-nbitq), 
to_sfixed(199907527.0/4294967296.0,1,-nbitq), 
to_sfixed(-705972799.0/4294967296.0,1,-nbitq), 
to_sfixed(207341870.0/4294967296.0,1,-nbitq), 
to_sfixed(-263554735.0/4294967296.0,1,-nbitq), 
to_sfixed(265851483.0/4294967296.0,1,-nbitq), 
to_sfixed(43682959.0/4294967296.0,1,-nbitq), 
to_sfixed(44908754.0/4294967296.0,1,-nbitq), 
to_sfixed(846748873.0/4294967296.0,1,-nbitq), 
to_sfixed(-328612012.0/4294967296.0,1,-nbitq), 
to_sfixed(-359608935.0/4294967296.0,1,-nbitq), 
to_sfixed(-361181216.0/4294967296.0,1,-nbitq), 
to_sfixed(-311194196.0/4294967296.0,1,-nbitq), 
to_sfixed(134803672.0/4294967296.0,1,-nbitq), 
to_sfixed(187459788.0/4294967296.0,1,-nbitq), 
to_sfixed(291587407.0/4294967296.0,1,-nbitq), 
to_sfixed(-455595988.0/4294967296.0,1,-nbitq), 
to_sfixed(223782114.0/4294967296.0,1,-nbitq), 
to_sfixed(-547045039.0/4294967296.0,1,-nbitq), 
to_sfixed(-712251437.0/4294967296.0,1,-nbitq), 
to_sfixed(-735285337.0/4294967296.0,1,-nbitq), 
to_sfixed(-811648096.0/4294967296.0,1,-nbitq), 
to_sfixed(220660924.0/4294967296.0,1,-nbitq), 
to_sfixed(-78400081.0/4294967296.0,1,-nbitq), 
to_sfixed(613241308.0/4294967296.0,1,-nbitq), 
to_sfixed(1053650107.0/4294967296.0,1,-nbitq), 
to_sfixed(189698892.0/4294967296.0,1,-nbitq), 
to_sfixed(1357148524.0/4294967296.0,1,-nbitq), 
to_sfixed(-332324084.0/4294967296.0,1,-nbitq), 
to_sfixed(-293186874.0/4294967296.0,1,-nbitq), 
to_sfixed(56487063.0/4294967296.0,1,-nbitq), 
to_sfixed(-817281759.0/4294967296.0,1,-nbitq), 
to_sfixed(837239105.0/4294967296.0,1,-nbitq), 
to_sfixed(960486969.0/4294967296.0,1,-nbitq), 
to_sfixed(193577486.0/4294967296.0,1,-nbitq), 
to_sfixed(171678608.0/4294967296.0,1,-nbitq), 
to_sfixed(68507900.0/4294967296.0,1,-nbitq), 
to_sfixed(835124734.0/4294967296.0,1,-nbitq), 
to_sfixed(-588191410.0/4294967296.0,1,-nbitq), 
to_sfixed(1038491348.0/4294967296.0,1,-nbitq), 
to_sfixed(-431630844.0/4294967296.0,1,-nbitq), 
to_sfixed(-244868304.0/4294967296.0,1,-nbitq), 
to_sfixed(-379473050.0/4294967296.0,1,-nbitq), 
to_sfixed(796506430.0/4294967296.0,1,-nbitq), 
to_sfixed(1407536664.0/4294967296.0,1,-nbitq), 
to_sfixed(-296176193.0/4294967296.0,1,-nbitq), 
to_sfixed(-284194977.0/4294967296.0,1,-nbitq), 
to_sfixed(-1161717807.0/4294967296.0,1,-nbitq), 
to_sfixed(211716761.0/4294967296.0,1,-nbitq), 
to_sfixed(-321257188.0/4294967296.0,1,-nbitq), 
to_sfixed(-338114252.0/4294967296.0,1,-nbitq), 
to_sfixed(1001279483.0/4294967296.0,1,-nbitq), 
to_sfixed(-952125303.0/4294967296.0,1,-nbitq), 
to_sfixed(-607220059.0/4294967296.0,1,-nbitq), 
to_sfixed(-447068375.0/4294967296.0,1,-nbitq), 
to_sfixed(26329998.0/4294967296.0,1,-nbitq), 
to_sfixed(-712526983.0/4294967296.0,1,-nbitq), 
to_sfixed(1534659398.0/4294967296.0,1,-nbitq), 
to_sfixed(205908842.0/4294967296.0,1,-nbitq), 
to_sfixed(-222296761.0/4294967296.0,1,-nbitq), 
to_sfixed(22809226.0/4294967296.0,1,-nbitq), 
to_sfixed(-316744292.0/4294967296.0,1,-nbitq), 
to_sfixed(-187916971.0/4294967296.0,1,-nbitq), 
to_sfixed(122572457.0/4294967296.0,1,-nbitq), 
to_sfixed(-29775891.0/4294967296.0,1,-nbitq), 
to_sfixed(522206859.0/4294967296.0,1,-nbitq), 
to_sfixed(300529806.0/4294967296.0,1,-nbitq), 
to_sfixed(-240151234.0/4294967296.0,1,-nbitq), 
to_sfixed(340244411.0/4294967296.0,1,-nbitq), 
to_sfixed(351347843.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(759853724.0/4294967296.0,1,-nbitq), 
to_sfixed(-737086606.0/4294967296.0,1,-nbitq), 
to_sfixed(-278149745.0/4294967296.0,1,-nbitq), 
to_sfixed(-93644776.0/4294967296.0,1,-nbitq), 
to_sfixed(-380387390.0/4294967296.0,1,-nbitq), 
to_sfixed(318395131.0/4294967296.0,1,-nbitq), 
to_sfixed(295114326.0/4294967296.0,1,-nbitq), 
to_sfixed(-213156335.0/4294967296.0,1,-nbitq), 
to_sfixed(-451017108.0/4294967296.0,1,-nbitq), 
to_sfixed(-180223388.0/4294967296.0,1,-nbitq), 
to_sfixed(75889337.0/4294967296.0,1,-nbitq), 
to_sfixed(278312554.0/4294967296.0,1,-nbitq), 
to_sfixed(-777206814.0/4294967296.0,1,-nbitq), 
to_sfixed(514173470.0/4294967296.0,1,-nbitq), 
to_sfixed(117846662.0/4294967296.0,1,-nbitq), 
to_sfixed(74118251.0/4294967296.0,1,-nbitq), 
to_sfixed(-248826517.0/4294967296.0,1,-nbitq), 
to_sfixed(390483792.0/4294967296.0,1,-nbitq), 
to_sfixed(930140304.0/4294967296.0,1,-nbitq), 
to_sfixed(139988708.0/4294967296.0,1,-nbitq), 
to_sfixed(329755694.0/4294967296.0,1,-nbitq), 
to_sfixed(-848179401.0/4294967296.0,1,-nbitq), 
to_sfixed(-383741948.0/4294967296.0,1,-nbitq), 
to_sfixed(354119119.0/4294967296.0,1,-nbitq), 
to_sfixed(-39973783.0/4294967296.0,1,-nbitq), 
to_sfixed(617414326.0/4294967296.0,1,-nbitq), 
to_sfixed(-225535857.0/4294967296.0,1,-nbitq), 
to_sfixed(-46439583.0/4294967296.0,1,-nbitq), 
to_sfixed(-109529222.0/4294967296.0,1,-nbitq), 
to_sfixed(117671722.0/4294967296.0,1,-nbitq), 
to_sfixed(-350707689.0/4294967296.0,1,-nbitq), 
to_sfixed(-1076065271.0/4294967296.0,1,-nbitq), 
to_sfixed(60060409.0/4294967296.0,1,-nbitq), 
to_sfixed(-211620614.0/4294967296.0,1,-nbitq), 
to_sfixed(-54045452.0/4294967296.0,1,-nbitq), 
to_sfixed(946732053.0/4294967296.0,1,-nbitq), 
to_sfixed(-4255729.0/4294967296.0,1,-nbitq), 
to_sfixed(771486676.0/4294967296.0,1,-nbitq), 
to_sfixed(499977937.0/4294967296.0,1,-nbitq), 
to_sfixed(219890155.0/4294967296.0,1,-nbitq), 
to_sfixed(783044865.0/4294967296.0,1,-nbitq), 
to_sfixed(-169935967.0/4294967296.0,1,-nbitq), 
to_sfixed(413887357.0/4294967296.0,1,-nbitq), 
to_sfixed(526366680.0/4294967296.0,1,-nbitq), 
to_sfixed(289202637.0/4294967296.0,1,-nbitq), 
to_sfixed(-94484380.0/4294967296.0,1,-nbitq), 
to_sfixed(114045957.0/4294967296.0,1,-nbitq), 
to_sfixed(632115169.0/4294967296.0,1,-nbitq), 
to_sfixed(-413476755.0/4294967296.0,1,-nbitq), 
to_sfixed(187339796.0/4294967296.0,1,-nbitq), 
to_sfixed(-92019581.0/4294967296.0,1,-nbitq), 
to_sfixed(645485727.0/4294967296.0,1,-nbitq), 
to_sfixed(-382435394.0/4294967296.0,1,-nbitq), 
to_sfixed(296935641.0/4294967296.0,1,-nbitq), 
to_sfixed(660376841.0/4294967296.0,1,-nbitq), 
to_sfixed(-259834466.0/4294967296.0,1,-nbitq), 
to_sfixed(-50316030.0/4294967296.0,1,-nbitq), 
to_sfixed(-974600001.0/4294967296.0,1,-nbitq), 
to_sfixed(454970312.0/4294967296.0,1,-nbitq), 
to_sfixed(359845090.0/4294967296.0,1,-nbitq), 
to_sfixed(329027192.0/4294967296.0,1,-nbitq), 
to_sfixed(722323499.0/4294967296.0,1,-nbitq), 
to_sfixed(-1075147963.0/4294967296.0,1,-nbitq), 
to_sfixed(-486043507.0/4294967296.0,1,-nbitq), 
to_sfixed(-191806841.0/4294967296.0,1,-nbitq), 
to_sfixed(300707752.0/4294967296.0,1,-nbitq), 
to_sfixed(-619430681.0/4294967296.0,1,-nbitq), 
to_sfixed(1393842937.0/4294967296.0,1,-nbitq), 
to_sfixed(-264624972.0/4294967296.0,1,-nbitq), 
to_sfixed(-697356696.0/4294967296.0,1,-nbitq), 
to_sfixed(641778201.0/4294967296.0,1,-nbitq), 
to_sfixed(4692.0/4294967296.0,1,-nbitq), 
to_sfixed(195088105.0/4294967296.0,1,-nbitq), 
to_sfixed(376750572.0/4294967296.0,1,-nbitq), 
to_sfixed(-224671449.0/4294967296.0,1,-nbitq), 
to_sfixed(-108031415.0/4294967296.0,1,-nbitq), 
to_sfixed(-63341416.0/4294967296.0,1,-nbitq), 
to_sfixed(65324534.0/4294967296.0,1,-nbitq), 
to_sfixed(90018901.0/4294967296.0,1,-nbitq), 
to_sfixed(-20637294.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-106106765.0/4294967296.0,1,-nbitq), 
to_sfixed(19951193.0/4294967296.0,1,-nbitq), 
to_sfixed(279841566.0/4294967296.0,1,-nbitq), 
to_sfixed(-465501010.0/4294967296.0,1,-nbitq), 
to_sfixed(-479224505.0/4294967296.0,1,-nbitq), 
to_sfixed(-111613287.0/4294967296.0,1,-nbitq), 
to_sfixed(-276087987.0/4294967296.0,1,-nbitq), 
to_sfixed(-115682885.0/4294967296.0,1,-nbitq), 
to_sfixed(-259703253.0/4294967296.0,1,-nbitq), 
to_sfixed(-299310244.0/4294967296.0,1,-nbitq), 
to_sfixed(-14422487.0/4294967296.0,1,-nbitq), 
to_sfixed(-599812109.0/4294967296.0,1,-nbitq), 
to_sfixed(-706610231.0/4294967296.0,1,-nbitq), 
to_sfixed(880816402.0/4294967296.0,1,-nbitq), 
to_sfixed(-201234008.0/4294967296.0,1,-nbitq), 
to_sfixed(-512746598.0/4294967296.0,1,-nbitq), 
to_sfixed(-400242920.0/4294967296.0,1,-nbitq), 
to_sfixed(-153178895.0/4294967296.0,1,-nbitq), 
to_sfixed(1082642049.0/4294967296.0,1,-nbitq), 
to_sfixed(-442358692.0/4294967296.0,1,-nbitq), 
to_sfixed(-273339311.0/4294967296.0,1,-nbitq), 
to_sfixed(-489548052.0/4294967296.0,1,-nbitq), 
to_sfixed(-670465833.0/4294967296.0,1,-nbitq), 
to_sfixed(536801516.0/4294967296.0,1,-nbitq), 
to_sfixed(278383951.0/4294967296.0,1,-nbitq), 
to_sfixed(-471372381.0/4294967296.0,1,-nbitq), 
to_sfixed(-697001288.0/4294967296.0,1,-nbitq), 
to_sfixed(611100908.0/4294967296.0,1,-nbitq), 
to_sfixed(223457903.0/4294967296.0,1,-nbitq), 
to_sfixed(-422086957.0/4294967296.0,1,-nbitq), 
to_sfixed(182251718.0/4294967296.0,1,-nbitq), 
to_sfixed(-615377787.0/4294967296.0,1,-nbitq), 
to_sfixed(-436746330.0/4294967296.0,1,-nbitq), 
to_sfixed(-651842931.0/4294967296.0,1,-nbitq), 
to_sfixed(498423506.0/4294967296.0,1,-nbitq), 
to_sfixed(166820853.0/4294967296.0,1,-nbitq), 
to_sfixed(-29662140.0/4294967296.0,1,-nbitq), 
to_sfixed(392951870.0/4294967296.0,1,-nbitq), 
to_sfixed(75379609.0/4294967296.0,1,-nbitq), 
to_sfixed(240434041.0/4294967296.0,1,-nbitq), 
to_sfixed(521091457.0/4294967296.0,1,-nbitq), 
to_sfixed(-355554845.0/4294967296.0,1,-nbitq), 
to_sfixed(-56788992.0/4294967296.0,1,-nbitq), 
to_sfixed(1137038314.0/4294967296.0,1,-nbitq), 
to_sfixed(98854226.0/4294967296.0,1,-nbitq), 
to_sfixed(511289205.0/4294967296.0,1,-nbitq), 
to_sfixed(286670497.0/4294967296.0,1,-nbitq), 
to_sfixed(758360293.0/4294967296.0,1,-nbitq), 
to_sfixed(-340052156.0/4294967296.0,1,-nbitq), 
to_sfixed(456816073.0/4294967296.0,1,-nbitq), 
to_sfixed(160241864.0/4294967296.0,1,-nbitq), 
to_sfixed(34378569.0/4294967296.0,1,-nbitq), 
to_sfixed(-664579766.0/4294967296.0,1,-nbitq), 
to_sfixed(385934439.0/4294967296.0,1,-nbitq), 
to_sfixed(-101599028.0/4294967296.0,1,-nbitq), 
to_sfixed(40460868.0/4294967296.0,1,-nbitq), 
to_sfixed(253306930.0/4294967296.0,1,-nbitq), 
to_sfixed(-1115382318.0/4294967296.0,1,-nbitq), 
to_sfixed(415262573.0/4294967296.0,1,-nbitq), 
to_sfixed(-147365904.0/4294967296.0,1,-nbitq), 
to_sfixed(-262052014.0/4294967296.0,1,-nbitq), 
to_sfixed(526976526.0/4294967296.0,1,-nbitq), 
to_sfixed(-511325851.0/4294967296.0,1,-nbitq), 
to_sfixed(-321788801.0/4294967296.0,1,-nbitq), 
to_sfixed(382962800.0/4294967296.0,1,-nbitq), 
to_sfixed(231477671.0/4294967296.0,1,-nbitq), 
to_sfixed(-85863304.0/4294967296.0,1,-nbitq), 
to_sfixed(1342722258.0/4294967296.0,1,-nbitq), 
to_sfixed(-217577143.0/4294967296.0,1,-nbitq), 
to_sfixed(-406728989.0/4294967296.0,1,-nbitq), 
to_sfixed(-121214201.0/4294967296.0,1,-nbitq), 
to_sfixed(-205591214.0/4294967296.0,1,-nbitq), 
to_sfixed(624596654.0/4294967296.0,1,-nbitq), 
to_sfixed(-9725920.0/4294967296.0,1,-nbitq), 
to_sfixed(475826217.0/4294967296.0,1,-nbitq), 
to_sfixed(604747767.0/4294967296.0,1,-nbitq), 
to_sfixed(-592825749.0/4294967296.0,1,-nbitq), 
to_sfixed(143270714.0/4294967296.0,1,-nbitq), 
to_sfixed(-137936297.0/4294967296.0,1,-nbitq), 
to_sfixed(-312644467.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-154012322.0/4294967296.0,1,-nbitq), 
to_sfixed(132827952.0/4294967296.0,1,-nbitq), 
to_sfixed(-325888148.0/4294967296.0,1,-nbitq), 
to_sfixed(79434999.0/4294967296.0,1,-nbitq), 
to_sfixed(-457625052.0/4294967296.0,1,-nbitq), 
to_sfixed(344303870.0/4294967296.0,1,-nbitq), 
to_sfixed(320669699.0/4294967296.0,1,-nbitq), 
to_sfixed(-250722732.0/4294967296.0,1,-nbitq), 
to_sfixed(795954946.0/4294967296.0,1,-nbitq), 
to_sfixed(212869172.0/4294967296.0,1,-nbitq), 
to_sfixed(358298105.0/4294967296.0,1,-nbitq), 
to_sfixed(-45275642.0/4294967296.0,1,-nbitq), 
to_sfixed(318162426.0/4294967296.0,1,-nbitq), 
to_sfixed(960878227.0/4294967296.0,1,-nbitq), 
to_sfixed(-87108082.0/4294967296.0,1,-nbitq), 
to_sfixed(84363794.0/4294967296.0,1,-nbitq), 
to_sfixed(-377649628.0/4294967296.0,1,-nbitq), 
to_sfixed(371209775.0/4294967296.0,1,-nbitq), 
to_sfixed(-210289501.0/4294967296.0,1,-nbitq), 
to_sfixed(-188584059.0/4294967296.0,1,-nbitq), 
to_sfixed(-60565642.0/4294967296.0,1,-nbitq), 
to_sfixed(-423344340.0/4294967296.0,1,-nbitq), 
to_sfixed(-719596788.0/4294967296.0,1,-nbitq), 
to_sfixed(-239335809.0/4294967296.0,1,-nbitq), 
to_sfixed(202186203.0/4294967296.0,1,-nbitq), 
to_sfixed(-519201148.0/4294967296.0,1,-nbitq), 
to_sfixed(-570369615.0/4294967296.0,1,-nbitq), 
to_sfixed(840709962.0/4294967296.0,1,-nbitq), 
to_sfixed(-46554393.0/4294967296.0,1,-nbitq), 
to_sfixed(-518508124.0/4294967296.0,1,-nbitq), 
to_sfixed(289285243.0/4294967296.0,1,-nbitq), 
to_sfixed(-420273015.0/4294967296.0,1,-nbitq), 
to_sfixed(-134550417.0/4294967296.0,1,-nbitq), 
to_sfixed(-559834132.0/4294967296.0,1,-nbitq), 
to_sfixed(-156798333.0/4294967296.0,1,-nbitq), 
to_sfixed(134899965.0/4294967296.0,1,-nbitq), 
to_sfixed(-55747467.0/4294967296.0,1,-nbitq), 
to_sfixed(-275873388.0/4294967296.0,1,-nbitq), 
to_sfixed(329938625.0/4294967296.0,1,-nbitq), 
to_sfixed(44363166.0/4294967296.0,1,-nbitq), 
to_sfixed(727603556.0/4294967296.0,1,-nbitq), 
to_sfixed(430966102.0/4294967296.0,1,-nbitq), 
to_sfixed(-147327488.0/4294967296.0,1,-nbitq), 
to_sfixed(674500168.0/4294967296.0,1,-nbitq), 
to_sfixed(379003528.0/4294967296.0,1,-nbitq), 
to_sfixed(278946749.0/4294967296.0,1,-nbitq), 
to_sfixed(-261308588.0/4294967296.0,1,-nbitq), 
to_sfixed(466071120.0/4294967296.0,1,-nbitq), 
to_sfixed(-191430559.0/4294967296.0,1,-nbitq), 
to_sfixed(595827973.0/4294967296.0,1,-nbitq), 
to_sfixed(24838214.0/4294967296.0,1,-nbitq), 
to_sfixed(267873390.0/4294967296.0,1,-nbitq), 
to_sfixed(-466546042.0/4294967296.0,1,-nbitq), 
to_sfixed(401353387.0/4294967296.0,1,-nbitq), 
to_sfixed(450792146.0/4294967296.0,1,-nbitq), 
to_sfixed(750134268.0/4294967296.0,1,-nbitq), 
to_sfixed(221347138.0/4294967296.0,1,-nbitq), 
to_sfixed(-919667573.0/4294967296.0,1,-nbitq), 
to_sfixed(378115259.0/4294967296.0,1,-nbitq), 
to_sfixed(-376631016.0/4294967296.0,1,-nbitq), 
to_sfixed(463147958.0/4294967296.0,1,-nbitq), 
to_sfixed(290133119.0/4294967296.0,1,-nbitq), 
to_sfixed(-380446912.0/4294967296.0,1,-nbitq), 
to_sfixed(-252710429.0/4294967296.0,1,-nbitq), 
to_sfixed(-7771692.0/4294967296.0,1,-nbitq), 
to_sfixed(-285571227.0/4294967296.0,1,-nbitq), 
to_sfixed(75208751.0/4294967296.0,1,-nbitq), 
to_sfixed(562845382.0/4294967296.0,1,-nbitq), 
to_sfixed(252257035.0/4294967296.0,1,-nbitq), 
to_sfixed(114119737.0/4294967296.0,1,-nbitq), 
to_sfixed(-649917819.0/4294967296.0,1,-nbitq), 
to_sfixed(-33046432.0/4294967296.0,1,-nbitq), 
to_sfixed(201862590.0/4294967296.0,1,-nbitq), 
to_sfixed(61561842.0/4294967296.0,1,-nbitq), 
to_sfixed(134258926.0/4294967296.0,1,-nbitq), 
to_sfixed(628995027.0/4294967296.0,1,-nbitq), 
to_sfixed(-370265507.0/4294967296.0,1,-nbitq), 
to_sfixed(83406066.0/4294967296.0,1,-nbitq), 
to_sfixed(286586548.0/4294967296.0,1,-nbitq), 
to_sfixed(37490385.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-109354944.0/4294967296.0,1,-nbitq), 
to_sfixed(-468938975.0/4294967296.0,1,-nbitq), 
to_sfixed(267353797.0/4294967296.0,1,-nbitq), 
to_sfixed(33399002.0/4294967296.0,1,-nbitq), 
to_sfixed(-595477228.0/4294967296.0,1,-nbitq), 
to_sfixed(645685855.0/4294967296.0,1,-nbitq), 
to_sfixed(169824275.0/4294967296.0,1,-nbitq), 
to_sfixed(-452811588.0/4294967296.0,1,-nbitq), 
to_sfixed(467788563.0/4294967296.0,1,-nbitq), 
to_sfixed(-215036206.0/4294967296.0,1,-nbitq), 
to_sfixed(-304615791.0/4294967296.0,1,-nbitq), 
to_sfixed(263103455.0/4294967296.0,1,-nbitq), 
to_sfixed(173709322.0/4294967296.0,1,-nbitq), 
to_sfixed(1260633357.0/4294967296.0,1,-nbitq), 
to_sfixed(-397233000.0/4294967296.0,1,-nbitq), 
to_sfixed(-97509858.0/4294967296.0,1,-nbitq), 
to_sfixed(-406628707.0/4294967296.0,1,-nbitq), 
to_sfixed(5695382.0/4294967296.0,1,-nbitq), 
to_sfixed(-313673578.0/4294967296.0,1,-nbitq), 
to_sfixed(319194319.0/4294967296.0,1,-nbitq), 
to_sfixed(336584012.0/4294967296.0,1,-nbitq), 
to_sfixed(292048507.0/4294967296.0,1,-nbitq), 
to_sfixed(-366389507.0/4294967296.0,1,-nbitq), 
to_sfixed(-381849955.0/4294967296.0,1,-nbitq), 
to_sfixed(-341434604.0/4294967296.0,1,-nbitq), 
to_sfixed(-15910506.0/4294967296.0,1,-nbitq), 
to_sfixed(76205013.0/4294967296.0,1,-nbitq), 
to_sfixed(692274512.0/4294967296.0,1,-nbitq), 
to_sfixed(-444137783.0/4294967296.0,1,-nbitq), 
to_sfixed(-118214805.0/4294967296.0,1,-nbitq), 
to_sfixed(320604082.0/4294967296.0,1,-nbitq), 
to_sfixed(-136193356.0/4294967296.0,1,-nbitq), 
to_sfixed(-823073771.0/4294967296.0,1,-nbitq), 
to_sfixed(-426699500.0/4294967296.0,1,-nbitq), 
to_sfixed(261788420.0/4294967296.0,1,-nbitq), 
to_sfixed(81732882.0/4294967296.0,1,-nbitq), 
to_sfixed(487271549.0/4294967296.0,1,-nbitq), 
to_sfixed(-593885981.0/4294967296.0,1,-nbitq), 
to_sfixed(-9035367.0/4294967296.0,1,-nbitq), 
to_sfixed(80750377.0/4294967296.0,1,-nbitq), 
to_sfixed(262991085.0/4294967296.0,1,-nbitq), 
to_sfixed(150731199.0/4294967296.0,1,-nbitq), 
to_sfixed(47611648.0/4294967296.0,1,-nbitq), 
to_sfixed(949153633.0/4294967296.0,1,-nbitq), 
to_sfixed(382196144.0/4294967296.0,1,-nbitq), 
to_sfixed(65746430.0/4294967296.0,1,-nbitq), 
to_sfixed(247022536.0/4294967296.0,1,-nbitq), 
to_sfixed(259300267.0/4294967296.0,1,-nbitq), 
to_sfixed(-275660804.0/4294967296.0,1,-nbitq), 
to_sfixed(41580388.0/4294967296.0,1,-nbitq), 
to_sfixed(55838830.0/4294967296.0,1,-nbitq), 
to_sfixed(-356208338.0/4294967296.0,1,-nbitq), 
to_sfixed(4447385.0/4294967296.0,1,-nbitq), 
to_sfixed(103169688.0/4294967296.0,1,-nbitq), 
to_sfixed(-340510400.0/4294967296.0,1,-nbitq), 
to_sfixed(496231591.0/4294967296.0,1,-nbitq), 
to_sfixed(33680314.0/4294967296.0,1,-nbitq), 
to_sfixed(-1142314161.0/4294967296.0,1,-nbitq), 
to_sfixed(-89914023.0/4294967296.0,1,-nbitq), 
to_sfixed(25273226.0/4294967296.0,1,-nbitq), 
to_sfixed(296766871.0/4294967296.0,1,-nbitq), 
to_sfixed(-305481989.0/4294967296.0,1,-nbitq), 
to_sfixed(-503771582.0/4294967296.0,1,-nbitq), 
to_sfixed(-176480350.0/4294967296.0,1,-nbitq), 
to_sfixed(203972614.0/4294967296.0,1,-nbitq), 
to_sfixed(-8317566.0/4294967296.0,1,-nbitq), 
to_sfixed(-35065751.0/4294967296.0,1,-nbitq), 
to_sfixed(-459147320.0/4294967296.0,1,-nbitq), 
to_sfixed(-165460511.0/4294967296.0,1,-nbitq), 
to_sfixed(-165723709.0/4294967296.0,1,-nbitq), 
to_sfixed(-476367257.0/4294967296.0,1,-nbitq), 
to_sfixed(414073930.0/4294967296.0,1,-nbitq), 
to_sfixed(-428256007.0/4294967296.0,1,-nbitq), 
to_sfixed(145553070.0/4294967296.0,1,-nbitq), 
to_sfixed(52847573.0/4294967296.0,1,-nbitq), 
to_sfixed(67429397.0/4294967296.0,1,-nbitq), 
to_sfixed(-512708360.0/4294967296.0,1,-nbitq), 
to_sfixed(-2990577.0/4294967296.0,1,-nbitq), 
to_sfixed(694600018.0/4294967296.0,1,-nbitq), 
to_sfixed(146517515.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-82898881.0/4294967296.0,1,-nbitq), 
to_sfixed(-157028366.0/4294967296.0,1,-nbitq), 
to_sfixed(611037251.0/4294967296.0,1,-nbitq), 
to_sfixed(493942234.0/4294967296.0,1,-nbitq), 
to_sfixed(-220852214.0/4294967296.0,1,-nbitq), 
to_sfixed(992022846.0/4294967296.0,1,-nbitq), 
to_sfixed(-8982417.0/4294967296.0,1,-nbitq), 
to_sfixed(122496522.0/4294967296.0,1,-nbitq), 
to_sfixed(467396168.0/4294967296.0,1,-nbitq), 
to_sfixed(-230525971.0/4294967296.0,1,-nbitq), 
to_sfixed(189373912.0/4294967296.0,1,-nbitq), 
to_sfixed(566349235.0/4294967296.0,1,-nbitq), 
to_sfixed(192926749.0/4294967296.0,1,-nbitq), 
to_sfixed(238293521.0/4294967296.0,1,-nbitq), 
to_sfixed(122339397.0/4294967296.0,1,-nbitq), 
to_sfixed(528811540.0/4294967296.0,1,-nbitq), 
to_sfixed(-144417953.0/4294967296.0,1,-nbitq), 
to_sfixed(38017418.0/4294967296.0,1,-nbitq), 
to_sfixed(-151248688.0/4294967296.0,1,-nbitq), 
to_sfixed(-177350339.0/4294967296.0,1,-nbitq), 
to_sfixed(-269917635.0/4294967296.0,1,-nbitq), 
to_sfixed(1120706296.0/4294967296.0,1,-nbitq), 
to_sfixed(-187445874.0/4294967296.0,1,-nbitq), 
to_sfixed(197501829.0/4294967296.0,1,-nbitq), 
to_sfixed(-67985737.0/4294967296.0,1,-nbitq), 
to_sfixed(-180008269.0/4294967296.0,1,-nbitq), 
to_sfixed(279359292.0/4294967296.0,1,-nbitq), 
to_sfixed(674227718.0/4294967296.0,1,-nbitq), 
to_sfixed(287757303.0/4294967296.0,1,-nbitq), 
to_sfixed(-179826869.0/4294967296.0,1,-nbitq), 
to_sfixed(547581021.0/4294967296.0,1,-nbitq), 
to_sfixed(-85038666.0/4294967296.0,1,-nbitq), 
to_sfixed(-136317245.0/4294967296.0,1,-nbitq), 
to_sfixed(-149328687.0/4294967296.0,1,-nbitq), 
to_sfixed(128969687.0/4294967296.0,1,-nbitq), 
to_sfixed(378658266.0/4294967296.0,1,-nbitq), 
to_sfixed(628177443.0/4294967296.0,1,-nbitq), 
to_sfixed(-98180544.0/4294967296.0,1,-nbitq), 
to_sfixed(395784903.0/4294967296.0,1,-nbitq), 
to_sfixed(458947913.0/4294967296.0,1,-nbitq), 
to_sfixed(-285980538.0/4294967296.0,1,-nbitq), 
to_sfixed(650292165.0/4294967296.0,1,-nbitq), 
to_sfixed(-119181722.0/4294967296.0,1,-nbitq), 
to_sfixed(202178105.0/4294967296.0,1,-nbitq), 
to_sfixed(27164309.0/4294967296.0,1,-nbitq), 
to_sfixed(421239112.0/4294967296.0,1,-nbitq), 
to_sfixed(-423311806.0/4294967296.0,1,-nbitq), 
to_sfixed(-31675955.0/4294967296.0,1,-nbitq), 
to_sfixed(170064912.0/4294967296.0,1,-nbitq), 
to_sfixed(-252895325.0/4294967296.0,1,-nbitq), 
to_sfixed(515393227.0/4294967296.0,1,-nbitq), 
to_sfixed(155116225.0/4294967296.0,1,-nbitq), 
to_sfixed(62332253.0/4294967296.0,1,-nbitq), 
to_sfixed(270597122.0/4294967296.0,1,-nbitq), 
to_sfixed(-733592933.0/4294967296.0,1,-nbitq), 
to_sfixed(466403781.0/4294967296.0,1,-nbitq), 
to_sfixed(407606030.0/4294967296.0,1,-nbitq), 
to_sfixed(-1145826303.0/4294967296.0,1,-nbitq), 
to_sfixed(394391427.0/4294967296.0,1,-nbitq), 
to_sfixed(-248206065.0/4294967296.0,1,-nbitq), 
to_sfixed(316661691.0/4294967296.0,1,-nbitq), 
to_sfixed(-190457800.0/4294967296.0,1,-nbitq), 
to_sfixed(-259131401.0/4294967296.0,1,-nbitq), 
to_sfixed(-757115342.0/4294967296.0,1,-nbitq), 
to_sfixed(137581772.0/4294967296.0,1,-nbitq), 
to_sfixed(259270747.0/4294967296.0,1,-nbitq), 
to_sfixed(-243315125.0/4294967296.0,1,-nbitq), 
to_sfixed(361031977.0/4294967296.0,1,-nbitq), 
to_sfixed(67740804.0/4294967296.0,1,-nbitq), 
to_sfixed(-149271883.0/4294967296.0,1,-nbitq), 
to_sfixed(-725169267.0/4294967296.0,1,-nbitq), 
to_sfixed(421466480.0/4294967296.0,1,-nbitq), 
to_sfixed(-179845967.0/4294967296.0,1,-nbitq), 
to_sfixed(309571047.0/4294967296.0,1,-nbitq), 
to_sfixed(-480281897.0/4294967296.0,1,-nbitq), 
to_sfixed(283520570.0/4294967296.0,1,-nbitq), 
to_sfixed(298087752.0/4294967296.0,1,-nbitq), 
to_sfixed(456465216.0/4294967296.0,1,-nbitq), 
to_sfixed(-140286344.0/4294967296.0,1,-nbitq), 
to_sfixed(328009761.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-320176807.0/4294967296.0,1,-nbitq), 
to_sfixed(-24861650.0/4294967296.0,1,-nbitq), 
to_sfixed(865303700.0/4294967296.0,1,-nbitq), 
to_sfixed(-137721442.0/4294967296.0,1,-nbitq), 
to_sfixed(-83434564.0/4294967296.0,1,-nbitq), 
to_sfixed(106918938.0/4294967296.0,1,-nbitq), 
to_sfixed(-144164986.0/4294967296.0,1,-nbitq), 
to_sfixed(505142906.0/4294967296.0,1,-nbitq), 
to_sfixed(187047086.0/4294967296.0,1,-nbitq), 
to_sfixed(-359651478.0/4294967296.0,1,-nbitq), 
to_sfixed(-158940995.0/4294967296.0,1,-nbitq), 
to_sfixed(-52952093.0/4294967296.0,1,-nbitq), 
to_sfixed(-79532683.0/4294967296.0,1,-nbitq), 
to_sfixed(170482254.0/4294967296.0,1,-nbitq), 
to_sfixed(271622691.0/4294967296.0,1,-nbitq), 
to_sfixed(209627502.0/4294967296.0,1,-nbitq), 
to_sfixed(201539467.0/4294967296.0,1,-nbitq), 
to_sfixed(-24665013.0/4294967296.0,1,-nbitq), 
to_sfixed(-349392291.0/4294967296.0,1,-nbitq), 
to_sfixed(-156255828.0/4294967296.0,1,-nbitq), 
to_sfixed(-214468619.0/4294967296.0,1,-nbitq), 
to_sfixed(642799542.0/4294967296.0,1,-nbitq), 
to_sfixed(-258092458.0/4294967296.0,1,-nbitq), 
to_sfixed(458178342.0/4294967296.0,1,-nbitq), 
to_sfixed(388298510.0/4294967296.0,1,-nbitq), 
to_sfixed(-433393685.0/4294967296.0,1,-nbitq), 
to_sfixed(531579154.0/4294967296.0,1,-nbitq), 
to_sfixed(166106060.0/4294967296.0,1,-nbitq), 
to_sfixed(204665668.0/4294967296.0,1,-nbitq), 
to_sfixed(123641554.0/4294967296.0,1,-nbitq), 
to_sfixed(8801069.0/4294967296.0,1,-nbitq), 
to_sfixed(-82484210.0/4294967296.0,1,-nbitq), 
to_sfixed(-145362997.0/4294967296.0,1,-nbitq), 
to_sfixed(104645838.0/4294967296.0,1,-nbitq), 
to_sfixed(-63100192.0/4294967296.0,1,-nbitq), 
to_sfixed(8821770.0/4294967296.0,1,-nbitq), 
to_sfixed(455222586.0/4294967296.0,1,-nbitq), 
to_sfixed(-563342339.0/4294967296.0,1,-nbitq), 
to_sfixed(138432289.0/4294967296.0,1,-nbitq), 
to_sfixed(419162.0/4294967296.0,1,-nbitq), 
to_sfixed(-215188146.0/4294967296.0,1,-nbitq), 
to_sfixed(139537372.0/4294967296.0,1,-nbitq), 
to_sfixed(99079273.0/4294967296.0,1,-nbitq), 
to_sfixed(-107390606.0/4294967296.0,1,-nbitq), 
to_sfixed(-163964659.0/4294967296.0,1,-nbitq), 
to_sfixed(-434129174.0/4294967296.0,1,-nbitq), 
to_sfixed(155769148.0/4294967296.0,1,-nbitq), 
to_sfixed(-332720888.0/4294967296.0,1,-nbitq), 
to_sfixed(-243325043.0/4294967296.0,1,-nbitq), 
to_sfixed(-616836023.0/4294967296.0,1,-nbitq), 
to_sfixed(320672603.0/4294967296.0,1,-nbitq), 
to_sfixed(-114537081.0/4294967296.0,1,-nbitq), 
to_sfixed(-275347740.0/4294967296.0,1,-nbitq), 
to_sfixed(247783252.0/4294967296.0,1,-nbitq), 
to_sfixed(-629720906.0/4294967296.0,1,-nbitq), 
to_sfixed(256681968.0/4294967296.0,1,-nbitq), 
to_sfixed(285005164.0/4294967296.0,1,-nbitq), 
to_sfixed(108358743.0/4294967296.0,1,-nbitq), 
to_sfixed(101249380.0/4294967296.0,1,-nbitq), 
to_sfixed(18863333.0/4294967296.0,1,-nbitq), 
to_sfixed(-187588879.0/4294967296.0,1,-nbitq), 
to_sfixed(-263839072.0/4294967296.0,1,-nbitq), 
to_sfixed(-174229903.0/4294967296.0,1,-nbitq), 
to_sfixed(-83410229.0/4294967296.0,1,-nbitq), 
to_sfixed(-45270790.0/4294967296.0,1,-nbitq), 
to_sfixed(-248034838.0/4294967296.0,1,-nbitq), 
to_sfixed(80609863.0/4294967296.0,1,-nbitq), 
to_sfixed(376632225.0/4294967296.0,1,-nbitq), 
to_sfixed(326769467.0/4294967296.0,1,-nbitq), 
to_sfixed(110192047.0/4294967296.0,1,-nbitq), 
to_sfixed(-397106312.0/4294967296.0,1,-nbitq), 
to_sfixed(437841208.0/4294967296.0,1,-nbitq), 
to_sfixed(9463994.0/4294967296.0,1,-nbitq), 
to_sfixed(422870461.0/4294967296.0,1,-nbitq), 
to_sfixed(248175685.0/4294967296.0,1,-nbitq), 
to_sfixed(118158939.0/4294967296.0,1,-nbitq), 
to_sfixed(47942038.0/4294967296.0,1,-nbitq), 
to_sfixed(-126776248.0/4294967296.0,1,-nbitq), 
to_sfixed(307413665.0/4294967296.0,1,-nbitq), 
to_sfixed(222039696.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(182358789.0/4294967296.0,1,-nbitq), 
to_sfixed(-200667910.0/4294967296.0,1,-nbitq), 
to_sfixed(1039915583.0/4294967296.0,1,-nbitq), 
to_sfixed(155734102.0/4294967296.0,1,-nbitq), 
to_sfixed(-280234104.0/4294967296.0,1,-nbitq), 
to_sfixed(-571533624.0/4294967296.0,1,-nbitq), 
to_sfixed(290714526.0/4294967296.0,1,-nbitq), 
to_sfixed(160455693.0/4294967296.0,1,-nbitq), 
to_sfixed(-447829007.0/4294967296.0,1,-nbitq), 
to_sfixed(8767016.0/4294967296.0,1,-nbitq), 
to_sfixed(281470966.0/4294967296.0,1,-nbitq), 
to_sfixed(279203934.0/4294967296.0,1,-nbitq), 
to_sfixed(-224464123.0/4294967296.0,1,-nbitq), 
to_sfixed(447427607.0/4294967296.0,1,-nbitq), 
to_sfixed(21102987.0/4294967296.0,1,-nbitq), 
to_sfixed(382113648.0/4294967296.0,1,-nbitq), 
to_sfixed(25070154.0/4294967296.0,1,-nbitq), 
to_sfixed(-23818341.0/4294967296.0,1,-nbitq), 
to_sfixed(4610828.0/4294967296.0,1,-nbitq), 
to_sfixed(-375367529.0/4294967296.0,1,-nbitq), 
to_sfixed(-46937447.0/4294967296.0,1,-nbitq), 
to_sfixed(573483568.0/4294967296.0,1,-nbitq), 
to_sfixed(-304250045.0/4294967296.0,1,-nbitq), 
to_sfixed(-133766516.0/4294967296.0,1,-nbitq), 
to_sfixed(400299944.0/4294967296.0,1,-nbitq), 
to_sfixed(-103699617.0/4294967296.0,1,-nbitq), 
to_sfixed(412691683.0/4294967296.0,1,-nbitq), 
to_sfixed(147714847.0/4294967296.0,1,-nbitq), 
to_sfixed(288566987.0/4294967296.0,1,-nbitq), 
to_sfixed(30092552.0/4294967296.0,1,-nbitq), 
to_sfixed(-83321316.0/4294967296.0,1,-nbitq), 
to_sfixed(-170263221.0/4294967296.0,1,-nbitq), 
to_sfixed(16545132.0/4294967296.0,1,-nbitq), 
to_sfixed(166670483.0/4294967296.0,1,-nbitq), 
to_sfixed(-219428106.0/4294967296.0,1,-nbitq), 
to_sfixed(-283501078.0/4294967296.0,1,-nbitq), 
to_sfixed(356854642.0/4294967296.0,1,-nbitq), 
to_sfixed(-433993435.0/4294967296.0,1,-nbitq), 
to_sfixed(-247967966.0/4294967296.0,1,-nbitq), 
to_sfixed(130153981.0/4294967296.0,1,-nbitq), 
to_sfixed(-389629480.0/4294967296.0,1,-nbitq), 
to_sfixed(549046583.0/4294967296.0,1,-nbitq), 
to_sfixed(-252825565.0/4294967296.0,1,-nbitq), 
to_sfixed(-107313704.0/4294967296.0,1,-nbitq), 
to_sfixed(-196212698.0/4294967296.0,1,-nbitq), 
to_sfixed(-216568778.0/4294967296.0,1,-nbitq), 
to_sfixed(-355196804.0/4294967296.0,1,-nbitq), 
to_sfixed(-502526399.0/4294967296.0,1,-nbitq), 
to_sfixed(225802432.0/4294967296.0,1,-nbitq), 
to_sfixed(-561219210.0/4294967296.0,1,-nbitq), 
to_sfixed(-113443900.0/4294967296.0,1,-nbitq), 
to_sfixed(291586944.0/4294967296.0,1,-nbitq), 
to_sfixed(18528975.0/4294967296.0,1,-nbitq), 
to_sfixed(122298971.0/4294967296.0,1,-nbitq), 
to_sfixed(-232557955.0/4294967296.0,1,-nbitq), 
to_sfixed(378331653.0/4294967296.0,1,-nbitq), 
to_sfixed(-292821695.0/4294967296.0,1,-nbitq), 
to_sfixed(-505519696.0/4294967296.0,1,-nbitq), 
to_sfixed(168752883.0/4294967296.0,1,-nbitq), 
to_sfixed(-5326044.0/4294967296.0,1,-nbitq), 
to_sfixed(-147420015.0/4294967296.0,1,-nbitq), 
to_sfixed(62014494.0/4294967296.0,1,-nbitq), 
to_sfixed(-89299083.0/4294967296.0,1,-nbitq), 
to_sfixed(99491514.0/4294967296.0,1,-nbitq), 
to_sfixed(192075615.0/4294967296.0,1,-nbitq), 
to_sfixed(153972389.0/4294967296.0,1,-nbitq), 
to_sfixed(83903199.0/4294967296.0,1,-nbitq), 
to_sfixed(126564991.0/4294967296.0,1,-nbitq), 
to_sfixed(-176711468.0/4294967296.0,1,-nbitq), 
to_sfixed(396109882.0/4294967296.0,1,-nbitq), 
to_sfixed(-439469638.0/4294967296.0,1,-nbitq), 
to_sfixed(244462178.0/4294967296.0,1,-nbitq), 
to_sfixed(-628229391.0/4294967296.0,1,-nbitq), 
to_sfixed(166688221.0/4294967296.0,1,-nbitq), 
to_sfixed(202384996.0/4294967296.0,1,-nbitq), 
to_sfixed(316707187.0/4294967296.0,1,-nbitq), 
to_sfixed(-359733292.0/4294967296.0,1,-nbitq), 
to_sfixed(-424023088.0/4294967296.0,1,-nbitq), 
to_sfixed(-206963089.0/4294967296.0,1,-nbitq), 
to_sfixed(-237964313.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-99413256.0/4294967296.0,1,-nbitq), 
to_sfixed(58382902.0/4294967296.0,1,-nbitq), 
to_sfixed(749315447.0/4294967296.0,1,-nbitq), 
to_sfixed(169571879.0/4294967296.0,1,-nbitq), 
to_sfixed(-86914851.0/4294967296.0,1,-nbitq), 
to_sfixed(3874473.0/4294967296.0,1,-nbitq), 
to_sfixed(364718791.0/4294967296.0,1,-nbitq), 
to_sfixed(4569059.0/4294967296.0,1,-nbitq), 
to_sfixed(190807115.0/4294967296.0,1,-nbitq), 
to_sfixed(77340776.0/4294967296.0,1,-nbitq), 
to_sfixed(91038513.0/4294967296.0,1,-nbitq), 
to_sfixed(156452503.0/4294967296.0,1,-nbitq), 
to_sfixed(-592571589.0/4294967296.0,1,-nbitq), 
to_sfixed(84667275.0/4294967296.0,1,-nbitq), 
to_sfixed(-440331232.0/4294967296.0,1,-nbitq), 
to_sfixed(548770149.0/4294967296.0,1,-nbitq), 
to_sfixed(377125100.0/4294967296.0,1,-nbitq), 
to_sfixed(-60059453.0/4294967296.0,1,-nbitq), 
to_sfixed(-465367898.0/4294967296.0,1,-nbitq), 
to_sfixed(-274170170.0/4294967296.0,1,-nbitq), 
to_sfixed(-229876370.0/4294967296.0,1,-nbitq), 
to_sfixed(461880419.0/4294967296.0,1,-nbitq), 
to_sfixed(386061289.0/4294967296.0,1,-nbitq), 
to_sfixed(306439505.0/4294967296.0,1,-nbitq), 
to_sfixed(377015462.0/4294967296.0,1,-nbitq), 
to_sfixed(351518566.0/4294967296.0,1,-nbitq), 
to_sfixed(11902783.0/4294967296.0,1,-nbitq), 
to_sfixed(111778493.0/4294967296.0,1,-nbitq), 
to_sfixed(-140850054.0/4294967296.0,1,-nbitq), 
to_sfixed(349568896.0/4294967296.0,1,-nbitq), 
to_sfixed(-4766730.0/4294967296.0,1,-nbitq), 
to_sfixed(-224847670.0/4294967296.0,1,-nbitq), 
to_sfixed(-242366080.0/4294967296.0,1,-nbitq), 
to_sfixed(-211057035.0/4294967296.0,1,-nbitq), 
to_sfixed(261066051.0/4294967296.0,1,-nbitq), 
to_sfixed(195392635.0/4294967296.0,1,-nbitq), 
to_sfixed(23736555.0/4294967296.0,1,-nbitq), 
to_sfixed(-261248079.0/4294967296.0,1,-nbitq), 
to_sfixed(5904598.0/4294967296.0,1,-nbitq), 
to_sfixed(-97455311.0/4294967296.0,1,-nbitq), 
to_sfixed(-410237835.0/4294967296.0,1,-nbitq), 
to_sfixed(490143748.0/4294967296.0,1,-nbitq), 
to_sfixed(247117171.0/4294967296.0,1,-nbitq), 
to_sfixed(352951040.0/4294967296.0,1,-nbitq), 
to_sfixed(466608802.0/4294967296.0,1,-nbitq), 
to_sfixed(-343429505.0/4294967296.0,1,-nbitq), 
to_sfixed(-400767618.0/4294967296.0,1,-nbitq), 
to_sfixed(62527542.0/4294967296.0,1,-nbitq), 
to_sfixed(-253231744.0/4294967296.0,1,-nbitq), 
to_sfixed(-338305949.0/4294967296.0,1,-nbitq), 
to_sfixed(-38147872.0/4294967296.0,1,-nbitq), 
to_sfixed(528089179.0/4294967296.0,1,-nbitq), 
to_sfixed(44934782.0/4294967296.0,1,-nbitq), 
to_sfixed(-196024079.0/4294967296.0,1,-nbitq), 
to_sfixed(-286448870.0/4294967296.0,1,-nbitq), 
to_sfixed(17215948.0/4294967296.0,1,-nbitq), 
to_sfixed(-43341584.0/4294967296.0,1,-nbitq), 
to_sfixed(-77338155.0/4294967296.0,1,-nbitq), 
to_sfixed(300600456.0/4294967296.0,1,-nbitq), 
to_sfixed(154590979.0/4294967296.0,1,-nbitq), 
to_sfixed(296356697.0/4294967296.0,1,-nbitq), 
to_sfixed(433277926.0/4294967296.0,1,-nbitq), 
to_sfixed(123565586.0/4294967296.0,1,-nbitq), 
to_sfixed(-146452205.0/4294967296.0,1,-nbitq), 
to_sfixed(-355589107.0/4294967296.0,1,-nbitq), 
to_sfixed(-392881924.0/4294967296.0,1,-nbitq), 
to_sfixed(580362793.0/4294967296.0,1,-nbitq), 
to_sfixed(-150196182.0/4294967296.0,1,-nbitq), 
to_sfixed(-284559509.0/4294967296.0,1,-nbitq), 
to_sfixed(-1034508.0/4294967296.0,1,-nbitq), 
to_sfixed(-402402671.0/4294967296.0,1,-nbitq), 
to_sfixed(-6852528.0/4294967296.0,1,-nbitq), 
to_sfixed(-143350768.0/4294967296.0,1,-nbitq), 
to_sfixed(334473238.0/4294967296.0,1,-nbitq), 
to_sfixed(382429198.0/4294967296.0,1,-nbitq), 
to_sfixed(-466310745.0/4294967296.0,1,-nbitq), 
to_sfixed(-245040162.0/4294967296.0,1,-nbitq), 
to_sfixed(177725500.0/4294967296.0,1,-nbitq), 
to_sfixed(-154878896.0/4294967296.0,1,-nbitq), 
to_sfixed(-262824448.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(247233223.0/4294967296.0,1,-nbitq), 
to_sfixed(172882208.0/4294967296.0,1,-nbitq), 
to_sfixed(50500278.0/4294967296.0,1,-nbitq), 
to_sfixed(-317187631.0/4294967296.0,1,-nbitq), 
to_sfixed(412123258.0/4294967296.0,1,-nbitq), 
to_sfixed(43728912.0/4294967296.0,1,-nbitq), 
to_sfixed(-329049839.0/4294967296.0,1,-nbitq), 
to_sfixed(-390755548.0/4294967296.0,1,-nbitq), 
to_sfixed(79089144.0/4294967296.0,1,-nbitq), 
to_sfixed(-24583110.0/4294967296.0,1,-nbitq), 
to_sfixed(-49727179.0/4294967296.0,1,-nbitq), 
to_sfixed(556003374.0/4294967296.0,1,-nbitq), 
to_sfixed(-60271865.0/4294967296.0,1,-nbitq), 
to_sfixed(165593975.0/4294967296.0,1,-nbitq), 
to_sfixed(12375130.0/4294967296.0,1,-nbitq), 
to_sfixed(125775924.0/4294967296.0,1,-nbitq), 
to_sfixed(-349249183.0/4294967296.0,1,-nbitq), 
to_sfixed(399838606.0/4294967296.0,1,-nbitq), 
to_sfixed(-233720000.0/4294967296.0,1,-nbitq), 
to_sfixed(246437495.0/4294967296.0,1,-nbitq), 
to_sfixed(-151378573.0/4294967296.0,1,-nbitq), 
to_sfixed(210621365.0/4294967296.0,1,-nbitq), 
to_sfixed(415988276.0/4294967296.0,1,-nbitq), 
to_sfixed(28510265.0/4294967296.0,1,-nbitq), 
to_sfixed(-36121990.0/4294967296.0,1,-nbitq), 
to_sfixed(-185566887.0/4294967296.0,1,-nbitq), 
to_sfixed(143922572.0/4294967296.0,1,-nbitq), 
to_sfixed(-446971784.0/4294967296.0,1,-nbitq), 
to_sfixed(477120143.0/4294967296.0,1,-nbitq), 
to_sfixed(-98148290.0/4294967296.0,1,-nbitq), 
to_sfixed(-187054215.0/4294967296.0,1,-nbitq), 
to_sfixed(75827825.0/4294967296.0,1,-nbitq), 
to_sfixed(492529280.0/4294967296.0,1,-nbitq), 
to_sfixed(-460042334.0/4294967296.0,1,-nbitq), 
to_sfixed(-266318575.0/4294967296.0,1,-nbitq), 
to_sfixed(184755307.0/4294967296.0,1,-nbitq), 
to_sfixed(-238842560.0/4294967296.0,1,-nbitq), 
to_sfixed(-104100460.0/4294967296.0,1,-nbitq), 
to_sfixed(-388236854.0/4294967296.0,1,-nbitq), 
to_sfixed(376427544.0/4294967296.0,1,-nbitq), 
to_sfixed(-427738978.0/4294967296.0,1,-nbitq), 
to_sfixed(31567085.0/4294967296.0,1,-nbitq), 
to_sfixed(48301093.0/4294967296.0,1,-nbitq), 
to_sfixed(-83812270.0/4294967296.0,1,-nbitq), 
to_sfixed(409188473.0/4294967296.0,1,-nbitq), 
to_sfixed(360044134.0/4294967296.0,1,-nbitq), 
to_sfixed(-369574824.0/4294967296.0,1,-nbitq), 
to_sfixed(-518093804.0/4294967296.0,1,-nbitq), 
to_sfixed(-183763818.0/4294967296.0,1,-nbitq), 
to_sfixed(50365236.0/4294967296.0,1,-nbitq), 
to_sfixed(208579707.0/4294967296.0,1,-nbitq), 
to_sfixed(240469533.0/4294967296.0,1,-nbitq), 
to_sfixed(-192352799.0/4294967296.0,1,-nbitq), 
to_sfixed(2320757.0/4294967296.0,1,-nbitq), 
to_sfixed(320271267.0/4294967296.0,1,-nbitq), 
to_sfixed(295258564.0/4294967296.0,1,-nbitq), 
to_sfixed(-55960211.0/4294967296.0,1,-nbitq), 
to_sfixed(71422354.0/4294967296.0,1,-nbitq), 
to_sfixed(-127091733.0/4294967296.0,1,-nbitq), 
to_sfixed(413015744.0/4294967296.0,1,-nbitq), 
to_sfixed(-406541390.0/4294967296.0,1,-nbitq), 
to_sfixed(445166920.0/4294967296.0,1,-nbitq), 
to_sfixed(282764350.0/4294967296.0,1,-nbitq), 
to_sfixed(213339749.0/4294967296.0,1,-nbitq), 
to_sfixed(25698944.0/4294967296.0,1,-nbitq), 
to_sfixed(-194612965.0/4294967296.0,1,-nbitq), 
to_sfixed(509874660.0/4294967296.0,1,-nbitq), 
to_sfixed(-274596430.0/4294967296.0,1,-nbitq), 
to_sfixed(323526508.0/4294967296.0,1,-nbitq), 
to_sfixed(-103197600.0/4294967296.0,1,-nbitq), 
to_sfixed(-156138507.0/4294967296.0,1,-nbitq), 
to_sfixed(-329838288.0/4294967296.0,1,-nbitq), 
to_sfixed(173203983.0/4294967296.0,1,-nbitq), 
to_sfixed(2697585.0/4294967296.0,1,-nbitq), 
to_sfixed(320961389.0/4294967296.0,1,-nbitq), 
to_sfixed(-422457476.0/4294967296.0,1,-nbitq), 
to_sfixed(133398761.0/4294967296.0,1,-nbitq), 
to_sfixed(-219582783.0/4294967296.0,1,-nbitq), 
to_sfixed(-270391885.0/4294967296.0,1,-nbitq), 
to_sfixed(395598321.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-207751832.0/4294967296.0,1,-nbitq), 
to_sfixed(133999019.0/4294967296.0,1,-nbitq), 
to_sfixed(353555112.0/4294967296.0,1,-nbitq), 
to_sfixed(-560443.0/4294967296.0,1,-nbitq), 
to_sfixed(-110632834.0/4294967296.0,1,-nbitq), 
to_sfixed(309867418.0/4294967296.0,1,-nbitq), 
to_sfixed(-94637094.0/4294967296.0,1,-nbitq), 
to_sfixed(40544880.0/4294967296.0,1,-nbitq), 
to_sfixed(-170698139.0/4294967296.0,1,-nbitq), 
to_sfixed(-1044094.0/4294967296.0,1,-nbitq), 
to_sfixed(-158929461.0/4294967296.0,1,-nbitq), 
to_sfixed(99174295.0/4294967296.0,1,-nbitq), 
to_sfixed(-182106791.0/4294967296.0,1,-nbitq), 
to_sfixed(318972071.0/4294967296.0,1,-nbitq), 
to_sfixed(313908901.0/4294967296.0,1,-nbitq), 
to_sfixed(-269517626.0/4294967296.0,1,-nbitq), 
to_sfixed(-259519496.0/4294967296.0,1,-nbitq), 
to_sfixed(392760459.0/4294967296.0,1,-nbitq), 
to_sfixed(-203639296.0/4294967296.0,1,-nbitq), 
to_sfixed(-15831734.0/4294967296.0,1,-nbitq), 
to_sfixed(78181783.0/4294967296.0,1,-nbitq), 
to_sfixed(515248171.0/4294967296.0,1,-nbitq), 
to_sfixed(73298855.0/4294967296.0,1,-nbitq), 
to_sfixed(249573613.0/4294967296.0,1,-nbitq), 
to_sfixed(-216200928.0/4294967296.0,1,-nbitq), 
to_sfixed(-126791961.0/4294967296.0,1,-nbitq), 
to_sfixed(-316111838.0/4294967296.0,1,-nbitq), 
to_sfixed(-212325620.0/4294967296.0,1,-nbitq), 
to_sfixed(454720729.0/4294967296.0,1,-nbitq), 
to_sfixed(-177034381.0/4294967296.0,1,-nbitq), 
to_sfixed(140873748.0/4294967296.0,1,-nbitq), 
to_sfixed(-40515428.0/4294967296.0,1,-nbitq), 
to_sfixed(-62608329.0/4294967296.0,1,-nbitq), 
to_sfixed(-515363836.0/4294967296.0,1,-nbitq), 
to_sfixed(54782954.0/4294967296.0,1,-nbitq), 
to_sfixed(384778132.0/4294967296.0,1,-nbitq), 
to_sfixed(-286108498.0/4294967296.0,1,-nbitq), 
to_sfixed(235126274.0/4294967296.0,1,-nbitq), 
to_sfixed(-272781624.0/4294967296.0,1,-nbitq), 
to_sfixed(-63739802.0/4294967296.0,1,-nbitq), 
to_sfixed(-133901019.0/4294967296.0,1,-nbitq), 
to_sfixed(-205805002.0/4294967296.0,1,-nbitq), 
to_sfixed(113258283.0/4294967296.0,1,-nbitq), 
to_sfixed(90742983.0/4294967296.0,1,-nbitq), 
to_sfixed(377832391.0/4294967296.0,1,-nbitq), 
to_sfixed(118085913.0/4294967296.0,1,-nbitq), 
to_sfixed(328829420.0/4294967296.0,1,-nbitq), 
to_sfixed(99982928.0/4294967296.0,1,-nbitq), 
to_sfixed(236154631.0/4294967296.0,1,-nbitq), 
to_sfixed(357540018.0/4294967296.0,1,-nbitq), 
to_sfixed(-259448523.0/4294967296.0,1,-nbitq), 
to_sfixed(-202353678.0/4294967296.0,1,-nbitq), 
to_sfixed(-601750753.0/4294967296.0,1,-nbitq), 
to_sfixed(361889923.0/4294967296.0,1,-nbitq), 
to_sfixed(532193298.0/4294967296.0,1,-nbitq), 
to_sfixed(-343692749.0/4294967296.0,1,-nbitq), 
to_sfixed(28875418.0/4294967296.0,1,-nbitq), 
to_sfixed(66817586.0/4294967296.0,1,-nbitq), 
to_sfixed(270576543.0/4294967296.0,1,-nbitq), 
to_sfixed(-332429601.0/4294967296.0,1,-nbitq), 
to_sfixed(260725394.0/4294967296.0,1,-nbitq), 
to_sfixed(-163615097.0/4294967296.0,1,-nbitq), 
to_sfixed(-371895686.0/4294967296.0,1,-nbitq), 
to_sfixed(-70522032.0/4294967296.0,1,-nbitq), 
to_sfixed(381855951.0/4294967296.0,1,-nbitq), 
to_sfixed(-443523224.0/4294967296.0,1,-nbitq), 
to_sfixed(101367289.0/4294967296.0,1,-nbitq), 
to_sfixed(-72020947.0/4294967296.0,1,-nbitq), 
to_sfixed(-197597007.0/4294967296.0,1,-nbitq), 
to_sfixed(23871973.0/4294967296.0,1,-nbitq), 
to_sfixed(188702705.0/4294967296.0,1,-nbitq), 
to_sfixed(-275458522.0/4294967296.0,1,-nbitq), 
to_sfixed(-81966227.0/4294967296.0,1,-nbitq), 
to_sfixed(-202751247.0/4294967296.0,1,-nbitq), 
to_sfixed(463634619.0/4294967296.0,1,-nbitq), 
to_sfixed(-524274532.0/4294967296.0,1,-nbitq), 
to_sfixed(-393507747.0/4294967296.0,1,-nbitq), 
to_sfixed(-305441552.0/4294967296.0,1,-nbitq), 
to_sfixed(181116974.0/4294967296.0,1,-nbitq), 
to_sfixed(149449295.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(80855962.0/4294967296.0,1,-nbitq), 
to_sfixed(-146563392.0/4294967296.0,1,-nbitq), 
to_sfixed(165914765.0/4294967296.0,1,-nbitq), 
to_sfixed(267408250.0/4294967296.0,1,-nbitq), 
to_sfixed(28817984.0/4294967296.0,1,-nbitq), 
to_sfixed(36147649.0/4294967296.0,1,-nbitq), 
to_sfixed(-182385445.0/4294967296.0,1,-nbitq), 
to_sfixed(54016485.0/4294967296.0,1,-nbitq), 
to_sfixed(176423696.0/4294967296.0,1,-nbitq), 
to_sfixed(-34490363.0/4294967296.0,1,-nbitq), 
to_sfixed(245205719.0/4294967296.0,1,-nbitq), 
to_sfixed(-107587593.0/4294967296.0,1,-nbitq), 
to_sfixed(-327110179.0/4294967296.0,1,-nbitq), 
to_sfixed(431952886.0/4294967296.0,1,-nbitq), 
to_sfixed(-44788271.0/4294967296.0,1,-nbitq), 
to_sfixed(328012531.0/4294967296.0,1,-nbitq), 
to_sfixed(374493963.0/4294967296.0,1,-nbitq), 
to_sfixed(-265879863.0/4294967296.0,1,-nbitq), 
to_sfixed(-154244869.0/4294967296.0,1,-nbitq), 
to_sfixed(-321799261.0/4294967296.0,1,-nbitq), 
to_sfixed(-21284304.0/4294967296.0,1,-nbitq), 
to_sfixed(311858517.0/4294967296.0,1,-nbitq), 
to_sfixed(-97265314.0/4294967296.0,1,-nbitq), 
to_sfixed(305267932.0/4294967296.0,1,-nbitq), 
to_sfixed(413322159.0/4294967296.0,1,-nbitq), 
to_sfixed(242439848.0/4294967296.0,1,-nbitq), 
to_sfixed(188846765.0/4294967296.0,1,-nbitq), 
to_sfixed(101973973.0/4294967296.0,1,-nbitq), 
to_sfixed(225053054.0/4294967296.0,1,-nbitq), 
to_sfixed(345702112.0/4294967296.0,1,-nbitq), 
to_sfixed(-456973988.0/4294967296.0,1,-nbitq), 
to_sfixed(-95552574.0/4294967296.0,1,-nbitq), 
to_sfixed(90813234.0/4294967296.0,1,-nbitq), 
to_sfixed(219116340.0/4294967296.0,1,-nbitq), 
to_sfixed(57712933.0/4294967296.0,1,-nbitq), 
to_sfixed(-180573950.0/4294967296.0,1,-nbitq), 
to_sfixed(439445646.0/4294967296.0,1,-nbitq), 
to_sfixed(174076412.0/4294967296.0,1,-nbitq), 
to_sfixed(-92641925.0/4294967296.0,1,-nbitq), 
to_sfixed(-154202682.0/4294967296.0,1,-nbitq), 
to_sfixed(-209556420.0/4294967296.0,1,-nbitq), 
to_sfixed(-31149706.0/4294967296.0,1,-nbitq), 
to_sfixed(226369469.0/4294967296.0,1,-nbitq), 
to_sfixed(-236997589.0/4294967296.0,1,-nbitq), 
to_sfixed(327875207.0/4294967296.0,1,-nbitq), 
to_sfixed(-27115150.0/4294967296.0,1,-nbitq), 
to_sfixed(-346748908.0/4294967296.0,1,-nbitq), 
to_sfixed(-328153419.0/4294967296.0,1,-nbitq), 
to_sfixed(241255327.0/4294967296.0,1,-nbitq), 
to_sfixed(180105950.0/4294967296.0,1,-nbitq), 
to_sfixed(-147167001.0/4294967296.0,1,-nbitq), 
to_sfixed(-118171436.0/4294967296.0,1,-nbitq), 
to_sfixed(-189690574.0/4294967296.0,1,-nbitq), 
to_sfixed(-286368802.0/4294967296.0,1,-nbitq), 
to_sfixed(190406221.0/4294967296.0,1,-nbitq), 
to_sfixed(-241038496.0/4294967296.0,1,-nbitq), 
to_sfixed(-178927835.0/4294967296.0,1,-nbitq), 
to_sfixed(-208292774.0/4294967296.0,1,-nbitq), 
to_sfixed(-194469039.0/4294967296.0,1,-nbitq), 
to_sfixed(151679838.0/4294967296.0,1,-nbitq), 
to_sfixed(117030302.0/4294967296.0,1,-nbitq), 
to_sfixed(-205978780.0/4294967296.0,1,-nbitq), 
to_sfixed(-152415713.0/4294967296.0,1,-nbitq), 
to_sfixed(348982886.0/4294967296.0,1,-nbitq), 
to_sfixed(306458596.0/4294967296.0,1,-nbitq), 
to_sfixed(-109656237.0/4294967296.0,1,-nbitq), 
to_sfixed(471380361.0/4294967296.0,1,-nbitq), 
to_sfixed(-316534337.0/4294967296.0,1,-nbitq), 
to_sfixed(-325465039.0/4294967296.0,1,-nbitq), 
to_sfixed(-27413724.0/4294967296.0,1,-nbitq), 
to_sfixed(-75665794.0/4294967296.0,1,-nbitq), 
to_sfixed(-91472134.0/4294967296.0,1,-nbitq), 
to_sfixed(-214937870.0/4294967296.0,1,-nbitq), 
to_sfixed(-109085905.0/4294967296.0,1,-nbitq), 
to_sfixed(107572698.0/4294967296.0,1,-nbitq), 
to_sfixed(-488319781.0/4294967296.0,1,-nbitq), 
to_sfixed(-314266763.0/4294967296.0,1,-nbitq), 
to_sfixed(-143861070.0/4294967296.0,1,-nbitq), 
to_sfixed(-135111921.0/4294967296.0,1,-nbitq), 
to_sfixed(68812203.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-237204751.0/4294967296.0,1,-nbitq), 
to_sfixed(187313715.0/4294967296.0,1,-nbitq), 
to_sfixed(-166858611.0/4294967296.0,1,-nbitq), 
to_sfixed(198812195.0/4294967296.0,1,-nbitq), 
to_sfixed(-173671143.0/4294967296.0,1,-nbitq), 
to_sfixed(-345607174.0/4294967296.0,1,-nbitq), 
to_sfixed(136049079.0/4294967296.0,1,-nbitq), 
to_sfixed(-406531777.0/4294967296.0,1,-nbitq), 
to_sfixed(9482560.0/4294967296.0,1,-nbitq), 
to_sfixed(19589993.0/4294967296.0,1,-nbitq), 
to_sfixed(-30379555.0/4294967296.0,1,-nbitq), 
to_sfixed(131929662.0/4294967296.0,1,-nbitq), 
to_sfixed(-375557967.0/4294967296.0,1,-nbitq), 
to_sfixed(335499928.0/4294967296.0,1,-nbitq), 
to_sfixed(196241775.0/4294967296.0,1,-nbitq), 
to_sfixed(162053539.0/4294967296.0,1,-nbitq), 
to_sfixed(-428543163.0/4294967296.0,1,-nbitq), 
to_sfixed(222849223.0/4294967296.0,1,-nbitq), 
to_sfixed(-199467828.0/4294967296.0,1,-nbitq), 
to_sfixed(32884352.0/4294967296.0,1,-nbitq), 
to_sfixed(-241427014.0/4294967296.0,1,-nbitq), 
to_sfixed(-25631372.0/4294967296.0,1,-nbitq), 
to_sfixed(495461493.0/4294967296.0,1,-nbitq), 
to_sfixed(-47195122.0/4294967296.0,1,-nbitq), 
to_sfixed(385080676.0/4294967296.0,1,-nbitq), 
to_sfixed(343998703.0/4294967296.0,1,-nbitq), 
to_sfixed(-203840349.0/4294967296.0,1,-nbitq), 
to_sfixed(57101867.0/4294967296.0,1,-nbitq), 
to_sfixed(329436434.0/4294967296.0,1,-nbitq), 
to_sfixed(-227467817.0/4294967296.0,1,-nbitq), 
to_sfixed(-3435317.0/4294967296.0,1,-nbitq), 
to_sfixed(153896794.0/4294967296.0,1,-nbitq), 
to_sfixed(188811915.0/4294967296.0,1,-nbitq), 
to_sfixed(241046529.0/4294967296.0,1,-nbitq), 
to_sfixed(512381987.0/4294967296.0,1,-nbitq), 
to_sfixed(-47626657.0/4294967296.0,1,-nbitq), 
to_sfixed(456476384.0/4294967296.0,1,-nbitq), 
to_sfixed(342581233.0/4294967296.0,1,-nbitq), 
to_sfixed(155229945.0/4294967296.0,1,-nbitq), 
to_sfixed(370161118.0/4294967296.0,1,-nbitq), 
to_sfixed(-355172480.0/4294967296.0,1,-nbitq), 
to_sfixed(512759145.0/4294967296.0,1,-nbitq), 
to_sfixed(382982840.0/4294967296.0,1,-nbitq), 
to_sfixed(357417799.0/4294967296.0,1,-nbitq), 
to_sfixed(-377728473.0/4294967296.0,1,-nbitq), 
to_sfixed(-217564068.0/4294967296.0,1,-nbitq), 
to_sfixed(20928300.0/4294967296.0,1,-nbitq), 
to_sfixed(-294564994.0/4294967296.0,1,-nbitq), 
to_sfixed(-77478435.0/4294967296.0,1,-nbitq), 
to_sfixed(250868742.0/4294967296.0,1,-nbitq), 
to_sfixed(229183909.0/4294967296.0,1,-nbitq), 
to_sfixed(-116827717.0/4294967296.0,1,-nbitq), 
to_sfixed(63834416.0/4294967296.0,1,-nbitq), 
to_sfixed(339266298.0/4294967296.0,1,-nbitq), 
to_sfixed(296613865.0/4294967296.0,1,-nbitq), 
to_sfixed(-198288676.0/4294967296.0,1,-nbitq), 
to_sfixed(-205298284.0/4294967296.0,1,-nbitq), 
to_sfixed(-252232548.0/4294967296.0,1,-nbitq), 
to_sfixed(40487671.0/4294967296.0,1,-nbitq), 
to_sfixed(253918059.0/4294967296.0,1,-nbitq), 
to_sfixed(-207321936.0/4294967296.0,1,-nbitq), 
to_sfixed(336727376.0/4294967296.0,1,-nbitq), 
to_sfixed(222094262.0/4294967296.0,1,-nbitq), 
to_sfixed(321371271.0/4294967296.0,1,-nbitq), 
to_sfixed(33560382.0/4294967296.0,1,-nbitq), 
to_sfixed(-72147522.0/4294967296.0,1,-nbitq), 
to_sfixed(354116684.0/4294967296.0,1,-nbitq), 
to_sfixed(-453529880.0/4294967296.0,1,-nbitq), 
to_sfixed(91588694.0/4294967296.0,1,-nbitq), 
to_sfixed(11453940.0/4294967296.0,1,-nbitq), 
to_sfixed(-94428350.0/4294967296.0,1,-nbitq), 
to_sfixed(70815770.0/4294967296.0,1,-nbitq), 
to_sfixed(-284350420.0/4294967296.0,1,-nbitq), 
to_sfixed(96492364.0/4294967296.0,1,-nbitq), 
to_sfixed(320155119.0/4294967296.0,1,-nbitq), 
to_sfixed(-485640243.0/4294967296.0,1,-nbitq), 
to_sfixed(-317182896.0/4294967296.0,1,-nbitq), 
to_sfixed(111944755.0/4294967296.0,1,-nbitq), 
to_sfixed(121726897.0/4294967296.0,1,-nbitq), 
to_sfixed(-92108893.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(336199753.0/4294967296.0,1,-nbitq), 
to_sfixed(-134692055.0/4294967296.0,1,-nbitq), 
to_sfixed(-505083563.0/4294967296.0,1,-nbitq), 
to_sfixed(310046803.0/4294967296.0,1,-nbitq), 
to_sfixed(890338812.0/4294967296.0,1,-nbitq), 
to_sfixed(37088653.0/4294967296.0,1,-nbitq), 
to_sfixed(-185382084.0/4294967296.0,1,-nbitq), 
to_sfixed(284851177.0/4294967296.0,1,-nbitq), 
to_sfixed(-160207016.0/4294967296.0,1,-nbitq), 
to_sfixed(213842433.0/4294967296.0,1,-nbitq), 
to_sfixed(302314252.0/4294967296.0,1,-nbitq), 
to_sfixed(446583767.0/4294967296.0,1,-nbitq), 
to_sfixed(101922259.0/4294967296.0,1,-nbitq), 
to_sfixed(-571506278.0/4294967296.0,1,-nbitq), 
to_sfixed(-390814528.0/4294967296.0,1,-nbitq), 
to_sfixed(9320216.0/4294967296.0,1,-nbitq), 
to_sfixed(14986684.0/4294967296.0,1,-nbitq), 
to_sfixed(76902754.0/4294967296.0,1,-nbitq), 
to_sfixed(-651304230.0/4294967296.0,1,-nbitq), 
to_sfixed(-145809242.0/4294967296.0,1,-nbitq), 
to_sfixed(184856938.0/4294967296.0,1,-nbitq), 
to_sfixed(403443298.0/4294967296.0,1,-nbitq), 
to_sfixed(182278575.0/4294967296.0,1,-nbitq), 
to_sfixed(-363271048.0/4294967296.0,1,-nbitq), 
to_sfixed(193521671.0/4294967296.0,1,-nbitq), 
to_sfixed(-198010319.0/4294967296.0,1,-nbitq), 
to_sfixed(-417137144.0/4294967296.0,1,-nbitq), 
to_sfixed(21302585.0/4294967296.0,1,-nbitq), 
to_sfixed(88526022.0/4294967296.0,1,-nbitq), 
to_sfixed(-277512128.0/4294967296.0,1,-nbitq), 
to_sfixed(-1202855.0/4294967296.0,1,-nbitq), 
to_sfixed(-602667034.0/4294967296.0,1,-nbitq), 
to_sfixed(-71554439.0/4294967296.0,1,-nbitq), 
to_sfixed(230794317.0/4294967296.0,1,-nbitq), 
to_sfixed(136547538.0/4294967296.0,1,-nbitq), 
to_sfixed(143151266.0/4294967296.0,1,-nbitq), 
to_sfixed(-10471546.0/4294967296.0,1,-nbitq), 
to_sfixed(104028182.0/4294967296.0,1,-nbitq), 
to_sfixed(136687221.0/4294967296.0,1,-nbitq), 
to_sfixed(-75429863.0/4294967296.0,1,-nbitq), 
to_sfixed(-70870182.0/4294967296.0,1,-nbitq), 
to_sfixed(-235863904.0/4294967296.0,1,-nbitq), 
to_sfixed(203197702.0/4294967296.0,1,-nbitq), 
to_sfixed(289917504.0/4294967296.0,1,-nbitq), 
to_sfixed(-371418023.0/4294967296.0,1,-nbitq), 
to_sfixed(355019866.0/4294967296.0,1,-nbitq), 
to_sfixed(-10164726.0/4294967296.0,1,-nbitq), 
to_sfixed(-35870543.0/4294967296.0,1,-nbitq), 
to_sfixed(285484416.0/4294967296.0,1,-nbitq), 
to_sfixed(380866426.0/4294967296.0,1,-nbitq), 
to_sfixed(-271425490.0/4294967296.0,1,-nbitq), 
to_sfixed(19656442.0/4294967296.0,1,-nbitq), 
to_sfixed(-57752479.0/4294967296.0,1,-nbitq), 
to_sfixed(325339203.0/4294967296.0,1,-nbitq), 
to_sfixed(509232831.0/4294967296.0,1,-nbitq), 
to_sfixed(169716460.0/4294967296.0,1,-nbitq), 
to_sfixed(5696256.0/4294967296.0,1,-nbitq), 
to_sfixed(-147541145.0/4294967296.0,1,-nbitq), 
to_sfixed(-72712741.0/4294967296.0,1,-nbitq), 
to_sfixed(252881817.0/4294967296.0,1,-nbitq), 
to_sfixed(-65454130.0/4294967296.0,1,-nbitq), 
to_sfixed(474719075.0/4294967296.0,1,-nbitq), 
to_sfixed(-452195408.0/4294967296.0,1,-nbitq), 
to_sfixed(149300024.0/4294967296.0,1,-nbitq), 
to_sfixed(-143421173.0/4294967296.0,1,-nbitq), 
to_sfixed(-121335130.0/4294967296.0,1,-nbitq), 
to_sfixed(-55765000.0/4294967296.0,1,-nbitq), 
to_sfixed(99923278.0/4294967296.0,1,-nbitq), 
to_sfixed(-324565811.0/4294967296.0,1,-nbitq), 
to_sfixed(241936395.0/4294967296.0,1,-nbitq), 
to_sfixed(139245216.0/4294967296.0,1,-nbitq), 
to_sfixed(108614419.0/4294967296.0,1,-nbitq), 
to_sfixed(131065086.0/4294967296.0,1,-nbitq), 
to_sfixed(125755168.0/4294967296.0,1,-nbitq), 
to_sfixed(268319027.0/4294967296.0,1,-nbitq), 
to_sfixed(-200936243.0/4294967296.0,1,-nbitq), 
to_sfixed(-164141217.0/4294967296.0,1,-nbitq), 
to_sfixed(-265603078.0/4294967296.0,1,-nbitq), 
to_sfixed(25863947.0/4294967296.0,1,-nbitq), 
to_sfixed(-61084398.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(279508423.0/4294967296.0,1,-nbitq), 
to_sfixed(-718673908.0/4294967296.0,1,-nbitq), 
to_sfixed(-612871738.0/4294967296.0,1,-nbitq), 
to_sfixed(118375824.0/4294967296.0,1,-nbitq), 
to_sfixed(1113011955.0/4294967296.0,1,-nbitq), 
to_sfixed(560960395.0/4294967296.0,1,-nbitq), 
to_sfixed(222775871.0/4294967296.0,1,-nbitq), 
to_sfixed(194705347.0/4294967296.0,1,-nbitq), 
to_sfixed(188897855.0/4294967296.0,1,-nbitq), 
to_sfixed(-47751525.0/4294967296.0,1,-nbitq), 
to_sfixed(-182235682.0/4294967296.0,1,-nbitq), 
to_sfixed(600014945.0/4294967296.0,1,-nbitq), 
to_sfixed(-521557529.0/4294967296.0,1,-nbitq), 
to_sfixed(-545010188.0/4294967296.0,1,-nbitq), 
to_sfixed(-247065795.0/4294967296.0,1,-nbitq), 
to_sfixed(41689758.0/4294967296.0,1,-nbitq), 
to_sfixed(272172346.0/4294967296.0,1,-nbitq), 
to_sfixed(81943303.0/4294967296.0,1,-nbitq), 
to_sfixed(-528797789.0/4294967296.0,1,-nbitq), 
to_sfixed(234495688.0/4294967296.0,1,-nbitq), 
to_sfixed(152327708.0/4294967296.0,1,-nbitq), 
to_sfixed(-251794906.0/4294967296.0,1,-nbitq), 
to_sfixed(-200363696.0/4294967296.0,1,-nbitq), 
to_sfixed(74784365.0/4294967296.0,1,-nbitq), 
to_sfixed(-97483917.0/4294967296.0,1,-nbitq), 
to_sfixed(-239084562.0/4294967296.0,1,-nbitq), 
to_sfixed(376230188.0/4294967296.0,1,-nbitq), 
to_sfixed(100648341.0/4294967296.0,1,-nbitq), 
to_sfixed(-737909013.0/4294967296.0,1,-nbitq), 
to_sfixed(-420076980.0/4294967296.0,1,-nbitq), 
to_sfixed(-342434882.0/4294967296.0,1,-nbitq), 
to_sfixed(-646565143.0/4294967296.0,1,-nbitq), 
to_sfixed(16385160.0/4294967296.0,1,-nbitq), 
to_sfixed(-8279482.0/4294967296.0,1,-nbitq), 
to_sfixed(-143009815.0/4294967296.0,1,-nbitq), 
to_sfixed(-108868822.0/4294967296.0,1,-nbitq), 
to_sfixed(629189825.0/4294967296.0,1,-nbitq), 
to_sfixed(772538934.0/4294967296.0,1,-nbitq), 
to_sfixed(116066102.0/4294967296.0,1,-nbitq), 
to_sfixed(-280401670.0/4294967296.0,1,-nbitq), 
to_sfixed(34598532.0/4294967296.0,1,-nbitq), 
to_sfixed(-323724811.0/4294967296.0,1,-nbitq), 
to_sfixed(-187344036.0/4294967296.0,1,-nbitq), 
to_sfixed(30158827.0/4294967296.0,1,-nbitq), 
to_sfixed(-180807252.0/4294967296.0,1,-nbitq), 
to_sfixed(379572956.0/4294967296.0,1,-nbitq), 
to_sfixed(-332326704.0/4294967296.0,1,-nbitq), 
to_sfixed(71963260.0/4294967296.0,1,-nbitq), 
to_sfixed(-396393876.0/4294967296.0,1,-nbitq), 
to_sfixed(-294325588.0/4294967296.0,1,-nbitq), 
to_sfixed(269841830.0/4294967296.0,1,-nbitq), 
to_sfixed(200941636.0/4294967296.0,1,-nbitq), 
to_sfixed(33595764.0/4294967296.0,1,-nbitq), 
to_sfixed(155445728.0/4294967296.0,1,-nbitq), 
to_sfixed(597232090.0/4294967296.0,1,-nbitq), 
to_sfixed(219689936.0/4294967296.0,1,-nbitq), 
to_sfixed(-212801476.0/4294967296.0,1,-nbitq), 
to_sfixed(-557353222.0/4294967296.0,1,-nbitq), 
to_sfixed(-20320830.0/4294967296.0,1,-nbitq), 
to_sfixed(-354748437.0/4294967296.0,1,-nbitq), 
to_sfixed(234981610.0/4294967296.0,1,-nbitq), 
to_sfixed(100179812.0/4294967296.0,1,-nbitq), 
to_sfixed(166653505.0/4294967296.0,1,-nbitq), 
to_sfixed(301070363.0/4294967296.0,1,-nbitq), 
to_sfixed(-25800606.0/4294967296.0,1,-nbitq), 
to_sfixed(-313944215.0/4294967296.0,1,-nbitq), 
to_sfixed(-427098617.0/4294967296.0,1,-nbitq), 
to_sfixed(-233975178.0/4294967296.0,1,-nbitq), 
to_sfixed(-48669797.0/4294967296.0,1,-nbitq), 
to_sfixed(-94328741.0/4294967296.0,1,-nbitq), 
to_sfixed(54658735.0/4294967296.0,1,-nbitq), 
to_sfixed(261948059.0/4294967296.0,1,-nbitq), 
to_sfixed(210099775.0/4294967296.0,1,-nbitq), 
to_sfixed(120090077.0/4294967296.0,1,-nbitq), 
to_sfixed(349681646.0/4294967296.0,1,-nbitq), 
to_sfixed(493374671.0/4294967296.0,1,-nbitq), 
to_sfixed(217156343.0/4294967296.0,1,-nbitq), 
to_sfixed(-17305159.0/4294967296.0,1,-nbitq), 
to_sfixed(-233715772.0/4294967296.0,1,-nbitq), 
to_sfixed(-178673956.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(75480187.0/4294967296.0,1,-nbitq), 
to_sfixed(-505083827.0/4294967296.0,1,-nbitq), 
to_sfixed(-46946568.0/4294967296.0,1,-nbitq), 
to_sfixed(278102983.0/4294967296.0,1,-nbitq), 
to_sfixed(416260840.0/4294967296.0,1,-nbitq), 
to_sfixed(410691127.0/4294967296.0,1,-nbitq), 
to_sfixed(-105693788.0/4294967296.0,1,-nbitq), 
to_sfixed(56341319.0/4294967296.0,1,-nbitq), 
to_sfixed(319428476.0/4294967296.0,1,-nbitq), 
to_sfixed(-168383414.0/4294967296.0,1,-nbitq), 
to_sfixed(-104152722.0/4294967296.0,1,-nbitq), 
to_sfixed(133816725.0/4294967296.0,1,-nbitq), 
to_sfixed(-96816737.0/4294967296.0,1,-nbitq), 
to_sfixed(-641170516.0/4294967296.0,1,-nbitq), 
to_sfixed(10045388.0/4294967296.0,1,-nbitq), 
to_sfixed(541215808.0/4294967296.0,1,-nbitq), 
to_sfixed(-332518955.0/4294967296.0,1,-nbitq), 
to_sfixed(-156008334.0/4294967296.0,1,-nbitq), 
to_sfixed(-655560257.0/4294967296.0,1,-nbitq), 
to_sfixed(104192841.0/4294967296.0,1,-nbitq), 
to_sfixed(-85140755.0/4294967296.0,1,-nbitq), 
to_sfixed(-346274234.0/4294967296.0,1,-nbitq), 
to_sfixed(-170443503.0/4294967296.0,1,-nbitq), 
to_sfixed(127752096.0/4294967296.0,1,-nbitq), 
to_sfixed(57637397.0/4294967296.0,1,-nbitq), 
to_sfixed(-660263193.0/4294967296.0,1,-nbitq), 
to_sfixed(519345089.0/4294967296.0,1,-nbitq), 
to_sfixed(-93729280.0/4294967296.0,1,-nbitq), 
to_sfixed(-63081471.0/4294967296.0,1,-nbitq), 
to_sfixed(-1179547981.0/4294967296.0,1,-nbitq), 
to_sfixed(351009218.0/4294967296.0,1,-nbitq), 
to_sfixed(-89800533.0/4294967296.0,1,-nbitq), 
to_sfixed(264434128.0/4294967296.0,1,-nbitq), 
to_sfixed(-163119193.0/4294967296.0,1,-nbitq), 
to_sfixed(-324081287.0/4294967296.0,1,-nbitq), 
to_sfixed(-317249830.0/4294967296.0,1,-nbitq), 
to_sfixed(797155445.0/4294967296.0,1,-nbitq), 
to_sfixed(459505807.0/4294967296.0,1,-nbitq), 
to_sfixed(12631980.0/4294967296.0,1,-nbitq), 
to_sfixed(60327325.0/4294967296.0,1,-nbitq), 
to_sfixed(94992448.0/4294967296.0,1,-nbitq), 
to_sfixed(-573969665.0/4294967296.0,1,-nbitq), 
to_sfixed(254974601.0/4294967296.0,1,-nbitq), 
to_sfixed(108317959.0/4294967296.0,1,-nbitq), 
to_sfixed(-89214519.0/4294967296.0,1,-nbitq), 
to_sfixed(-149920567.0/4294967296.0,1,-nbitq), 
to_sfixed(-284698613.0/4294967296.0,1,-nbitq), 
to_sfixed(-39331927.0/4294967296.0,1,-nbitq), 
to_sfixed(-122801880.0/4294967296.0,1,-nbitq), 
to_sfixed(-448861304.0/4294967296.0,1,-nbitq), 
to_sfixed(-311555006.0/4294967296.0,1,-nbitq), 
to_sfixed(892588985.0/4294967296.0,1,-nbitq), 
to_sfixed(143527858.0/4294967296.0,1,-nbitq), 
to_sfixed(400870728.0/4294967296.0,1,-nbitq), 
to_sfixed(-107940805.0/4294967296.0,1,-nbitq), 
to_sfixed(231701096.0/4294967296.0,1,-nbitq), 
to_sfixed(388951792.0/4294967296.0,1,-nbitq), 
to_sfixed(-65165815.0/4294967296.0,1,-nbitq), 
to_sfixed(111564633.0/4294967296.0,1,-nbitq), 
to_sfixed(407971527.0/4294967296.0,1,-nbitq), 
to_sfixed(188803635.0/4294967296.0,1,-nbitq), 
to_sfixed(-562721381.0/4294967296.0,1,-nbitq), 
to_sfixed(713965104.0/4294967296.0,1,-nbitq), 
to_sfixed(296248661.0/4294967296.0,1,-nbitq), 
to_sfixed(300264502.0/4294967296.0,1,-nbitq), 
to_sfixed(262254511.0/4294967296.0,1,-nbitq), 
to_sfixed(-638691802.0/4294967296.0,1,-nbitq), 
to_sfixed(-691264693.0/4294967296.0,1,-nbitq), 
to_sfixed(-275225811.0/4294967296.0,1,-nbitq), 
to_sfixed(209073779.0/4294967296.0,1,-nbitq), 
to_sfixed(-53601858.0/4294967296.0,1,-nbitq), 
to_sfixed(106334255.0/4294967296.0,1,-nbitq), 
to_sfixed(31178635.0/4294967296.0,1,-nbitq), 
to_sfixed(-109361808.0/4294967296.0,1,-nbitq), 
to_sfixed(116185764.0/4294967296.0,1,-nbitq), 
to_sfixed(640777895.0/4294967296.0,1,-nbitq), 
to_sfixed(265878356.0/4294967296.0,1,-nbitq), 
to_sfixed(154577426.0/4294967296.0,1,-nbitq), 
to_sfixed(-463201536.0/4294967296.0,1,-nbitq), 
to_sfixed(186593581.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(381398835.0/4294967296.0,1,-nbitq), 
to_sfixed(-266279813.0/4294967296.0,1,-nbitq), 
to_sfixed(3574165.0/4294967296.0,1,-nbitq), 
to_sfixed(293333806.0/4294967296.0,1,-nbitq), 
to_sfixed(-105534127.0/4294967296.0,1,-nbitq), 
to_sfixed(529244035.0/4294967296.0,1,-nbitq), 
to_sfixed(75560142.0/4294967296.0,1,-nbitq), 
to_sfixed(213181177.0/4294967296.0,1,-nbitq), 
to_sfixed(972567613.0/4294967296.0,1,-nbitq), 
to_sfixed(-364322197.0/4294967296.0,1,-nbitq), 
to_sfixed(46125067.0/4294967296.0,1,-nbitq), 
to_sfixed(-503195885.0/4294967296.0,1,-nbitq), 
to_sfixed(-126875633.0/4294967296.0,1,-nbitq), 
to_sfixed(-462540547.0/4294967296.0,1,-nbitq), 
to_sfixed(194624656.0/4294967296.0,1,-nbitq), 
to_sfixed(102425417.0/4294967296.0,1,-nbitq), 
to_sfixed(2273386.0/4294967296.0,1,-nbitq), 
to_sfixed(-261512770.0/4294967296.0,1,-nbitq), 
to_sfixed(-795732328.0/4294967296.0,1,-nbitq), 
to_sfixed(157586217.0/4294967296.0,1,-nbitq), 
to_sfixed(-136139449.0/4294967296.0,1,-nbitq), 
to_sfixed(-45494127.0/4294967296.0,1,-nbitq), 
to_sfixed(-136357310.0/4294967296.0,1,-nbitq), 
to_sfixed(293799228.0/4294967296.0,1,-nbitq), 
to_sfixed(9618546.0/4294967296.0,1,-nbitq), 
to_sfixed(-844909128.0/4294967296.0,1,-nbitq), 
to_sfixed(406335378.0/4294967296.0,1,-nbitq), 
to_sfixed(248770807.0/4294967296.0,1,-nbitq), 
to_sfixed(-309964307.0/4294967296.0,1,-nbitq), 
to_sfixed(-687130348.0/4294967296.0,1,-nbitq), 
to_sfixed(223607741.0/4294967296.0,1,-nbitq), 
to_sfixed(-567137007.0/4294967296.0,1,-nbitq), 
to_sfixed(774763337.0/4294967296.0,1,-nbitq), 
to_sfixed(508570183.0/4294967296.0,1,-nbitq), 
to_sfixed(-415244350.0/4294967296.0,1,-nbitq), 
to_sfixed(129333147.0/4294967296.0,1,-nbitq), 
to_sfixed(445313802.0/4294967296.0,1,-nbitq), 
to_sfixed(-63892692.0/4294967296.0,1,-nbitq), 
to_sfixed(-332297221.0/4294967296.0,1,-nbitq), 
to_sfixed(402213399.0/4294967296.0,1,-nbitq), 
to_sfixed(826269588.0/4294967296.0,1,-nbitq), 
to_sfixed(-781662821.0/4294967296.0,1,-nbitq), 
to_sfixed(-172418579.0/4294967296.0,1,-nbitq), 
to_sfixed(-129080668.0/4294967296.0,1,-nbitq), 
to_sfixed(481434451.0/4294967296.0,1,-nbitq), 
to_sfixed(102652201.0/4294967296.0,1,-nbitq), 
to_sfixed(-38249946.0/4294967296.0,1,-nbitq), 
to_sfixed(504952799.0/4294967296.0,1,-nbitq), 
to_sfixed(-164100432.0/4294967296.0,1,-nbitq), 
to_sfixed(-111975874.0/4294967296.0,1,-nbitq), 
to_sfixed(-393788977.0/4294967296.0,1,-nbitq), 
to_sfixed(808313680.0/4294967296.0,1,-nbitq), 
to_sfixed(181508195.0/4294967296.0,1,-nbitq), 
to_sfixed(-444831771.0/4294967296.0,1,-nbitq), 
to_sfixed(-597971721.0/4294967296.0,1,-nbitq), 
to_sfixed(1134297605.0/4294967296.0,1,-nbitq), 
to_sfixed(-125107833.0/4294967296.0,1,-nbitq), 
to_sfixed(44967089.0/4294967296.0,1,-nbitq), 
to_sfixed(81433412.0/4294967296.0,1,-nbitq), 
to_sfixed(188747.0/4294967296.0,1,-nbitq), 
to_sfixed(262220655.0/4294967296.0,1,-nbitq), 
to_sfixed(-776115467.0/4294967296.0,1,-nbitq), 
to_sfixed(-214509786.0/4294967296.0,1,-nbitq), 
to_sfixed(-53017537.0/4294967296.0,1,-nbitq), 
to_sfixed(-162354247.0/4294967296.0,1,-nbitq), 
to_sfixed(240194479.0/4294967296.0,1,-nbitq), 
to_sfixed(-1667960188.0/4294967296.0,1,-nbitq), 
to_sfixed(-881222092.0/4294967296.0,1,-nbitq), 
to_sfixed(-17473671.0/4294967296.0,1,-nbitq), 
to_sfixed(181758929.0/4294967296.0,1,-nbitq), 
to_sfixed(-751751011.0/4294967296.0,1,-nbitq), 
to_sfixed(-11489874.0/4294967296.0,1,-nbitq), 
to_sfixed(401995174.0/4294967296.0,1,-nbitq), 
to_sfixed(-306406572.0/4294967296.0,1,-nbitq), 
to_sfixed(98908989.0/4294967296.0,1,-nbitq), 
to_sfixed(351983892.0/4294967296.0,1,-nbitq), 
to_sfixed(-43468569.0/4294967296.0,1,-nbitq), 
to_sfixed(356293094.0/4294967296.0,1,-nbitq), 
to_sfixed(-1072562454.0/4294967296.0,1,-nbitq), 
to_sfixed(-325795798.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(275148201.0/4294967296.0,1,-nbitq), 
to_sfixed(-579790557.0/4294967296.0,1,-nbitq), 
to_sfixed(380680377.0/4294967296.0,1,-nbitq), 
to_sfixed(428842237.0/4294967296.0,1,-nbitq), 
to_sfixed(155180040.0/4294967296.0,1,-nbitq), 
to_sfixed(150504538.0/4294967296.0,1,-nbitq), 
to_sfixed(-226959988.0/4294967296.0,1,-nbitq), 
to_sfixed(487952377.0/4294967296.0,1,-nbitq), 
to_sfixed(877863260.0/4294967296.0,1,-nbitq), 
to_sfixed(-23252412.0/4294967296.0,1,-nbitq), 
to_sfixed(-580325238.0/4294967296.0,1,-nbitq), 
to_sfixed(196882611.0/4294967296.0,1,-nbitq), 
to_sfixed(223112844.0/4294967296.0,1,-nbitq), 
to_sfixed(-408458217.0/4294967296.0,1,-nbitq), 
to_sfixed(-281806901.0/4294967296.0,1,-nbitq), 
to_sfixed(391560250.0/4294967296.0,1,-nbitq), 
to_sfixed(243725430.0/4294967296.0,1,-nbitq), 
to_sfixed(346011326.0/4294967296.0,1,-nbitq), 
to_sfixed(-595435560.0/4294967296.0,1,-nbitq), 
to_sfixed(213338026.0/4294967296.0,1,-nbitq), 
to_sfixed(-98816422.0/4294967296.0,1,-nbitq), 
to_sfixed(291311994.0/4294967296.0,1,-nbitq), 
to_sfixed(235816391.0/4294967296.0,1,-nbitq), 
to_sfixed(234657248.0/4294967296.0,1,-nbitq), 
to_sfixed(-252679354.0/4294967296.0,1,-nbitq), 
to_sfixed(-320388332.0/4294967296.0,1,-nbitq), 
to_sfixed(238560261.0/4294967296.0,1,-nbitq), 
to_sfixed(1518266.0/4294967296.0,1,-nbitq), 
to_sfixed(218891604.0/4294967296.0,1,-nbitq), 
to_sfixed(-1068520202.0/4294967296.0,1,-nbitq), 
to_sfixed(546956981.0/4294967296.0,1,-nbitq), 
to_sfixed(150036514.0/4294967296.0,1,-nbitq), 
to_sfixed(422099619.0/4294967296.0,1,-nbitq), 
to_sfixed(530901004.0/4294967296.0,1,-nbitq), 
to_sfixed(-915285693.0/4294967296.0,1,-nbitq), 
to_sfixed(-517995887.0/4294967296.0,1,-nbitq), 
to_sfixed(437642113.0/4294967296.0,1,-nbitq), 
to_sfixed(-249374675.0/4294967296.0,1,-nbitq), 
to_sfixed(284218243.0/4294967296.0,1,-nbitq), 
to_sfixed(247696102.0/4294967296.0,1,-nbitq), 
to_sfixed(321462407.0/4294967296.0,1,-nbitq), 
to_sfixed(-708688796.0/4294967296.0,1,-nbitq), 
to_sfixed(129261041.0/4294967296.0,1,-nbitq), 
to_sfixed(-406667718.0/4294967296.0,1,-nbitq), 
to_sfixed(-408556930.0/4294967296.0,1,-nbitq), 
to_sfixed(-433539452.0/4294967296.0,1,-nbitq), 
to_sfixed(325788788.0/4294967296.0,1,-nbitq), 
to_sfixed(136181898.0/4294967296.0,1,-nbitq), 
to_sfixed(-187718310.0/4294967296.0,1,-nbitq), 
to_sfixed(-298744403.0/4294967296.0,1,-nbitq), 
to_sfixed(-669739000.0/4294967296.0,1,-nbitq), 
to_sfixed(1247181457.0/4294967296.0,1,-nbitq), 
to_sfixed(336644879.0/4294967296.0,1,-nbitq), 
to_sfixed(-235588315.0/4294967296.0,1,-nbitq), 
to_sfixed(-605384806.0/4294967296.0,1,-nbitq), 
to_sfixed(419052549.0/4294967296.0,1,-nbitq), 
to_sfixed(-486063577.0/4294967296.0,1,-nbitq), 
to_sfixed(272154838.0/4294967296.0,1,-nbitq), 
to_sfixed(99942790.0/4294967296.0,1,-nbitq), 
to_sfixed(-276798693.0/4294967296.0,1,-nbitq), 
to_sfixed(-309205595.0/4294967296.0,1,-nbitq), 
to_sfixed(-249091189.0/4294967296.0,1,-nbitq), 
to_sfixed(218880408.0/4294967296.0,1,-nbitq), 
to_sfixed(-81039152.0/4294967296.0,1,-nbitq), 
to_sfixed(-580575296.0/4294967296.0,1,-nbitq), 
to_sfixed(47909911.0/4294967296.0,1,-nbitq), 
to_sfixed(-1226491141.0/4294967296.0,1,-nbitq), 
to_sfixed(-413830759.0/4294967296.0,1,-nbitq), 
to_sfixed(-115442591.0/4294967296.0,1,-nbitq), 
to_sfixed(557039575.0/4294967296.0,1,-nbitq), 
to_sfixed(-480964535.0/4294967296.0,1,-nbitq), 
to_sfixed(-50614127.0/4294967296.0,1,-nbitq), 
to_sfixed(264336039.0/4294967296.0,1,-nbitq), 
to_sfixed(-232380063.0/4294967296.0,1,-nbitq), 
to_sfixed(384858444.0/4294967296.0,1,-nbitq), 
to_sfixed(-74088237.0/4294967296.0,1,-nbitq), 
to_sfixed(45194685.0/4294967296.0,1,-nbitq), 
to_sfixed(-481942850.0/4294967296.0,1,-nbitq), 
to_sfixed(-630970410.0/4294967296.0,1,-nbitq), 
to_sfixed(-356064624.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-82953614.0/4294967296.0,1,-nbitq), 
to_sfixed(-207097696.0/4294967296.0,1,-nbitq), 
to_sfixed(280885353.0/4294967296.0,1,-nbitq), 
to_sfixed(225302100.0/4294967296.0,1,-nbitq), 
to_sfixed(-53453939.0/4294967296.0,1,-nbitq), 
to_sfixed(177191942.0/4294967296.0,1,-nbitq), 
to_sfixed(-120984465.0/4294967296.0,1,-nbitq), 
to_sfixed(304742550.0/4294967296.0,1,-nbitq), 
to_sfixed(1108904976.0/4294967296.0,1,-nbitq), 
to_sfixed(158313320.0/4294967296.0,1,-nbitq), 
to_sfixed(-815805786.0/4294967296.0,1,-nbitq), 
to_sfixed(732850484.0/4294967296.0,1,-nbitq), 
to_sfixed(-192247514.0/4294967296.0,1,-nbitq), 
to_sfixed(-135203012.0/4294967296.0,1,-nbitq), 
to_sfixed(-191912163.0/4294967296.0,1,-nbitq), 
to_sfixed(86784894.0/4294967296.0,1,-nbitq), 
to_sfixed(53337585.0/4294967296.0,1,-nbitq), 
to_sfixed(414855180.0/4294967296.0,1,-nbitq), 
to_sfixed(-206056899.0/4294967296.0,1,-nbitq), 
to_sfixed(-160516529.0/4294967296.0,1,-nbitq), 
to_sfixed(-395569434.0/4294967296.0,1,-nbitq), 
to_sfixed(-144073155.0/4294967296.0,1,-nbitq), 
to_sfixed(642274703.0/4294967296.0,1,-nbitq), 
to_sfixed(796221188.0/4294967296.0,1,-nbitq), 
to_sfixed(-249368574.0/4294967296.0,1,-nbitq), 
to_sfixed(478613803.0/4294967296.0,1,-nbitq), 
to_sfixed(-495545626.0/4294967296.0,1,-nbitq), 
to_sfixed(-209729219.0/4294967296.0,1,-nbitq), 
to_sfixed(57340141.0/4294967296.0,1,-nbitq), 
to_sfixed(-835104909.0/4294967296.0,1,-nbitq), 
to_sfixed(573465041.0/4294967296.0,1,-nbitq), 
to_sfixed(-141205314.0/4294967296.0,1,-nbitq), 
to_sfixed(519484923.0/4294967296.0,1,-nbitq), 
to_sfixed(202438220.0/4294967296.0,1,-nbitq), 
to_sfixed(-1115126281.0/4294967296.0,1,-nbitq), 
to_sfixed(-714361181.0/4294967296.0,1,-nbitq), 
to_sfixed(940736300.0/4294967296.0,1,-nbitq), 
to_sfixed(-184441234.0/4294967296.0,1,-nbitq), 
to_sfixed(-59911432.0/4294967296.0,1,-nbitq), 
to_sfixed(-342477609.0/4294967296.0,1,-nbitq), 
to_sfixed(483032047.0/4294967296.0,1,-nbitq), 
to_sfixed(-515813798.0/4294967296.0,1,-nbitq), 
to_sfixed(-4281926.0/4294967296.0,1,-nbitq), 
to_sfixed(-81792609.0/4294967296.0,1,-nbitq), 
to_sfixed(-150412281.0/4294967296.0,1,-nbitq), 
to_sfixed(-556110974.0/4294967296.0,1,-nbitq), 
to_sfixed(106587122.0/4294967296.0,1,-nbitq), 
to_sfixed(565656654.0/4294967296.0,1,-nbitq), 
to_sfixed(-20314870.0/4294967296.0,1,-nbitq), 
to_sfixed(-605476122.0/4294967296.0,1,-nbitq), 
to_sfixed(-383292010.0/4294967296.0,1,-nbitq), 
to_sfixed(894600196.0/4294967296.0,1,-nbitq), 
to_sfixed(-710128295.0/4294967296.0,1,-nbitq), 
to_sfixed(146990547.0/4294967296.0,1,-nbitq), 
to_sfixed(-217883222.0/4294967296.0,1,-nbitq), 
to_sfixed(979030883.0/4294967296.0,1,-nbitq), 
to_sfixed(-388259957.0/4294967296.0,1,-nbitq), 
to_sfixed(472182604.0/4294967296.0,1,-nbitq), 
to_sfixed(173608138.0/4294967296.0,1,-nbitq), 
to_sfixed(309492076.0/4294967296.0,1,-nbitq), 
to_sfixed(-209942906.0/4294967296.0,1,-nbitq), 
to_sfixed(-933891700.0/4294967296.0,1,-nbitq), 
to_sfixed(-439098293.0/4294967296.0,1,-nbitq), 
to_sfixed(-608572231.0/4294967296.0,1,-nbitq), 
to_sfixed(-15100301.0/4294967296.0,1,-nbitq), 
to_sfixed(-102117349.0/4294967296.0,1,-nbitq), 
to_sfixed(-1064659497.0/4294967296.0,1,-nbitq), 
to_sfixed(-545528997.0/4294967296.0,1,-nbitq), 
to_sfixed(178158692.0/4294967296.0,1,-nbitq), 
to_sfixed(466535029.0/4294967296.0,1,-nbitq), 
to_sfixed(-748185592.0/4294967296.0,1,-nbitq), 
to_sfixed(575912681.0/4294967296.0,1,-nbitq), 
to_sfixed(695453575.0/4294967296.0,1,-nbitq), 
to_sfixed(-273687098.0/4294967296.0,1,-nbitq), 
to_sfixed(26613911.0/4294967296.0,1,-nbitq), 
to_sfixed(-490221540.0/4294967296.0,1,-nbitq), 
to_sfixed(359383885.0/4294967296.0,1,-nbitq), 
to_sfixed(-688279178.0/4294967296.0,1,-nbitq), 
to_sfixed(137923284.0/4294967296.0,1,-nbitq), 
to_sfixed(-84580947.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(368360097.0/4294967296.0,1,-nbitq), 
to_sfixed(-151731785.0/4294967296.0,1,-nbitq), 
to_sfixed(-468190016.0/4294967296.0,1,-nbitq), 
to_sfixed(530570506.0/4294967296.0,1,-nbitq), 
to_sfixed(-234309004.0/4294967296.0,1,-nbitq), 
to_sfixed(-260481481.0/4294967296.0,1,-nbitq), 
to_sfixed(41067932.0/4294967296.0,1,-nbitq), 
to_sfixed(997535587.0/4294967296.0,1,-nbitq), 
to_sfixed(1041351881.0/4294967296.0,1,-nbitq), 
to_sfixed(317276007.0/4294967296.0,1,-nbitq), 
to_sfixed(-1175631757.0/4294967296.0,1,-nbitq), 
to_sfixed(626534651.0/4294967296.0,1,-nbitq), 
to_sfixed(-282562824.0/4294967296.0,1,-nbitq), 
to_sfixed(-165028891.0/4294967296.0,1,-nbitq), 
to_sfixed(481438372.0/4294967296.0,1,-nbitq), 
to_sfixed(-282628047.0/4294967296.0,1,-nbitq), 
to_sfixed(-431141670.0/4294967296.0,1,-nbitq), 
to_sfixed(-128701359.0/4294967296.0,1,-nbitq), 
to_sfixed(-78608934.0/4294967296.0,1,-nbitq), 
to_sfixed(-126297420.0/4294967296.0,1,-nbitq), 
to_sfixed(174456297.0/4294967296.0,1,-nbitq), 
to_sfixed(-513930140.0/4294967296.0,1,-nbitq), 
to_sfixed(742404148.0/4294967296.0,1,-nbitq), 
to_sfixed(594317450.0/4294967296.0,1,-nbitq), 
to_sfixed(129643963.0/4294967296.0,1,-nbitq), 
to_sfixed(-527909272.0/4294967296.0,1,-nbitq), 
to_sfixed(-734716780.0/4294967296.0,1,-nbitq), 
to_sfixed(126246285.0/4294967296.0,1,-nbitq), 
to_sfixed(230691277.0/4294967296.0,1,-nbitq), 
to_sfixed(-655751238.0/4294967296.0,1,-nbitq), 
to_sfixed(797740180.0/4294967296.0,1,-nbitq), 
to_sfixed(493487943.0/4294967296.0,1,-nbitq), 
to_sfixed(256451531.0/4294967296.0,1,-nbitq), 
to_sfixed(-491464558.0/4294967296.0,1,-nbitq), 
to_sfixed(-955455206.0/4294967296.0,1,-nbitq), 
to_sfixed(-1642475131.0/4294967296.0,1,-nbitq), 
to_sfixed(661227118.0/4294967296.0,1,-nbitq), 
to_sfixed(-549641784.0/4294967296.0,1,-nbitq), 
to_sfixed(-64608814.0/4294967296.0,1,-nbitq), 
to_sfixed(191969214.0/4294967296.0,1,-nbitq), 
to_sfixed(343429394.0/4294967296.0,1,-nbitq), 
to_sfixed(-578910331.0/4294967296.0,1,-nbitq), 
to_sfixed(-336388268.0/4294967296.0,1,-nbitq), 
to_sfixed(621433801.0/4294967296.0,1,-nbitq), 
to_sfixed(-185384203.0/4294967296.0,1,-nbitq), 
to_sfixed(-960506081.0/4294967296.0,1,-nbitq), 
to_sfixed(290184492.0/4294967296.0,1,-nbitq), 
to_sfixed(135473674.0/4294967296.0,1,-nbitq), 
to_sfixed(-551900370.0/4294967296.0,1,-nbitq), 
to_sfixed(-864237888.0/4294967296.0,1,-nbitq), 
to_sfixed(6793895.0/4294967296.0,1,-nbitq), 
to_sfixed(1010347678.0/4294967296.0,1,-nbitq), 
to_sfixed(-549352654.0/4294967296.0,1,-nbitq), 
to_sfixed(634483272.0/4294967296.0,1,-nbitq), 
to_sfixed(-444300435.0/4294967296.0,1,-nbitq), 
to_sfixed(868797252.0/4294967296.0,1,-nbitq), 
to_sfixed(-465292375.0/4294967296.0,1,-nbitq), 
to_sfixed(223005544.0/4294967296.0,1,-nbitq), 
to_sfixed(-368182490.0/4294967296.0,1,-nbitq), 
to_sfixed(241617462.0/4294967296.0,1,-nbitq), 
to_sfixed(272875492.0/4294967296.0,1,-nbitq), 
to_sfixed(-604638335.0/4294967296.0,1,-nbitq), 
to_sfixed(-606236311.0/4294967296.0,1,-nbitq), 
to_sfixed(-625793754.0/4294967296.0,1,-nbitq), 
to_sfixed(-219110864.0/4294967296.0,1,-nbitq), 
to_sfixed(359155857.0/4294967296.0,1,-nbitq), 
to_sfixed(-200708783.0/4294967296.0,1,-nbitq), 
to_sfixed(-398279819.0/4294967296.0,1,-nbitq), 
to_sfixed(224852687.0/4294967296.0,1,-nbitq), 
to_sfixed(174870821.0/4294967296.0,1,-nbitq), 
to_sfixed(-1524954584.0/4294967296.0,1,-nbitq), 
to_sfixed(637337581.0/4294967296.0,1,-nbitq), 
to_sfixed(682811793.0/4294967296.0,1,-nbitq), 
to_sfixed(167465913.0/4294967296.0,1,-nbitq), 
to_sfixed(-30785647.0/4294967296.0,1,-nbitq), 
to_sfixed(-811540653.0/4294967296.0,1,-nbitq), 
to_sfixed(-123102115.0/4294967296.0,1,-nbitq), 
to_sfixed(-552254275.0/4294967296.0,1,-nbitq), 
to_sfixed(101131448.0/4294967296.0,1,-nbitq), 
to_sfixed(185828050.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(384139767.0/4294967296.0,1,-nbitq), 
to_sfixed(-480789344.0/4294967296.0,1,-nbitq), 
to_sfixed(-113049351.0/4294967296.0,1,-nbitq), 
to_sfixed(933038369.0/4294967296.0,1,-nbitq), 
to_sfixed(-947438049.0/4294967296.0,1,-nbitq), 
to_sfixed(-636169597.0/4294967296.0,1,-nbitq), 
to_sfixed(94856993.0/4294967296.0,1,-nbitq), 
to_sfixed(269471965.0/4294967296.0,1,-nbitq), 
to_sfixed(720937414.0/4294967296.0,1,-nbitq), 
to_sfixed(170946017.0/4294967296.0,1,-nbitq), 
to_sfixed(-294082761.0/4294967296.0,1,-nbitq), 
to_sfixed(538442035.0/4294967296.0,1,-nbitq), 
to_sfixed(-20205905.0/4294967296.0,1,-nbitq), 
to_sfixed(-398994242.0/4294967296.0,1,-nbitq), 
to_sfixed(-108943362.0/4294967296.0,1,-nbitq), 
to_sfixed(-318938199.0/4294967296.0,1,-nbitq), 
to_sfixed(-303570696.0/4294967296.0,1,-nbitq), 
to_sfixed(46589262.0/4294967296.0,1,-nbitq), 
to_sfixed(-609906452.0/4294967296.0,1,-nbitq), 
to_sfixed(-543232585.0/4294967296.0,1,-nbitq), 
to_sfixed(171378089.0/4294967296.0,1,-nbitq), 
to_sfixed(-71018595.0/4294967296.0,1,-nbitq), 
to_sfixed(150735467.0/4294967296.0,1,-nbitq), 
to_sfixed(56200754.0/4294967296.0,1,-nbitq), 
to_sfixed(-161811969.0/4294967296.0,1,-nbitq), 
to_sfixed(-898309117.0/4294967296.0,1,-nbitq), 
to_sfixed(-172623745.0/4294967296.0,1,-nbitq), 
to_sfixed(253086517.0/4294967296.0,1,-nbitq), 
to_sfixed(-212502471.0/4294967296.0,1,-nbitq), 
to_sfixed(-1347268388.0/4294967296.0,1,-nbitq), 
to_sfixed(1048467564.0/4294967296.0,1,-nbitq), 
to_sfixed(-996988.0/4294967296.0,1,-nbitq), 
to_sfixed(519297739.0/4294967296.0,1,-nbitq), 
to_sfixed(-1200779903.0/4294967296.0,1,-nbitq), 
to_sfixed(-772242546.0/4294967296.0,1,-nbitq), 
to_sfixed(-1416766738.0/4294967296.0,1,-nbitq), 
to_sfixed(247574663.0/4294967296.0,1,-nbitq), 
to_sfixed(-490947077.0/4294967296.0,1,-nbitq), 
to_sfixed(-20913866.0/4294967296.0,1,-nbitq), 
to_sfixed(100192455.0/4294967296.0,1,-nbitq), 
to_sfixed(387434547.0/4294967296.0,1,-nbitq), 
to_sfixed(-615236424.0/4294967296.0,1,-nbitq), 
to_sfixed(665810216.0/4294967296.0,1,-nbitq), 
to_sfixed(845523823.0/4294967296.0,1,-nbitq), 
to_sfixed(-227669014.0/4294967296.0,1,-nbitq), 
to_sfixed(-212884417.0/4294967296.0,1,-nbitq), 
to_sfixed(-442112274.0/4294967296.0,1,-nbitq), 
to_sfixed(143025697.0/4294967296.0,1,-nbitq), 
to_sfixed(-302142172.0/4294967296.0,1,-nbitq), 
to_sfixed(-525039241.0/4294967296.0,1,-nbitq), 
to_sfixed(-252706003.0/4294967296.0,1,-nbitq), 
to_sfixed(539610520.0/4294967296.0,1,-nbitq), 
to_sfixed(-1317727356.0/4294967296.0,1,-nbitq), 
to_sfixed(404470150.0/4294967296.0,1,-nbitq), 
to_sfixed(-1263493836.0/4294967296.0,1,-nbitq), 
to_sfixed(614531128.0/4294967296.0,1,-nbitq), 
to_sfixed(-366340054.0/4294967296.0,1,-nbitq), 
to_sfixed(38636247.0/4294967296.0,1,-nbitq), 
to_sfixed(4267834.0/4294967296.0,1,-nbitq), 
to_sfixed(167342857.0/4294967296.0,1,-nbitq), 
to_sfixed(271279228.0/4294967296.0,1,-nbitq), 
to_sfixed(-1053931550.0/4294967296.0,1,-nbitq), 
to_sfixed(-874309082.0/4294967296.0,1,-nbitq), 
to_sfixed(-534484470.0/4294967296.0,1,-nbitq), 
to_sfixed(40272380.0/4294967296.0,1,-nbitq), 
to_sfixed(16036359.0/4294967296.0,1,-nbitq), 
to_sfixed(987045178.0/4294967296.0,1,-nbitq), 
to_sfixed(-842334392.0/4294967296.0,1,-nbitq), 
to_sfixed(-173571884.0/4294967296.0,1,-nbitq), 
to_sfixed(19633901.0/4294967296.0,1,-nbitq), 
to_sfixed(-2471646923.0/4294967296.0,1,-nbitq), 
to_sfixed(-124958489.0/4294967296.0,1,-nbitq), 
to_sfixed(1252243240.0/4294967296.0,1,-nbitq), 
to_sfixed(22583639.0/4294967296.0,1,-nbitq), 
to_sfixed(332811572.0/4294967296.0,1,-nbitq), 
to_sfixed(328374436.0/4294967296.0,1,-nbitq), 
to_sfixed(-685689793.0/4294967296.0,1,-nbitq), 
to_sfixed(-118931592.0/4294967296.0,1,-nbitq), 
to_sfixed(290243865.0/4294967296.0,1,-nbitq), 
to_sfixed(-256770986.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(282496701.0/4294967296.0,1,-nbitq), 
to_sfixed(-1383922454.0/4294967296.0,1,-nbitq), 
to_sfixed(-797822662.0/4294967296.0,1,-nbitq), 
to_sfixed(1362325183.0/4294967296.0,1,-nbitq), 
to_sfixed(-1299052976.0/4294967296.0,1,-nbitq), 
to_sfixed(-511229248.0/4294967296.0,1,-nbitq), 
to_sfixed(386207624.0/4294967296.0,1,-nbitq), 
to_sfixed(-704784100.0/4294967296.0,1,-nbitq), 
to_sfixed(685721697.0/4294967296.0,1,-nbitq), 
to_sfixed(388136743.0/4294967296.0,1,-nbitq), 
to_sfixed(-876475120.0/4294967296.0,1,-nbitq), 
to_sfixed(488226647.0/4294967296.0,1,-nbitq), 
to_sfixed(140310547.0/4294967296.0,1,-nbitq), 
to_sfixed(-803507658.0/4294967296.0,1,-nbitq), 
to_sfixed(239842796.0/4294967296.0,1,-nbitq), 
to_sfixed(-472355571.0/4294967296.0,1,-nbitq), 
to_sfixed(67978942.0/4294967296.0,1,-nbitq), 
to_sfixed(65869704.0/4294967296.0,1,-nbitq), 
to_sfixed(60196931.0/4294967296.0,1,-nbitq), 
to_sfixed(-679877408.0/4294967296.0,1,-nbitq), 
to_sfixed(196151785.0/4294967296.0,1,-nbitq), 
to_sfixed(168614618.0/4294967296.0,1,-nbitq), 
to_sfixed(490734263.0/4294967296.0,1,-nbitq), 
to_sfixed(480735552.0/4294967296.0,1,-nbitq), 
to_sfixed(-364007565.0/4294967296.0,1,-nbitq), 
to_sfixed(694587409.0/4294967296.0,1,-nbitq), 
to_sfixed(-281424067.0/4294967296.0,1,-nbitq), 
to_sfixed(-400683721.0/4294967296.0,1,-nbitq), 
to_sfixed(-117964663.0/4294967296.0,1,-nbitq), 
to_sfixed(-477823958.0/4294967296.0,1,-nbitq), 
to_sfixed(941757363.0/4294967296.0,1,-nbitq), 
to_sfixed(-59220255.0/4294967296.0,1,-nbitq), 
to_sfixed(726936369.0/4294967296.0,1,-nbitq), 
to_sfixed(-671975119.0/4294967296.0,1,-nbitq), 
to_sfixed(98891756.0/4294967296.0,1,-nbitq), 
to_sfixed(741506020.0/4294967296.0,1,-nbitq), 
to_sfixed(1108576923.0/4294967296.0,1,-nbitq), 
to_sfixed(-630771409.0/4294967296.0,1,-nbitq), 
to_sfixed(-270833405.0/4294967296.0,1,-nbitq), 
to_sfixed(317682771.0/4294967296.0,1,-nbitq), 
to_sfixed(163082288.0/4294967296.0,1,-nbitq), 
to_sfixed(187743105.0/4294967296.0,1,-nbitq), 
to_sfixed(1846709785.0/4294967296.0,1,-nbitq), 
to_sfixed(420209969.0/4294967296.0,1,-nbitq), 
to_sfixed(-279147795.0/4294967296.0,1,-nbitq), 
to_sfixed(-318553243.0/4294967296.0,1,-nbitq), 
to_sfixed(321841712.0/4294967296.0,1,-nbitq), 
to_sfixed(204096282.0/4294967296.0,1,-nbitq), 
to_sfixed(-312078890.0/4294967296.0,1,-nbitq), 
to_sfixed(-269814961.0/4294967296.0,1,-nbitq), 
to_sfixed(-447199494.0/4294967296.0,1,-nbitq), 
to_sfixed(739121999.0/4294967296.0,1,-nbitq), 
to_sfixed(-856137660.0/4294967296.0,1,-nbitq), 
to_sfixed(-82222458.0/4294967296.0,1,-nbitq), 
to_sfixed(494818259.0/4294967296.0,1,-nbitq), 
to_sfixed(-572323390.0/4294967296.0,1,-nbitq), 
to_sfixed(-546402145.0/4294967296.0,1,-nbitq), 
to_sfixed(-94789247.0/4294967296.0,1,-nbitq), 
to_sfixed(-71810704.0/4294967296.0,1,-nbitq), 
to_sfixed(-206371959.0/4294967296.0,1,-nbitq), 
to_sfixed(160488604.0/4294967296.0,1,-nbitq), 
to_sfixed(-395304419.0/4294967296.0,1,-nbitq), 
to_sfixed(-1212235473.0/4294967296.0,1,-nbitq), 
to_sfixed(259246119.0/4294967296.0,1,-nbitq), 
to_sfixed(373612175.0/4294967296.0,1,-nbitq), 
to_sfixed(-128546111.0/4294967296.0,1,-nbitq), 
to_sfixed(1050659061.0/4294967296.0,1,-nbitq), 
to_sfixed(371889546.0/4294967296.0,1,-nbitq), 
to_sfixed(-38138326.0/4294967296.0,1,-nbitq), 
to_sfixed(18837260.0/4294967296.0,1,-nbitq), 
to_sfixed(-1571371749.0/4294967296.0,1,-nbitq), 
to_sfixed(29333606.0/4294967296.0,1,-nbitq), 
to_sfixed(679731078.0/4294967296.0,1,-nbitq), 
to_sfixed(-118817994.0/4294967296.0,1,-nbitq), 
to_sfixed(251512540.0/4294967296.0,1,-nbitq), 
to_sfixed(489163716.0/4294967296.0,1,-nbitq), 
to_sfixed(-337573689.0/4294967296.0,1,-nbitq), 
to_sfixed(-198251716.0/4294967296.0,1,-nbitq), 
to_sfixed(-119573822.0/4294967296.0,1,-nbitq), 
to_sfixed(-275092296.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-204264735.0/4294967296.0,1,-nbitq), 
to_sfixed(-588669416.0/4294967296.0,1,-nbitq), 
to_sfixed(-1102992030.0/4294967296.0,1,-nbitq), 
to_sfixed(790242034.0/4294967296.0,1,-nbitq), 
to_sfixed(-1356256578.0/4294967296.0,1,-nbitq), 
to_sfixed(-1028545209.0/4294967296.0,1,-nbitq), 
to_sfixed(572812979.0/4294967296.0,1,-nbitq), 
to_sfixed(-934344487.0/4294967296.0,1,-nbitq), 
to_sfixed(-13586702.0/4294967296.0,1,-nbitq), 
to_sfixed(213885150.0/4294967296.0,1,-nbitq), 
to_sfixed(-989045751.0/4294967296.0,1,-nbitq), 
to_sfixed(666928860.0/4294967296.0,1,-nbitq), 
to_sfixed(-276418236.0/4294967296.0,1,-nbitq), 
to_sfixed(254729887.0/4294967296.0,1,-nbitq), 
to_sfixed(153529542.0/4294967296.0,1,-nbitq), 
to_sfixed(610045209.0/4294967296.0,1,-nbitq), 
to_sfixed(23691862.0/4294967296.0,1,-nbitq), 
to_sfixed(-285871311.0/4294967296.0,1,-nbitq), 
to_sfixed(1380302633.0/4294967296.0,1,-nbitq), 
to_sfixed(-837975257.0/4294967296.0,1,-nbitq), 
to_sfixed(158069192.0/4294967296.0,1,-nbitq), 
to_sfixed(-462965276.0/4294967296.0,1,-nbitq), 
to_sfixed(978295148.0/4294967296.0,1,-nbitq), 
to_sfixed(415691632.0/4294967296.0,1,-nbitq), 
to_sfixed(-137644504.0/4294967296.0,1,-nbitq), 
to_sfixed(509887021.0/4294967296.0,1,-nbitq), 
to_sfixed(150478753.0/4294967296.0,1,-nbitq), 
to_sfixed(-1628625786.0/4294967296.0,1,-nbitq), 
to_sfixed(-496054779.0/4294967296.0,1,-nbitq), 
to_sfixed(-870238538.0/4294967296.0,1,-nbitq), 
to_sfixed(921960420.0/4294967296.0,1,-nbitq), 
to_sfixed(-1025021079.0/4294967296.0,1,-nbitq), 
to_sfixed(797752963.0/4294967296.0,1,-nbitq), 
to_sfixed(-932844722.0/4294967296.0,1,-nbitq), 
to_sfixed(616014286.0/4294967296.0,1,-nbitq), 
to_sfixed(999447655.0/4294967296.0,1,-nbitq), 
to_sfixed(200897051.0/4294967296.0,1,-nbitq), 
to_sfixed(-1059831588.0/4294967296.0,1,-nbitq), 
to_sfixed(-126173442.0/4294967296.0,1,-nbitq), 
to_sfixed(572114007.0/4294967296.0,1,-nbitq), 
to_sfixed(-340642302.0/4294967296.0,1,-nbitq), 
to_sfixed(-342574478.0/4294967296.0,1,-nbitq), 
to_sfixed(1406762253.0/4294967296.0,1,-nbitq), 
to_sfixed(314560952.0/4294967296.0,1,-nbitq), 
to_sfixed(233401019.0/4294967296.0,1,-nbitq), 
to_sfixed(-195059598.0/4294967296.0,1,-nbitq), 
to_sfixed(-127753247.0/4294967296.0,1,-nbitq), 
to_sfixed(380178340.0/4294967296.0,1,-nbitq), 
to_sfixed(-186061724.0/4294967296.0,1,-nbitq), 
to_sfixed(211884199.0/4294967296.0,1,-nbitq), 
to_sfixed(-375286336.0/4294967296.0,1,-nbitq), 
to_sfixed(1178262067.0/4294967296.0,1,-nbitq), 
to_sfixed(-706038793.0/4294967296.0,1,-nbitq), 
to_sfixed(-730115210.0/4294967296.0,1,-nbitq), 
to_sfixed(-270797675.0/4294967296.0,1,-nbitq), 
to_sfixed(-106629334.0/4294967296.0,1,-nbitq), 
to_sfixed(-21785766.0/4294967296.0,1,-nbitq), 
to_sfixed(42028713.0/4294967296.0,1,-nbitq), 
to_sfixed(-102800691.0/4294967296.0,1,-nbitq), 
to_sfixed(208683750.0/4294967296.0,1,-nbitq), 
to_sfixed(-108897144.0/4294967296.0,1,-nbitq), 
to_sfixed(151008452.0/4294967296.0,1,-nbitq), 
to_sfixed(-105044608.0/4294967296.0,1,-nbitq), 
to_sfixed(-157754051.0/4294967296.0,1,-nbitq), 
to_sfixed(245916842.0/4294967296.0,1,-nbitq), 
to_sfixed(91184242.0/4294967296.0,1,-nbitq), 
to_sfixed(-178598805.0/4294967296.0,1,-nbitq), 
to_sfixed(292054327.0/4294967296.0,1,-nbitq), 
to_sfixed(-118441287.0/4294967296.0,1,-nbitq), 
to_sfixed(-459712862.0/4294967296.0,1,-nbitq), 
to_sfixed(-1433214090.0/4294967296.0,1,-nbitq), 
to_sfixed(327334469.0/4294967296.0,1,-nbitq), 
to_sfixed(-165943951.0/4294967296.0,1,-nbitq), 
to_sfixed(49075356.0/4294967296.0,1,-nbitq), 
to_sfixed(-4381039.0/4294967296.0,1,-nbitq), 
to_sfixed(818874583.0/4294967296.0,1,-nbitq), 
to_sfixed(-343234104.0/4294967296.0,1,-nbitq), 
to_sfixed(397829680.0/4294967296.0,1,-nbitq), 
to_sfixed(73657422.0/4294967296.0,1,-nbitq), 
to_sfixed(-175008274.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-487613649.0/4294967296.0,1,-nbitq), 
to_sfixed(395195958.0/4294967296.0,1,-nbitq), 
to_sfixed(-1098404628.0/4294967296.0,1,-nbitq), 
to_sfixed(70025949.0/4294967296.0,1,-nbitq), 
to_sfixed(-530238188.0/4294967296.0,1,-nbitq), 
to_sfixed(-953249405.0/4294967296.0,1,-nbitq), 
to_sfixed(150932804.0/4294967296.0,1,-nbitq), 
to_sfixed(-214988153.0/4294967296.0,1,-nbitq), 
to_sfixed(1058540352.0/4294967296.0,1,-nbitq), 
to_sfixed(-134881905.0/4294967296.0,1,-nbitq), 
to_sfixed(-976963762.0/4294967296.0,1,-nbitq), 
to_sfixed(-287910962.0/4294967296.0,1,-nbitq), 
to_sfixed(-1068989623.0/4294967296.0,1,-nbitq), 
to_sfixed(640419681.0/4294967296.0,1,-nbitq), 
to_sfixed(-120527719.0/4294967296.0,1,-nbitq), 
to_sfixed(269439654.0/4294967296.0,1,-nbitq), 
to_sfixed(-13682384.0/4294967296.0,1,-nbitq), 
to_sfixed(171921177.0/4294967296.0,1,-nbitq), 
to_sfixed(995514374.0/4294967296.0,1,-nbitq), 
to_sfixed(-700158813.0/4294967296.0,1,-nbitq), 
to_sfixed(-91413396.0/4294967296.0,1,-nbitq), 
to_sfixed(-714773340.0/4294967296.0,1,-nbitq), 
to_sfixed(282577991.0/4294967296.0,1,-nbitq), 
to_sfixed(404487912.0/4294967296.0,1,-nbitq), 
to_sfixed(347223907.0/4294967296.0,1,-nbitq), 
to_sfixed(-545341067.0/4294967296.0,1,-nbitq), 
to_sfixed(-246722552.0/4294967296.0,1,-nbitq), 
to_sfixed(-1254626966.0/4294967296.0,1,-nbitq), 
to_sfixed(-797221891.0/4294967296.0,1,-nbitq), 
to_sfixed(-381802637.0/4294967296.0,1,-nbitq), 
to_sfixed(-530796062.0/4294967296.0,1,-nbitq), 
to_sfixed(-88548876.0/4294967296.0,1,-nbitq), 
to_sfixed(-309544067.0/4294967296.0,1,-nbitq), 
to_sfixed(21588561.0/4294967296.0,1,-nbitq), 
to_sfixed(828134316.0/4294967296.0,1,-nbitq), 
to_sfixed(1017470453.0/4294967296.0,1,-nbitq), 
to_sfixed(1034274025.0/4294967296.0,1,-nbitq), 
to_sfixed(-754507002.0/4294967296.0,1,-nbitq), 
to_sfixed(-280244103.0/4294967296.0,1,-nbitq), 
to_sfixed(-22683461.0/4294967296.0,1,-nbitq), 
to_sfixed(-177563475.0/4294967296.0,1,-nbitq), 
to_sfixed(-611113258.0/4294967296.0,1,-nbitq), 
to_sfixed(676303218.0/4294967296.0,1,-nbitq), 
to_sfixed(105026302.0/4294967296.0,1,-nbitq), 
to_sfixed(-167136406.0/4294967296.0,1,-nbitq), 
to_sfixed(127397820.0/4294967296.0,1,-nbitq), 
to_sfixed(-35767726.0/4294967296.0,1,-nbitq), 
to_sfixed(650052263.0/4294967296.0,1,-nbitq), 
to_sfixed(-137877126.0/4294967296.0,1,-nbitq), 
to_sfixed(242902347.0/4294967296.0,1,-nbitq), 
to_sfixed(-671520419.0/4294967296.0,1,-nbitq), 
to_sfixed(-78957186.0/4294967296.0,1,-nbitq), 
to_sfixed(404254087.0/4294967296.0,1,-nbitq), 
to_sfixed(-772207875.0/4294967296.0,1,-nbitq), 
to_sfixed(735346267.0/4294967296.0,1,-nbitq), 
to_sfixed(-167341070.0/4294967296.0,1,-nbitq), 
to_sfixed(-789292685.0/4294967296.0,1,-nbitq), 
to_sfixed(-7319548.0/4294967296.0,1,-nbitq), 
to_sfixed(-330816644.0/4294967296.0,1,-nbitq), 
to_sfixed(112001896.0/4294967296.0,1,-nbitq), 
to_sfixed(-245259165.0/4294967296.0,1,-nbitq), 
to_sfixed(67524443.0/4294967296.0,1,-nbitq), 
to_sfixed(118742397.0/4294967296.0,1,-nbitq), 
to_sfixed(-322226023.0/4294967296.0,1,-nbitq), 
to_sfixed(154578493.0/4294967296.0,1,-nbitq), 
to_sfixed(-70259775.0/4294967296.0,1,-nbitq), 
to_sfixed(127632860.0/4294967296.0,1,-nbitq), 
to_sfixed(1083552812.0/4294967296.0,1,-nbitq), 
to_sfixed(-229653678.0/4294967296.0,1,-nbitq), 
to_sfixed(-86175254.0/4294967296.0,1,-nbitq), 
to_sfixed(-817083088.0/4294967296.0,1,-nbitq), 
to_sfixed(190732788.0/4294967296.0,1,-nbitq), 
to_sfixed(128647215.0/4294967296.0,1,-nbitq), 
to_sfixed(-303083345.0/4294967296.0,1,-nbitq), 
to_sfixed(324395691.0/4294967296.0,1,-nbitq), 
to_sfixed(985118296.0/4294967296.0,1,-nbitq), 
to_sfixed(-1164748041.0/4294967296.0,1,-nbitq), 
to_sfixed(676813265.0/4294967296.0,1,-nbitq), 
to_sfixed(188173785.0/4294967296.0,1,-nbitq), 
to_sfixed(-218847079.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(312155843.0/4294967296.0,1,-nbitq), 
to_sfixed(-923319676.0/4294967296.0,1,-nbitq), 
to_sfixed(656939964.0/4294967296.0,1,-nbitq), 
to_sfixed(731503622.0/4294967296.0,1,-nbitq), 
to_sfixed(-243766730.0/4294967296.0,1,-nbitq), 
to_sfixed(-376720260.0/4294967296.0,1,-nbitq), 
to_sfixed(516822222.0/4294967296.0,1,-nbitq), 
to_sfixed(-368539003.0/4294967296.0,1,-nbitq), 
to_sfixed(116903517.0/4294967296.0,1,-nbitq), 
to_sfixed(300562152.0/4294967296.0,1,-nbitq), 
to_sfixed(-132990032.0/4294967296.0,1,-nbitq), 
to_sfixed(783267984.0/4294967296.0,1,-nbitq), 
to_sfixed(-645376894.0/4294967296.0,1,-nbitq), 
to_sfixed(62281295.0/4294967296.0,1,-nbitq), 
to_sfixed(361096943.0/4294967296.0,1,-nbitq), 
to_sfixed(659816775.0/4294967296.0,1,-nbitq), 
to_sfixed(-363904924.0/4294967296.0,1,-nbitq), 
to_sfixed(57135392.0/4294967296.0,1,-nbitq), 
to_sfixed(206388004.0/4294967296.0,1,-nbitq), 
to_sfixed(-260871429.0/4294967296.0,1,-nbitq), 
to_sfixed(-72500340.0/4294967296.0,1,-nbitq), 
to_sfixed(10786132.0/4294967296.0,1,-nbitq), 
to_sfixed(-210539484.0/4294967296.0,1,-nbitq), 
to_sfixed(-220712974.0/4294967296.0,1,-nbitq), 
to_sfixed(-288855751.0/4294967296.0,1,-nbitq), 
to_sfixed(-241745990.0/4294967296.0,1,-nbitq), 
to_sfixed(-1130241835.0/4294967296.0,1,-nbitq), 
to_sfixed(-918612097.0/4294967296.0,1,-nbitq), 
to_sfixed(111746578.0/4294967296.0,1,-nbitq), 
to_sfixed(-137372351.0/4294967296.0,1,-nbitq), 
to_sfixed(-699162873.0/4294967296.0,1,-nbitq), 
to_sfixed(-465240256.0/4294967296.0,1,-nbitq), 
to_sfixed(-874459008.0/4294967296.0,1,-nbitq), 
to_sfixed(296194353.0/4294967296.0,1,-nbitq), 
to_sfixed(1244570815.0/4294967296.0,1,-nbitq), 
to_sfixed(365413504.0/4294967296.0,1,-nbitq), 
to_sfixed(1008332135.0/4294967296.0,1,-nbitq), 
to_sfixed(523665797.0/4294967296.0,1,-nbitq), 
to_sfixed(-344751974.0/4294967296.0,1,-nbitq), 
to_sfixed(21194154.0/4294967296.0,1,-nbitq), 
to_sfixed(77361900.0/4294967296.0,1,-nbitq), 
to_sfixed(-362533809.0/4294967296.0,1,-nbitq), 
to_sfixed(237292382.0/4294967296.0,1,-nbitq), 
to_sfixed(353710631.0/4294967296.0,1,-nbitq), 
to_sfixed(258453675.0/4294967296.0,1,-nbitq), 
to_sfixed(466309036.0/4294967296.0,1,-nbitq), 
to_sfixed(-262447886.0/4294967296.0,1,-nbitq), 
to_sfixed(727891518.0/4294967296.0,1,-nbitq), 
to_sfixed(-318847760.0/4294967296.0,1,-nbitq), 
to_sfixed(912345945.0/4294967296.0,1,-nbitq), 
to_sfixed(-462077329.0/4294967296.0,1,-nbitq), 
to_sfixed(759844591.0/4294967296.0,1,-nbitq), 
to_sfixed(-188918302.0/4294967296.0,1,-nbitq), 
to_sfixed(-305305986.0/4294967296.0,1,-nbitq), 
to_sfixed(633377828.0/4294967296.0,1,-nbitq), 
to_sfixed(869640378.0/4294967296.0,1,-nbitq), 
to_sfixed(-725009699.0/4294967296.0,1,-nbitq), 
to_sfixed(-19142454.0/4294967296.0,1,-nbitq), 
to_sfixed(423093654.0/4294967296.0,1,-nbitq), 
to_sfixed(282322927.0/4294967296.0,1,-nbitq), 
to_sfixed(-283760210.0/4294967296.0,1,-nbitq), 
to_sfixed(240168954.0/4294967296.0,1,-nbitq), 
to_sfixed(-551360882.0/4294967296.0,1,-nbitq), 
to_sfixed(399875445.0/4294967296.0,1,-nbitq), 
to_sfixed(-52829542.0/4294967296.0,1,-nbitq), 
to_sfixed(361122591.0/4294967296.0,1,-nbitq), 
to_sfixed(-652378236.0/4294967296.0,1,-nbitq), 
to_sfixed(604419171.0/4294967296.0,1,-nbitq), 
to_sfixed(64674546.0/4294967296.0,1,-nbitq), 
to_sfixed(12283639.0/4294967296.0,1,-nbitq), 
to_sfixed(-1012132345.0/4294967296.0,1,-nbitq), 
to_sfixed(-292679949.0/4294967296.0,1,-nbitq), 
to_sfixed(-38634071.0/4294967296.0,1,-nbitq), 
to_sfixed(-179015046.0/4294967296.0,1,-nbitq), 
to_sfixed(418728020.0/4294967296.0,1,-nbitq), 
to_sfixed(490849443.0/4294967296.0,1,-nbitq), 
to_sfixed(-148677997.0/4294967296.0,1,-nbitq), 
to_sfixed(-45311374.0/4294967296.0,1,-nbitq), 
to_sfixed(489934098.0/4294967296.0,1,-nbitq), 
to_sfixed(-372333538.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(552662699.0/4294967296.0,1,-nbitq), 
to_sfixed(-994551249.0/4294967296.0,1,-nbitq), 
to_sfixed(314975502.0/4294967296.0,1,-nbitq), 
to_sfixed(-287417983.0/4294967296.0,1,-nbitq), 
to_sfixed(-578935513.0/4294967296.0,1,-nbitq), 
to_sfixed(141128109.0/4294967296.0,1,-nbitq), 
to_sfixed(87048595.0/4294967296.0,1,-nbitq), 
to_sfixed(-187734966.0/4294967296.0,1,-nbitq), 
to_sfixed(88741310.0/4294967296.0,1,-nbitq), 
to_sfixed(294482638.0/4294967296.0,1,-nbitq), 
to_sfixed(-634544814.0/4294967296.0,1,-nbitq), 
to_sfixed(395883355.0/4294967296.0,1,-nbitq), 
to_sfixed(-97299679.0/4294967296.0,1,-nbitq), 
to_sfixed(1434658327.0/4294967296.0,1,-nbitq), 
to_sfixed(-327045799.0/4294967296.0,1,-nbitq), 
to_sfixed(850230807.0/4294967296.0,1,-nbitq), 
to_sfixed(-73830224.0/4294967296.0,1,-nbitq), 
to_sfixed(219994284.0/4294967296.0,1,-nbitq), 
to_sfixed(210258360.0/4294967296.0,1,-nbitq), 
to_sfixed(-405802697.0/4294967296.0,1,-nbitq), 
to_sfixed(323841755.0/4294967296.0,1,-nbitq), 
to_sfixed(-453604622.0/4294967296.0,1,-nbitq), 
to_sfixed(-154039884.0/4294967296.0,1,-nbitq), 
to_sfixed(494158861.0/4294967296.0,1,-nbitq), 
to_sfixed(100724538.0/4294967296.0,1,-nbitq), 
to_sfixed(1112126086.0/4294967296.0,1,-nbitq), 
to_sfixed(-317312187.0/4294967296.0,1,-nbitq), 
to_sfixed(-696739756.0/4294967296.0,1,-nbitq), 
to_sfixed(156447297.0/4294967296.0,1,-nbitq), 
to_sfixed(-324464344.0/4294967296.0,1,-nbitq), 
to_sfixed(-370085909.0/4294967296.0,1,-nbitq), 
to_sfixed(-1103821665.0/4294967296.0,1,-nbitq), 
to_sfixed(-1604904064.0/4294967296.0,1,-nbitq), 
to_sfixed(-13303834.0/4294967296.0,1,-nbitq), 
to_sfixed(690455292.0/4294967296.0,1,-nbitq), 
to_sfixed(534304190.0/4294967296.0,1,-nbitq), 
to_sfixed(564769016.0/4294967296.0,1,-nbitq), 
to_sfixed(387966093.0/4294967296.0,1,-nbitq), 
to_sfixed(-627543644.0/4294967296.0,1,-nbitq), 
to_sfixed(594480755.0/4294967296.0,1,-nbitq), 
to_sfixed(66690807.0/4294967296.0,1,-nbitq), 
to_sfixed(21050458.0/4294967296.0,1,-nbitq), 
to_sfixed(91543578.0/4294967296.0,1,-nbitq), 
to_sfixed(1029885073.0/4294967296.0,1,-nbitq), 
to_sfixed(764483453.0/4294967296.0,1,-nbitq), 
to_sfixed(514000478.0/4294967296.0,1,-nbitq), 
to_sfixed(241999381.0/4294967296.0,1,-nbitq), 
to_sfixed(326432676.0/4294967296.0,1,-nbitq), 
to_sfixed(-542603529.0/4294967296.0,1,-nbitq), 
to_sfixed(945705128.0/4294967296.0,1,-nbitq), 
to_sfixed(-96360889.0/4294967296.0,1,-nbitq), 
to_sfixed(1420495.0/4294967296.0,1,-nbitq), 
to_sfixed(-1434937122.0/4294967296.0,1,-nbitq), 
to_sfixed(576785059.0/4294967296.0,1,-nbitq), 
to_sfixed(447482111.0/4294967296.0,1,-nbitq), 
to_sfixed(396511679.0/4294967296.0,1,-nbitq), 
to_sfixed(101579276.0/4294967296.0,1,-nbitq), 
to_sfixed(-1621022631.0/4294967296.0,1,-nbitq), 
to_sfixed(-288398067.0/4294967296.0,1,-nbitq), 
to_sfixed(357119778.0/4294967296.0,1,-nbitq), 
to_sfixed(149705562.0/4294967296.0,1,-nbitq), 
to_sfixed(594171328.0/4294967296.0,1,-nbitq), 
to_sfixed(-910698467.0/4294967296.0,1,-nbitq), 
to_sfixed(-177597689.0/4294967296.0,1,-nbitq), 
to_sfixed(-745409219.0/4294967296.0,1,-nbitq), 
to_sfixed(-61752524.0/4294967296.0,1,-nbitq), 
to_sfixed(-1691296738.0/4294967296.0,1,-nbitq), 
to_sfixed(939371158.0/4294967296.0,1,-nbitq), 
to_sfixed(-311183380.0/4294967296.0,1,-nbitq), 
to_sfixed(13659594.0/4294967296.0,1,-nbitq), 
to_sfixed(-96220910.0/4294967296.0,1,-nbitq), 
to_sfixed(-180866336.0/4294967296.0,1,-nbitq), 
to_sfixed(-564726263.0/4294967296.0,1,-nbitq), 
to_sfixed(-218555094.0/4294967296.0,1,-nbitq), 
to_sfixed(191680385.0/4294967296.0,1,-nbitq), 
to_sfixed(510855700.0/4294967296.0,1,-nbitq), 
to_sfixed(-35542657.0/4294967296.0,1,-nbitq), 
to_sfixed(294231736.0/4294967296.0,1,-nbitq), 
to_sfixed(665539318.0/4294967296.0,1,-nbitq), 
to_sfixed(192741039.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(183767751.0/4294967296.0,1,-nbitq), 
to_sfixed(-436726777.0/4294967296.0,1,-nbitq), 
to_sfixed(512535993.0/4294967296.0,1,-nbitq), 
to_sfixed(-430961184.0/4294967296.0,1,-nbitq), 
to_sfixed(-106924874.0/4294967296.0,1,-nbitq), 
to_sfixed(-460174750.0/4294967296.0,1,-nbitq), 
to_sfixed(89128609.0/4294967296.0,1,-nbitq), 
to_sfixed(87876648.0/4294967296.0,1,-nbitq), 
to_sfixed(202439343.0/4294967296.0,1,-nbitq), 
to_sfixed(-312185632.0/4294967296.0,1,-nbitq), 
to_sfixed(-281046264.0/4294967296.0,1,-nbitq), 
to_sfixed(681663361.0/4294967296.0,1,-nbitq), 
to_sfixed(-106006200.0/4294967296.0,1,-nbitq), 
to_sfixed(691760606.0/4294967296.0,1,-nbitq), 
to_sfixed(351625935.0/4294967296.0,1,-nbitq), 
to_sfixed(355219913.0/4294967296.0,1,-nbitq), 
to_sfixed(-158125993.0/4294967296.0,1,-nbitq), 
to_sfixed(387228644.0/4294967296.0,1,-nbitq), 
to_sfixed(64298839.0/4294967296.0,1,-nbitq), 
to_sfixed(-147095645.0/4294967296.0,1,-nbitq), 
to_sfixed(-371611624.0/4294967296.0,1,-nbitq), 
to_sfixed(-401976726.0/4294967296.0,1,-nbitq), 
to_sfixed(-1036176713.0/4294967296.0,1,-nbitq), 
to_sfixed(105414709.0/4294967296.0,1,-nbitq), 
to_sfixed(445600157.0/4294967296.0,1,-nbitq), 
to_sfixed(824580021.0/4294967296.0,1,-nbitq), 
to_sfixed(-166407320.0/4294967296.0,1,-nbitq), 
to_sfixed(478439274.0/4294967296.0,1,-nbitq), 
to_sfixed(-231797393.0/4294967296.0,1,-nbitq), 
to_sfixed(-266427811.0/4294967296.0,1,-nbitq), 
to_sfixed(-61588855.0/4294967296.0,1,-nbitq), 
to_sfixed(-809554911.0/4294967296.0,1,-nbitq), 
to_sfixed(-987332752.0/4294967296.0,1,-nbitq), 
to_sfixed(79537820.0/4294967296.0,1,-nbitq), 
to_sfixed(479593407.0/4294967296.0,1,-nbitq), 
to_sfixed(1300751783.0/4294967296.0,1,-nbitq), 
to_sfixed(852459430.0/4294967296.0,1,-nbitq), 
to_sfixed(638353832.0/4294967296.0,1,-nbitq), 
to_sfixed(-122398088.0/4294967296.0,1,-nbitq), 
to_sfixed(-75130308.0/4294967296.0,1,-nbitq), 
to_sfixed(528642891.0/4294967296.0,1,-nbitq), 
to_sfixed(60085131.0/4294967296.0,1,-nbitq), 
to_sfixed(38976518.0/4294967296.0,1,-nbitq), 
to_sfixed(1585983204.0/4294967296.0,1,-nbitq), 
to_sfixed(222699352.0/4294967296.0,1,-nbitq), 
to_sfixed(1893309948.0/4294967296.0,1,-nbitq), 
to_sfixed(374700211.0/4294967296.0,1,-nbitq), 
to_sfixed(322433089.0/4294967296.0,1,-nbitq), 
to_sfixed(76223874.0/4294967296.0,1,-nbitq), 
to_sfixed(261243710.0/4294967296.0,1,-nbitq), 
to_sfixed(-162628235.0/4294967296.0,1,-nbitq), 
to_sfixed(-48566811.0/4294967296.0,1,-nbitq), 
to_sfixed(-881024652.0/4294967296.0,1,-nbitq), 
to_sfixed(1430555263.0/4294967296.0,1,-nbitq), 
to_sfixed(-6880780.0/4294967296.0,1,-nbitq), 
to_sfixed(86204243.0/4294967296.0,1,-nbitq), 
to_sfixed(1099330512.0/4294967296.0,1,-nbitq), 
to_sfixed(-1705020884.0/4294967296.0,1,-nbitq), 
to_sfixed(140835021.0/4294967296.0,1,-nbitq), 
to_sfixed(-37146565.0/4294967296.0,1,-nbitq), 
to_sfixed(188418003.0/4294967296.0,1,-nbitq), 
to_sfixed(8831546.0/4294967296.0,1,-nbitq), 
to_sfixed(-1485042062.0/4294967296.0,1,-nbitq), 
to_sfixed(-42897936.0/4294967296.0,1,-nbitq), 
to_sfixed(162316951.0/4294967296.0,1,-nbitq), 
to_sfixed(-332547924.0/4294967296.0,1,-nbitq), 
to_sfixed(-761643162.0/4294967296.0,1,-nbitq), 
to_sfixed(1016561219.0/4294967296.0,1,-nbitq), 
to_sfixed(-226870901.0/4294967296.0,1,-nbitq), 
to_sfixed(-342636415.0/4294967296.0,1,-nbitq), 
to_sfixed(587000095.0/4294967296.0,1,-nbitq), 
to_sfixed(-44394576.0/4294967296.0,1,-nbitq), 
to_sfixed(241425659.0/4294967296.0,1,-nbitq), 
to_sfixed(-194738702.0/4294967296.0,1,-nbitq), 
to_sfixed(-86773182.0/4294967296.0,1,-nbitq), 
to_sfixed(393274403.0/4294967296.0,1,-nbitq), 
to_sfixed(-178387473.0/4294967296.0,1,-nbitq), 
to_sfixed(363926110.0/4294967296.0,1,-nbitq), 
to_sfixed(555903843.0/4294967296.0,1,-nbitq), 
to_sfixed(175314323.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-31753070.0/4294967296.0,1,-nbitq), 
to_sfixed(-32414575.0/4294967296.0,1,-nbitq), 
to_sfixed(-8620960.0/4294967296.0,1,-nbitq), 
to_sfixed(-468390914.0/4294967296.0,1,-nbitq), 
to_sfixed(-579335241.0/4294967296.0,1,-nbitq), 
to_sfixed(-534005324.0/4294967296.0,1,-nbitq), 
to_sfixed(-58216676.0/4294967296.0,1,-nbitq), 
to_sfixed(-586322923.0/4294967296.0,1,-nbitq), 
to_sfixed(-429091337.0/4294967296.0,1,-nbitq), 
to_sfixed(-165821184.0/4294967296.0,1,-nbitq), 
to_sfixed(-160019657.0/4294967296.0,1,-nbitq), 
to_sfixed(551200639.0/4294967296.0,1,-nbitq), 
to_sfixed(-129370373.0/4294967296.0,1,-nbitq), 
to_sfixed(1211213054.0/4294967296.0,1,-nbitq), 
to_sfixed(-213325749.0/4294967296.0,1,-nbitq), 
to_sfixed(375803753.0/4294967296.0,1,-nbitq), 
to_sfixed(194788405.0/4294967296.0,1,-nbitq), 
to_sfixed(83349135.0/4294967296.0,1,-nbitq), 
to_sfixed(152951046.0/4294967296.0,1,-nbitq), 
to_sfixed(-345664161.0/4294967296.0,1,-nbitq), 
to_sfixed(107642421.0/4294967296.0,1,-nbitq), 
to_sfixed(-734477786.0/4294967296.0,1,-nbitq), 
to_sfixed(-844380671.0/4294967296.0,1,-nbitq), 
to_sfixed(3212509.0/4294967296.0,1,-nbitq), 
to_sfixed(-83150193.0/4294967296.0,1,-nbitq), 
to_sfixed(282719812.0/4294967296.0,1,-nbitq), 
to_sfixed(-453994098.0/4294967296.0,1,-nbitq), 
to_sfixed(556399702.0/4294967296.0,1,-nbitq), 
to_sfixed(407978627.0/4294967296.0,1,-nbitq), 
to_sfixed(-56193784.0/4294967296.0,1,-nbitq), 
to_sfixed(838347729.0/4294967296.0,1,-nbitq), 
to_sfixed(-894276290.0/4294967296.0,1,-nbitq), 
to_sfixed(-966495286.0/4294967296.0,1,-nbitq), 
to_sfixed(-145096160.0/4294967296.0,1,-nbitq), 
to_sfixed(493113514.0/4294967296.0,1,-nbitq), 
to_sfixed(506494382.0/4294967296.0,1,-nbitq), 
to_sfixed(488704338.0/4294967296.0,1,-nbitq), 
to_sfixed(543327667.0/4294967296.0,1,-nbitq), 
to_sfixed(-48005527.0/4294967296.0,1,-nbitq), 
to_sfixed(92368119.0/4294967296.0,1,-nbitq), 
to_sfixed(645573484.0/4294967296.0,1,-nbitq), 
to_sfixed(1177046006.0/4294967296.0,1,-nbitq), 
to_sfixed(-1133377967.0/4294967296.0,1,-nbitq), 
to_sfixed(1479121462.0/4294967296.0,1,-nbitq), 
to_sfixed(-101447882.0/4294967296.0,1,-nbitq), 
to_sfixed(1355762816.0/4294967296.0,1,-nbitq), 
to_sfixed(361900276.0/4294967296.0,1,-nbitq), 
to_sfixed(268559468.0/4294967296.0,1,-nbitq), 
to_sfixed(-311898510.0/4294967296.0,1,-nbitq), 
to_sfixed(-115945003.0/4294967296.0,1,-nbitq), 
to_sfixed(-457227174.0/4294967296.0,1,-nbitq), 
to_sfixed(472659396.0/4294967296.0,1,-nbitq), 
to_sfixed(-1048073437.0/4294967296.0,1,-nbitq), 
to_sfixed(624942073.0/4294967296.0,1,-nbitq), 
to_sfixed(28628573.0/4294967296.0,1,-nbitq), 
to_sfixed(402935524.0/4294967296.0,1,-nbitq), 
to_sfixed(458662756.0/4294967296.0,1,-nbitq), 
to_sfixed(-1182739729.0/4294967296.0,1,-nbitq), 
to_sfixed(159205220.0/4294967296.0,1,-nbitq), 
to_sfixed(232996238.0/4294967296.0,1,-nbitq), 
to_sfixed(45331608.0/4294967296.0,1,-nbitq), 
to_sfixed(652861879.0/4294967296.0,1,-nbitq), 
to_sfixed(-960381843.0/4294967296.0,1,-nbitq), 
to_sfixed(-272080287.0/4294967296.0,1,-nbitq), 
to_sfixed(-73949412.0/4294967296.0,1,-nbitq), 
to_sfixed(236933419.0/4294967296.0,1,-nbitq), 
to_sfixed(-154813588.0/4294967296.0,1,-nbitq), 
to_sfixed(1098759566.0/4294967296.0,1,-nbitq), 
to_sfixed(329089321.0/4294967296.0,1,-nbitq), 
to_sfixed(-1169467787.0/4294967296.0,1,-nbitq), 
to_sfixed(686487089.0/4294967296.0,1,-nbitq), 
to_sfixed(-94992905.0/4294967296.0,1,-nbitq), 
to_sfixed(-455570980.0/4294967296.0,1,-nbitq), 
to_sfixed(-294452204.0/4294967296.0,1,-nbitq), 
to_sfixed(-217273973.0/4294967296.0,1,-nbitq), 
to_sfixed(-53821867.0/4294967296.0,1,-nbitq), 
to_sfixed(-668359552.0/4294967296.0,1,-nbitq), 
to_sfixed(111883496.0/4294967296.0,1,-nbitq), 
to_sfixed(162556465.0/4294967296.0,1,-nbitq), 
to_sfixed(-241419768.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-60135925.0/4294967296.0,1,-nbitq), 
to_sfixed(488389504.0/4294967296.0,1,-nbitq), 
to_sfixed(435837779.0/4294967296.0,1,-nbitq), 
to_sfixed(-195825953.0/4294967296.0,1,-nbitq), 
to_sfixed(-514826154.0/4294967296.0,1,-nbitq), 
to_sfixed(-680735705.0/4294967296.0,1,-nbitq), 
to_sfixed(-367694063.0/4294967296.0,1,-nbitq), 
to_sfixed(-507977399.0/4294967296.0,1,-nbitq), 
to_sfixed(-226792992.0/4294967296.0,1,-nbitq), 
to_sfixed(368953867.0/4294967296.0,1,-nbitq), 
to_sfixed(-256413000.0/4294967296.0,1,-nbitq), 
to_sfixed(375431477.0/4294967296.0,1,-nbitq), 
to_sfixed(-760831234.0/4294967296.0,1,-nbitq), 
to_sfixed(1156042382.0/4294967296.0,1,-nbitq), 
to_sfixed(324447025.0/4294967296.0,1,-nbitq), 
to_sfixed(202059340.0/4294967296.0,1,-nbitq), 
to_sfixed(-133713301.0/4294967296.0,1,-nbitq), 
to_sfixed(-80735316.0/4294967296.0,1,-nbitq), 
to_sfixed(-361067935.0/4294967296.0,1,-nbitq), 
to_sfixed(-110440332.0/4294967296.0,1,-nbitq), 
to_sfixed(362004203.0/4294967296.0,1,-nbitq), 
to_sfixed(-68454462.0/4294967296.0,1,-nbitq), 
to_sfixed(-895119701.0/4294967296.0,1,-nbitq), 
to_sfixed(514929071.0/4294967296.0,1,-nbitq), 
to_sfixed(-87236801.0/4294967296.0,1,-nbitq), 
to_sfixed(-1131349524.0/4294967296.0,1,-nbitq), 
to_sfixed(-638359288.0/4294967296.0,1,-nbitq), 
to_sfixed(786643847.0/4294967296.0,1,-nbitq), 
to_sfixed(-44574848.0/4294967296.0,1,-nbitq), 
to_sfixed(-648261180.0/4294967296.0,1,-nbitq), 
to_sfixed(1325998368.0/4294967296.0,1,-nbitq), 
to_sfixed(-723146987.0/4294967296.0,1,-nbitq), 
to_sfixed(-767923850.0/4294967296.0,1,-nbitq), 
to_sfixed(-671069817.0/4294967296.0,1,-nbitq), 
to_sfixed(454209484.0/4294967296.0,1,-nbitq), 
to_sfixed(497006511.0/4294967296.0,1,-nbitq), 
to_sfixed(363197021.0/4294967296.0,1,-nbitq), 
to_sfixed(101849610.0/4294967296.0,1,-nbitq), 
to_sfixed(593221129.0/4294967296.0,1,-nbitq), 
to_sfixed(5795499.0/4294967296.0,1,-nbitq), 
to_sfixed(208945369.0/4294967296.0,1,-nbitq), 
to_sfixed(638148620.0/4294967296.0,1,-nbitq), 
to_sfixed(-339296132.0/4294967296.0,1,-nbitq), 
to_sfixed(1307738371.0/4294967296.0,1,-nbitq), 
to_sfixed(-125899013.0/4294967296.0,1,-nbitq), 
to_sfixed(826806276.0/4294967296.0,1,-nbitq), 
to_sfixed(320455936.0/4294967296.0,1,-nbitq), 
to_sfixed(-522966142.0/4294967296.0,1,-nbitq), 
to_sfixed(-401287364.0/4294967296.0,1,-nbitq), 
to_sfixed(-496160556.0/4294967296.0,1,-nbitq), 
to_sfixed(355523745.0/4294967296.0,1,-nbitq), 
to_sfixed(-109851584.0/4294967296.0,1,-nbitq), 
to_sfixed(-244442972.0/4294967296.0,1,-nbitq), 
to_sfixed(359969407.0/4294967296.0,1,-nbitq), 
to_sfixed(-273029451.0/4294967296.0,1,-nbitq), 
to_sfixed(-88277492.0/4294967296.0,1,-nbitq), 
to_sfixed(-83679598.0/4294967296.0,1,-nbitq), 
to_sfixed(-303472629.0/4294967296.0,1,-nbitq), 
to_sfixed(-311388144.0/4294967296.0,1,-nbitq), 
to_sfixed(-115143393.0/4294967296.0,1,-nbitq), 
to_sfixed(-307803272.0/4294967296.0,1,-nbitq), 
to_sfixed(245476439.0/4294967296.0,1,-nbitq), 
to_sfixed(173650768.0/4294967296.0,1,-nbitq), 
to_sfixed(-185271483.0/4294967296.0,1,-nbitq), 
to_sfixed(166437919.0/4294967296.0,1,-nbitq), 
to_sfixed(-244154640.0/4294967296.0,1,-nbitq), 
to_sfixed(-445469372.0/4294967296.0,1,-nbitq), 
to_sfixed(392210839.0/4294967296.0,1,-nbitq), 
to_sfixed(181140724.0/4294967296.0,1,-nbitq), 
to_sfixed(-701603952.0/4294967296.0,1,-nbitq), 
to_sfixed(-560943231.0/4294967296.0,1,-nbitq), 
to_sfixed(180159270.0/4294967296.0,1,-nbitq), 
to_sfixed(-39277108.0/4294967296.0,1,-nbitq), 
to_sfixed(-130639743.0/4294967296.0,1,-nbitq), 
to_sfixed(-234324248.0/4294967296.0,1,-nbitq), 
to_sfixed(459151219.0/4294967296.0,1,-nbitq), 
to_sfixed(-311995933.0/4294967296.0,1,-nbitq), 
to_sfixed(385941437.0/4294967296.0,1,-nbitq), 
to_sfixed(486177956.0/4294967296.0,1,-nbitq), 
to_sfixed(293852584.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-529879715.0/4294967296.0,1,-nbitq), 
to_sfixed(23584059.0/4294967296.0,1,-nbitq), 
to_sfixed(-781937881.0/4294967296.0,1,-nbitq), 
to_sfixed(-401599897.0/4294967296.0,1,-nbitq), 
to_sfixed(-330656306.0/4294967296.0,1,-nbitq), 
to_sfixed(76088939.0/4294967296.0,1,-nbitq), 
to_sfixed(-200533398.0/4294967296.0,1,-nbitq), 
to_sfixed(-426790051.0/4294967296.0,1,-nbitq), 
to_sfixed(-194840351.0/4294967296.0,1,-nbitq), 
to_sfixed(-31259506.0/4294967296.0,1,-nbitq), 
to_sfixed(-118084489.0/4294967296.0,1,-nbitq), 
to_sfixed(3263031.0/4294967296.0,1,-nbitq), 
to_sfixed(-183427006.0/4294967296.0,1,-nbitq), 
to_sfixed(843890363.0/4294967296.0,1,-nbitq), 
to_sfixed(266239541.0/4294967296.0,1,-nbitq), 
to_sfixed(222171415.0/4294967296.0,1,-nbitq), 
to_sfixed(190663576.0/4294967296.0,1,-nbitq), 
to_sfixed(-73344188.0/4294967296.0,1,-nbitq), 
to_sfixed(-1222243266.0/4294967296.0,1,-nbitq), 
to_sfixed(78781675.0/4294967296.0,1,-nbitq), 
to_sfixed(170353209.0/4294967296.0,1,-nbitq), 
to_sfixed(-635751177.0/4294967296.0,1,-nbitq), 
to_sfixed(-895081621.0/4294967296.0,1,-nbitq), 
to_sfixed(376076015.0/4294967296.0,1,-nbitq), 
to_sfixed(258930359.0/4294967296.0,1,-nbitq), 
to_sfixed(-826828161.0/4294967296.0,1,-nbitq), 
to_sfixed(340177379.0/4294967296.0,1,-nbitq), 
to_sfixed(433651262.0/4294967296.0,1,-nbitq), 
to_sfixed(-332138901.0/4294967296.0,1,-nbitq), 
to_sfixed(-412293689.0/4294967296.0,1,-nbitq), 
to_sfixed(509893973.0/4294967296.0,1,-nbitq), 
to_sfixed(-501501207.0/4294967296.0,1,-nbitq), 
to_sfixed(-634069094.0/4294967296.0,1,-nbitq), 
to_sfixed(-397195618.0/4294967296.0,1,-nbitq), 
to_sfixed(581802434.0/4294967296.0,1,-nbitq), 
to_sfixed(720249330.0/4294967296.0,1,-nbitq), 
to_sfixed(-75443998.0/4294967296.0,1,-nbitq), 
to_sfixed(486159290.0/4294967296.0,1,-nbitq), 
to_sfixed(96234991.0/4294967296.0,1,-nbitq), 
to_sfixed(27111943.0/4294967296.0,1,-nbitq), 
to_sfixed(334149273.0/4294967296.0,1,-nbitq), 
to_sfixed(97225443.0/4294967296.0,1,-nbitq), 
to_sfixed(-729431454.0/4294967296.0,1,-nbitq), 
to_sfixed(598718534.0/4294967296.0,1,-nbitq), 
to_sfixed(19119423.0/4294967296.0,1,-nbitq), 
to_sfixed(-24020955.0/4294967296.0,1,-nbitq), 
to_sfixed(135286231.0/4294967296.0,1,-nbitq), 
to_sfixed(-262904154.0/4294967296.0,1,-nbitq), 
to_sfixed(-46645477.0/4294967296.0,1,-nbitq), 
to_sfixed(-17451644.0/4294967296.0,1,-nbitq), 
to_sfixed(90548891.0/4294967296.0,1,-nbitq), 
to_sfixed(-101274331.0/4294967296.0,1,-nbitq), 
to_sfixed(298802920.0/4294967296.0,1,-nbitq), 
to_sfixed(-461775394.0/4294967296.0,1,-nbitq), 
to_sfixed(-739025703.0/4294967296.0,1,-nbitq), 
to_sfixed(357402290.0/4294967296.0,1,-nbitq), 
to_sfixed(366457433.0/4294967296.0,1,-nbitq), 
to_sfixed(-752646239.0/4294967296.0,1,-nbitq), 
to_sfixed(366838013.0/4294967296.0,1,-nbitq), 
to_sfixed(-355234172.0/4294967296.0,1,-nbitq), 
to_sfixed(-260511181.0/4294967296.0,1,-nbitq), 
to_sfixed(-550832486.0/4294967296.0,1,-nbitq), 
to_sfixed(-45220777.0/4294967296.0,1,-nbitq), 
to_sfixed(-101402859.0/4294967296.0,1,-nbitq), 
to_sfixed(533863535.0/4294967296.0,1,-nbitq), 
to_sfixed(235611896.0/4294967296.0,1,-nbitq), 
to_sfixed(58999655.0/4294967296.0,1,-nbitq), 
to_sfixed(-137952353.0/4294967296.0,1,-nbitq), 
to_sfixed(153359045.0/4294967296.0,1,-nbitq), 
to_sfixed(238403230.0/4294967296.0,1,-nbitq), 
to_sfixed(-62809716.0/4294967296.0,1,-nbitq), 
to_sfixed(-267137165.0/4294967296.0,1,-nbitq), 
to_sfixed(469804709.0/4294967296.0,1,-nbitq), 
to_sfixed(153823726.0/4294967296.0,1,-nbitq), 
to_sfixed(-260833351.0/4294967296.0,1,-nbitq), 
to_sfixed(619067400.0/4294967296.0,1,-nbitq), 
to_sfixed(-850603404.0/4294967296.0,1,-nbitq), 
to_sfixed(354305070.0/4294967296.0,1,-nbitq), 
to_sfixed(565223426.0/4294967296.0,1,-nbitq), 
to_sfixed(-80120439.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-85307950.0/4294967296.0,1,-nbitq), 
to_sfixed(-578673220.0/4294967296.0,1,-nbitq), 
to_sfixed(485083640.0/4294967296.0,1,-nbitq), 
to_sfixed(533854659.0/4294967296.0,1,-nbitq), 
to_sfixed(-630721583.0/4294967296.0,1,-nbitq), 
to_sfixed(250772645.0/4294967296.0,1,-nbitq), 
to_sfixed(227747901.0/4294967296.0,1,-nbitq), 
to_sfixed(-128837746.0/4294967296.0,1,-nbitq), 
to_sfixed(310439975.0/4294967296.0,1,-nbitq), 
to_sfixed(399599234.0/4294967296.0,1,-nbitq), 
to_sfixed(-412254185.0/4294967296.0,1,-nbitq), 
to_sfixed(625676056.0/4294967296.0,1,-nbitq), 
to_sfixed(-560460548.0/4294967296.0,1,-nbitq), 
to_sfixed(331095523.0/4294967296.0,1,-nbitq), 
to_sfixed(49813915.0/4294967296.0,1,-nbitq), 
to_sfixed(-29457688.0/4294967296.0,1,-nbitq), 
to_sfixed(-307140786.0/4294967296.0,1,-nbitq), 
to_sfixed(331825116.0/4294967296.0,1,-nbitq), 
to_sfixed(-877128368.0/4294967296.0,1,-nbitq), 
to_sfixed(230831982.0/4294967296.0,1,-nbitq), 
to_sfixed(-156365573.0/4294967296.0,1,-nbitq), 
to_sfixed(805323125.0/4294967296.0,1,-nbitq), 
to_sfixed(195363996.0/4294967296.0,1,-nbitq), 
to_sfixed(750754911.0/4294967296.0,1,-nbitq), 
to_sfixed(237733122.0/4294967296.0,1,-nbitq), 
to_sfixed(161662404.0/4294967296.0,1,-nbitq), 
to_sfixed(444014618.0/4294967296.0,1,-nbitq), 
to_sfixed(811162414.0/4294967296.0,1,-nbitq), 
to_sfixed(-430064304.0/4294967296.0,1,-nbitq), 
to_sfixed(-573979988.0/4294967296.0,1,-nbitq), 
to_sfixed(777499495.0/4294967296.0,1,-nbitq), 
to_sfixed(-141540957.0/4294967296.0,1,-nbitq), 
to_sfixed(-629497805.0/4294967296.0,1,-nbitq), 
to_sfixed(-257692285.0/4294967296.0,1,-nbitq), 
to_sfixed(1405161.0/4294967296.0,1,-nbitq), 
to_sfixed(601006567.0/4294967296.0,1,-nbitq), 
to_sfixed(17175909.0/4294967296.0,1,-nbitq), 
to_sfixed(112957327.0/4294967296.0,1,-nbitq), 
to_sfixed(496360624.0/4294967296.0,1,-nbitq), 
to_sfixed(-12697474.0/4294967296.0,1,-nbitq), 
to_sfixed(-248823661.0/4294967296.0,1,-nbitq), 
to_sfixed(572898446.0/4294967296.0,1,-nbitq), 
to_sfixed(42274938.0/4294967296.0,1,-nbitq), 
to_sfixed(235346302.0/4294967296.0,1,-nbitq), 
to_sfixed(338724436.0/4294967296.0,1,-nbitq), 
to_sfixed(81508708.0/4294967296.0,1,-nbitq), 
to_sfixed(10746297.0/4294967296.0,1,-nbitq), 
to_sfixed(-387613830.0/4294967296.0,1,-nbitq), 
to_sfixed(281129516.0/4294967296.0,1,-nbitq), 
to_sfixed(-271230321.0/4294967296.0,1,-nbitq), 
to_sfixed(-102798773.0/4294967296.0,1,-nbitq), 
to_sfixed(146278180.0/4294967296.0,1,-nbitq), 
to_sfixed(40039992.0/4294967296.0,1,-nbitq), 
to_sfixed(20534518.0/4294967296.0,1,-nbitq), 
to_sfixed(-1043479394.0/4294967296.0,1,-nbitq), 
to_sfixed(814790045.0/4294967296.0,1,-nbitq), 
to_sfixed(135661272.0/4294967296.0,1,-nbitq), 
to_sfixed(-1185372429.0/4294967296.0,1,-nbitq), 
to_sfixed(216491755.0/4294967296.0,1,-nbitq), 
to_sfixed(241168176.0/4294967296.0,1,-nbitq), 
to_sfixed(-107353259.0/4294967296.0,1,-nbitq), 
to_sfixed(-295410805.0/4294967296.0,1,-nbitq), 
to_sfixed(-137144506.0/4294967296.0,1,-nbitq), 
to_sfixed(-278118214.0/4294967296.0,1,-nbitq), 
to_sfixed(148947215.0/4294967296.0,1,-nbitq), 
to_sfixed(-336466169.0/4294967296.0,1,-nbitq), 
to_sfixed(272544901.0/4294967296.0,1,-nbitq), 
to_sfixed(156271242.0/4294967296.0,1,-nbitq), 
to_sfixed(255847868.0/4294967296.0,1,-nbitq), 
to_sfixed(-535814324.0/4294967296.0,1,-nbitq), 
to_sfixed(-427851567.0/4294967296.0,1,-nbitq), 
to_sfixed(24057121.0/4294967296.0,1,-nbitq), 
to_sfixed(50125035.0/4294967296.0,1,-nbitq), 
to_sfixed(-297132735.0/4294967296.0,1,-nbitq), 
to_sfixed(187418907.0/4294967296.0,1,-nbitq), 
to_sfixed(233725061.0/4294967296.0,1,-nbitq), 
to_sfixed(-171582097.0/4294967296.0,1,-nbitq), 
to_sfixed(514910365.0/4294967296.0,1,-nbitq), 
to_sfixed(338129159.0/4294967296.0,1,-nbitq), 
to_sfixed(28699729.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-224606294.0/4294967296.0,1,-nbitq), 
to_sfixed(-463502192.0/4294967296.0,1,-nbitq), 
to_sfixed(351278273.0/4294967296.0,1,-nbitq), 
to_sfixed(95953444.0/4294967296.0,1,-nbitq), 
to_sfixed(-490295061.0/4294967296.0,1,-nbitq), 
to_sfixed(151874917.0/4294967296.0,1,-nbitq), 
to_sfixed(-179538998.0/4294967296.0,1,-nbitq), 
to_sfixed(726011781.0/4294967296.0,1,-nbitq), 
to_sfixed(-94845993.0/4294967296.0,1,-nbitq), 
to_sfixed(-126203923.0/4294967296.0,1,-nbitq), 
to_sfixed(454725929.0/4294967296.0,1,-nbitq), 
to_sfixed(937153749.0/4294967296.0,1,-nbitq), 
to_sfixed(-188211515.0/4294967296.0,1,-nbitq), 
to_sfixed(-554040080.0/4294967296.0,1,-nbitq), 
to_sfixed(-260673649.0/4294967296.0,1,-nbitq), 
to_sfixed(-258455749.0/4294967296.0,1,-nbitq), 
to_sfixed(198173637.0/4294967296.0,1,-nbitq), 
to_sfixed(293438314.0/4294967296.0,1,-nbitq), 
to_sfixed(-831480234.0/4294967296.0,1,-nbitq), 
to_sfixed(102711948.0/4294967296.0,1,-nbitq), 
to_sfixed(-142062693.0/4294967296.0,1,-nbitq), 
to_sfixed(467562126.0/4294967296.0,1,-nbitq), 
to_sfixed(70839684.0/4294967296.0,1,-nbitq), 
to_sfixed(433552086.0/4294967296.0,1,-nbitq), 
to_sfixed(219471623.0/4294967296.0,1,-nbitq), 
to_sfixed(-670866282.0/4294967296.0,1,-nbitq), 
to_sfixed(614525370.0/4294967296.0,1,-nbitq), 
to_sfixed(507358756.0/4294967296.0,1,-nbitq), 
to_sfixed(-187747623.0/4294967296.0,1,-nbitq), 
to_sfixed(-493153845.0/4294967296.0,1,-nbitq), 
to_sfixed(773488741.0/4294967296.0,1,-nbitq), 
to_sfixed(-112935494.0/4294967296.0,1,-nbitq), 
to_sfixed(-208495222.0/4294967296.0,1,-nbitq), 
to_sfixed(45383013.0/4294967296.0,1,-nbitq), 
to_sfixed(-267474609.0/4294967296.0,1,-nbitq), 
to_sfixed(431796274.0/4294967296.0,1,-nbitq), 
to_sfixed(-212845822.0/4294967296.0,1,-nbitq), 
to_sfixed(-549708724.0/4294967296.0,1,-nbitq), 
to_sfixed(147188681.0/4294967296.0,1,-nbitq), 
to_sfixed(-97333680.0/4294967296.0,1,-nbitq), 
to_sfixed(-76824959.0/4294967296.0,1,-nbitq), 
to_sfixed(557326861.0/4294967296.0,1,-nbitq), 
to_sfixed(-123374137.0/4294967296.0,1,-nbitq), 
to_sfixed(15727820.0/4294967296.0,1,-nbitq), 
to_sfixed(332493163.0/4294967296.0,1,-nbitq), 
to_sfixed(-141375531.0/4294967296.0,1,-nbitq), 
to_sfixed(81075873.0/4294967296.0,1,-nbitq), 
to_sfixed(-143862435.0/4294967296.0,1,-nbitq), 
to_sfixed(382983678.0/4294967296.0,1,-nbitq), 
to_sfixed(-970564708.0/4294967296.0,1,-nbitq), 
to_sfixed(494906355.0/4294967296.0,1,-nbitq), 
to_sfixed(-178588702.0/4294967296.0,1,-nbitq), 
to_sfixed(-563803440.0/4294967296.0,1,-nbitq), 
to_sfixed(27958416.0/4294967296.0,1,-nbitq), 
to_sfixed(-1185729686.0/4294967296.0,1,-nbitq), 
to_sfixed(213782436.0/4294967296.0,1,-nbitq), 
to_sfixed(43109690.0/4294967296.0,1,-nbitq), 
to_sfixed(-510380318.0/4294967296.0,1,-nbitq), 
to_sfixed(91065774.0/4294967296.0,1,-nbitq), 
to_sfixed(299508426.0/4294967296.0,1,-nbitq), 
to_sfixed(-340405885.0/4294967296.0,1,-nbitq), 
to_sfixed(-154283751.0/4294967296.0,1,-nbitq), 
to_sfixed(-11002161.0/4294967296.0,1,-nbitq), 
to_sfixed(-431519188.0/4294967296.0,1,-nbitq), 
to_sfixed(-250214245.0/4294967296.0,1,-nbitq), 
to_sfixed(-93385913.0/4294967296.0,1,-nbitq), 
to_sfixed(-231319292.0/4294967296.0,1,-nbitq), 
to_sfixed(-157636953.0/4294967296.0,1,-nbitq), 
to_sfixed(101656466.0/4294967296.0,1,-nbitq), 
to_sfixed(-416296428.0/4294967296.0,1,-nbitq), 
to_sfixed(-442634127.0/4294967296.0,1,-nbitq), 
to_sfixed(293896603.0/4294967296.0,1,-nbitq), 
to_sfixed(282900873.0/4294967296.0,1,-nbitq), 
to_sfixed(-64135534.0/4294967296.0,1,-nbitq), 
to_sfixed(163347086.0/4294967296.0,1,-nbitq), 
to_sfixed(54976546.0/4294967296.0,1,-nbitq), 
to_sfixed(53739353.0/4294967296.0,1,-nbitq), 
to_sfixed(420616190.0/4294967296.0,1,-nbitq), 
to_sfixed(28630314.0/4294967296.0,1,-nbitq), 
to_sfixed(-359024248.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-126781972.0/4294967296.0,1,-nbitq), 
to_sfixed(-40555723.0/4294967296.0,1,-nbitq), 
to_sfixed(1093377350.0/4294967296.0,1,-nbitq), 
to_sfixed(-224692691.0/4294967296.0,1,-nbitq), 
to_sfixed(80323138.0/4294967296.0,1,-nbitq), 
to_sfixed(-340325640.0/4294967296.0,1,-nbitq), 
to_sfixed(-271411477.0/4294967296.0,1,-nbitq), 
to_sfixed(61443072.0/4294967296.0,1,-nbitq), 
to_sfixed(-197382153.0/4294967296.0,1,-nbitq), 
to_sfixed(301417454.0/4294967296.0,1,-nbitq), 
to_sfixed(-195840962.0/4294967296.0,1,-nbitq), 
to_sfixed(109933315.0/4294967296.0,1,-nbitq), 
to_sfixed(-699975059.0/4294967296.0,1,-nbitq), 
to_sfixed(523221973.0/4294967296.0,1,-nbitq), 
to_sfixed(-343241418.0/4294967296.0,1,-nbitq), 
to_sfixed(521737144.0/4294967296.0,1,-nbitq), 
to_sfixed(-109352235.0/4294967296.0,1,-nbitq), 
to_sfixed(234258718.0/4294967296.0,1,-nbitq), 
to_sfixed(-130349531.0/4294967296.0,1,-nbitq), 
to_sfixed(-319505946.0/4294967296.0,1,-nbitq), 
to_sfixed(-85663590.0/4294967296.0,1,-nbitq), 
to_sfixed(232778780.0/4294967296.0,1,-nbitq), 
to_sfixed(-120557150.0/4294967296.0,1,-nbitq), 
to_sfixed(426635998.0/4294967296.0,1,-nbitq), 
to_sfixed(-301906633.0/4294967296.0,1,-nbitq), 
to_sfixed(-158726738.0/4294967296.0,1,-nbitq), 
to_sfixed(402404887.0/4294967296.0,1,-nbitq), 
to_sfixed(-35468411.0/4294967296.0,1,-nbitq), 
to_sfixed(-7869124.0/4294967296.0,1,-nbitq), 
to_sfixed(136068861.0/4294967296.0,1,-nbitq), 
to_sfixed(467732518.0/4294967296.0,1,-nbitq), 
to_sfixed(-35887505.0/4294967296.0,1,-nbitq), 
to_sfixed(51908451.0/4294967296.0,1,-nbitq), 
to_sfixed(-289391037.0/4294967296.0,1,-nbitq), 
to_sfixed(-405771576.0/4294967296.0,1,-nbitq), 
to_sfixed(-401556158.0/4294967296.0,1,-nbitq), 
to_sfixed(385175929.0/4294967296.0,1,-nbitq), 
to_sfixed(-294663795.0/4294967296.0,1,-nbitq), 
to_sfixed(393861180.0/4294967296.0,1,-nbitq), 
to_sfixed(283843004.0/4294967296.0,1,-nbitq), 
to_sfixed(-302922434.0/4294967296.0,1,-nbitq), 
to_sfixed(435261887.0/4294967296.0,1,-nbitq), 
to_sfixed(207739398.0/4294967296.0,1,-nbitq), 
to_sfixed(241156004.0/4294967296.0,1,-nbitq), 
to_sfixed(63065343.0/4294967296.0,1,-nbitq), 
to_sfixed(-127155856.0/4294967296.0,1,-nbitq), 
to_sfixed(166160057.0/4294967296.0,1,-nbitq), 
to_sfixed(-133732663.0/4294967296.0,1,-nbitq), 
to_sfixed(209672725.0/4294967296.0,1,-nbitq), 
to_sfixed(-872369330.0/4294967296.0,1,-nbitq), 
to_sfixed(-209463465.0/4294967296.0,1,-nbitq), 
to_sfixed(317795596.0/4294967296.0,1,-nbitq), 
to_sfixed(-68663328.0/4294967296.0,1,-nbitq), 
to_sfixed(-284606905.0/4294967296.0,1,-nbitq), 
to_sfixed(-560351886.0/4294967296.0,1,-nbitq), 
to_sfixed(316734522.0/4294967296.0,1,-nbitq), 
to_sfixed(211907479.0/4294967296.0,1,-nbitq), 
to_sfixed(-173881878.0/4294967296.0,1,-nbitq), 
to_sfixed(-276039507.0/4294967296.0,1,-nbitq), 
to_sfixed(123136017.0/4294967296.0,1,-nbitq), 
to_sfixed(64820769.0/4294967296.0,1,-nbitq), 
to_sfixed(3934461.0/4294967296.0,1,-nbitq), 
to_sfixed(-10286051.0/4294967296.0,1,-nbitq), 
to_sfixed(-245095550.0/4294967296.0,1,-nbitq), 
to_sfixed(-43219999.0/4294967296.0,1,-nbitq), 
to_sfixed(-202468399.0/4294967296.0,1,-nbitq), 
to_sfixed(538417893.0/4294967296.0,1,-nbitq), 
to_sfixed(-332165948.0/4294967296.0,1,-nbitq), 
to_sfixed(341932721.0/4294967296.0,1,-nbitq), 
to_sfixed(458971684.0/4294967296.0,1,-nbitq), 
to_sfixed(83497140.0/4294967296.0,1,-nbitq), 
to_sfixed(-106703138.0/4294967296.0,1,-nbitq), 
to_sfixed(-308474896.0/4294967296.0,1,-nbitq), 
to_sfixed(247230144.0/4294967296.0,1,-nbitq), 
to_sfixed(234544798.0/4294967296.0,1,-nbitq), 
to_sfixed(-42070176.0/4294967296.0,1,-nbitq), 
to_sfixed(-41630129.0/4294967296.0,1,-nbitq), 
to_sfixed(-101432251.0/4294967296.0,1,-nbitq), 
to_sfixed(205854894.0/4294967296.0,1,-nbitq), 
to_sfixed(60118204.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-175123583.0/4294967296.0,1,-nbitq), 
to_sfixed(-5146816.0/4294967296.0,1,-nbitq), 
to_sfixed(1207051960.0/4294967296.0,1,-nbitq), 
to_sfixed(-306341333.0/4294967296.0,1,-nbitq), 
to_sfixed(-445553039.0/4294967296.0,1,-nbitq), 
to_sfixed(-675898086.0/4294967296.0,1,-nbitq), 
to_sfixed(-283011243.0/4294967296.0,1,-nbitq), 
to_sfixed(508479821.0/4294967296.0,1,-nbitq), 
to_sfixed(306415573.0/4294967296.0,1,-nbitq), 
to_sfixed(281906494.0/4294967296.0,1,-nbitq), 
to_sfixed(472312721.0/4294967296.0,1,-nbitq), 
to_sfixed(162212654.0/4294967296.0,1,-nbitq), 
to_sfixed(261784689.0/4294967296.0,1,-nbitq), 
to_sfixed(178484860.0/4294967296.0,1,-nbitq), 
to_sfixed(34392943.0/4294967296.0,1,-nbitq), 
to_sfixed(26767648.0/4294967296.0,1,-nbitq), 
to_sfixed(202942014.0/4294967296.0,1,-nbitq), 
to_sfixed(-321547919.0/4294967296.0,1,-nbitq), 
to_sfixed(-125935139.0/4294967296.0,1,-nbitq), 
to_sfixed(57028848.0/4294967296.0,1,-nbitq), 
to_sfixed(193184153.0/4294967296.0,1,-nbitq), 
to_sfixed(332597538.0/4294967296.0,1,-nbitq), 
to_sfixed(-257384034.0/4294967296.0,1,-nbitq), 
to_sfixed(166701222.0/4294967296.0,1,-nbitq), 
to_sfixed(-274926392.0/4294967296.0,1,-nbitq), 
to_sfixed(-228062510.0/4294967296.0,1,-nbitq), 
to_sfixed(-75432078.0/4294967296.0,1,-nbitq), 
to_sfixed(119365065.0/4294967296.0,1,-nbitq), 
to_sfixed(546538918.0/4294967296.0,1,-nbitq), 
to_sfixed(253476168.0/4294967296.0,1,-nbitq), 
to_sfixed(-69328089.0/4294967296.0,1,-nbitq), 
to_sfixed(-439003970.0/4294967296.0,1,-nbitq), 
to_sfixed(248754329.0/4294967296.0,1,-nbitq), 
to_sfixed(-281198081.0/4294967296.0,1,-nbitq), 
to_sfixed(-50964381.0/4294967296.0,1,-nbitq), 
to_sfixed(-473626356.0/4294967296.0,1,-nbitq), 
to_sfixed(-18921557.0/4294967296.0,1,-nbitq), 
to_sfixed(-445482452.0/4294967296.0,1,-nbitq), 
to_sfixed(67789036.0/4294967296.0,1,-nbitq), 
to_sfixed(280570076.0/4294967296.0,1,-nbitq), 
to_sfixed(-376363529.0/4294967296.0,1,-nbitq), 
to_sfixed(-8091318.0/4294967296.0,1,-nbitq), 
to_sfixed(241176631.0/4294967296.0,1,-nbitq), 
to_sfixed(34547463.0/4294967296.0,1,-nbitq), 
to_sfixed(289350047.0/4294967296.0,1,-nbitq), 
to_sfixed(-87040319.0/4294967296.0,1,-nbitq), 
to_sfixed(26771832.0/4294967296.0,1,-nbitq), 
to_sfixed(-359941366.0/4294967296.0,1,-nbitq), 
to_sfixed(-13685313.0/4294967296.0,1,-nbitq), 
to_sfixed(-75200570.0/4294967296.0,1,-nbitq), 
to_sfixed(-145969582.0/4294967296.0,1,-nbitq), 
to_sfixed(351452160.0/4294967296.0,1,-nbitq), 
to_sfixed(168259240.0/4294967296.0,1,-nbitq), 
to_sfixed(122874548.0/4294967296.0,1,-nbitq), 
to_sfixed(-17450110.0/4294967296.0,1,-nbitq), 
to_sfixed(211293130.0/4294967296.0,1,-nbitq), 
to_sfixed(237351881.0/4294967296.0,1,-nbitq), 
to_sfixed(-375674210.0/4294967296.0,1,-nbitq), 
to_sfixed(127007200.0/4294967296.0,1,-nbitq), 
to_sfixed(427140371.0/4294967296.0,1,-nbitq), 
to_sfixed(-323222240.0/4294967296.0,1,-nbitq), 
to_sfixed(-221806461.0/4294967296.0,1,-nbitq), 
to_sfixed(-248784486.0/4294967296.0,1,-nbitq), 
to_sfixed(-263563291.0/4294967296.0,1,-nbitq), 
to_sfixed(54008620.0/4294967296.0,1,-nbitq), 
to_sfixed(344942454.0/4294967296.0,1,-nbitq), 
to_sfixed(457929655.0/4294967296.0,1,-nbitq), 
to_sfixed(-308195896.0/4294967296.0,1,-nbitq), 
to_sfixed(-3680760.0/4294967296.0,1,-nbitq), 
to_sfixed(628967606.0/4294967296.0,1,-nbitq), 
to_sfixed(-2895030.0/4294967296.0,1,-nbitq), 
to_sfixed(172250065.0/4294967296.0,1,-nbitq), 
to_sfixed(-64543797.0/4294967296.0,1,-nbitq), 
to_sfixed(150541008.0/4294967296.0,1,-nbitq), 
to_sfixed(323592622.0/4294967296.0,1,-nbitq), 
to_sfixed(253500844.0/4294967296.0,1,-nbitq), 
to_sfixed(68744070.0/4294967296.0,1,-nbitq), 
to_sfixed(51225904.0/4294967296.0,1,-nbitq), 
to_sfixed(-25487997.0/4294967296.0,1,-nbitq), 
to_sfixed(-101199156.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(383459414.0/4294967296.0,1,-nbitq), 
to_sfixed(-265183694.0/4294967296.0,1,-nbitq), 
to_sfixed(775435325.0/4294967296.0,1,-nbitq), 
to_sfixed(205723082.0/4294967296.0,1,-nbitq), 
to_sfixed(219685679.0/4294967296.0,1,-nbitq), 
to_sfixed(-535830189.0/4294967296.0,1,-nbitq), 
to_sfixed(-10394036.0/4294967296.0,1,-nbitq), 
to_sfixed(55476564.0/4294967296.0,1,-nbitq), 
to_sfixed(289144330.0/4294967296.0,1,-nbitq), 
to_sfixed(-33477359.0/4294967296.0,1,-nbitq), 
to_sfixed(107221916.0/4294967296.0,1,-nbitq), 
to_sfixed(40409417.0/4294967296.0,1,-nbitq), 
to_sfixed(-423055569.0/4294967296.0,1,-nbitq), 
to_sfixed(129134693.0/4294967296.0,1,-nbitq), 
to_sfixed(-40282098.0/4294967296.0,1,-nbitq), 
to_sfixed(360975757.0/4294967296.0,1,-nbitq), 
to_sfixed(91844611.0/4294967296.0,1,-nbitq), 
to_sfixed(-165627354.0/4294967296.0,1,-nbitq), 
to_sfixed(-111342758.0/4294967296.0,1,-nbitq), 
to_sfixed(-309164886.0/4294967296.0,1,-nbitq), 
to_sfixed(-247895866.0/4294967296.0,1,-nbitq), 
to_sfixed(-178323685.0/4294967296.0,1,-nbitq), 
to_sfixed(-4910105.0/4294967296.0,1,-nbitq), 
to_sfixed(-55676973.0/4294967296.0,1,-nbitq), 
to_sfixed(104200852.0/4294967296.0,1,-nbitq), 
to_sfixed(184941529.0/4294967296.0,1,-nbitq), 
to_sfixed(72342114.0/4294967296.0,1,-nbitq), 
to_sfixed(202475821.0/4294967296.0,1,-nbitq), 
to_sfixed(553281692.0/4294967296.0,1,-nbitq), 
to_sfixed(-149298472.0/4294967296.0,1,-nbitq), 
to_sfixed(-91539677.0/4294967296.0,1,-nbitq), 
to_sfixed(-51521858.0/4294967296.0,1,-nbitq), 
to_sfixed(-198586791.0/4294967296.0,1,-nbitq), 
to_sfixed(-165403379.0/4294967296.0,1,-nbitq), 
to_sfixed(24494779.0/4294967296.0,1,-nbitq), 
to_sfixed(-185343701.0/4294967296.0,1,-nbitq), 
to_sfixed(-228441327.0/4294967296.0,1,-nbitq), 
to_sfixed(151102702.0/4294967296.0,1,-nbitq), 
to_sfixed(103850919.0/4294967296.0,1,-nbitq), 
to_sfixed(41033348.0/4294967296.0,1,-nbitq), 
to_sfixed(-328479578.0/4294967296.0,1,-nbitq), 
to_sfixed(-362931500.0/4294967296.0,1,-nbitq), 
to_sfixed(21747136.0/4294967296.0,1,-nbitq), 
to_sfixed(-133498619.0/4294967296.0,1,-nbitq), 
to_sfixed(224622262.0/4294967296.0,1,-nbitq), 
to_sfixed(-378112543.0/4294967296.0,1,-nbitq), 
to_sfixed(123553487.0/4294967296.0,1,-nbitq), 
to_sfixed(-75441648.0/4294967296.0,1,-nbitq), 
to_sfixed(135514171.0/4294967296.0,1,-nbitq), 
to_sfixed(-105982918.0/4294967296.0,1,-nbitq), 
to_sfixed(65696765.0/4294967296.0,1,-nbitq), 
to_sfixed(-305339593.0/4294967296.0,1,-nbitq), 
to_sfixed(-351509307.0/4294967296.0,1,-nbitq), 
to_sfixed(-292409570.0/4294967296.0,1,-nbitq), 
to_sfixed(-62780727.0/4294967296.0,1,-nbitq), 
to_sfixed(-361260071.0/4294967296.0,1,-nbitq), 
to_sfixed(-276411488.0/4294967296.0,1,-nbitq), 
to_sfixed(-125415519.0/4294967296.0,1,-nbitq), 
to_sfixed(160210776.0/4294967296.0,1,-nbitq), 
to_sfixed(353848090.0/4294967296.0,1,-nbitq), 
to_sfixed(-3031056.0/4294967296.0,1,-nbitq), 
to_sfixed(154750337.0/4294967296.0,1,-nbitq), 
to_sfixed(-236694809.0/4294967296.0,1,-nbitq), 
to_sfixed(353319865.0/4294967296.0,1,-nbitq), 
to_sfixed(-263512455.0/4294967296.0,1,-nbitq), 
to_sfixed(73442737.0/4294967296.0,1,-nbitq), 
to_sfixed(433516874.0/4294967296.0,1,-nbitq), 
to_sfixed(-264036962.0/4294967296.0,1,-nbitq), 
to_sfixed(-316307647.0/4294967296.0,1,-nbitq), 
to_sfixed(529764899.0/4294967296.0,1,-nbitq), 
to_sfixed(55743101.0/4294967296.0,1,-nbitq), 
to_sfixed(358655898.0/4294967296.0,1,-nbitq), 
to_sfixed(185248006.0/4294967296.0,1,-nbitq), 
to_sfixed(-95581218.0/4294967296.0,1,-nbitq), 
to_sfixed(177819332.0/4294967296.0,1,-nbitq), 
to_sfixed(40873227.0/4294967296.0,1,-nbitq), 
to_sfixed(-61170994.0/4294967296.0,1,-nbitq), 
to_sfixed(-164901729.0/4294967296.0,1,-nbitq), 
to_sfixed(-233009290.0/4294967296.0,1,-nbitq), 
to_sfixed(372219487.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-27761352.0/4294967296.0,1,-nbitq), 
to_sfixed(238382307.0/4294967296.0,1,-nbitq), 
to_sfixed(-112477338.0/4294967296.0,1,-nbitq), 
to_sfixed(-366267328.0/4294967296.0,1,-nbitq), 
to_sfixed(135454452.0/4294967296.0,1,-nbitq), 
to_sfixed(-37451240.0/4294967296.0,1,-nbitq), 
to_sfixed(-6481827.0/4294967296.0,1,-nbitq), 
to_sfixed(-400072928.0/4294967296.0,1,-nbitq), 
to_sfixed(-182298652.0/4294967296.0,1,-nbitq), 
to_sfixed(356924106.0/4294967296.0,1,-nbitq), 
to_sfixed(-367646880.0/4294967296.0,1,-nbitq), 
to_sfixed(-285754058.0/4294967296.0,1,-nbitq), 
to_sfixed(-292943667.0/4294967296.0,1,-nbitq), 
to_sfixed(203851351.0/4294967296.0,1,-nbitq), 
to_sfixed(-59835472.0/4294967296.0,1,-nbitq), 
to_sfixed(47695368.0/4294967296.0,1,-nbitq), 
to_sfixed(347282404.0/4294967296.0,1,-nbitq), 
to_sfixed(193766686.0/4294967296.0,1,-nbitq), 
to_sfixed(408401236.0/4294967296.0,1,-nbitq), 
to_sfixed(52672485.0/4294967296.0,1,-nbitq), 
to_sfixed(-169150496.0/4294967296.0,1,-nbitq), 
to_sfixed(-172376226.0/4294967296.0,1,-nbitq), 
to_sfixed(-94565829.0/4294967296.0,1,-nbitq), 
to_sfixed(-290778281.0/4294967296.0,1,-nbitq), 
to_sfixed(-274151266.0/4294967296.0,1,-nbitq), 
to_sfixed(94855502.0/4294967296.0,1,-nbitq), 
to_sfixed(22514967.0/4294967296.0,1,-nbitq), 
to_sfixed(-404912704.0/4294967296.0,1,-nbitq), 
to_sfixed(-351103941.0/4294967296.0,1,-nbitq), 
to_sfixed(-87264384.0/4294967296.0,1,-nbitq), 
to_sfixed(-379910569.0/4294967296.0,1,-nbitq), 
to_sfixed(-72824218.0/4294967296.0,1,-nbitq), 
to_sfixed(-264281865.0/4294967296.0,1,-nbitq), 
to_sfixed(-318806502.0/4294967296.0,1,-nbitq), 
to_sfixed(-178919075.0/4294967296.0,1,-nbitq), 
to_sfixed(-156519040.0/4294967296.0,1,-nbitq), 
to_sfixed(33661023.0/4294967296.0,1,-nbitq), 
to_sfixed(-230146024.0/4294967296.0,1,-nbitq), 
to_sfixed(136580857.0/4294967296.0,1,-nbitq), 
to_sfixed(400675201.0/4294967296.0,1,-nbitq), 
to_sfixed(-146126746.0/4294967296.0,1,-nbitq), 
to_sfixed(-149158872.0/4294967296.0,1,-nbitq), 
to_sfixed(197055156.0/4294967296.0,1,-nbitq), 
to_sfixed(-394216887.0/4294967296.0,1,-nbitq), 
to_sfixed(120730229.0/4294967296.0,1,-nbitq), 
to_sfixed(211653508.0/4294967296.0,1,-nbitq), 
to_sfixed(91026509.0/4294967296.0,1,-nbitq), 
to_sfixed(-176950635.0/4294967296.0,1,-nbitq), 
to_sfixed(-353804382.0/4294967296.0,1,-nbitq), 
to_sfixed(531373865.0/4294967296.0,1,-nbitq), 
to_sfixed(124652393.0/4294967296.0,1,-nbitq), 
to_sfixed(-301461313.0/4294967296.0,1,-nbitq), 
to_sfixed(209033531.0/4294967296.0,1,-nbitq), 
to_sfixed(355919816.0/4294967296.0,1,-nbitq), 
to_sfixed(70667413.0/4294967296.0,1,-nbitq), 
to_sfixed(155521170.0/4294967296.0,1,-nbitq), 
to_sfixed(-255852203.0/4294967296.0,1,-nbitq), 
to_sfixed(76764223.0/4294967296.0,1,-nbitq), 
to_sfixed(439337512.0/4294967296.0,1,-nbitq), 
to_sfixed(-195170328.0/4294967296.0,1,-nbitq), 
to_sfixed(-397168257.0/4294967296.0,1,-nbitq), 
to_sfixed(503846781.0/4294967296.0,1,-nbitq), 
to_sfixed(270071688.0/4294967296.0,1,-nbitq), 
to_sfixed(29864854.0/4294967296.0,1,-nbitq), 
to_sfixed(172901698.0/4294967296.0,1,-nbitq), 
to_sfixed(-116152108.0/4294967296.0,1,-nbitq), 
to_sfixed(866799050.0/4294967296.0,1,-nbitq), 
to_sfixed(53459540.0/4294967296.0,1,-nbitq), 
to_sfixed(-291938718.0/4294967296.0,1,-nbitq), 
to_sfixed(492196532.0/4294967296.0,1,-nbitq), 
to_sfixed(273011175.0/4294967296.0,1,-nbitq), 
to_sfixed(-130102375.0/4294967296.0,1,-nbitq), 
to_sfixed(-312842561.0/4294967296.0,1,-nbitq), 
to_sfixed(219452279.0/4294967296.0,1,-nbitq), 
to_sfixed(26494.0/4294967296.0,1,-nbitq), 
to_sfixed(-451131435.0/4294967296.0,1,-nbitq), 
to_sfixed(-429278551.0/4294967296.0,1,-nbitq), 
to_sfixed(-174119085.0/4294967296.0,1,-nbitq), 
to_sfixed(-298193588.0/4294967296.0,1,-nbitq), 
to_sfixed(-61568207.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-275915401.0/4294967296.0,1,-nbitq), 
to_sfixed(-204970883.0/4294967296.0,1,-nbitq), 
to_sfixed(277511757.0/4294967296.0,1,-nbitq), 
to_sfixed(-157231153.0/4294967296.0,1,-nbitq), 
to_sfixed(155936085.0/4294967296.0,1,-nbitq), 
to_sfixed(169183489.0/4294967296.0,1,-nbitq), 
to_sfixed(-344156331.0/4294967296.0,1,-nbitq), 
to_sfixed(-202827370.0/4294967296.0,1,-nbitq), 
to_sfixed(184335575.0/4294967296.0,1,-nbitq), 
to_sfixed(-144426198.0/4294967296.0,1,-nbitq), 
to_sfixed(-352027306.0/4294967296.0,1,-nbitq), 
to_sfixed(261741751.0/4294967296.0,1,-nbitq), 
to_sfixed(-352405392.0/4294967296.0,1,-nbitq), 
to_sfixed(-110776481.0/4294967296.0,1,-nbitq), 
to_sfixed(-381448615.0/4294967296.0,1,-nbitq), 
to_sfixed(256240640.0/4294967296.0,1,-nbitq), 
to_sfixed(105456392.0/4294967296.0,1,-nbitq), 
to_sfixed(-9120180.0/4294967296.0,1,-nbitq), 
to_sfixed(408192896.0/4294967296.0,1,-nbitq), 
to_sfixed(309437507.0/4294967296.0,1,-nbitq), 
to_sfixed(-226054256.0/4294967296.0,1,-nbitq), 
to_sfixed(-157732933.0/4294967296.0,1,-nbitq), 
to_sfixed(320303344.0/4294967296.0,1,-nbitq), 
to_sfixed(-23855574.0/4294967296.0,1,-nbitq), 
to_sfixed(-337858961.0/4294967296.0,1,-nbitq), 
to_sfixed(61623047.0/4294967296.0,1,-nbitq), 
to_sfixed(-155952290.0/4294967296.0,1,-nbitq), 
to_sfixed(-328689887.0/4294967296.0,1,-nbitq), 
to_sfixed(181205883.0/4294967296.0,1,-nbitq), 
to_sfixed(314810311.0/4294967296.0,1,-nbitq), 
to_sfixed(-472820791.0/4294967296.0,1,-nbitq), 
to_sfixed(-151310276.0/4294967296.0,1,-nbitq), 
to_sfixed(161857572.0/4294967296.0,1,-nbitq), 
to_sfixed(-286521836.0/4294967296.0,1,-nbitq), 
to_sfixed(423738813.0/4294967296.0,1,-nbitq), 
to_sfixed(-260178099.0/4294967296.0,1,-nbitq), 
to_sfixed(386923782.0/4294967296.0,1,-nbitq), 
to_sfixed(473959773.0/4294967296.0,1,-nbitq), 
to_sfixed(170974478.0/4294967296.0,1,-nbitq), 
to_sfixed(-71458113.0/4294967296.0,1,-nbitq), 
to_sfixed(-110629635.0/4294967296.0,1,-nbitq), 
to_sfixed(-152007037.0/4294967296.0,1,-nbitq), 
to_sfixed(406405817.0/4294967296.0,1,-nbitq), 
to_sfixed(435564783.0/4294967296.0,1,-nbitq), 
to_sfixed(-224365496.0/4294967296.0,1,-nbitq), 
to_sfixed(243582612.0/4294967296.0,1,-nbitq), 
to_sfixed(80530257.0/4294967296.0,1,-nbitq), 
to_sfixed(-460100665.0/4294967296.0,1,-nbitq), 
to_sfixed(23400782.0/4294967296.0,1,-nbitq), 
to_sfixed(223814545.0/4294967296.0,1,-nbitq), 
to_sfixed(-163689069.0/4294967296.0,1,-nbitq), 
to_sfixed(143567051.0/4294967296.0,1,-nbitq), 
to_sfixed(-294061552.0/4294967296.0,1,-nbitq), 
to_sfixed(149992034.0/4294967296.0,1,-nbitq), 
to_sfixed(611158786.0/4294967296.0,1,-nbitq), 
to_sfixed(230118921.0/4294967296.0,1,-nbitq), 
to_sfixed(-49448165.0/4294967296.0,1,-nbitq), 
to_sfixed(-33804573.0/4294967296.0,1,-nbitq), 
to_sfixed(-101997288.0/4294967296.0,1,-nbitq), 
to_sfixed(73275045.0/4294967296.0,1,-nbitq), 
to_sfixed(354227886.0/4294967296.0,1,-nbitq), 
to_sfixed(186487766.0/4294967296.0,1,-nbitq), 
to_sfixed(365750109.0/4294967296.0,1,-nbitq), 
to_sfixed(366063042.0/4294967296.0,1,-nbitq), 
to_sfixed(-140116346.0/4294967296.0,1,-nbitq), 
to_sfixed(295683719.0/4294967296.0,1,-nbitq), 
to_sfixed(644889562.0/4294967296.0,1,-nbitq), 
to_sfixed(-147469958.0/4294967296.0,1,-nbitq), 
to_sfixed(-27981230.0/4294967296.0,1,-nbitq), 
to_sfixed(-54313356.0/4294967296.0,1,-nbitq), 
to_sfixed(-444464566.0/4294967296.0,1,-nbitq), 
to_sfixed(-188411329.0/4294967296.0,1,-nbitq), 
to_sfixed(-16453039.0/4294967296.0,1,-nbitq), 
to_sfixed(-257532460.0/4294967296.0,1,-nbitq), 
to_sfixed(466879901.0/4294967296.0,1,-nbitq), 
to_sfixed(-234696589.0/4294967296.0,1,-nbitq), 
to_sfixed(81831868.0/4294967296.0,1,-nbitq), 
to_sfixed(-294156418.0/4294967296.0,1,-nbitq), 
to_sfixed(-348524606.0/4294967296.0,1,-nbitq), 
to_sfixed(81738221.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-322473792.0/4294967296.0,1,-nbitq), 
to_sfixed(-127155786.0/4294967296.0,1,-nbitq), 
to_sfixed(66651553.0/4294967296.0,1,-nbitq), 
to_sfixed(444193441.0/4294967296.0,1,-nbitq), 
to_sfixed(575179319.0/4294967296.0,1,-nbitq), 
to_sfixed(-170138251.0/4294967296.0,1,-nbitq), 
to_sfixed(-116207192.0/4294967296.0,1,-nbitq), 
to_sfixed(-301235820.0/4294967296.0,1,-nbitq), 
to_sfixed(323972909.0/4294967296.0,1,-nbitq), 
to_sfixed(196413764.0/4294967296.0,1,-nbitq), 
to_sfixed(-275555197.0/4294967296.0,1,-nbitq), 
to_sfixed(379019396.0/4294967296.0,1,-nbitq), 
to_sfixed(326175887.0/4294967296.0,1,-nbitq), 
to_sfixed(360625550.0/4294967296.0,1,-nbitq), 
to_sfixed(95233282.0/4294967296.0,1,-nbitq), 
to_sfixed(267673674.0/4294967296.0,1,-nbitq), 
to_sfixed(-351584459.0/4294967296.0,1,-nbitq), 
to_sfixed(-83599848.0/4294967296.0,1,-nbitq), 
to_sfixed(-65877745.0/4294967296.0,1,-nbitq), 
to_sfixed(287837306.0/4294967296.0,1,-nbitq), 
to_sfixed(-342009604.0/4294967296.0,1,-nbitq), 
to_sfixed(-89678613.0/4294967296.0,1,-nbitq), 
to_sfixed(345527021.0/4294967296.0,1,-nbitq), 
to_sfixed(-245110567.0/4294967296.0,1,-nbitq), 
to_sfixed(353800159.0/4294967296.0,1,-nbitq), 
to_sfixed(99954726.0/4294967296.0,1,-nbitq), 
to_sfixed(-105244184.0/4294967296.0,1,-nbitq), 
to_sfixed(-551630710.0/4294967296.0,1,-nbitq), 
to_sfixed(-49297283.0/4294967296.0,1,-nbitq), 
to_sfixed(188741445.0/4294967296.0,1,-nbitq), 
to_sfixed(-480503446.0/4294967296.0,1,-nbitq), 
to_sfixed(-186068758.0/4294967296.0,1,-nbitq), 
to_sfixed(283401298.0/4294967296.0,1,-nbitq), 
to_sfixed(143647479.0/4294967296.0,1,-nbitq), 
to_sfixed(543506602.0/4294967296.0,1,-nbitq), 
to_sfixed(310897497.0/4294967296.0,1,-nbitq), 
to_sfixed(-252401931.0/4294967296.0,1,-nbitq), 
to_sfixed(693818516.0/4294967296.0,1,-nbitq), 
to_sfixed(-438376045.0/4294967296.0,1,-nbitq), 
to_sfixed(286012559.0/4294967296.0,1,-nbitq), 
to_sfixed(145418669.0/4294967296.0,1,-nbitq), 
to_sfixed(211082713.0/4294967296.0,1,-nbitq), 
to_sfixed(-98845429.0/4294967296.0,1,-nbitq), 
to_sfixed(-159475583.0/4294967296.0,1,-nbitq), 
to_sfixed(-90649450.0/4294967296.0,1,-nbitq), 
to_sfixed(-127228330.0/4294967296.0,1,-nbitq), 
to_sfixed(-408500755.0/4294967296.0,1,-nbitq), 
to_sfixed(-20725197.0/4294967296.0,1,-nbitq), 
to_sfixed(205539264.0/4294967296.0,1,-nbitq), 
to_sfixed(-171720162.0/4294967296.0,1,-nbitq), 
to_sfixed(132647855.0/4294967296.0,1,-nbitq), 
to_sfixed(33233253.0/4294967296.0,1,-nbitq), 
to_sfixed(-339169378.0/4294967296.0,1,-nbitq), 
to_sfixed(358861443.0/4294967296.0,1,-nbitq), 
to_sfixed(596496054.0/4294967296.0,1,-nbitq), 
to_sfixed(339622783.0/4294967296.0,1,-nbitq), 
to_sfixed(-125404199.0/4294967296.0,1,-nbitq), 
to_sfixed(-309522152.0/4294967296.0,1,-nbitq), 
to_sfixed(-155422002.0/4294967296.0,1,-nbitq), 
to_sfixed(-326006531.0/4294967296.0,1,-nbitq), 
to_sfixed(1663861.0/4294967296.0,1,-nbitq), 
to_sfixed(503805048.0/4294967296.0,1,-nbitq), 
to_sfixed(213503756.0/4294967296.0,1,-nbitq), 
to_sfixed(296291626.0/4294967296.0,1,-nbitq), 
to_sfixed(366031489.0/4294967296.0,1,-nbitq), 
to_sfixed(601603.0/4294967296.0,1,-nbitq), 
to_sfixed(602353583.0/4294967296.0,1,-nbitq), 
to_sfixed(-234512750.0/4294967296.0,1,-nbitq), 
to_sfixed(350340039.0/4294967296.0,1,-nbitq), 
to_sfixed(61519534.0/4294967296.0,1,-nbitq), 
to_sfixed(-317151089.0/4294967296.0,1,-nbitq), 
to_sfixed(-152607559.0/4294967296.0,1,-nbitq), 
to_sfixed(-366945464.0/4294967296.0,1,-nbitq), 
to_sfixed(16409819.0/4294967296.0,1,-nbitq), 
to_sfixed(-208264617.0/4294967296.0,1,-nbitq), 
to_sfixed(-439476526.0/4294967296.0,1,-nbitq), 
to_sfixed(37832861.0/4294967296.0,1,-nbitq), 
to_sfixed(-88044635.0/4294967296.0,1,-nbitq), 
to_sfixed(29209936.0/4294967296.0,1,-nbitq), 
to_sfixed(-89465556.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(370983947.0/4294967296.0,1,-nbitq), 
to_sfixed(-359072296.0/4294967296.0,1,-nbitq), 
to_sfixed(305777741.0/4294967296.0,1,-nbitq), 
to_sfixed(-169391288.0/4294967296.0,1,-nbitq), 
to_sfixed(572808620.0/4294967296.0,1,-nbitq), 
to_sfixed(106203480.0/4294967296.0,1,-nbitq), 
to_sfixed(-38823043.0/4294967296.0,1,-nbitq), 
to_sfixed(244517752.0/4294967296.0,1,-nbitq), 
to_sfixed(175709770.0/4294967296.0,1,-nbitq), 
to_sfixed(-324807413.0/4294967296.0,1,-nbitq), 
to_sfixed(-94608458.0/4294967296.0,1,-nbitq), 
to_sfixed(-128454474.0/4294967296.0,1,-nbitq), 
to_sfixed(218019257.0/4294967296.0,1,-nbitq), 
to_sfixed(128819761.0/4294967296.0,1,-nbitq), 
to_sfixed(363833528.0/4294967296.0,1,-nbitq), 
to_sfixed(136200529.0/4294967296.0,1,-nbitq), 
to_sfixed(-6140543.0/4294967296.0,1,-nbitq), 
to_sfixed(314953546.0/4294967296.0,1,-nbitq), 
to_sfixed(137534347.0/4294967296.0,1,-nbitq), 
to_sfixed(308860986.0/4294967296.0,1,-nbitq), 
to_sfixed(249578103.0/4294967296.0,1,-nbitq), 
to_sfixed(384232418.0/4294967296.0,1,-nbitq), 
to_sfixed(-392671678.0/4294967296.0,1,-nbitq), 
to_sfixed(277133715.0/4294967296.0,1,-nbitq), 
to_sfixed(-232064320.0/4294967296.0,1,-nbitq), 
to_sfixed(-360111082.0/4294967296.0,1,-nbitq), 
to_sfixed(254959269.0/4294967296.0,1,-nbitq), 
to_sfixed(139468488.0/4294967296.0,1,-nbitq), 
to_sfixed(-74259491.0/4294967296.0,1,-nbitq), 
to_sfixed(-189137064.0/4294967296.0,1,-nbitq), 
to_sfixed(240536557.0/4294967296.0,1,-nbitq), 
to_sfixed(-662654768.0/4294967296.0,1,-nbitq), 
to_sfixed(-66328193.0/4294967296.0,1,-nbitq), 
to_sfixed(-14184436.0/4294967296.0,1,-nbitq), 
to_sfixed(30469893.0/4294967296.0,1,-nbitq), 
to_sfixed(399486129.0/4294967296.0,1,-nbitq), 
to_sfixed(122377341.0/4294967296.0,1,-nbitq), 
to_sfixed(468509533.0/4294967296.0,1,-nbitq), 
to_sfixed(99101683.0/4294967296.0,1,-nbitq), 
to_sfixed(9175053.0/4294967296.0,1,-nbitq), 
to_sfixed(-192042985.0/4294967296.0,1,-nbitq), 
to_sfixed(-265785933.0/4294967296.0,1,-nbitq), 
to_sfixed(13490288.0/4294967296.0,1,-nbitq), 
to_sfixed(-203546798.0/4294967296.0,1,-nbitq), 
to_sfixed(-566350961.0/4294967296.0,1,-nbitq), 
to_sfixed(383328976.0/4294967296.0,1,-nbitq), 
to_sfixed(305499795.0/4294967296.0,1,-nbitq), 
to_sfixed(170461239.0/4294967296.0,1,-nbitq), 
to_sfixed(137065889.0/4294967296.0,1,-nbitq), 
to_sfixed(-352509521.0/4294967296.0,1,-nbitq), 
to_sfixed(86513906.0/4294967296.0,1,-nbitq), 
to_sfixed(443136452.0/4294967296.0,1,-nbitq), 
to_sfixed(-73694294.0/4294967296.0,1,-nbitq), 
to_sfixed(423547571.0/4294967296.0,1,-nbitq), 
to_sfixed(113436425.0/4294967296.0,1,-nbitq), 
to_sfixed(-233801091.0/4294967296.0,1,-nbitq), 
to_sfixed(-192011070.0/4294967296.0,1,-nbitq), 
to_sfixed(-285671409.0/4294967296.0,1,-nbitq), 
to_sfixed(-59964348.0/4294967296.0,1,-nbitq), 
to_sfixed(-27500993.0/4294967296.0,1,-nbitq), 
to_sfixed(90322962.0/4294967296.0,1,-nbitq), 
to_sfixed(163194868.0/4294967296.0,1,-nbitq), 
to_sfixed(321564636.0/4294967296.0,1,-nbitq), 
to_sfixed(-196005008.0/4294967296.0,1,-nbitq), 
to_sfixed(-244266786.0/4294967296.0,1,-nbitq), 
to_sfixed(307227654.0/4294967296.0,1,-nbitq), 
to_sfixed(-282692473.0/4294967296.0,1,-nbitq), 
to_sfixed(-291107309.0/4294967296.0,1,-nbitq), 
to_sfixed(-158213816.0/4294967296.0,1,-nbitq), 
to_sfixed(563341480.0/4294967296.0,1,-nbitq), 
to_sfixed(293774046.0/4294967296.0,1,-nbitq), 
to_sfixed(-197603022.0/4294967296.0,1,-nbitq), 
to_sfixed(296774845.0/4294967296.0,1,-nbitq), 
to_sfixed(9230256.0/4294967296.0,1,-nbitq), 
to_sfixed(-2230594.0/4294967296.0,1,-nbitq), 
to_sfixed(-132604940.0/4294967296.0,1,-nbitq), 
to_sfixed(273751014.0/4294967296.0,1,-nbitq), 
to_sfixed(175696977.0/4294967296.0,1,-nbitq), 
to_sfixed(-114300953.0/4294967296.0,1,-nbitq), 
to_sfixed(375727650.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-286232853.0/4294967296.0,1,-nbitq), 
to_sfixed(-339519976.0/4294967296.0,1,-nbitq), 
to_sfixed(-160368277.0/4294967296.0,1,-nbitq), 
to_sfixed(169002225.0/4294967296.0,1,-nbitq), 
to_sfixed(-117170968.0/4294967296.0,1,-nbitq), 
to_sfixed(275349052.0/4294967296.0,1,-nbitq), 
to_sfixed(390425453.0/4294967296.0,1,-nbitq), 
to_sfixed(90261011.0/4294967296.0,1,-nbitq), 
to_sfixed(356698243.0/4294967296.0,1,-nbitq), 
to_sfixed(89039276.0/4294967296.0,1,-nbitq), 
to_sfixed(216156182.0/4294967296.0,1,-nbitq), 
to_sfixed(299203425.0/4294967296.0,1,-nbitq), 
to_sfixed(307882528.0/4294967296.0,1,-nbitq), 
to_sfixed(-562659871.0/4294967296.0,1,-nbitq), 
to_sfixed(130351298.0/4294967296.0,1,-nbitq), 
to_sfixed(251858696.0/4294967296.0,1,-nbitq), 
to_sfixed(-82859034.0/4294967296.0,1,-nbitq), 
to_sfixed(-267822600.0/4294967296.0,1,-nbitq), 
to_sfixed(-898520969.0/4294967296.0,1,-nbitq), 
to_sfixed(447456145.0/4294967296.0,1,-nbitq), 
to_sfixed(-101842315.0/4294967296.0,1,-nbitq), 
to_sfixed(121405667.0/4294967296.0,1,-nbitq), 
to_sfixed(-359990371.0/4294967296.0,1,-nbitq), 
to_sfixed(179306714.0/4294967296.0,1,-nbitq), 
to_sfixed(-234514301.0/4294967296.0,1,-nbitq), 
to_sfixed(-70391193.0/4294967296.0,1,-nbitq), 
to_sfixed(100326858.0/4294967296.0,1,-nbitq), 
to_sfixed(-64418207.0/4294967296.0,1,-nbitq), 
to_sfixed(-634964435.0/4294967296.0,1,-nbitq), 
to_sfixed(-672217470.0/4294967296.0,1,-nbitq), 
to_sfixed(329370169.0/4294967296.0,1,-nbitq), 
to_sfixed(-643473480.0/4294967296.0,1,-nbitq), 
to_sfixed(329518049.0/4294967296.0,1,-nbitq), 
to_sfixed(309154042.0/4294967296.0,1,-nbitq), 
to_sfixed(-207595394.0/4294967296.0,1,-nbitq), 
to_sfixed(608867266.0/4294967296.0,1,-nbitq), 
to_sfixed(313403120.0/4294967296.0,1,-nbitq), 
to_sfixed(6333168.0/4294967296.0,1,-nbitq), 
to_sfixed(-30744385.0/4294967296.0,1,-nbitq), 
to_sfixed(118570023.0/4294967296.0,1,-nbitq), 
to_sfixed(343933687.0/4294967296.0,1,-nbitq), 
to_sfixed(-539101079.0/4294967296.0,1,-nbitq), 
to_sfixed(-602337328.0/4294967296.0,1,-nbitq), 
to_sfixed(-737400498.0/4294967296.0,1,-nbitq), 
to_sfixed(-62762235.0/4294967296.0,1,-nbitq), 
to_sfixed(312906547.0/4294967296.0,1,-nbitq), 
to_sfixed(-52724094.0/4294967296.0,1,-nbitq), 
to_sfixed(-249330176.0/4294967296.0,1,-nbitq), 
to_sfixed(-23802074.0/4294967296.0,1,-nbitq), 
to_sfixed(-588193887.0/4294967296.0,1,-nbitq), 
to_sfixed(-98448648.0/4294967296.0,1,-nbitq), 
to_sfixed(725701952.0/4294967296.0,1,-nbitq), 
to_sfixed(350519868.0/4294967296.0,1,-nbitq), 
to_sfixed(-141281323.0/4294967296.0,1,-nbitq), 
to_sfixed(243623757.0/4294967296.0,1,-nbitq), 
to_sfixed(119038509.0/4294967296.0,1,-nbitq), 
to_sfixed(243445908.0/4294967296.0,1,-nbitq), 
to_sfixed(272255929.0/4294967296.0,1,-nbitq), 
to_sfixed(-8905044.0/4294967296.0,1,-nbitq), 
to_sfixed(-94519209.0/4294967296.0,1,-nbitq), 
to_sfixed(-185974257.0/4294967296.0,1,-nbitq), 
to_sfixed(-668205962.0/4294967296.0,1,-nbitq), 
to_sfixed(84026766.0/4294967296.0,1,-nbitq), 
to_sfixed(-141165132.0/4294967296.0,1,-nbitq), 
to_sfixed(-216691062.0/4294967296.0,1,-nbitq), 
to_sfixed(345603535.0/4294967296.0,1,-nbitq), 
to_sfixed(-446724237.0/4294967296.0,1,-nbitq), 
to_sfixed(141436814.0/4294967296.0,1,-nbitq), 
to_sfixed(40448552.0/4294967296.0,1,-nbitq), 
to_sfixed(579062828.0/4294967296.0,1,-nbitq), 
to_sfixed(-200840695.0/4294967296.0,1,-nbitq), 
to_sfixed(135154578.0/4294967296.0,1,-nbitq), 
to_sfixed(157669318.0/4294967296.0,1,-nbitq), 
to_sfixed(79824498.0/4294967296.0,1,-nbitq), 
to_sfixed(62714710.0/4294967296.0,1,-nbitq), 
to_sfixed(-357283879.0/4294967296.0,1,-nbitq), 
to_sfixed(-52925105.0/4294967296.0,1,-nbitq), 
to_sfixed(326171372.0/4294967296.0,1,-nbitq), 
to_sfixed(-45515234.0/4294967296.0,1,-nbitq), 
to_sfixed(-276094181.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-137941635.0/4294967296.0,1,-nbitq), 
to_sfixed(106827341.0/4294967296.0,1,-nbitq), 
to_sfixed(410891049.0/4294967296.0,1,-nbitq), 
to_sfixed(594839693.0/4294967296.0,1,-nbitq), 
to_sfixed(-267458016.0/4294967296.0,1,-nbitq), 
to_sfixed(357973901.0/4294967296.0,1,-nbitq), 
to_sfixed(361602281.0/4294967296.0,1,-nbitq), 
to_sfixed(-107737415.0/4294967296.0,1,-nbitq), 
to_sfixed(339698693.0/4294967296.0,1,-nbitq), 
to_sfixed(-53127271.0/4294967296.0,1,-nbitq), 
to_sfixed(-63028978.0/4294967296.0,1,-nbitq), 
to_sfixed(-810449005.0/4294967296.0,1,-nbitq), 
to_sfixed(-159224915.0/4294967296.0,1,-nbitq), 
to_sfixed(-861900492.0/4294967296.0,1,-nbitq), 
to_sfixed(361339685.0/4294967296.0,1,-nbitq), 
to_sfixed(486809907.0/4294967296.0,1,-nbitq), 
to_sfixed(-202655058.0/4294967296.0,1,-nbitq), 
to_sfixed(206323831.0/4294967296.0,1,-nbitq), 
to_sfixed(-907019409.0/4294967296.0,1,-nbitq), 
to_sfixed(353505833.0/4294967296.0,1,-nbitq), 
to_sfixed(-365640106.0/4294967296.0,1,-nbitq), 
to_sfixed(47196549.0/4294967296.0,1,-nbitq), 
to_sfixed(-583031350.0/4294967296.0,1,-nbitq), 
to_sfixed(244875076.0/4294967296.0,1,-nbitq), 
to_sfixed(-122363226.0/4294967296.0,1,-nbitq), 
to_sfixed(-545057140.0/4294967296.0,1,-nbitq), 
to_sfixed(552795020.0/4294967296.0,1,-nbitq), 
to_sfixed(61577948.0/4294967296.0,1,-nbitq), 
to_sfixed(-475858254.0/4294967296.0,1,-nbitq), 
to_sfixed(-1235210778.0/4294967296.0,1,-nbitq), 
to_sfixed(79754583.0/4294967296.0,1,-nbitq), 
to_sfixed(-237632245.0/4294967296.0,1,-nbitq), 
to_sfixed(778154956.0/4294967296.0,1,-nbitq), 
to_sfixed(638169486.0/4294967296.0,1,-nbitq), 
to_sfixed(-423674986.0/4294967296.0,1,-nbitq), 
to_sfixed(14697192.0/4294967296.0,1,-nbitq), 
to_sfixed(306238578.0/4294967296.0,1,-nbitq), 
to_sfixed(-474796965.0/4294967296.0,1,-nbitq), 
to_sfixed(231896560.0/4294967296.0,1,-nbitq), 
to_sfixed(-39447605.0/4294967296.0,1,-nbitq), 
to_sfixed(-121900528.0/4294967296.0,1,-nbitq), 
to_sfixed(-445884758.0/4294967296.0,1,-nbitq), 
to_sfixed(-546215240.0/4294967296.0,1,-nbitq), 
to_sfixed(-296823739.0/4294967296.0,1,-nbitq), 
to_sfixed(-228567989.0/4294967296.0,1,-nbitq), 
to_sfixed(-137293922.0/4294967296.0,1,-nbitq), 
to_sfixed(-388844206.0/4294967296.0,1,-nbitq), 
to_sfixed(-383487219.0/4294967296.0,1,-nbitq), 
to_sfixed(76753595.0/4294967296.0,1,-nbitq), 
to_sfixed(-131164567.0/4294967296.0,1,-nbitq), 
to_sfixed(-24891319.0/4294967296.0,1,-nbitq), 
to_sfixed(586313201.0/4294967296.0,1,-nbitq), 
to_sfixed(231375584.0/4294967296.0,1,-nbitq), 
to_sfixed(-302771623.0/4294967296.0,1,-nbitq), 
to_sfixed(-654292556.0/4294967296.0,1,-nbitq), 
to_sfixed(410179441.0/4294967296.0,1,-nbitq), 
to_sfixed(273906076.0/4294967296.0,1,-nbitq), 
to_sfixed(-247975048.0/4294967296.0,1,-nbitq), 
to_sfixed(-72109731.0/4294967296.0,1,-nbitq), 
to_sfixed(157291848.0/4294967296.0,1,-nbitq), 
to_sfixed(72927918.0/4294967296.0,1,-nbitq), 
to_sfixed(-671401866.0/4294967296.0,1,-nbitq), 
to_sfixed(162977053.0/4294967296.0,1,-nbitq), 
to_sfixed(-414022887.0/4294967296.0,1,-nbitq), 
to_sfixed(-153244728.0/4294967296.0,1,-nbitq), 
to_sfixed(-206339779.0/4294967296.0,1,-nbitq), 
to_sfixed(-1492428474.0/4294967296.0,1,-nbitq), 
to_sfixed(36290752.0/4294967296.0,1,-nbitq), 
to_sfixed(-185790045.0/4294967296.0,1,-nbitq), 
to_sfixed(277807658.0/4294967296.0,1,-nbitq), 
to_sfixed(-722822658.0/4294967296.0,1,-nbitq), 
to_sfixed(58306374.0/4294967296.0,1,-nbitq), 
to_sfixed(577990526.0/4294967296.0,1,-nbitq), 
to_sfixed(228317294.0/4294967296.0,1,-nbitq), 
to_sfixed(-144308099.0/4294967296.0,1,-nbitq), 
to_sfixed(87516221.0/4294967296.0,1,-nbitq), 
to_sfixed(95858639.0/4294967296.0,1,-nbitq), 
to_sfixed(-251725263.0/4294967296.0,1,-nbitq), 
to_sfixed(-1033073864.0/4294967296.0,1,-nbitq), 
to_sfixed(-109329830.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(432200575.0/4294967296.0,1,-nbitq), 
to_sfixed(-9105772.0/4294967296.0,1,-nbitq), 
to_sfixed(832081550.0/4294967296.0,1,-nbitq), 
to_sfixed(118212541.0/4294967296.0,1,-nbitq), 
to_sfixed(-248148695.0/4294967296.0,1,-nbitq), 
to_sfixed(717641943.0/4294967296.0,1,-nbitq), 
to_sfixed(-42108718.0/4294967296.0,1,-nbitq), 
to_sfixed(396893566.0/4294967296.0,1,-nbitq), 
to_sfixed(637268725.0/4294967296.0,1,-nbitq), 
to_sfixed(186354917.0/4294967296.0,1,-nbitq), 
to_sfixed(231885401.0/4294967296.0,1,-nbitq), 
to_sfixed(-271982148.0/4294967296.0,1,-nbitq), 
to_sfixed(-415717143.0/4294967296.0,1,-nbitq), 
to_sfixed(-495542692.0/4294967296.0,1,-nbitq), 
to_sfixed(371349211.0/4294967296.0,1,-nbitq), 
to_sfixed(431856753.0/4294967296.0,1,-nbitq), 
to_sfixed(315170313.0/4294967296.0,1,-nbitq), 
to_sfixed(407530946.0/4294967296.0,1,-nbitq), 
to_sfixed(-1010742356.0/4294967296.0,1,-nbitq), 
to_sfixed(7650096.0/4294967296.0,1,-nbitq), 
to_sfixed(-211548509.0/4294967296.0,1,-nbitq), 
to_sfixed(-210321603.0/4294967296.0,1,-nbitq), 
to_sfixed(-35018363.0/4294967296.0,1,-nbitq), 
to_sfixed(-46071113.0/4294967296.0,1,-nbitq), 
to_sfixed(218057163.0/4294967296.0,1,-nbitq), 
to_sfixed(-978699621.0/4294967296.0,1,-nbitq), 
to_sfixed(190496620.0/4294967296.0,1,-nbitq), 
to_sfixed(353106676.0/4294967296.0,1,-nbitq), 
to_sfixed(3713348.0/4294967296.0,1,-nbitq), 
to_sfixed(-907534293.0/4294967296.0,1,-nbitq), 
to_sfixed(501021578.0/4294967296.0,1,-nbitq), 
to_sfixed(24471709.0/4294967296.0,1,-nbitq), 
to_sfixed(536852566.0/4294967296.0,1,-nbitq), 
to_sfixed(600230826.0/4294967296.0,1,-nbitq), 
to_sfixed(-68509056.0/4294967296.0,1,-nbitq), 
to_sfixed(-682977127.0/4294967296.0,1,-nbitq), 
to_sfixed(296255672.0/4294967296.0,1,-nbitq), 
to_sfixed(248247182.0/4294967296.0,1,-nbitq), 
to_sfixed(119680167.0/4294967296.0,1,-nbitq), 
to_sfixed(122194874.0/4294967296.0,1,-nbitq), 
to_sfixed(511715501.0/4294967296.0,1,-nbitq), 
to_sfixed(-713408431.0/4294967296.0,1,-nbitq), 
to_sfixed(-339742438.0/4294967296.0,1,-nbitq), 
to_sfixed(-396671122.0/4294967296.0,1,-nbitq), 
to_sfixed(334645246.0/4294967296.0,1,-nbitq), 
to_sfixed(-282416434.0/4294967296.0,1,-nbitq), 
to_sfixed(307288810.0/4294967296.0,1,-nbitq), 
to_sfixed(253014133.0/4294967296.0,1,-nbitq), 
to_sfixed(93014041.0/4294967296.0,1,-nbitq), 
to_sfixed(-33113156.0/4294967296.0,1,-nbitq), 
to_sfixed(-383612181.0/4294967296.0,1,-nbitq), 
to_sfixed(574868599.0/4294967296.0,1,-nbitq), 
to_sfixed(622313023.0/4294967296.0,1,-nbitq), 
to_sfixed(-249418420.0/4294967296.0,1,-nbitq), 
to_sfixed(-1325799298.0/4294967296.0,1,-nbitq), 
to_sfixed(855422555.0/4294967296.0,1,-nbitq), 
to_sfixed(-108016738.0/4294967296.0,1,-nbitq), 
to_sfixed(273731462.0/4294967296.0,1,-nbitq), 
to_sfixed(8728635.0/4294967296.0,1,-nbitq), 
to_sfixed(-65223365.0/4294967296.0,1,-nbitq), 
to_sfixed(45274669.0/4294967296.0,1,-nbitq), 
to_sfixed(-30903443.0/4294967296.0,1,-nbitq), 
to_sfixed(81551526.0/4294967296.0,1,-nbitq), 
to_sfixed(-233644276.0/4294967296.0,1,-nbitq), 
to_sfixed(-111599488.0/4294967296.0,1,-nbitq), 
to_sfixed(140034768.0/4294967296.0,1,-nbitq), 
to_sfixed(-1327892258.0/4294967296.0,1,-nbitq), 
to_sfixed(-209904342.0/4294967296.0,1,-nbitq), 
to_sfixed(199219815.0/4294967296.0,1,-nbitq), 
to_sfixed(-43408123.0/4294967296.0,1,-nbitq), 
to_sfixed(-1181609681.0/4294967296.0,1,-nbitq), 
to_sfixed(-95730358.0/4294967296.0,1,-nbitq), 
to_sfixed(565317685.0/4294967296.0,1,-nbitq), 
to_sfixed(-39809401.0/4294967296.0,1,-nbitq), 
to_sfixed(108601814.0/4294967296.0,1,-nbitq), 
to_sfixed(472534491.0/4294967296.0,1,-nbitq), 
to_sfixed(-459553511.0/4294967296.0,1,-nbitq), 
to_sfixed(115375102.0/4294967296.0,1,-nbitq), 
to_sfixed(-851086073.0/4294967296.0,1,-nbitq), 
to_sfixed(-318544485.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-252308985.0/4294967296.0,1,-nbitq), 
to_sfixed(-4801313.0/4294967296.0,1,-nbitq), 
to_sfixed(931520752.0/4294967296.0,1,-nbitq), 
to_sfixed(800855025.0/4294967296.0,1,-nbitq), 
to_sfixed(-93542735.0/4294967296.0,1,-nbitq), 
to_sfixed(1129642583.0/4294967296.0,1,-nbitq), 
to_sfixed(-176958299.0/4294967296.0,1,-nbitq), 
to_sfixed(568723784.0/4294967296.0,1,-nbitq), 
to_sfixed(1293199340.0/4294967296.0,1,-nbitq), 
to_sfixed(259646463.0/4294967296.0,1,-nbitq), 
to_sfixed(-191519212.0/4294967296.0,1,-nbitq), 
to_sfixed(-42790345.0/4294967296.0,1,-nbitq), 
to_sfixed(-851053093.0/4294967296.0,1,-nbitq), 
to_sfixed(-970267139.0/4294967296.0,1,-nbitq), 
to_sfixed(-134568225.0/4294967296.0,1,-nbitq), 
to_sfixed(209303457.0/4294967296.0,1,-nbitq), 
to_sfixed(-17295991.0/4294967296.0,1,-nbitq), 
to_sfixed(395074082.0/4294967296.0,1,-nbitq), 
to_sfixed(-1032791322.0/4294967296.0,1,-nbitq), 
to_sfixed(-123169523.0/4294967296.0,1,-nbitq), 
to_sfixed(-353370567.0/4294967296.0,1,-nbitq), 
to_sfixed(-224902294.0/4294967296.0,1,-nbitq), 
to_sfixed(128798940.0/4294967296.0,1,-nbitq), 
to_sfixed(11059595.0/4294967296.0,1,-nbitq), 
to_sfixed(62581599.0/4294967296.0,1,-nbitq), 
to_sfixed(-992898718.0/4294967296.0,1,-nbitq), 
to_sfixed(235914931.0/4294967296.0,1,-nbitq), 
to_sfixed(468327521.0/4294967296.0,1,-nbitq), 
to_sfixed(226159969.0/4294967296.0,1,-nbitq), 
to_sfixed(-195701596.0/4294967296.0,1,-nbitq), 
to_sfixed(584008721.0/4294967296.0,1,-nbitq), 
to_sfixed(-191644816.0/4294967296.0,1,-nbitq), 
to_sfixed(755164302.0/4294967296.0,1,-nbitq), 
to_sfixed(1071367859.0/4294967296.0,1,-nbitq), 
to_sfixed(-662317719.0/4294967296.0,1,-nbitq), 
to_sfixed(-890001001.0/4294967296.0,1,-nbitq), 
to_sfixed(834353531.0/4294967296.0,1,-nbitq), 
to_sfixed(548500419.0/4294967296.0,1,-nbitq), 
to_sfixed(7300512.0/4294967296.0,1,-nbitq), 
to_sfixed(-120020377.0/4294967296.0,1,-nbitq), 
to_sfixed(123324744.0/4294967296.0,1,-nbitq), 
to_sfixed(-852185744.0/4294967296.0,1,-nbitq), 
to_sfixed(-188455222.0/4294967296.0,1,-nbitq), 
to_sfixed(-597752522.0/4294967296.0,1,-nbitq), 
to_sfixed(-347634339.0/4294967296.0,1,-nbitq), 
to_sfixed(-1162909193.0/4294967296.0,1,-nbitq), 
to_sfixed(-167570962.0/4294967296.0,1,-nbitq), 
to_sfixed(258666694.0/4294967296.0,1,-nbitq), 
to_sfixed(-345949390.0/4294967296.0,1,-nbitq), 
to_sfixed(-960587250.0/4294967296.0,1,-nbitq), 
to_sfixed(-271165560.0/4294967296.0,1,-nbitq), 
to_sfixed(284801938.0/4294967296.0,1,-nbitq), 
to_sfixed(380474419.0/4294967296.0,1,-nbitq), 
to_sfixed(-851514379.0/4294967296.0,1,-nbitq), 
to_sfixed(-922803421.0/4294967296.0,1,-nbitq), 
to_sfixed(642966927.0/4294967296.0,1,-nbitq), 
to_sfixed(-199390705.0/4294967296.0,1,-nbitq), 
to_sfixed(222709158.0/4294967296.0,1,-nbitq), 
to_sfixed(-125605876.0/4294967296.0,1,-nbitq), 
to_sfixed(420253316.0/4294967296.0,1,-nbitq), 
to_sfixed(-280548960.0/4294967296.0,1,-nbitq), 
to_sfixed(-366765151.0/4294967296.0,1,-nbitq), 
to_sfixed(-527835339.0/4294967296.0,1,-nbitq), 
to_sfixed(-423967129.0/4294967296.0,1,-nbitq), 
to_sfixed(-476433185.0/4294967296.0,1,-nbitq), 
to_sfixed(414761959.0/4294967296.0,1,-nbitq), 
to_sfixed(-1349304183.0/4294967296.0,1,-nbitq), 
to_sfixed(-985955529.0/4294967296.0,1,-nbitq), 
to_sfixed(-230539294.0/4294967296.0,1,-nbitq), 
to_sfixed(818041391.0/4294967296.0,1,-nbitq), 
to_sfixed(-478442394.0/4294967296.0,1,-nbitq), 
to_sfixed(67331604.0/4294967296.0,1,-nbitq), 
to_sfixed(-65551054.0/4294967296.0,1,-nbitq), 
to_sfixed(148007216.0/4294967296.0,1,-nbitq), 
to_sfixed(523288038.0/4294967296.0,1,-nbitq), 
to_sfixed(396531400.0/4294967296.0,1,-nbitq), 
to_sfixed(257218603.0/4294967296.0,1,-nbitq), 
to_sfixed(27028069.0/4294967296.0,1,-nbitq), 
to_sfixed(-962531427.0/4294967296.0,1,-nbitq), 
to_sfixed(14860341.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-115226225.0/4294967296.0,1,-nbitq), 
to_sfixed(513430823.0/4294967296.0,1,-nbitq), 
to_sfixed(1500974649.0/4294967296.0,1,-nbitq), 
to_sfixed(578994689.0/4294967296.0,1,-nbitq), 
to_sfixed(69020859.0/4294967296.0,1,-nbitq), 
to_sfixed(936123764.0/4294967296.0,1,-nbitq), 
to_sfixed(-362216274.0/4294967296.0,1,-nbitq), 
to_sfixed(133724805.0/4294967296.0,1,-nbitq), 
to_sfixed(589875815.0/4294967296.0,1,-nbitq), 
to_sfixed(-321312811.0/4294967296.0,1,-nbitq), 
to_sfixed(-83868034.0/4294967296.0,1,-nbitq), 
to_sfixed(418752158.0/4294967296.0,1,-nbitq), 
to_sfixed(-791041069.0/4294967296.0,1,-nbitq), 
to_sfixed(-877177547.0/4294967296.0,1,-nbitq), 
to_sfixed(270698663.0/4294967296.0,1,-nbitq), 
to_sfixed(367629864.0/4294967296.0,1,-nbitq), 
to_sfixed(-256801480.0/4294967296.0,1,-nbitq), 
to_sfixed(411982306.0/4294967296.0,1,-nbitq), 
to_sfixed(-270011181.0/4294967296.0,1,-nbitq), 
to_sfixed(209054277.0/4294967296.0,1,-nbitq), 
to_sfixed(-353235060.0/4294967296.0,1,-nbitq), 
to_sfixed(350703318.0/4294967296.0,1,-nbitq), 
to_sfixed(336917680.0/4294967296.0,1,-nbitq), 
to_sfixed(113272167.0/4294967296.0,1,-nbitq), 
to_sfixed(-148335328.0/4294967296.0,1,-nbitq), 
to_sfixed(209559168.0/4294967296.0,1,-nbitq), 
to_sfixed(-72808088.0/4294967296.0,1,-nbitq), 
to_sfixed(874375359.0/4294967296.0,1,-nbitq), 
to_sfixed(583623328.0/4294967296.0,1,-nbitq), 
to_sfixed(-149533948.0/4294967296.0,1,-nbitq), 
to_sfixed(626945390.0/4294967296.0,1,-nbitq), 
to_sfixed(-281955114.0/4294967296.0,1,-nbitq), 
to_sfixed(597515981.0/4294967296.0,1,-nbitq), 
to_sfixed(651204807.0/4294967296.0,1,-nbitq), 
to_sfixed(-1137797215.0/4294967296.0,1,-nbitq), 
to_sfixed(-619833219.0/4294967296.0,1,-nbitq), 
to_sfixed(721279866.0/4294967296.0,1,-nbitq), 
to_sfixed(-473537938.0/4294967296.0,1,-nbitq), 
to_sfixed(113737633.0/4294967296.0,1,-nbitq), 
to_sfixed(205568589.0/4294967296.0,1,-nbitq), 
to_sfixed(79394633.0/4294967296.0,1,-nbitq), 
to_sfixed(-271667291.0/4294967296.0,1,-nbitq), 
to_sfixed(-318965084.0/4294967296.0,1,-nbitq), 
to_sfixed(-399551613.0/4294967296.0,1,-nbitq), 
to_sfixed(-353744659.0/4294967296.0,1,-nbitq), 
to_sfixed(-1698747648.0/4294967296.0,1,-nbitq), 
to_sfixed(-253189872.0/4294967296.0,1,-nbitq), 
to_sfixed(749876659.0/4294967296.0,1,-nbitq), 
to_sfixed(-599404127.0/4294967296.0,1,-nbitq), 
to_sfixed(-1193799345.0/4294967296.0,1,-nbitq), 
to_sfixed(-834781109.0/4294967296.0,1,-nbitq), 
to_sfixed(880574674.0/4294967296.0,1,-nbitq), 
to_sfixed(-778717036.0/4294967296.0,1,-nbitq), 
to_sfixed(353415546.0/4294967296.0,1,-nbitq), 
to_sfixed(117876668.0/4294967296.0,1,-nbitq), 
to_sfixed(250732097.0/4294967296.0,1,-nbitq), 
to_sfixed(-345856554.0/4294967296.0,1,-nbitq), 
to_sfixed(699235656.0/4294967296.0,1,-nbitq), 
to_sfixed(-19819594.0/4294967296.0,1,-nbitq), 
to_sfixed(-164801356.0/4294967296.0,1,-nbitq), 
to_sfixed(43754735.0/4294967296.0,1,-nbitq), 
to_sfixed(-345227823.0/4294967296.0,1,-nbitq), 
to_sfixed(-665679149.0/4294967296.0,1,-nbitq), 
to_sfixed(-749522191.0/4294967296.0,1,-nbitq), 
to_sfixed(-354354445.0/4294967296.0,1,-nbitq), 
to_sfixed(213763490.0/4294967296.0,1,-nbitq), 
to_sfixed(-1200832963.0/4294967296.0,1,-nbitq), 
to_sfixed(-1195892737.0/4294967296.0,1,-nbitq), 
to_sfixed(-85928211.0/4294967296.0,1,-nbitq), 
to_sfixed(517116790.0/4294967296.0,1,-nbitq), 
to_sfixed(-1325521141.0/4294967296.0,1,-nbitq), 
to_sfixed(164697748.0/4294967296.0,1,-nbitq), 
to_sfixed(502590389.0/4294967296.0,1,-nbitq), 
to_sfixed(-108961024.0/4294967296.0,1,-nbitq), 
to_sfixed(-126507935.0/4294967296.0,1,-nbitq), 
to_sfixed(179265838.0/4294967296.0,1,-nbitq), 
to_sfixed(-11473558.0/4294967296.0,1,-nbitq), 
to_sfixed(-848429382.0/4294967296.0,1,-nbitq), 
to_sfixed(43922646.0/4294967296.0,1,-nbitq), 
to_sfixed(310076675.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-83472893.0/4294967296.0,1,-nbitq), 
to_sfixed(1202396015.0/4294967296.0,1,-nbitq), 
to_sfixed(683051288.0/4294967296.0,1,-nbitq), 
to_sfixed(996323433.0/4294967296.0,1,-nbitq), 
to_sfixed(467346578.0/4294967296.0,1,-nbitq), 
to_sfixed(-376857785.0/4294967296.0,1,-nbitq), 
to_sfixed(82043088.0/4294967296.0,1,-nbitq), 
to_sfixed(167734454.0/4294967296.0,1,-nbitq), 
to_sfixed(669263259.0/4294967296.0,1,-nbitq), 
to_sfixed(-287044501.0/4294967296.0,1,-nbitq), 
to_sfixed(-1251346399.0/4294967296.0,1,-nbitq), 
to_sfixed(259504543.0/4294967296.0,1,-nbitq), 
to_sfixed(-542867880.0/4294967296.0,1,-nbitq), 
to_sfixed(-967069128.0/4294967296.0,1,-nbitq), 
to_sfixed(492635567.0/4294967296.0,1,-nbitq), 
to_sfixed(-63341803.0/4294967296.0,1,-nbitq), 
to_sfixed(28495332.0/4294967296.0,1,-nbitq), 
to_sfixed(269655726.0/4294967296.0,1,-nbitq), 
to_sfixed(-546224343.0/4294967296.0,1,-nbitq), 
to_sfixed(-1106550946.0/4294967296.0,1,-nbitq), 
to_sfixed(-339188943.0/4294967296.0,1,-nbitq), 
to_sfixed(-258684268.0/4294967296.0,1,-nbitq), 
to_sfixed(352135941.0/4294967296.0,1,-nbitq), 
to_sfixed(-245430171.0/4294967296.0,1,-nbitq), 
to_sfixed(339167118.0/4294967296.0,1,-nbitq), 
to_sfixed(-343759998.0/4294967296.0,1,-nbitq), 
to_sfixed(-565738982.0/4294967296.0,1,-nbitq), 
to_sfixed(936120091.0/4294967296.0,1,-nbitq), 
to_sfixed(486484763.0/4294967296.0,1,-nbitq), 
to_sfixed(-804449284.0/4294967296.0,1,-nbitq), 
to_sfixed(461068810.0/4294967296.0,1,-nbitq), 
to_sfixed(-519364555.0/4294967296.0,1,-nbitq), 
to_sfixed(636549728.0/4294967296.0,1,-nbitq), 
to_sfixed(-425671498.0/4294967296.0,1,-nbitq), 
to_sfixed(-793497902.0/4294967296.0,1,-nbitq), 
to_sfixed(-1506120748.0/4294967296.0,1,-nbitq), 
to_sfixed(1063526333.0/4294967296.0,1,-nbitq), 
to_sfixed(-514399826.0/4294967296.0,1,-nbitq), 
to_sfixed(122389052.0/4294967296.0,1,-nbitq), 
to_sfixed(-181274605.0/4294967296.0,1,-nbitq), 
to_sfixed(-212545950.0/4294967296.0,1,-nbitq), 
to_sfixed(-976552514.0/4294967296.0,1,-nbitq), 
to_sfixed(29939544.0/4294967296.0,1,-nbitq), 
to_sfixed(388350100.0/4294967296.0,1,-nbitq), 
to_sfixed(2528562.0/4294967296.0,1,-nbitq), 
to_sfixed(-1715618166.0/4294967296.0,1,-nbitq), 
to_sfixed(-32793590.0/4294967296.0,1,-nbitq), 
to_sfixed(374217230.0/4294967296.0,1,-nbitq), 
to_sfixed(44484150.0/4294967296.0,1,-nbitq), 
to_sfixed(-941581579.0/4294967296.0,1,-nbitq), 
to_sfixed(-642463516.0/4294967296.0,1,-nbitq), 
to_sfixed(565051791.0/4294967296.0,1,-nbitq), 
to_sfixed(-1264868847.0/4294967296.0,1,-nbitq), 
to_sfixed(770379404.0/4294967296.0,1,-nbitq), 
to_sfixed(-213417932.0/4294967296.0,1,-nbitq), 
to_sfixed(-222473696.0/4294967296.0,1,-nbitq), 
to_sfixed(-772365471.0/4294967296.0,1,-nbitq), 
to_sfixed(91338853.0/4294967296.0,1,-nbitq), 
to_sfixed(115426965.0/4294967296.0,1,-nbitq), 
to_sfixed(347129058.0/4294967296.0,1,-nbitq), 
to_sfixed(413843637.0/4294967296.0,1,-nbitq), 
to_sfixed(-681262713.0/4294967296.0,1,-nbitq), 
to_sfixed(315300789.0/4294967296.0,1,-nbitq), 
to_sfixed(-110000919.0/4294967296.0,1,-nbitq), 
to_sfixed(-571770240.0/4294967296.0,1,-nbitq), 
to_sfixed(90171169.0/4294967296.0,1,-nbitq), 
to_sfixed(-539685851.0/4294967296.0,1,-nbitq), 
to_sfixed(-536001688.0/4294967296.0,1,-nbitq), 
to_sfixed(267271093.0/4294967296.0,1,-nbitq), 
to_sfixed(210713165.0/4294967296.0,1,-nbitq), 
to_sfixed(-1573267216.0/4294967296.0,1,-nbitq), 
to_sfixed(-219068370.0/4294967296.0,1,-nbitq), 
to_sfixed(555429893.0/4294967296.0,1,-nbitq), 
to_sfixed(273722364.0/4294967296.0,1,-nbitq), 
to_sfixed(-207908337.0/4294967296.0,1,-nbitq), 
to_sfixed(-417019583.0/4294967296.0,1,-nbitq), 
to_sfixed(-866438327.0/4294967296.0,1,-nbitq), 
to_sfixed(-739372833.0/4294967296.0,1,-nbitq), 
to_sfixed(311312940.0/4294967296.0,1,-nbitq), 
to_sfixed(-82883052.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-20406019.0/4294967296.0,1,-nbitq), 
to_sfixed(869755392.0/4294967296.0,1,-nbitq), 
to_sfixed(701982342.0/4294967296.0,1,-nbitq), 
to_sfixed(1306402919.0/4294967296.0,1,-nbitq), 
to_sfixed(-325961957.0/4294967296.0,1,-nbitq), 
to_sfixed(-365877484.0/4294967296.0,1,-nbitq), 
to_sfixed(-315248092.0/4294967296.0,1,-nbitq), 
to_sfixed(-514621274.0/4294967296.0,1,-nbitq), 
to_sfixed(782253423.0/4294967296.0,1,-nbitq), 
to_sfixed(120001360.0/4294967296.0,1,-nbitq), 
to_sfixed(-1209031964.0/4294967296.0,1,-nbitq), 
to_sfixed(33707775.0/4294967296.0,1,-nbitq), 
to_sfixed(-885714543.0/4294967296.0,1,-nbitq), 
to_sfixed(-943530299.0/4294967296.0,1,-nbitq), 
to_sfixed(-160520355.0/4294967296.0,1,-nbitq), 
to_sfixed(-243808959.0/4294967296.0,1,-nbitq), 
to_sfixed(-271033386.0/4294967296.0,1,-nbitq), 
to_sfixed(-71357395.0/4294967296.0,1,-nbitq), 
to_sfixed(-522363971.0/4294967296.0,1,-nbitq), 
to_sfixed(-1126588493.0/4294967296.0,1,-nbitq), 
to_sfixed(66529024.0/4294967296.0,1,-nbitq), 
to_sfixed(402085673.0/4294967296.0,1,-nbitq), 
to_sfixed(-2710180.0/4294967296.0,1,-nbitq), 
to_sfixed(973324992.0/4294967296.0,1,-nbitq), 
to_sfixed(347109750.0/4294967296.0,1,-nbitq), 
to_sfixed(-217659353.0/4294967296.0,1,-nbitq), 
to_sfixed(-624820177.0/4294967296.0,1,-nbitq), 
to_sfixed(878120879.0/4294967296.0,1,-nbitq), 
to_sfixed(1096706758.0/4294967296.0,1,-nbitq), 
to_sfixed(-1029399968.0/4294967296.0,1,-nbitq), 
to_sfixed(1083890010.0/4294967296.0,1,-nbitq), 
to_sfixed(-116345495.0/4294967296.0,1,-nbitq), 
to_sfixed(541808214.0/4294967296.0,1,-nbitq), 
to_sfixed(-827595590.0/4294967296.0,1,-nbitq), 
to_sfixed(-484711047.0/4294967296.0,1,-nbitq), 
to_sfixed(-1097122341.0/4294967296.0,1,-nbitq), 
to_sfixed(593549516.0/4294967296.0,1,-nbitq), 
to_sfixed(-928828806.0/4294967296.0,1,-nbitq), 
to_sfixed(58175937.0/4294967296.0,1,-nbitq), 
to_sfixed(353127803.0/4294967296.0,1,-nbitq), 
to_sfixed(725309620.0/4294967296.0,1,-nbitq), 
to_sfixed(-344934765.0/4294967296.0,1,-nbitq), 
to_sfixed(828479117.0/4294967296.0,1,-nbitq), 
to_sfixed(170993275.0/4294967296.0,1,-nbitq), 
to_sfixed(629633203.0/4294967296.0,1,-nbitq), 
to_sfixed(-795289762.0/4294967296.0,1,-nbitq), 
to_sfixed(275125689.0/4294967296.0,1,-nbitq), 
to_sfixed(276102775.0/4294967296.0,1,-nbitq), 
to_sfixed(-634352362.0/4294967296.0,1,-nbitq), 
to_sfixed(-963700669.0/4294967296.0,1,-nbitq), 
to_sfixed(-745626609.0/4294967296.0,1,-nbitq), 
to_sfixed(52626105.0/4294967296.0,1,-nbitq), 
to_sfixed(-1007351436.0/4294967296.0,1,-nbitq), 
to_sfixed(697177287.0/4294967296.0,1,-nbitq), 
to_sfixed(-285857057.0/4294967296.0,1,-nbitq), 
to_sfixed(63793316.0/4294967296.0,1,-nbitq), 
to_sfixed(-699076256.0/4294967296.0,1,-nbitq), 
to_sfixed(312705390.0/4294967296.0,1,-nbitq), 
to_sfixed(142218943.0/4294967296.0,1,-nbitq), 
to_sfixed(208342915.0/4294967296.0,1,-nbitq), 
to_sfixed(477695572.0/4294967296.0,1,-nbitq), 
to_sfixed(-710348742.0/4294967296.0,1,-nbitq), 
to_sfixed(496351889.0/4294967296.0,1,-nbitq), 
to_sfixed(-334980613.0/4294967296.0,1,-nbitq), 
to_sfixed(178564995.0/4294967296.0,1,-nbitq), 
to_sfixed(183237226.0/4294967296.0,1,-nbitq), 
to_sfixed(697166765.0/4294967296.0,1,-nbitq), 
to_sfixed(-175312422.0/4294967296.0,1,-nbitq), 
to_sfixed(-173665627.0/4294967296.0,1,-nbitq), 
to_sfixed(836530674.0/4294967296.0,1,-nbitq), 
to_sfixed(-2276532882.0/4294967296.0,1,-nbitq), 
to_sfixed(540625288.0/4294967296.0,1,-nbitq), 
to_sfixed(734126634.0/4294967296.0,1,-nbitq), 
to_sfixed(199472469.0/4294967296.0,1,-nbitq), 
to_sfixed(172299912.0/4294967296.0,1,-nbitq), 
to_sfixed(-680979099.0/4294967296.0,1,-nbitq), 
to_sfixed(-46485205.0/4294967296.0,1,-nbitq), 
to_sfixed(89568939.0/4294967296.0,1,-nbitq), 
to_sfixed(373600746.0/4294967296.0,1,-nbitq), 
to_sfixed(-216813286.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-314239399.0/4294967296.0,1,-nbitq), 
to_sfixed(-336138311.0/4294967296.0,1,-nbitq), 
to_sfixed(-1458256629.0/4294967296.0,1,-nbitq), 
to_sfixed(910926752.0/4294967296.0,1,-nbitq), 
to_sfixed(-654638734.0/4294967296.0,1,-nbitq), 
to_sfixed(229385868.0/4294967296.0,1,-nbitq), 
to_sfixed(-6748215.0/4294967296.0,1,-nbitq), 
to_sfixed(-888735755.0/4294967296.0,1,-nbitq), 
to_sfixed(333577037.0/4294967296.0,1,-nbitq), 
to_sfixed(-208883833.0/4294967296.0,1,-nbitq), 
to_sfixed(-947989877.0/4294967296.0,1,-nbitq), 
to_sfixed(1005735019.0/4294967296.0,1,-nbitq), 
to_sfixed(-221311334.0/4294967296.0,1,-nbitq), 
to_sfixed(-745421084.0/4294967296.0,1,-nbitq), 
to_sfixed(140583956.0/4294967296.0,1,-nbitq), 
to_sfixed(-484683330.0/4294967296.0,1,-nbitq), 
to_sfixed(-22839441.0/4294967296.0,1,-nbitq), 
to_sfixed(250598735.0/4294967296.0,1,-nbitq), 
to_sfixed(808627212.0/4294967296.0,1,-nbitq), 
to_sfixed(-849567972.0/4294967296.0,1,-nbitq), 
to_sfixed(-238708115.0/4294967296.0,1,-nbitq), 
to_sfixed(-180464286.0/4294967296.0,1,-nbitq), 
to_sfixed(1201398864.0/4294967296.0,1,-nbitq), 
to_sfixed(521129354.0/4294967296.0,1,-nbitq), 
to_sfixed(340139842.0/4294967296.0,1,-nbitq), 
to_sfixed(640979426.0/4294967296.0,1,-nbitq), 
to_sfixed(-469884287.0/4294967296.0,1,-nbitq), 
to_sfixed(430552907.0/4294967296.0,1,-nbitq), 
to_sfixed(-76284254.0/4294967296.0,1,-nbitq), 
to_sfixed(-853132488.0/4294967296.0,1,-nbitq), 
to_sfixed(1403767532.0/4294967296.0,1,-nbitq), 
to_sfixed(-292758572.0/4294967296.0,1,-nbitq), 
to_sfixed(662768449.0/4294967296.0,1,-nbitq), 
to_sfixed(-1192376911.0/4294967296.0,1,-nbitq), 
to_sfixed(-95833202.0/4294967296.0,1,-nbitq), 
to_sfixed(1200615407.0/4294967296.0,1,-nbitq), 
to_sfixed(7985730.0/4294967296.0,1,-nbitq), 
to_sfixed(-599022663.0/4294967296.0,1,-nbitq), 
to_sfixed(-343542701.0/4294967296.0,1,-nbitq), 
to_sfixed(118596014.0/4294967296.0,1,-nbitq), 
to_sfixed(215061169.0/4294967296.0,1,-nbitq), 
to_sfixed(377433934.0/4294967296.0,1,-nbitq), 
to_sfixed(831272270.0/4294967296.0,1,-nbitq), 
to_sfixed(-208653055.0/4294967296.0,1,-nbitq), 
to_sfixed(-76175250.0/4294967296.0,1,-nbitq), 
to_sfixed(-1464222189.0/4294967296.0,1,-nbitq), 
to_sfixed(-48885812.0/4294967296.0,1,-nbitq), 
to_sfixed(694751384.0/4294967296.0,1,-nbitq), 
to_sfixed(-448161055.0/4294967296.0,1,-nbitq), 
to_sfixed(-1004446983.0/4294967296.0,1,-nbitq), 
to_sfixed(-476314165.0/4294967296.0,1,-nbitq), 
to_sfixed(620573437.0/4294967296.0,1,-nbitq), 
to_sfixed(-1593630355.0/4294967296.0,1,-nbitq), 
to_sfixed(182946618.0/4294967296.0,1,-nbitq), 
to_sfixed(10156284.0/4294967296.0,1,-nbitq), 
to_sfixed(-763158152.0/4294967296.0,1,-nbitq), 
to_sfixed(-416561328.0/4294967296.0,1,-nbitq), 
to_sfixed(1140206126.0/4294967296.0,1,-nbitq), 
to_sfixed(55088142.0/4294967296.0,1,-nbitq), 
to_sfixed(-333610770.0/4294967296.0,1,-nbitq), 
to_sfixed(31989552.0/4294967296.0,1,-nbitq), 
to_sfixed(-985135838.0/4294967296.0,1,-nbitq), 
to_sfixed(40855802.0/4294967296.0,1,-nbitq), 
to_sfixed(-689114822.0/4294967296.0,1,-nbitq), 
to_sfixed(420738404.0/4294967296.0,1,-nbitq), 
to_sfixed(325738224.0/4294967296.0,1,-nbitq), 
to_sfixed(1790577902.0/4294967296.0,1,-nbitq), 
to_sfixed(-229757610.0/4294967296.0,1,-nbitq), 
to_sfixed(156465107.0/4294967296.0,1,-nbitq), 
to_sfixed(476670889.0/4294967296.0,1,-nbitq), 
to_sfixed(-1255116413.0/4294967296.0,1,-nbitq), 
to_sfixed(78320479.0/4294967296.0,1,-nbitq), 
to_sfixed(392150099.0/4294967296.0,1,-nbitq), 
to_sfixed(143563701.0/4294967296.0,1,-nbitq), 
to_sfixed(-167103937.0/4294967296.0,1,-nbitq), 
to_sfixed(-685016376.0/4294967296.0,1,-nbitq), 
to_sfixed(194534624.0/4294967296.0,1,-nbitq), 
to_sfixed(348289079.0/4294967296.0,1,-nbitq), 
to_sfixed(56776229.0/4294967296.0,1,-nbitq), 
to_sfixed(-55698979.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-266648836.0/4294967296.0,1,-nbitq), 
to_sfixed(-260502490.0/4294967296.0,1,-nbitq), 
to_sfixed(-1593856301.0/4294967296.0,1,-nbitq), 
to_sfixed(891307232.0/4294967296.0,1,-nbitq), 
to_sfixed(-1170046000.0/4294967296.0,1,-nbitq), 
to_sfixed(52614740.0/4294967296.0,1,-nbitq), 
to_sfixed(371203918.0/4294967296.0,1,-nbitq), 
to_sfixed(-1368571810.0/4294967296.0,1,-nbitq), 
to_sfixed(594315320.0/4294967296.0,1,-nbitq), 
to_sfixed(34232925.0/4294967296.0,1,-nbitq), 
to_sfixed(-1045114856.0/4294967296.0,1,-nbitq), 
to_sfixed(507736191.0/4294967296.0,1,-nbitq), 
to_sfixed(-365264661.0/4294967296.0,1,-nbitq), 
to_sfixed(-173123233.0/4294967296.0,1,-nbitq), 
to_sfixed(-250587758.0/4294967296.0,1,-nbitq), 
to_sfixed(-266598279.0/4294967296.0,1,-nbitq), 
to_sfixed(-245873141.0/4294967296.0,1,-nbitq), 
to_sfixed(290755166.0/4294967296.0,1,-nbitq), 
to_sfixed(2083002204.0/4294967296.0,1,-nbitq), 
to_sfixed(-1212284683.0/4294967296.0,1,-nbitq), 
to_sfixed(-291367746.0/4294967296.0,1,-nbitq), 
to_sfixed(-190865342.0/4294967296.0,1,-nbitq), 
to_sfixed(1139192776.0/4294967296.0,1,-nbitq), 
to_sfixed(306344277.0/4294967296.0,1,-nbitq), 
to_sfixed(-292109766.0/4294967296.0,1,-nbitq), 
to_sfixed(77995163.0/4294967296.0,1,-nbitq), 
to_sfixed(-127411475.0/4294967296.0,1,-nbitq), 
to_sfixed(-1045501361.0/4294967296.0,1,-nbitq), 
to_sfixed(-1345593187.0/4294967296.0,1,-nbitq), 
to_sfixed(-1290543305.0/4294967296.0,1,-nbitq), 
to_sfixed(1114331152.0/4294967296.0,1,-nbitq), 
to_sfixed(-1027741016.0/4294967296.0,1,-nbitq), 
to_sfixed(104167375.0/4294967296.0,1,-nbitq), 
to_sfixed(-1238179689.0/4294967296.0,1,-nbitq), 
to_sfixed(128868012.0/4294967296.0,1,-nbitq), 
to_sfixed(1021976414.0/4294967296.0,1,-nbitq), 
to_sfixed(143782781.0/4294967296.0,1,-nbitq), 
to_sfixed(-950507045.0/4294967296.0,1,-nbitq), 
to_sfixed(-614962012.0/4294967296.0,1,-nbitq), 
to_sfixed(-99053952.0/4294967296.0,1,-nbitq), 
to_sfixed(-274928604.0/4294967296.0,1,-nbitq), 
to_sfixed(126578389.0/4294967296.0,1,-nbitq), 
to_sfixed(1454918294.0/4294967296.0,1,-nbitq), 
to_sfixed(-171323856.0/4294967296.0,1,-nbitq), 
to_sfixed(128723115.0/4294967296.0,1,-nbitq), 
to_sfixed(-287330194.0/4294967296.0,1,-nbitq), 
to_sfixed(66054118.0/4294967296.0,1,-nbitq), 
to_sfixed(537304399.0/4294967296.0,1,-nbitq), 
to_sfixed(144836005.0/4294967296.0,1,-nbitq), 
to_sfixed(-773965175.0/4294967296.0,1,-nbitq), 
to_sfixed(-152515054.0/4294967296.0,1,-nbitq), 
to_sfixed(450025845.0/4294967296.0,1,-nbitq), 
to_sfixed(-1185641084.0/4294967296.0,1,-nbitq), 
to_sfixed(-347239948.0/4294967296.0,1,-nbitq), 
to_sfixed(-32663755.0/4294967296.0,1,-nbitq), 
to_sfixed(-939842686.0/4294967296.0,1,-nbitq), 
to_sfixed(-983217900.0/4294967296.0,1,-nbitq), 
to_sfixed(-156196378.0/4294967296.0,1,-nbitq), 
to_sfixed(-345846058.0/4294967296.0,1,-nbitq), 
to_sfixed(184556305.0/4294967296.0,1,-nbitq), 
to_sfixed(108904204.0/4294967296.0,1,-nbitq), 
to_sfixed(-640136190.0/4294967296.0,1,-nbitq), 
to_sfixed(-70869612.0/4294967296.0,1,-nbitq), 
to_sfixed(-362326274.0/4294967296.0,1,-nbitq), 
to_sfixed(200957231.0/4294967296.0,1,-nbitq), 
to_sfixed(80842952.0/4294967296.0,1,-nbitq), 
to_sfixed(-89177937.0/4294967296.0,1,-nbitq), 
to_sfixed(658441765.0/4294967296.0,1,-nbitq), 
to_sfixed(-381529057.0/4294967296.0,1,-nbitq), 
to_sfixed(-600493344.0/4294967296.0,1,-nbitq), 
to_sfixed(-1497208496.0/4294967296.0,1,-nbitq), 
to_sfixed(-203819438.0/4294967296.0,1,-nbitq), 
to_sfixed(142875037.0/4294967296.0,1,-nbitq), 
to_sfixed(-241696416.0/4294967296.0,1,-nbitq), 
to_sfixed(-61478203.0/4294967296.0,1,-nbitq), 
to_sfixed(322080862.0/4294967296.0,1,-nbitq), 
to_sfixed(-193151972.0/4294967296.0,1,-nbitq), 
to_sfixed(309463853.0/4294967296.0,1,-nbitq), 
to_sfixed(-142887290.0/4294967296.0,1,-nbitq), 
to_sfixed(390880458.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-598880761.0/4294967296.0,1,-nbitq), 
to_sfixed(106007983.0/4294967296.0,1,-nbitq), 
to_sfixed(-1332572623.0/4294967296.0,1,-nbitq), 
to_sfixed(150228704.0/4294967296.0,1,-nbitq), 
to_sfixed(-507015551.0/4294967296.0,1,-nbitq), 
to_sfixed(-251856362.0/4294967296.0,1,-nbitq), 
to_sfixed(301911269.0/4294967296.0,1,-nbitq), 
to_sfixed(-415568721.0/4294967296.0,1,-nbitq), 
to_sfixed(1219346475.0/4294967296.0,1,-nbitq), 
to_sfixed(108030592.0/4294967296.0,1,-nbitq), 
to_sfixed(-716068834.0/4294967296.0,1,-nbitq), 
to_sfixed(46844930.0/4294967296.0,1,-nbitq), 
to_sfixed(-770223352.0/4294967296.0,1,-nbitq), 
to_sfixed(-52251816.0/4294967296.0,1,-nbitq), 
to_sfixed(-226658798.0/4294967296.0,1,-nbitq), 
to_sfixed(42676340.0/4294967296.0,1,-nbitq), 
to_sfixed(-4383509.0/4294967296.0,1,-nbitq), 
to_sfixed(-69668741.0/4294967296.0,1,-nbitq), 
to_sfixed(653928107.0/4294967296.0,1,-nbitq), 
to_sfixed(-1125416907.0/4294967296.0,1,-nbitq), 
to_sfixed(67688104.0/4294967296.0,1,-nbitq), 
to_sfixed(-1016159507.0/4294967296.0,1,-nbitq), 
to_sfixed(801788630.0/4294967296.0,1,-nbitq), 
to_sfixed(887130087.0/4294967296.0,1,-nbitq), 
to_sfixed(248834475.0/4294967296.0,1,-nbitq), 
to_sfixed(-229659451.0/4294967296.0,1,-nbitq), 
to_sfixed(-878910032.0/4294967296.0,1,-nbitq), 
to_sfixed(-1261022318.0/4294967296.0,1,-nbitq), 
to_sfixed(-355328387.0/4294967296.0,1,-nbitq), 
to_sfixed(-482523647.0/4294967296.0,1,-nbitq), 
to_sfixed(-280345087.0/4294967296.0,1,-nbitq), 
to_sfixed(256500161.0/4294967296.0,1,-nbitq), 
to_sfixed(-1137022670.0/4294967296.0,1,-nbitq), 
to_sfixed(-313034274.0/4294967296.0,1,-nbitq), 
to_sfixed(-243563213.0/4294967296.0,1,-nbitq), 
to_sfixed(647511464.0/4294967296.0,1,-nbitq), 
to_sfixed(226718752.0/4294967296.0,1,-nbitq), 
to_sfixed(-635452016.0/4294967296.0,1,-nbitq), 
to_sfixed(-721864925.0/4294967296.0,1,-nbitq), 
to_sfixed(255727369.0/4294967296.0,1,-nbitq), 
to_sfixed(-99047537.0/4294967296.0,1,-nbitq), 
to_sfixed(-401396494.0/4294967296.0,1,-nbitq), 
to_sfixed(-2672305.0/4294967296.0,1,-nbitq), 
to_sfixed(-466630518.0/4294967296.0,1,-nbitq), 
to_sfixed(240412594.0/4294967296.0,1,-nbitq), 
to_sfixed(-443860228.0/4294967296.0,1,-nbitq), 
to_sfixed(316457129.0/4294967296.0,1,-nbitq), 
to_sfixed(652751394.0/4294967296.0,1,-nbitq), 
to_sfixed(93399578.0/4294967296.0,1,-nbitq), 
to_sfixed(41048270.0/4294967296.0,1,-nbitq), 
to_sfixed(204875966.0/4294967296.0,1,-nbitq), 
to_sfixed(-551701141.0/4294967296.0,1,-nbitq), 
to_sfixed(-456287666.0/4294967296.0,1,-nbitq), 
to_sfixed(-954554627.0/4294967296.0,1,-nbitq), 
to_sfixed(1301195036.0/4294967296.0,1,-nbitq), 
to_sfixed(-495437611.0/4294967296.0,1,-nbitq), 
to_sfixed(-557757464.0/4294967296.0,1,-nbitq), 
to_sfixed(-486092338.0/4294967296.0,1,-nbitq), 
to_sfixed(117504212.0/4294967296.0,1,-nbitq), 
to_sfixed(-245975513.0/4294967296.0,1,-nbitq), 
to_sfixed(289227436.0/4294967296.0,1,-nbitq), 
to_sfixed(-495259378.0/4294967296.0,1,-nbitq), 
to_sfixed(394144453.0/4294967296.0,1,-nbitq), 
to_sfixed(-123387299.0/4294967296.0,1,-nbitq), 
to_sfixed(-173129351.0/4294967296.0,1,-nbitq), 
to_sfixed(398843679.0/4294967296.0,1,-nbitq), 
to_sfixed(-549938973.0/4294967296.0,1,-nbitq), 
to_sfixed(33424587.0/4294967296.0,1,-nbitq), 
to_sfixed(143672623.0/4294967296.0,1,-nbitq), 
to_sfixed(63220618.0/4294967296.0,1,-nbitq), 
to_sfixed(-160407332.0/4294967296.0,1,-nbitq), 
to_sfixed(253491512.0/4294967296.0,1,-nbitq), 
to_sfixed(70896025.0/4294967296.0,1,-nbitq), 
to_sfixed(442945087.0/4294967296.0,1,-nbitq), 
to_sfixed(126645509.0/4294967296.0,1,-nbitq), 
to_sfixed(1228981295.0/4294967296.0,1,-nbitq), 
to_sfixed(-347070188.0/4294967296.0,1,-nbitq), 
to_sfixed(120279657.0/4294967296.0,1,-nbitq), 
to_sfixed(-345799821.0/4294967296.0,1,-nbitq), 
to_sfixed(-12657499.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(63923674.0/4294967296.0,1,-nbitq), 
to_sfixed(-237536445.0/4294967296.0,1,-nbitq), 
to_sfixed(147482251.0/4294967296.0,1,-nbitq), 
to_sfixed(-252372861.0/4294967296.0,1,-nbitq), 
to_sfixed(563582414.0/4294967296.0,1,-nbitq), 
to_sfixed(-42480446.0/4294967296.0,1,-nbitq), 
to_sfixed(579643678.0/4294967296.0,1,-nbitq), 
to_sfixed(-237709327.0/4294967296.0,1,-nbitq), 
to_sfixed(-8154900.0/4294967296.0,1,-nbitq), 
to_sfixed(-328184130.0/4294967296.0,1,-nbitq), 
to_sfixed(-423910284.0/4294967296.0,1,-nbitq), 
to_sfixed(599702524.0/4294967296.0,1,-nbitq), 
to_sfixed(-462291034.0/4294967296.0,1,-nbitq), 
to_sfixed(-27875394.0/4294967296.0,1,-nbitq), 
to_sfixed(-266058107.0/4294967296.0,1,-nbitq), 
to_sfixed(569487381.0/4294967296.0,1,-nbitq), 
to_sfixed(-309111526.0/4294967296.0,1,-nbitq), 
to_sfixed(-239923886.0/4294967296.0,1,-nbitq), 
to_sfixed(33529146.0/4294967296.0,1,-nbitq), 
to_sfixed(-661167932.0/4294967296.0,1,-nbitq), 
to_sfixed(55929106.0/4294967296.0,1,-nbitq), 
to_sfixed(-74190716.0/4294967296.0,1,-nbitq), 
to_sfixed(667751426.0/4294967296.0,1,-nbitq), 
to_sfixed(-136026217.0/4294967296.0,1,-nbitq), 
to_sfixed(-83230593.0/4294967296.0,1,-nbitq), 
to_sfixed(198934893.0/4294967296.0,1,-nbitq), 
to_sfixed(-580938846.0/4294967296.0,1,-nbitq), 
to_sfixed(-748193686.0/4294967296.0,1,-nbitq), 
to_sfixed(-111492730.0/4294967296.0,1,-nbitq), 
to_sfixed(-903892556.0/4294967296.0,1,-nbitq), 
to_sfixed(-355834038.0/4294967296.0,1,-nbitq), 
to_sfixed(130231484.0/4294967296.0,1,-nbitq), 
to_sfixed(-1241553288.0/4294967296.0,1,-nbitq), 
to_sfixed(530213573.0/4294967296.0,1,-nbitq), 
to_sfixed(843585532.0/4294967296.0,1,-nbitq), 
to_sfixed(46813475.0/4294967296.0,1,-nbitq), 
to_sfixed(-230737839.0/4294967296.0,1,-nbitq), 
to_sfixed(-285511939.0/4294967296.0,1,-nbitq), 
to_sfixed(-889564522.0/4294967296.0,1,-nbitq), 
to_sfixed(91100755.0/4294967296.0,1,-nbitq), 
to_sfixed(53247866.0/4294967296.0,1,-nbitq), 
to_sfixed(-330314596.0/4294967296.0,1,-nbitq), 
to_sfixed(-142301996.0/4294967296.0,1,-nbitq), 
to_sfixed(-175660467.0/4294967296.0,1,-nbitq), 
to_sfixed(414511041.0/4294967296.0,1,-nbitq), 
to_sfixed(-206814621.0/4294967296.0,1,-nbitq), 
to_sfixed(-105698860.0/4294967296.0,1,-nbitq), 
to_sfixed(343350863.0/4294967296.0,1,-nbitq), 
to_sfixed(-116646113.0/4294967296.0,1,-nbitq), 
to_sfixed(-447610172.0/4294967296.0,1,-nbitq), 
to_sfixed(309004892.0/4294967296.0,1,-nbitq), 
to_sfixed(-64065836.0/4294967296.0,1,-nbitq), 
to_sfixed(-578523316.0/4294967296.0,1,-nbitq), 
to_sfixed(-1088444175.0/4294967296.0,1,-nbitq), 
to_sfixed(1326517609.0/4294967296.0,1,-nbitq), 
to_sfixed(-69704112.0/4294967296.0,1,-nbitq), 
to_sfixed(-611845661.0/4294967296.0,1,-nbitq), 
to_sfixed(-528339649.0/4294967296.0,1,-nbitq), 
to_sfixed(-31459958.0/4294967296.0,1,-nbitq), 
to_sfixed(289900999.0/4294967296.0,1,-nbitq), 
to_sfixed(-148560005.0/4294967296.0,1,-nbitq), 
to_sfixed(-754377378.0/4294967296.0,1,-nbitq), 
to_sfixed(15887475.0/4294967296.0,1,-nbitq), 
to_sfixed(317675748.0/4294967296.0,1,-nbitq), 
to_sfixed(-67515356.0/4294967296.0,1,-nbitq), 
to_sfixed(-230591461.0/4294967296.0,1,-nbitq), 
to_sfixed(-661988661.0/4294967296.0,1,-nbitq), 
to_sfixed(470011588.0/4294967296.0,1,-nbitq), 
to_sfixed(-56969289.0/4294967296.0,1,-nbitq), 
to_sfixed(-92298090.0/4294967296.0,1,-nbitq), 
to_sfixed(-798341740.0/4294967296.0,1,-nbitq), 
to_sfixed(336578235.0/4294967296.0,1,-nbitq), 
to_sfixed(-638635093.0/4294967296.0,1,-nbitq), 
to_sfixed(-309608265.0/4294967296.0,1,-nbitq), 
to_sfixed(237563204.0/4294967296.0,1,-nbitq), 
to_sfixed(645998349.0/4294967296.0,1,-nbitq), 
to_sfixed(-169599103.0/4294967296.0,1,-nbitq), 
to_sfixed(302282324.0/4294967296.0,1,-nbitq), 
to_sfixed(723417603.0/4294967296.0,1,-nbitq), 
to_sfixed(-17316573.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-130407561.0/4294967296.0,1,-nbitq), 
to_sfixed(-427331414.0/4294967296.0,1,-nbitq), 
to_sfixed(209316289.0/4294967296.0,1,-nbitq), 
to_sfixed(-243647469.0/4294967296.0,1,-nbitq), 
to_sfixed(-191446564.0/4294967296.0,1,-nbitq), 
to_sfixed(-609284659.0/4294967296.0,1,-nbitq), 
to_sfixed(410759735.0/4294967296.0,1,-nbitq), 
to_sfixed(453768510.0/4294967296.0,1,-nbitq), 
to_sfixed(211536457.0/4294967296.0,1,-nbitq), 
to_sfixed(-245891299.0/4294967296.0,1,-nbitq), 
to_sfixed(-197662467.0/4294967296.0,1,-nbitq), 
to_sfixed(245547406.0/4294967296.0,1,-nbitq), 
to_sfixed(-275656461.0/4294967296.0,1,-nbitq), 
to_sfixed(996569939.0/4294967296.0,1,-nbitq), 
to_sfixed(-388670492.0/4294967296.0,1,-nbitq), 
to_sfixed(413680191.0/4294967296.0,1,-nbitq), 
to_sfixed(-191031006.0/4294967296.0,1,-nbitq), 
to_sfixed(311745820.0/4294967296.0,1,-nbitq), 
to_sfixed(-213162941.0/4294967296.0,1,-nbitq), 
to_sfixed(-490267932.0/4294967296.0,1,-nbitq), 
to_sfixed(-315940208.0/4294967296.0,1,-nbitq), 
to_sfixed(-455099135.0/4294967296.0,1,-nbitq), 
to_sfixed(158785090.0/4294967296.0,1,-nbitq), 
to_sfixed(146874423.0/4294967296.0,1,-nbitq), 
to_sfixed(225862583.0/4294967296.0,1,-nbitq), 
to_sfixed(867661730.0/4294967296.0,1,-nbitq), 
to_sfixed(-340495459.0/4294967296.0,1,-nbitq), 
to_sfixed(-529096904.0/4294967296.0,1,-nbitq), 
to_sfixed(544968848.0/4294967296.0,1,-nbitq), 
to_sfixed(-1202291432.0/4294967296.0,1,-nbitq), 
to_sfixed(-441950245.0/4294967296.0,1,-nbitq), 
to_sfixed(-675616129.0/4294967296.0,1,-nbitq), 
to_sfixed(-1660290272.0/4294967296.0,1,-nbitq), 
to_sfixed(558402841.0/4294967296.0,1,-nbitq), 
to_sfixed(636946195.0/4294967296.0,1,-nbitq), 
to_sfixed(984014081.0/4294967296.0,1,-nbitq), 
to_sfixed(47313422.0/4294967296.0,1,-nbitq), 
to_sfixed(-67472607.0/4294967296.0,1,-nbitq), 
to_sfixed(-284114603.0/4294967296.0,1,-nbitq), 
to_sfixed(147248110.0/4294967296.0,1,-nbitq), 
to_sfixed(602954021.0/4294967296.0,1,-nbitq), 
to_sfixed(-293205555.0/4294967296.0,1,-nbitq), 
to_sfixed(-346994192.0/4294967296.0,1,-nbitq), 
to_sfixed(325126379.0/4294967296.0,1,-nbitq), 
to_sfixed(232734019.0/4294967296.0,1,-nbitq), 
to_sfixed(667479526.0/4294967296.0,1,-nbitq), 
to_sfixed(271841003.0/4294967296.0,1,-nbitq), 
to_sfixed(-534898136.0/4294967296.0,1,-nbitq), 
to_sfixed(-300951506.0/4294967296.0,1,-nbitq), 
to_sfixed(917422098.0/4294967296.0,1,-nbitq), 
to_sfixed(182330739.0/4294967296.0,1,-nbitq), 
to_sfixed(-492508766.0/4294967296.0,1,-nbitq), 
to_sfixed(-966463331.0/4294967296.0,1,-nbitq), 
to_sfixed(-56853677.0/4294967296.0,1,-nbitq), 
to_sfixed(736727279.0/4294967296.0,1,-nbitq), 
to_sfixed(421526175.0/4294967296.0,1,-nbitq), 
to_sfixed(-350897656.0/4294967296.0,1,-nbitq), 
to_sfixed(-689321080.0/4294967296.0,1,-nbitq), 
to_sfixed(277605808.0/4294967296.0,1,-nbitq), 
to_sfixed(-60002467.0/4294967296.0,1,-nbitq), 
to_sfixed(-377671091.0/4294967296.0,1,-nbitq), 
to_sfixed(-503015228.0/4294967296.0,1,-nbitq), 
to_sfixed(-373762261.0/4294967296.0,1,-nbitq), 
to_sfixed(13930250.0/4294967296.0,1,-nbitq), 
to_sfixed(-800876922.0/4294967296.0,1,-nbitq), 
to_sfixed(-194068065.0/4294967296.0,1,-nbitq), 
to_sfixed(-1714601153.0/4294967296.0,1,-nbitq), 
to_sfixed(1175627813.0/4294967296.0,1,-nbitq), 
to_sfixed(-266781183.0/4294967296.0,1,-nbitq), 
to_sfixed(-292573031.0/4294967296.0,1,-nbitq), 
to_sfixed(361495645.0/4294967296.0,1,-nbitq), 
to_sfixed(-403914985.0/4294967296.0,1,-nbitq), 
to_sfixed(72450501.0/4294967296.0,1,-nbitq), 
to_sfixed(-172935879.0/4294967296.0,1,-nbitq), 
to_sfixed(380495154.0/4294967296.0,1,-nbitq), 
to_sfixed(432334006.0/4294967296.0,1,-nbitq), 
to_sfixed(-376361391.0/4294967296.0,1,-nbitq), 
to_sfixed(502598394.0/4294967296.0,1,-nbitq), 
to_sfixed(1108569052.0/4294967296.0,1,-nbitq), 
to_sfixed(57862829.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-124211279.0/4294967296.0,1,-nbitq), 
to_sfixed(118559546.0/4294967296.0,1,-nbitq), 
to_sfixed(1226931114.0/4294967296.0,1,-nbitq), 
to_sfixed(-292516008.0/4294967296.0,1,-nbitq), 
to_sfixed(119502342.0/4294967296.0,1,-nbitq), 
to_sfixed(-587982795.0/4294967296.0,1,-nbitq), 
to_sfixed(618835744.0/4294967296.0,1,-nbitq), 
to_sfixed(-121411685.0/4294967296.0,1,-nbitq), 
to_sfixed(621604398.0/4294967296.0,1,-nbitq), 
to_sfixed(-56760152.0/4294967296.0,1,-nbitq), 
to_sfixed(-199214704.0/4294967296.0,1,-nbitq), 
to_sfixed(-76588231.0/4294967296.0,1,-nbitq), 
to_sfixed(121419392.0/4294967296.0,1,-nbitq), 
to_sfixed(468371249.0/4294967296.0,1,-nbitq), 
to_sfixed(-112643198.0/4294967296.0,1,-nbitq), 
to_sfixed(597601105.0/4294967296.0,1,-nbitq), 
to_sfixed(357177036.0/4294967296.0,1,-nbitq), 
to_sfixed(77965676.0/4294967296.0,1,-nbitq), 
to_sfixed(-132046092.0/4294967296.0,1,-nbitq), 
to_sfixed(-318493658.0/4294967296.0,1,-nbitq), 
to_sfixed(225445092.0/4294967296.0,1,-nbitq), 
to_sfixed(-526083566.0/4294967296.0,1,-nbitq), 
to_sfixed(-873336112.0/4294967296.0,1,-nbitq), 
to_sfixed(-316001934.0/4294967296.0,1,-nbitq), 
to_sfixed(261965181.0/4294967296.0,1,-nbitq), 
to_sfixed(636538736.0/4294967296.0,1,-nbitq), 
to_sfixed(-1044525844.0/4294967296.0,1,-nbitq), 
to_sfixed(494115370.0/4294967296.0,1,-nbitq), 
to_sfixed(113066884.0/4294967296.0,1,-nbitq), 
to_sfixed(-818663252.0/4294967296.0,1,-nbitq), 
to_sfixed(-271536414.0/4294967296.0,1,-nbitq), 
to_sfixed(-725585010.0/4294967296.0,1,-nbitq), 
to_sfixed(-1598333910.0/4294967296.0,1,-nbitq), 
to_sfixed(207547010.0/4294967296.0,1,-nbitq), 
to_sfixed(93307884.0/4294967296.0,1,-nbitq), 
to_sfixed(1011069118.0/4294967296.0,1,-nbitq), 
to_sfixed(239280063.0/4294967296.0,1,-nbitq), 
to_sfixed(522105323.0/4294967296.0,1,-nbitq), 
to_sfixed(142404581.0/4294967296.0,1,-nbitq), 
to_sfixed(125480853.0/4294967296.0,1,-nbitq), 
to_sfixed(764256058.0/4294967296.0,1,-nbitq), 
to_sfixed(40934935.0/4294967296.0,1,-nbitq), 
to_sfixed(-399869862.0/4294967296.0,1,-nbitq), 
to_sfixed(1462693267.0/4294967296.0,1,-nbitq), 
to_sfixed(469625392.0/4294967296.0,1,-nbitq), 
to_sfixed(951180424.0/4294967296.0,1,-nbitq), 
to_sfixed(-128444042.0/4294967296.0,1,-nbitq), 
to_sfixed(-992047580.0/4294967296.0,1,-nbitq), 
to_sfixed(-603991127.0/4294967296.0,1,-nbitq), 
to_sfixed(726069175.0/4294967296.0,1,-nbitq), 
to_sfixed(132527806.0/4294967296.0,1,-nbitq), 
to_sfixed(302089095.0/4294967296.0,1,-nbitq), 
to_sfixed(-1367572339.0/4294967296.0,1,-nbitq), 
to_sfixed(1009373872.0/4294967296.0,1,-nbitq), 
to_sfixed(178990963.0/4294967296.0,1,-nbitq), 
to_sfixed(338861660.0/4294967296.0,1,-nbitq), 
to_sfixed(300355941.0/4294967296.0,1,-nbitq), 
to_sfixed(-594158381.0/4294967296.0,1,-nbitq), 
to_sfixed(192849367.0/4294967296.0,1,-nbitq), 
to_sfixed(373900984.0/4294967296.0,1,-nbitq), 
to_sfixed(-666134404.0/4294967296.0,1,-nbitq), 
to_sfixed(-268437728.0/4294967296.0,1,-nbitq), 
to_sfixed(-1563498097.0/4294967296.0,1,-nbitq), 
to_sfixed(46095414.0/4294967296.0,1,-nbitq), 
to_sfixed(-613418175.0/4294967296.0,1,-nbitq), 
to_sfixed(-426674246.0/4294967296.0,1,-nbitq), 
to_sfixed(-1132170714.0/4294967296.0,1,-nbitq), 
to_sfixed(458717764.0/4294967296.0,1,-nbitq), 
to_sfixed(-218356083.0/4294967296.0,1,-nbitq), 
to_sfixed(-264420140.0/4294967296.0,1,-nbitq), 
to_sfixed(660104846.0/4294967296.0,1,-nbitq), 
to_sfixed(-424181300.0/4294967296.0,1,-nbitq), 
to_sfixed(294485232.0/4294967296.0,1,-nbitq), 
to_sfixed(335675787.0/4294967296.0,1,-nbitq), 
to_sfixed(493076809.0/4294967296.0,1,-nbitq), 
to_sfixed(501025102.0/4294967296.0,1,-nbitq), 
to_sfixed(180681185.0/4294967296.0,1,-nbitq), 
to_sfixed(-186848986.0/4294967296.0,1,-nbitq), 
to_sfixed(906831498.0/4294967296.0,1,-nbitq), 
to_sfixed(-371154475.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(161781022.0/4294967296.0,1,-nbitq), 
to_sfixed(29568834.0/4294967296.0,1,-nbitq), 
to_sfixed(923196930.0/4294967296.0,1,-nbitq), 
to_sfixed(-660935403.0/4294967296.0,1,-nbitq), 
to_sfixed(-112723931.0/4294967296.0,1,-nbitq), 
to_sfixed(-723390214.0/4294967296.0,1,-nbitq), 
to_sfixed(413097035.0/4294967296.0,1,-nbitq), 
to_sfixed(460399306.0/4294967296.0,1,-nbitq), 
to_sfixed(617485225.0/4294967296.0,1,-nbitq), 
to_sfixed(270818131.0/4294967296.0,1,-nbitq), 
to_sfixed(-391301453.0/4294967296.0,1,-nbitq), 
to_sfixed(-341146635.0/4294967296.0,1,-nbitq), 
to_sfixed(132616195.0/4294967296.0,1,-nbitq), 
to_sfixed(678705324.0/4294967296.0,1,-nbitq), 
to_sfixed(-244188406.0/4294967296.0,1,-nbitq), 
to_sfixed(588078114.0/4294967296.0,1,-nbitq), 
to_sfixed(-351314921.0/4294967296.0,1,-nbitq), 
to_sfixed(344473788.0/4294967296.0,1,-nbitq), 
to_sfixed(-297768879.0/4294967296.0,1,-nbitq), 
to_sfixed(-931823184.0/4294967296.0,1,-nbitq), 
to_sfixed(-191958105.0/4294967296.0,1,-nbitq), 
to_sfixed(101618301.0/4294967296.0,1,-nbitq), 
to_sfixed(-453947238.0/4294967296.0,1,-nbitq), 
to_sfixed(530044598.0/4294967296.0,1,-nbitq), 
to_sfixed(173441793.0/4294967296.0,1,-nbitq), 
to_sfixed(254695297.0/4294967296.0,1,-nbitq), 
to_sfixed(-630680097.0/4294967296.0,1,-nbitq), 
to_sfixed(425609827.0/4294967296.0,1,-nbitq), 
to_sfixed(495621072.0/4294967296.0,1,-nbitq), 
to_sfixed(-97704279.0/4294967296.0,1,-nbitq), 
to_sfixed(-645322898.0/4294967296.0,1,-nbitq), 
to_sfixed(-649740987.0/4294967296.0,1,-nbitq), 
to_sfixed(-2078872522.0/4294967296.0,1,-nbitq), 
to_sfixed(468899878.0/4294967296.0,1,-nbitq), 
to_sfixed(200991338.0/4294967296.0,1,-nbitq), 
to_sfixed(370959608.0/4294967296.0,1,-nbitq), 
to_sfixed(776793297.0/4294967296.0,1,-nbitq), 
to_sfixed(975797111.0/4294967296.0,1,-nbitq), 
to_sfixed(645083089.0/4294967296.0,1,-nbitq), 
to_sfixed(64832531.0/4294967296.0,1,-nbitq), 
to_sfixed(516289001.0/4294967296.0,1,-nbitq), 
to_sfixed(839231972.0/4294967296.0,1,-nbitq), 
to_sfixed(-724826471.0/4294967296.0,1,-nbitq), 
to_sfixed(1291417959.0/4294967296.0,1,-nbitq), 
to_sfixed(380218086.0/4294967296.0,1,-nbitq), 
to_sfixed(739997948.0/4294967296.0,1,-nbitq), 
to_sfixed(-345064308.0/4294967296.0,1,-nbitq), 
to_sfixed(-385945347.0/4294967296.0,1,-nbitq), 
to_sfixed(-842724919.0/4294967296.0,1,-nbitq), 
to_sfixed(491164238.0/4294967296.0,1,-nbitq), 
to_sfixed(257639645.0/4294967296.0,1,-nbitq), 
to_sfixed(296941597.0/4294967296.0,1,-nbitq), 
to_sfixed(-2096069263.0/4294967296.0,1,-nbitq), 
to_sfixed(482358907.0/4294967296.0,1,-nbitq), 
to_sfixed(-309239278.0/4294967296.0,1,-nbitq), 
to_sfixed(553819947.0/4294967296.0,1,-nbitq), 
to_sfixed(679442920.0/4294967296.0,1,-nbitq), 
to_sfixed(-6389823.0/4294967296.0,1,-nbitq), 
to_sfixed(282864646.0/4294967296.0,1,-nbitq), 
to_sfixed(-14478401.0/4294967296.0,1,-nbitq), 
to_sfixed(-325222452.0/4294967296.0,1,-nbitq), 
to_sfixed(295134989.0/4294967296.0,1,-nbitq), 
to_sfixed(-1224005083.0/4294967296.0,1,-nbitq), 
to_sfixed(-185734147.0/4294967296.0,1,-nbitq), 
to_sfixed(-476349450.0/4294967296.0,1,-nbitq), 
to_sfixed(-251786199.0/4294967296.0,1,-nbitq), 
to_sfixed(-611266543.0/4294967296.0,1,-nbitq), 
to_sfixed(266402114.0/4294967296.0,1,-nbitq), 
to_sfixed(70351870.0/4294967296.0,1,-nbitq), 
to_sfixed(-7259885.0/4294967296.0,1,-nbitq), 
to_sfixed(-115370747.0/4294967296.0,1,-nbitq), 
to_sfixed(-138575807.0/4294967296.0,1,-nbitq), 
to_sfixed(-675406470.0/4294967296.0,1,-nbitq), 
to_sfixed(103938807.0/4294967296.0,1,-nbitq), 
to_sfixed(51464149.0/4294967296.0,1,-nbitq), 
to_sfixed(106661865.0/4294967296.0,1,-nbitq), 
to_sfixed(144811698.0/4294967296.0,1,-nbitq), 
to_sfixed(82528551.0/4294967296.0,1,-nbitq), 
to_sfixed(622468969.0/4294967296.0,1,-nbitq), 
to_sfixed(-292184288.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(196021210.0/4294967296.0,1,-nbitq), 
to_sfixed(-335340145.0/4294967296.0,1,-nbitq), 
to_sfixed(780795088.0/4294967296.0,1,-nbitq), 
to_sfixed(-948999700.0/4294967296.0,1,-nbitq), 
to_sfixed(-397392435.0/4294967296.0,1,-nbitq), 
to_sfixed(-443976642.0/4294967296.0,1,-nbitq), 
to_sfixed(-24662573.0/4294967296.0,1,-nbitq), 
to_sfixed(170971300.0/4294967296.0,1,-nbitq), 
to_sfixed(203820085.0/4294967296.0,1,-nbitq), 
to_sfixed(157386428.0/4294967296.0,1,-nbitq), 
to_sfixed(-344386911.0/4294967296.0,1,-nbitq), 
to_sfixed(-133660154.0/4294967296.0,1,-nbitq), 
to_sfixed(-176214750.0/4294967296.0,1,-nbitq), 
to_sfixed(1765104199.0/4294967296.0,1,-nbitq), 
to_sfixed(-312123210.0/4294967296.0,1,-nbitq), 
to_sfixed(246436418.0/4294967296.0,1,-nbitq), 
to_sfixed(-143807112.0/4294967296.0,1,-nbitq), 
to_sfixed(321092930.0/4294967296.0,1,-nbitq), 
to_sfixed(-479721489.0/4294967296.0,1,-nbitq), 
to_sfixed(-863590308.0/4294967296.0,1,-nbitq), 
to_sfixed(-162363134.0/4294967296.0,1,-nbitq), 
to_sfixed(42214604.0/4294967296.0,1,-nbitq), 
to_sfixed(-690539929.0/4294967296.0,1,-nbitq), 
to_sfixed(704712077.0/4294967296.0,1,-nbitq), 
to_sfixed(17446199.0/4294967296.0,1,-nbitq), 
to_sfixed(-91931645.0/4294967296.0,1,-nbitq), 
to_sfixed(-503191549.0/4294967296.0,1,-nbitq), 
to_sfixed(699498850.0/4294967296.0,1,-nbitq), 
to_sfixed(-14783654.0/4294967296.0,1,-nbitq), 
to_sfixed(153345993.0/4294967296.0,1,-nbitq), 
to_sfixed(846839973.0/4294967296.0,1,-nbitq), 
to_sfixed(-481806331.0/4294967296.0,1,-nbitq), 
to_sfixed(-1869786825.0/4294967296.0,1,-nbitq), 
to_sfixed(145788884.0/4294967296.0,1,-nbitq), 
to_sfixed(409217727.0/4294967296.0,1,-nbitq), 
to_sfixed(1132487448.0/4294967296.0,1,-nbitq), 
to_sfixed(618806776.0/4294967296.0,1,-nbitq), 
to_sfixed(302059650.0/4294967296.0,1,-nbitq), 
to_sfixed(434580813.0/4294967296.0,1,-nbitq), 
to_sfixed(281192257.0/4294967296.0,1,-nbitq), 
to_sfixed(452030067.0/4294967296.0,1,-nbitq), 
to_sfixed(758440930.0/4294967296.0,1,-nbitq), 
to_sfixed(-714306901.0/4294967296.0,1,-nbitq), 
to_sfixed(1835650295.0/4294967296.0,1,-nbitq), 
to_sfixed(-26787364.0/4294967296.0,1,-nbitq), 
to_sfixed(721040086.0/4294967296.0,1,-nbitq), 
to_sfixed(327463139.0/4294967296.0,1,-nbitq), 
to_sfixed(198807160.0/4294967296.0,1,-nbitq), 
to_sfixed(-1022699268.0/4294967296.0,1,-nbitq), 
to_sfixed(366429852.0/4294967296.0,1,-nbitq), 
to_sfixed(40911427.0/4294967296.0,1,-nbitq), 
to_sfixed(175635828.0/4294967296.0,1,-nbitq), 
to_sfixed(-587501253.0/4294967296.0,1,-nbitq), 
to_sfixed(-208203676.0/4294967296.0,1,-nbitq), 
to_sfixed(-503998901.0/4294967296.0,1,-nbitq), 
to_sfixed(457921166.0/4294967296.0,1,-nbitq), 
to_sfixed(772555905.0/4294967296.0,1,-nbitq), 
to_sfixed(465854979.0/4294967296.0,1,-nbitq), 
to_sfixed(201579223.0/4294967296.0,1,-nbitq), 
to_sfixed(-96645397.0/4294967296.0,1,-nbitq), 
to_sfixed(-119570002.0/4294967296.0,1,-nbitq), 
to_sfixed(-20114246.0/4294967296.0,1,-nbitq), 
to_sfixed(-482987686.0/4294967296.0,1,-nbitq), 
to_sfixed(10413616.0/4294967296.0,1,-nbitq), 
to_sfixed(471480665.0/4294967296.0,1,-nbitq), 
to_sfixed(-73435406.0/4294967296.0,1,-nbitq), 
to_sfixed(88174527.0/4294967296.0,1,-nbitq), 
to_sfixed(43947742.0/4294967296.0,1,-nbitq), 
to_sfixed(187967233.0/4294967296.0,1,-nbitq), 
to_sfixed(-275167867.0/4294967296.0,1,-nbitq), 
to_sfixed(-8302703.0/4294967296.0,1,-nbitq), 
to_sfixed(-268323721.0/4294967296.0,1,-nbitq), 
to_sfixed(-451924743.0/4294967296.0,1,-nbitq), 
to_sfixed(308516594.0/4294967296.0,1,-nbitq), 
to_sfixed(-227024876.0/4294967296.0,1,-nbitq), 
to_sfixed(417845298.0/4294967296.0,1,-nbitq), 
to_sfixed(69905311.0/4294967296.0,1,-nbitq), 
to_sfixed(270931327.0/4294967296.0,1,-nbitq), 
to_sfixed(331494682.0/4294967296.0,1,-nbitq), 
to_sfixed(-267190854.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(83786010.0/4294967296.0,1,-nbitq), 
to_sfixed(-335451532.0/4294967296.0,1,-nbitq), 
to_sfixed(129220818.0/4294967296.0,1,-nbitq), 
to_sfixed(-392769892.0/4294967296.0,1,-nbitq), 
to_sfixed(-632170702.0/4294967296.0,1,-nbitq), 
to_sfixed(-484708700.0/4294967296.0,1,-nbitq), 
to_sfixed(173311963.0/4294967296.0,1,-nbitq), 
to_sfixed(-3157503.0/4294967296.0,1,-nbitq), 
to_sfixed(675816361.0/4294967296.0,1,-nbitq), 
to_sfixed(-115797263.0/4294967296.0,1,-nbitq), 
to_sfixed(-607518614.0/4294967296.0,1,-nbitq), 
to_sfixed(644338201.0/4294967296.0,1,-nbitq), 
to_sfixed(280683493.0/4294967296.0,1,-nbitq), 
to_sfixed(500712345.0/4294967296.0,1,-nbitq), 
to_sfixed(-287261660.0/4294967296.0,1,-nbitq), 
to_sfixed(-20440297.0/4294967296.0,1,-nbitq), 
to_sfixed(-405308205.0/4294967296.0,1,-nbitq), 
to_sfixed(117488658.0/4294967296.0,1,-nbitq), 
to_sfixed(-1193711606.0/4294967296.0,1,-nbitq), 
to_sfixed(-112878144.0/4294967296.0,1,-nbitq), 
to_sfixed(222550821.0/4294967296.0,1,-nbitq), 
to_sfixed(95157441.0/4294967296.0,1,-nbitq), 
to_sfixed(-622361575.0/4294967296.0,1,-nbitq), 
to_sfixed(130024734.0/4294967296.0,1,-nbitq), 
to_sfixed(94662740.0/4294967296.0,1,-nbitq), 
to_sfixed(-250784808.0/4294967296.0,1,-nbitq), 
to_sfixed(623011591.0/4294967296.0,1,-nbitq), 
to_sfixed(513086073.0/4294967296.0,1,-nbitq), 
to_sfixed(140953820.0/4294967296.0,1,-nbitq), 
to_sfixed(793759813.0/4294967296.0,1,-nbitq), 
to_sfixed(551058131.0/4294967296.0,1,-nbitq), 
to_sfixed(-69747321.0/4294967296.0,1,-nbitq), 
to_sfixed(-952623284.0/4294967296.0,1,-nbitq), 
to_sfixed(-644895831.0/4294967296.0,1,-nbitq), 
to_sfixed(530988327.0/4294967296.0,1,-nbitq), 
to_sfixed(732009213.0/4294967296.0,1,-nbitq), 
to_sfixed(64989784.0/4294967296.0,1,-nbitq), 
to_sfixed(170772332.0/4294967296.0,1,-nbitq), 
to_sfixed(-5614585.0/4294967296.0,1,-nbitq), 
to_sfixed(61035969.0/4294967296.0,1,-nbitq), 
to_sfixed(324400493.0/4294967296.0,1,-nbitq), 
to_sfixed(201265498.0/4294967296.0,1,-nbitq), 
to_sfixed(-959591351.0/4294967296.0,1,-nbitq), 
to_sfixed(783926825.0/4294967296.0,1,-nbitq), 
to_sfixed(-28037798.0/4294967296.0,1,-nbitq), 
to_sfixed(388399267.0/4294967296.0,1,-nbitq), 
to_sfixed(-275486776.0/4294967296.0,1,-nbitq), 
to_sfixed(-606013363.0/4294967296.0,1,-nbitq), 
to_sfixed(-535751318.0/4294967296.0,1,-nbitq), 
to_sfixed(-92787511.0/4294967296.0,1,-nbitq), 
to_sfixed(362268155.0/4294967296.0,1,-nbitq), 
to_sfixed(100817938.0/4294967296.0,1,-nbitq), 
to_sfixed(13752128.0/4294967296.0,1,-nbitq), 
to_sfixed(-156237004.0/4294967296.0,1,-nbitq), 
to_sfixed(-1090838331.0/4294967296.0,1,-nbitq), 
to_sfixed(571079429.0/4294967296.0,1,-nbitq), 
to_sfixed(-153115928.0/4294967296.0,1,-nbitq), 
to_sfixed(142209592.0/4294967296.0,1,-nbitq), 
to_sfixed(-95885047.0/4294967296.0,1,-nbitq), 
to_sfixed(96367479.0/4294967296.0,1,-nbitq), 
to_sfixed(19285563.0/4294967296.0,1,-nbitq), 
to_sfixed(-426204035.0/4294967296.0,1,-nbitq), 
to_sfixed(-146349155.0/4294967296.0,1,-nbitq), 
to_sfixed(-488648053.0/4294967296.0,1,-nbitq), 
to_sfixed(416437309.0/4294967296.0,1,-nbitq), 
to_sfixed(331727356.0/4294967296.0,1,-nbitq), 
to_sfixed(285499215.0/4294967296.0,1,-nbitq), 
to_sfixed(241545841.0/4294967296.0,1,-nbitq), 
to_sfixed(-206896097.0/4294967296.0,1,-nbitq), 
to_sfixed(255320032.0/4294967296.0,1,-nbitq), 
to_sfixed(244388731.0/4294967296.0,1,-nbitq), 
to_sfixed(143755517.0/4294967296.0,1,-nbitq), 
to_sfixed(197416694.0/4294967296.0,1,-nbitq), 
to_sfixed(237710420.0/4294967296.0,1,-nbitq), 
to_sfixed(183095870.0/4294967296.0,1,-nbitq), 
to_sfixed(112955112.0/4294967296.0,1,-nbitq), 
to_sfixed(-478536262.0/4294967296.0,1,-nbitq), 
to_sfixed(-165078506.0/4294967296.0,1,-nbitq), 
to_sfixed(597503544.0/4294967296.0,1,-nbitq), 
to_sfixed(-134963144.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-428297573.0/4294967296.0,1,-nbitq), 
to_sfixed(-355635181.0/4294967296.0,1,-nbitq), 
to_sfixed(276158691.0/4294967296.0,1,-nbitq), 
to_sfixed(53396475.0/4294967296.0,1,-nbitq), 
to_sfixed(-489248534.0/4294967296.0,1,-nbitq), 
to_sfixed(-265888178.0/4294967296.0,1,-nbitq), 
to_sfixed(-43457580.0/4294967296.0,1,-nbitq), 
to_sfixed(380160608.0/4294967296.0,1,-nbitq), 
to_sfixed(556892960.0/4294967296.0,1,-nbitq), 
to_sfixed(-157607112.0/4294967296.0,1,-nbitq), 
to_sfixed(20158415.0/4294967296.0,1,-nbitq), 
to_sfixed(-71231554.0/4294967296.0,1,-nbitq), 
to_sfixed(-115203250.0/4294967296.0,1,-nbitq), 
to_sfixed(1156502017.0/4294967296.0,1,-nbitq), 
to_sfixed(206896218.0/4294967296.0,1,-nbitq), 
to_sfixed(312960089.0/4294967296.0,1,-nbitq), 
to_sfixed(287690926.0/4294967296.0,1,-nbitq), 
to_sfixed(-197337254.0/4294967296.0,1,-nbitq), 
to_sfixed(-651813146.0/4294967296.0,1,-nbitq), 
to_sfixed(248185011.0/4294967296.0,1,-nbitq), 
to_sfixed(184788251.0/4294967296.0,1,-nbitq), 
to_sfixed(486630161.0/4294967296.0,1,-nbitq), 
to_sfixed(-368613818.0/4294967296.0,1,-nbitq), 
to_sfixed(1481275745.0/4294967296.0,1,-nbitq), 
to_sfixed(198098269.0/4294967296.0,1,-nbitq), 
to_sfixed(-83991316.0/4294967296.0,1,-nbitq), 
to_sfixed(524342942.0/4294967296.0,1,-nbitq), 
to_sfixed(171748367.0/4294967296.0,1,-nbitq), 
to_sfixed(381927044.0/4294967296.0,1,-nbitq), 
to_sfixed(9407436.0/4294967296.0,1,-nbitq), 
to_sfixed(1194416069.0/4294967296.0,1,-nbitq), 
to_sfixed(311085539.0/4294967296.0,1,-nbitq), 
to_sfixed(-975908254.0/4294967296.0,1,-nbitq), 
to_sfixed(104251096.0/4294967296.0,1,-nbitq), 
to_sfixed(624476497.0/4294967296.0,1,-nbitq), 
to_sfixed(360770762.0/4294967296.0,1,-nbitq), 
to_sfixed(279998799.0/4294967296.0,1,-nbitq), 
to_sfixed(558632047.0/4294967296.0,1,-nbitq), 
to_sfixed(177669622.0/4294967296.0,1,-nbitq), 
to_sfixed(-120921068.0/4294967296.0,1,-nbitq), 
to_sfixed(93052089.0/4294967296.0,1,-nbitq), 
to_sfixed(-330107324.0/4294967296.0,1,-nbitq), 
to_sfixed(37882811.0/4294967296.0,1,-nbitq), 
to_sfixed(297798170.0/4294967296.0,1,-nbitq), 
to_sfixed(162999468.0/4294967296.0,1,-nbitq), 
to_sfixed(-228352066.0/4294967296.0,1,-nbitq), 
to_sfixed(37958023.0/4294967296.0,1,-nbitq), 
to_sfixed(-313168560.0/4294967296.0,1,-nbitq), 
to_sfixed(-393685056.0/4294967296.0,1,-nbitq), 
to_sfixed(-314888909.0/4294967296.0,1,-nbitq), 
to_sfixed(-1445720.0/4294967296.0,1,-nbitq), 
to_sfixed(194640081.0/4294967296.0,1,-nbitq), 
to_sfixed(-217518699.0/4294967296.0,1,-nbitq), 
to_sfixed(-570156218.0/4294967296.0,1,-nbitq), 
to_sfixed(-2014006906.0/4294967296.0,1,-nbitq), 
to_sfixed(166945292.0/4294967296.0,1,-nbitq), 
to_sfixed(16748403.0/4294967296.0,1,-nbitq), 
to_sfixed(-384963569.0/4294967296.0,1,-nbitq), 
to_sfixed(-410213558.0/4294967296.0,1,-nbitq), 
to_sfixed(-321587931.0/4294967296.0,1,-nbitq), 
to_sfixed(-485475828.0/4294967296.0,1,-nbitq), 
to_sfixed(-800010521.0/4294967296.0,1,-nbitq), 
to_sfixed(97310579.0/4294967296.0,1,-nbitq), 
to_sfixed(185754834.0/4294967296.0,1,-nbitq), 
to_sfixed(-34930016.0/4294967296.0,1,-nbitq), 
to_sfixed(-287434242.0/4294967296.0,1,-nbitq), 
to_sfixed(717993845.0/4294967296.0,1,-nbitq), 
to_sfixed(86591030.0/4294967296.0,1,-nbitq), 
to_sfixed(-228294282.0/4294967296.0,1,-nbitq), 
to_sfixed(182053750.0/4294967296.0,1,-nbitq), 
to_sfixed(209679480.0/4294967296.0,1,-nbitq), 
to_sfixed(-10363645.0/4294967296.0,1,-nbitq), 
to_sfixed(563682027.0/4294967296.0,1,-nbitq), 
to_sfixed(-50267664.0/4294967296.0,1,-nbitq), 
to_sfixed(52569688.0/4294967296.0,1,-nbitq), 
to_sfixed(-465760505.0/4294967296.0,1,-nbitq), 
to_sfixed(309336153.0/4294967296.0,1,-nbitq), 
to_sfixed(-271787248.0/4294967296.0,1,-nbitq), 
to_sfixed(24067576.0/4294967296.0,1,-nbitq), 
to_sfixed(66986252.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-280015081.0/4294967296.0,1,-nbitq), 
to_sfixed(-956318844.0/4294967296.0,1,-nbitq), 
to_sfixed(1216020526.0/4294967296.0,1,-nbitq), 
to_sfixed(-51170488.0/4294967296.0,1,-nbitq), 
to_sfixed(-250731029.0/4294967296.0,1,-nbitq), 
to_sfixed(64707969.0/4294967296.0,1,-nbitq), 
to_sfixed(253069967.0/4294967296.0,1,-nbitq), 
to_sfixed(376908604.0/4294967296.0,1,-nbitq), 
to_sfixed(317809375.0/4294967296.0,1,-nbitq), 
to_sfixed(48286604.0/4294967296.0,1,-nbitq), 
to_sfixed(-252289813.0/4294967296.0,1,-nbitq), 
to_sfixed(390951222.0/4294967296.0,1,-nbitq), 
to_sfixed(92338099.0/4294967296.0,1,-nbitq), 
to_sfixed(212320466.0/4294967296.0,1,-nbitq), 
to_sfixed(-61820023.0/4294967296.0,1,-nbitq), 
to_sfixed(237253263.0/4294967296.0,1,-nbitq), 
to_sfixed(317323522.0/4294967296.0,1,-nbitq), 
to_sfixed(-159501652.0/4294967296.0,1,-nbitq), 
to_sfixed(-590923823.0/4294967296.0,1,-nbitq), 
to_sfixed(108427320.0/4294967296.0,1,-nbitq), 
to_sfixed(-255758124.0/4294967296.0,1,-nbitq), 
to_sfixed(743873808.0/4294967296.0,1,-nbitq), 
to_sfixed(-545984501.0/4294967296.0,1,-nbitq), 
to_sfixed(-22438636.0/4294967296.0,1,-nbitq), 
to_sfixed(-118974501.0/4294967296.0,1,-nbitq), 
to_sfixed(-841539230.0/4294967296.0,1,-nbitq), 
to_sfixed(269757337.0/4294967296.0,1,-nbitq), 
to_sfixed(64492733.0/4294967296.0,1,-nbitq), 
to_sfixed(202954969.0/4294967296.0,1,-nbitq), 
to_sfixed(283790018.0/4294967296.0,1,-nbitq), 
to_sfixed(894802011.0/4294967296.0,1,-nbitq), 
to_sfixed(233832308.0/4294967296.0,1,-nbitq), 
to_sfixed(-126110656.0/4294967296.0,1,-nbitq), 
to_sfixed(-206199354.0/4294967296.0,1,-nbitq), 
to_sfixed(-196017572.0/4294967296.0,1,-nbitq), 
to_sfixed(473393376.0/4294967296.0,1,-nbitq), 
to_sfixed(-292440543.0/4294967296.0,1,-nbitq), 
to_sfixed(422016812.0/4294967296.0,1,-nbitq), 
to_sfixed(-135904245.0/4294967296.0,1,-nbitq), 
to_sfixed(-88468111.0/4294967296.0,1,-nbitq), 
to_sfixed(231767414.0/4294967296.0,1,-nbitq), 
to_sfixed(-75392944.0/4294967296.0,1,-nbitq), 
to_sfixed(-320257558.0/4294967296.0,1,-nbitq), 
to_sfixed(-408951347.0/4294967296.0,1,-nbitq), 
to_sfixed(264944609.0/4294967296.0,1,-nbitq), 
to_sfixed(596904344.0/4294967296.0,1,-nbitq), 
to_sfixed(-405515234.0/4294967296.0,1,-nbitq), 
to_sfixed(-110105868.0/4294967296.0,1,-nbitq), 
to_sfixed(157306693.0/4294967296.0,1,-nbitq), 
to_sfixed(-1185867818.0/4294967296.0,1,-nbitq), 
to_sfixed(402251944.0/4294967296.0,1,-nbitq), 
to_sfixed(703109071.0/4294967296.0,1,-nbitq), 
to_sfixed(160342552.0/4294967296.0,1,-nbitq), 
to_sfixed(-270696993.0/4294967296.0,1,-nbitq), 
to_sfixed(-1229255378.0/4294967296.0,1,-nbitq), 
to_sfixed(534750749.0/4294967296.0,1,-nbitq), 
to_sfixed(416721468.0/4294967296.0,1,-nbitq), 
to_sfixed(445325794.0/4294967296.0,1,-nbitq), 
to_sfixed(240687647.0/4294967296.0,1,-nbitq), 
to_sfixed(275507257.0/4294967296.0,1,-nbitq), 
to_sfixed(101345391.0/4294967296.0,1,-nbitq), 
to_sfixed(-26324668.0/4294967296.0,1,-nbitq), 
to_sfixed(-141564784.0/4294967296.0,1,-nbitq), 
to_sfixed(28467908.0/4294967296.0,1,-nbitq), 
to_sfixed(448981207.0/4294967296.0,1,-nbitq), 
to_sfixed(234715525.0/4294967296.0,1,-nbitq), 
to_sfixed(277872201.0/4294967296.0,1,-nbitq), 
to_sfixed(-46539503.0/4294967296.0,1,-nbitq), 
to_sfixed(-173721421.0/4294967296.0,1,-nbitq), 
to_sfixed(366853702.0/4294967296.0,1,-nbitq), 
to_sfixed(-58068948.0/4294967296.0,1,-nbitq), 
to_sfixed(206917627.0/4294967296.0,1,-nbitq), 
to_sfixed(-8285640.0/4294967296.0,1,-nbitq), 
to_sfixed(256796774.0/4294967296.0,1,-nbitq), 
to_sfixed(168390833.0/4294967296.0,1,-nbitq), 
to_sfixed(-210917442.0/4294967296.0,1,-nbitq), 
to_sfixed(355708800.0/4294967296.0,1,-nbitq), 
to_sfixed(552301818.0/4294967296.0,1,-nbitq), 
to_sfixed(42926090.0/4294967296.0,1,-nbitq), 
to_sfixed(276376080.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(240061753.0/4294967296.0,1,-nbitq), 
to_sfixed(-1057177634.0/4294967296.0,1,-nbitq), 
to_sfixed(1011239136.0/4294967296.0,1,-nbitq), 
to_sfixed(77897320.0/4294967296.0,1,-nbitq), 
to_sfixed(-475270520.0/4294967296.0,1,-nbitq), 
to_sfixed(180780275.0/4294967296.0,1,-nbitq), 
to_sfixed(-373441193.0/4294967296.0,1,-nbitq), 
to_sfixed(699734531.0/4294967296.0,1,-nbitq), 
to_sfixed(-40986636.0/4294967296.0,1,-nbitq), 
to_sfixed(-299245846.0/4294967296.0,1,-nbitq), 
to_sfixed(-200713794.0/4294967296.0,1,-nbitq), 
to_sfixed(615246751.0/4294967296.0,1,-nbitq), 
to_sfixed(2678030.0/4294967296.0,1,-nbitq), 
to_sfixed(331708973.0/4294967296.0,1,-nbitq), 
to_sfixed(-241929492.0/4294967296.0,1,-nbitq), 
to_sfixed(519137555.0/4294967296.0,1,-nbitq), 
to_sfixed(-338800366.0/4294967296.0,1,-nbitq), 
to_sfixed(82965283.0/4294967296.0,1,-nbitq), 
to_sfixed(-304058822.0/4294967296.0,1,-nbitq), 
to_sfixed(198749754.0/4294967296.0,1,-nbitq), 
to_sfixed(-123605403.0/4294967296.0,1,-nbitq), 
to_sfixed(460215339.0/4294967296.0,1,-nbitq), 
to_sfixed(-5710633.0/4294967296.0,1,-nbitq), 
to_sfixed(-414197289.0/4294967296.0,1,-nbitq), 
to_sfixed(355830789.0/4294967296.0,1,-nbitq), 
to_sfixed(-325686428.0/4294967296.0,1,-nbitq), 
to_sfixed(404157930.0/4294967296.0,1,-nbitq), 
to_sfixed(-59830693.0/4294967296.0,1,-nbitq), 
to_sfixed(-330664800.0/4294967296.0,1,-nbitq), 
to_sfixed(560097721.0/4294967296.0,1,-nbitq), 
to_sfixed(128925352.0/4294967296.0,1,-nbitq), 
to_sfixed(-311809209.0/4294967296.0,1,-nbitq), 
to_sfixed(-236109532.0/4294967296.0,1,-nbitq), 
to_sfixed(320057416.0/4294967296.0,1,-nbitq), 
to_sfixed(-411706262.0/4294967296.0,1,-nbitq), 
to_sfixed(155003828.0/4294967296.0,1,-nbitq), 
to_sfixed(359287366.0/4294967296.0,1,-nbitq), 
to_sfixed(150884494.0/4294967296.0,1,-nbitq), 
to_sfixed(-84284147.0/4294967296.0,1,-nbitq), 
to_sfixed(-150261467.0/4294967296.0,1,-nbitq), 
to_sfixed(-301602122.0/4294967296.0,1,-nbitq), 
to_sfixed(167963769.0/4294967296.0,1,-nbitq), 
to_sfixed(-137251417.0/4294967296.0,1,-nbitq), 
to_sfixed(-387134106.0/4294967296.0,1,-nbitq), 
to_sfixed(-7139473.0/4294967296.0,1,-nbitq), 
to_sfixed(222198702.0/4294967296.0,1,-nbitq), 
to_sfixed(159764526.0/4294967296.0,1,-nbitq), 
to_sfixed(-285889360.0/4294967296.0,1,-nbitq), 
to_sfixed(-151121036.0/4294967296.0,1,-nbitq), 
to_sfixed(-176496752.0/4294967296.0,1,-nbitq), 
to_sfixed(391078760.0/4294967296.0,1,-nbitq), 
to_sfixed(-75164853.0/4294967296.0,1,-nbitq), 
to_sfixed(794564897.0/4294967296.0,1,-nbitq), 
to_sfixed(-180413572.0/4294967296.0,1,-nbitq), 
to_sfixed(-409688681.0/4294967296.0,1,-nbitq), 
to_sfixed(347423625.0/4294967296.0,1,-nbitq), 
to_sfixed(-50200742.0/4294967296.0,1,-nbitq), 
to_sfixed(164663753.0/4294967296.0,1,-nbitq), 
to_sfixed(-203274500.0/4294967296.0,1,-nbitq), 
to_sfixed(-131850558.0/4294967296.0,1,-nbitq), 
to_sfixed(243423737.0/4294967296.0,1,-nbitq), 
to_sfixed(-363574975.0/4294967296.0,1,-nbitq), 
to_sfixed(-95334335.0/4294967296.0,1,-nbitq), 
to_sfixed(35897550.0/4294967296.0,1,-nbitq), 
to_sfixed(-180933746.0/4294967296.0,1,-nbitq), 
to_sfixed(-91712567.0/4294967296.0,1,-nbitq), 
to_sfixed(278675802.0/4294967296.0,1,-nbitq), 
to_sfixed(-268495408.0/4294967296.0,1,-nbitq), 
to_sfixed(116769377.0/4294967296.0,1,-nbitq), 
to_sfixed(636094072.0/4294967296.0,1,-nbitq), 
to_sfixed(-154985152.0/4294967296.0,1,-nbitq), 
to_sfixed(2387841.0/4294967296.0,1,-nbitq), 
to_sfixed(-148159711.0/4294967296.0,1,-nbitq), 
to_sfixed(211923524.0/4294967296.0,1,-nbitq), 
to_sfixed(-239929078.0/4294967296.0,1,-nbitq), 
to_sfixed(-311397651.0/4294967296.0,1,-nbitq), 
to_sfixed(330977104.0/4294967296.0,1,-nbitq), 
to_sfixed(405022689.0/4294967296.0,1,-nbitq), 
to_sfixed(420129731.0/4294967296.0,1,-nbitq), 
to_sfixed(226073664.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(75523484.0/4294967296.0,1,-nbitq), 
to_sfixed(43766501.0/4294967296.0,1,-nbitq), 
to_sfixed(771773619.0/4294967296.0,1,-nbitq), 
to_sfixed(43797293.0/4294967296.0,1,-nbitq), 
to_sfixed(-50811258.0/4294967296.0,1,-nbitq), 
to_sfixed(-239511543.0/4294967296.0,1,-nbitq), 
to_sfixed(-162576993.0/4294967296.0,1,-nbitq), 
to_sfixed(560540476.0/4294967296.0,1,-nbitq), 
to_sfixed(-277608308.0/4294967296.0,1,-nbitq), 
to_sfixed(157792675.0/4294967296.0,1,-nbitq), 
to_sfixed(-1730571.0/4294967296.0,1,-nbitq), 
to_sfixed(152911842.0/4294967296.0,1,-nbitq), 
to_sfixed(-35739595.0/4294967296.0,1,-nbitq), 
to_sfixed(285920976.0/4294967296.0,1,-nbitq), 
to_sfixed(-130521364.0/4294967296.0,1,-nbitq), 
to_sfixed(527506751.0/4294967296.0,1,-nbitq), 
to_sfixed(196849342.0/4294967296.0,1,-nbitq), 
to_sfixed(242124888.0/4294967296.0,1,-nbitq), 
to_sfixed(90809701.0/4294967296.0,1,-nbitq), 
to_sfixed(363527203.0/4294967296.0,1,-nbitq), 
to_sfixed(278037310.0/4294967296.0,1,-nbitq), 
to_sfixed(457891044.0/4294967296.0,1,-nbitq), 
to_sfixed(-305537082.0/4294967296.0,1,-nbitq), 
to_sfixed(91660975.0/4294967296.0,1,-nbitq), 
to_sfixed(437210268.0/4294967296.0,1,-nbitq), 
to_sfixed(-416649389.0/4294967296.0,1,-nbitq), 
to_sfixed(243745957.0/4294967296.0,1,-nbitq), 
to_sfixed(-146964490.0/4294967296.0,1,-nbitq), 
to_sfixed(538988565.0/4294967296.0,1,-nbitq), 
to_sfixed(586359382.0/4294967296.0,1,-nbitq), 
to_sfixed(-213005448.0/4294967296.0,1,-nbitq), 
to_sfixed(-180331683.0/4294967296.0,1,-nbitq), 
to_sfixed(-136013726.0/4294967296.0,1,-nbitq), 
to_sfixed(-457944364.0/4294967296.0,1,-nbitq), 
to_sfixed(-78284863.0/4294967296.0,1,-nbitq), 
to_sfixed(-362082087.0/4294967296.0,1,-nbitq), 
to_sfixed(-185969874.0/4294967296.0,1,-nbitq), 
to_sfixed(-101917409.0/4294967296.0,1,-nbitq), 
to_sfixed(144942365.0/4294967296.0,1,-nbitq), 
to_sfixed(466500101.0/4294967296.0,1,-nbitq), 
to_sfixed(205467229.0/4294967296.0,1,-nbitq), 
to_sfixed(-903701.0/4294967296.0,1,-nbitq), 
to_sfixed(-288055299.0/4294967296.0,1,-nbitq), 
to_sfixed(-85750624.0/4294967296.0,1,-nbitq), 
to_sfixed(199138788.0/4294967296.0,1,-nbitq), 
to_sfixed(-304087575.0/4294967296.0,1,-nbitq), 
to_sfixed(176379501.0/4294967296.0,1,-nbitq), 
to_sfixed(-95361480.0/4294967296.0,1,-nbitq), 
to_sfixed(-182956506.0/4294967296.0,1,-nbitq), 
to_sfixed(-588816106.0/4294967296.0,1,-nbitq), 
to_sfixed(396754661.0/4294967296.0,1,-nbitq), 
to_sfixed(374458724.0/4294967296.0,1,-nbitq), 
to_sfixed(-196990117.0/4294967296.0,1,-nbitq), 
to_sfixed(447703549.0/4294967296.0,1,-nbitq), 
to_sfixed(-356579779.0/4294967296.0,1,-nbitq), 
to_sfixed(-307009412.0/4294967296.0,1,-nbitq), 
to_sfixed(-198389667.0/4294967296.0,1,-nbitq), 
to_sfixed(396019892.0/4294967296.0,1,-nbitq), 
to_sfixed(-29463974.0/4294967296.0,1,-nbitq), 
to_sfixed(-4599097.0/4294967296.0,1,-nbitq), 
to_sfixed(159840627.0/4294967296.0,1,-nbitq), 
to_sfixed(-279320290.0/4294967296.0,1,-nbitq), 
to_sfixed(-229655158.0/4294967296.0,1,-nbitq), 
to_sfixed(-442986928.0/4294967296.0,1,-nbitq), 
to_sfixed(-186881604.0/4294967296.0,1,-nbitq), 
to_sfixed(-331210937.0/4294967296.0,1,-nbitq), 
to_sfixed(366487210.0/4294967296.0,1,-nbitq), 
to_sfixed(208442949.0/4294967296.0,1,-nbitq), 
to_sfixed(98582802.0/4294967296.0,1,-nbitq), 
to_sfixed(558114251.0/4294967296.0,1,-nbitq), 
to_sfixed(-371569118.0/4294967296.0,1,-nbitq), 
to_sfixed(70366638.0/4294967296.0,1,-nbitq), 
to_sfixed(131173754.0/4294967296.0,1,-nbitq), 
to_sfixed(-271444213.0/4294967296.0,1,-nbitq), 
to_sfixed(136970326.0/4294967296.0,1,-nbitq), 
to_sfixed(-423664848.0/4294967296.0,1,-nbitq), 
to_sfixed(-388007205.0/4294967296.0,1,-nbitq), 
to_sfixed(-65166367.0/4294967296.0,1,-nbitq), 
to_sfixed(-16483574.0/4294967296.0,1,-nbitq), 
to_sfixed(338604651.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-379884289.0/4294967296.0,1,-nbitq), 
to_sfixed(22876699.0/4294967296.0,1,-nbitq), 
to_sfixed(705472579.0/4294967296.0,1,-nbitq), 
to_sfixed(-197857753.0/4294967296.0,1,-nbitq), 
to_sfixed(-160625140.0/4294967296.0,1,-nbitq), 
to_sfixed(-642651304.0/4294967296.0,1,-nbitq), 
to_sfixed(182006667.0/4294967296.0,1,-nbitq), 
to_sfixed(-250047428.0/4294967296.0,1,-nbitq), 
to_sfixed(-530603836.0/4294967296.0,1,-nbitq), 
to_sfixed(-60112616.0/4294967296.0,1,-nbitq), 
to_sfixed(244778231.0/4294967296.0,1,-nbitq), 
to_sfixed(451979759.0/4294967296.0,1,-nbitq), 
to_sfixed(-305022222.0/4294967296.0,1,-nbitq), 
to_sfixed(349402526.0/4294967296.0,1,-nbitq), 
to_sfixed(314784449.0/4294967296.0,1,-nbitq), 
to_sfixed(-103732998.0/4294967296.0,1,-nbitq), 
to_sfixed(-279168083.0/4294967296.0,1,-nbitq), 
to_sfixed(133397182.0/4294967296.0,1,-nbitq), 
to_sfixed(33582872.0/4294967296.0,1,-nbitq), 
to_sfixed(-314410976.0/4294967296.0,1,-nbitq), 
to_sfixed(363843696.0/4294967296.0,1,-nbitq), 
to_sfixed(-96784032.0/4294967296.0,1,-nbitq), 
to_sfixed(140119296.0/4294967296.0,1,-nbitq), 
to_sfixed(576971893.0/4294967296.0,1,-nbitq), 
to_sfixed(338216973.0/4294967296.0,1,-nbitq), 
to_sfixed(-14393758.0/4294967296.0,1,-nbitq), 
to_sfixed(-114012078.0/4294967296.0,1,-nbitq), 
to_sfixed(173851560.0/4294967296.0,1,-nbitq), 
to_sfixed(308886356.0/4294967296.0,1,-nbitq), 
to_sfixed(495917117.0/4294967296.0,1,-nbitq), 
to_sfixed(-450664815.0/4294967296.0,1,-nbitq), 
to_sfixed(-344777588.0/4294967296.0,1,-nbitq), 
to_sfixed(-205297714.0/4294967296.0,1,-nbitq), 
to_sfixed(215773223.0/4294967296.0,1,-nbitq), 
to_sfixed(-399682978.0/4294967296.0,1,-nbitq), 
to_sfixed(205275960.0/4294967296.0,1,-nbitq), 
to_sfixed(-477915199.0/4294967296.0,1,-nbitq), 
to_sfixed(67644888.0/4294967296.0,1,-nbitq), 
to_sfixed(358668208.0/4294967296.0,1,-nbitq), 
to_sfixed(-3378061.0/4294967296.0,1,-nbitq), 
to_sfixed(-65647506.0/4294967296.0,1,-nbitq), 
to_sfixed(371402773.0/4294967296.0,1,-nbitq), 
to_sfixed(-140392567.0/4294967296.0,1,-nbitq), 
to_sfixed(-203105283.0/4294967296.0,1,-nbitq), 
to_sfixed(171118683.0/4294967296.0,1,-nbitq), 
to_sfixed(-50195639.0/4294967296.0,1,-nbitq), 
to_sfixed(266868178.0/4294967296.0,1,-nbitq), 
to_sfixed(-315496718.0/4294967296.0,1,-nbitq), 
to_sfixed(-20637765.0/4294967296.0,1,-nbitq), 
to_sfixed(290626487.0/4294967296.0,1,-nbitq), 
to_sfixed(-162384974.0/4294967296.0,1,-nbitq), 
to_sfixed(-64579.0/4294967296.0,1,-nbitq), 
to_sfixed(-437084292.0/4294967296.0,1,-nbitq), 
to_sfixed(188408208.0/4294967296.0,1,-nbitq), 
to_sfixed(69878467.0/4294967296.0,1,-nbitq), 
to_sfixed(260542839.0/4294967296.0,1,-nbitq), 
to_sfixed(266438102.0/4294967296.0,1,-nbitq), 
to_sfixed(358327335.0/4294967296.0,1,-nbitq), 
to_sfixed(-62197457.0/4294967296.0,1,-nbitq), 
to_sfixed(170471762.0/4294967296.0,1,-nbitq), 
to_sfixed(-123905982.0/4294967296.0,1,-nbitq), 
to_sfixed(-114321310.0/4294967296.0,1,-nbitq), 
to_sfixed(402118931.0/4294967296.0,1,-nbitq), 
to_sfixed(164032148.0/4294967296.0,1,-nbitq), 
to_sfixed(263206254.0/4294967296.0,1,-nbitq), 
to_sfixed(226690120.0/4294967296.0,1,-nbitq), 
to_sfixed(301887274.0/4294967296.0,1,-nbitq), 
to_sfixed(-408966897.0/4294967296.0,1,-nbitq), 
to_sfixed(-75421818.0/4294967296.0,1,-nbitq), 
to_sfixed(532889338.0/4294967296.0,1,-nbitq), 
to_sfixed(-435865204.0/4294967296.0,1,-nbitq), 
to_sfixed(-305493398.0/4294967296.0,1,-nbitq), 
to_sfixed(184153262.0/4294967296.0,1,-nbitq), 
to_sfixed(180778127.0/4294967296.0,1,-nbitq), 
to_sfixed(288475218.0/4294967296.0,1,-nbitq), 
to_sfixed(25173678.0/4294967296.0,1,-nbitq), 
to_sfixed(-79729648.0/4294967296.0,1,-nbitq), 
to_sfixed(-159124152.0/4294967296.0,1,-nbitq), 
to_sfixed(-268871511.0/4294967296.0,1,-nbitq), 
to_sfixed(-257275324.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-283116665.0/4294967296.0,1,-nbitq), 
to_sfixed(-430229397.0/4294967296.0,1,-nbitq), 
to_sfixed(421132214.0/4294967296.0,1,-nbitq), 
to_sfixed(81243568.0/4294967296.0,1,-nbitq), 
to_sfixed(267282317.0/4294967296.0,1,-nbitq), 
to_sfixed(-57111647.0/4294967296.0,1,-nbitq), 
to_sfixed(-91928689.0/4294967296.0,1,-nbitq), 
to_sfixed(-77660017.0/4294967296.0,1,-nbitq), 
to_sfixed(-460413969.0/4294967296.0,1,-nbitq), 
to_sfixed(303645898.0/4294967296.0,1,-nbitq), 
to_sfixed(246101135.0/4294967296.0,1,-nbitq), 
to_sfixed(407959730.0/4294967296.0,1,-nbitq), 
to_sfixed(208251227.0/4294967296.0,1,-nbitq), 
to_sfixed(36564690.0/4294967296.0,1,-nbitq), 
to_sfixed(-339244010.0/4294967296.0,1,-nbitq), 
to_sfixed(306869995.0/4294967296.0,1,-nbitq), 
to_sfixed(-72435228.0/4294967296.0,1,-nbitq), 
to_sfixed(390145174.0/4294967296.0,1,-nbitq), 
to_sfixed(-219131132.0/4294967296.0,1,-nbitq), 
to_sfixed(-146109107.0/4294967296.0,1,-nbitq), 
to_sfixed(-296236429.0/4294967296.0,1,-nbitq), 
to_sfixed(-60548620.0/4294967296.0,1,-nbitq), 
to_sfixed(-43583428.0/4294967296.0,1,-nbitq), 
to_sfixed(479873210.0/4294967296.0,1,-nbitq), 
to_sfixed(-265084243.0/4294967296.0,1,-nbitq), 
to_sfixed(-401135232.0/4294967296.0,1,-nbitq), 
to_sfixed(99036339.0/4294967296.0,1,-nbitq), 
to_sfixed(-125173073.0/4294967296.0,1,-nbitq), 
to_sfixed(-51091511.0/4294967296.0,1,-nbitq), 
to_sfixed(329621227.0/4294967296.0,1,-nbitq), 
to_sfixed(-634031569.0/4294967296.0,1,-nbitq), 
to_sfixed(-156706939.0/4294967296.0,1,-nbitq), 
to_sfixed(268257476.0/4294967296.0,1,-nbitq), 
to_sfixed(62138708.0/4294967296.0,1,-nbitq), 
to_sfixed(-49007761.0/4294967296.0,1,-nbitq), 
to_sfixed(-506343717.0/4294967296.0,1,-nbitq), 
to_sfixed(-77761155.0/4294967296.0,1,-nbitq), 
to_sfixed(282534230.0/4294967296.0,1,-nbitq), 
to_sfixed(-264227223.0/4294967296.0,1,-nbitq), 
to_sfixed(5862112.0/4294967296.0,1,-nbitq), 
to_sfixed(-265862451.0/4294967296.0,1,-nbitq), 
to_sfixed(-203641984.0/4294967296.0,1,-nbitq), 
to_sfixed(-25103843.0/4294967296.0,1,-nbitq), 
to_sfixed(269637102.0/4294967296.0,1,-nbitq), 
to_sfixed(-137026888.0/4294967296.0,1,-nbitq), 
to_sfixed(-213125287.0/4294967296.0,1,-nbitq), 
to_sfixed(-301495993.0/4294967296.0,1,-nbitq), 
to_sfixed(-514156386.0/4294967296.0,1,-nbitq), 
to_sfixed(-15160011.0/4294967296.0,1,-nbitq), 
to_sfixed(33176647.0/4294967296.0,1,-nbitq), 
to_sfixed(-134647976.0/4294967296.0,1,-nbitq), 
to_sfixed(-213406197.0/4294967296.0,1,-nbitq), 
to_sfixed(146760113.0/4294967296.0,1,-nbitq), 
to_sfixed(197585430.0/4294967296.0,1,-nbitq), 
to_sfixed(441508011.0/4294967296.0,1,-nbitq), 
to_sfixed(-360853462.0/4294967296.0,1,-nbitq), 
to_sfixed(471444952.0/4294967296.0,1,-nbitq), 
to_sfixed(-340162431.0/4294967296.0,1,-nbitq), 
to_sfixed(236025337.0/4294967296.0,1,-nbitq), 
to_sfixed(395560604.0/4294967296.0,1,-nbitq), 
to_sfixed(109090148.0/4294967296.0,1,-nbitq), 
to_sfixed(67827863.0/4294967296.0,1,-nbitq), 
to_sfixed(317770436.0/4294967296.0,1,-nbitq), 
to_sfixed(-60866791.0/4294967296.0,1,-nbitq), 
to_sfixed(-376172555.0/4294967296.0,1,-nbitq), 
to_sfixed(-338327508.0/4294967296.0,1,-nbitq), 
to_sfixed(654146983.0/4294967296.0,1,-nbitq), 
to_sfixed(78048424.0/4294967296.0,1,-nbitq), 
to_sfixed(141053493.0/4294967296.0,1,-nbitq), 
to_sfixed(136669618.0/4294967296.0,1,-nbitq), 
to_sfixed(164467866.0/4294967296.0,1,-nbitq), 
to_sfixed(9853356.0/4294967296.0,1,-nbitq), 
to_sfixed(-205427711.0/4294967296.0,1,-nbitq), 
to_sfixed(-224685604.0/4294967296.0,1,-nbitq), 
to_sfixed(180197708.0/4294967296.0,1,-nbitq), 
to_sfixed(55456512.0/4294967296.0,1,-nbitq), 
to_sfixed(195038886.0/4294967296.0,1,-nbitq), 
to_sfixed(21106201.0/4294967296.0,1,-nbitq), 
to_sfixed(258622462.0/4294967296.0,1,-nbitq), 
to_sfixed(144873873.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-2951743.0/4294967296.0,1,-nbitq), 
to_sfixed(-343259540.0/4294967296.0,1,-nbitq), 
to_sfixed(445983058.0/4294967296.0,1,-nbitq), 
to_sfixed(-299487842.0/4294967296.0,1,-nbitq), 
to_sfixed(-54796873.0/4294967296.0,1,-nbitq), 
to_sfixed(174579686.0/4294967296.0,1,-nbitq), 
to_sfixed(-49501777.0/4294967296.0,1,-nbitq), 
to_sfixed(-262449579.0/4294967296.0,1,-nbitq), 
to_sfixed(82672443.0/4294967296.0,1,-nbitq), 
to_sfixed(147912528.0/4294967296.0,1,-nbitq), 
to_sfixed(339631827.0/4294967296.0,1,-nbitq), 
to_sfixed(310289450.0/4294967296.0,1,-nbitq), 
to_sfixed(-213158180.0/4294967296.0,1,-nbitq), 
to_sfixed(289834235.0/4294967296.0,1,-nbitq), 
to_sfixed(-85206764.0/4294967296.0,1,-nbitq), 
to_sfixed(-405551548.0/4294967296.0,1,-nbitq), 
to_sfixed(-355795250.0/4294967296.0,1,-nbitq), 
to_sfixed(311589231.0/4294967296.0,1,-nbitq), 
to_sfixed(-103471360.0/4294967296.0,1,-nbitq), 
to_sfixed(302134045.0/4294967296.0,1,-nbitq), 
to_sfixed(-110672090.0/4294967296.0,1,-nbitq), 
to_sfixed(446994078.0/4294967296.0,1,-nbitq), 
to_sfixed(-77470707.0/4294967296.0,1,-nbitq), 
to_sfixed(-361865153.0/4294967296.0,1,-nbitq), 
to_sfixed(-141998055.0/4294967296.0,1,-nbitq), 
to_sfixed(525446293.0/4294967296.0,1,-nbitq), 
to_sfixed(193212455.0/4294967296.0,1,-nbitq), 
to_sfixed(-386951879.0/4294967296.0,1,-nbitq), 
to_sfixed(-60614622.0/4294967296.0,1,-nbitq), 
to_sfixed(-23297356.0/4294967296.0,1,-nbitq), 
to_sfixed(37801179.0/4294967296.0,1,-nbitq), 
to_sfixed(-166113929.0/4294967296.0,1,-nbitq), 
to_sfixed(105373242.0/4294967296.0,1,-nbitq), 
to_sfixed(53433213.0/4294967296.0,1,-nbitq), 
to_sfixed(285272384.0/4294967296.0,1,-nbitq), 
to_sfixed(-188024039.0/4294967296.0,1,-nbitq), 
to_sfixed(-42302681.0/4294967296.0,1,-nbitq), 
to_sfixed(169728449.0/4294967296.0,1,-nbitq), 
to_sfixed(51950160.0/4294967296.0,1,-nbitq), 
to_sfixed(-66636891.0/4294967296.0,1,-nbitq), 
to_sfixed(-25183511.0/4294967296.0,1,-nbitq), 
to_sfixed(409509441.0/4294967296.0,1,-nbitq), 
to_sfixed(-192874782.0/4294967296.0,1,-nbitq), 
to_sfixed(-5732666.0/4294967296.0,1,-nbitq), 
to_sfixed(322317792.0/4294967296.0,1,-nbitq), 
to_sfixed(196706126.0/4294967296.0,1,-nbitq), 
to_sfixed(-61325780.0/4294967296.0,1,-nbitq), 
to_sfixed(-85704717.0/4294967296.0,1,-nbitq), 
to_sfixed(55774641.0/4294967296.0,1,-nbitq), 
to_sfixed(530240419.0/4294967296.0,1,-nbitq), 
to_sfixed(373092540.0/4294967296.0,1,-nbitq), 
to_sfixed(-304146620.0/4294967296.0,1,-nbitq), 
to_sfixed(-113656595.0/4294967296.0,1,-nbitq), 
to_sfixed(92454241.0/4294967296.0,1,-nbitq), 
to_sfixed(-60498914.0/4294967296.0,1,-nbitq), 
to_sfixed(37881419.0/4294967296.0,1,-nbitq), 
to_sfixed(8998735.0/4294967296.0,1,-nbitq), 
to_sfixed(157583567.0/4294967296.0,1,-nbitq), 
to_sfixed(-173815722.0/4294967296.0,1,-nbitq), 
to_sfixed(76187633.0/4294967296.0,1,-nbitq), 
to_sfixed(-109174550.0/4294967296.0,1,-nbitq), 
to_sfixed(-267962181.0/4294967296.0,1,-nbitq), 
to_sfixed(115906615.0/4294967296.0,1,-nbitq), 
to_sfixed(-66623961.0/4294967296.0,1,-nbitq), 
to_sfixed(-186625934.0/4294967296.0,1,-nbitq), 
to_sfixed(-256304046.0/4294967296.0,1,-nbitq), 
to_sfixed(619429474.0/4294967296.0,1,-nbitq), 
to_sfixed(342197586.0/4294967296.0,1,-nbitq), 
to_sfixed(-228396039.0/4294967296.0,1,-nbitq), 
to_sfixed(63317720.0/4294967296.0,1,-nbitq), 
to_sfixed(51688851.0/4294967296.0,1,-nbitq), 
to_sfixed(-156038051.0/4294967296.0,1,-nbitq), 
to_sfixed(154785237.0/4294967296.0,1,-nbitq), 
to_sfixed(246035493.0/4294967296.0,1,-nbitq), 
to_sfixed(263590118.0/4294967296.0,1,-nbitq), 
to_sfixed(-104562810.0/4294967296.0,1,-nbitq), 
to_sfixed(-41267888.0/4294967296.0,1,-nbitq), 
to_sfixed(134030834.0/4294967296.0,1,-nbitq), 
to_sfixed(81697503.0/4294967296.0,1,-nbitq), 
to_sfixed(-265615301.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-288932648.0/4294967296.0,1,-nbitq), 
to_sfixed(-334420016.0/4294967296.0,1,-nbitq), 
to_sfixed(-19006245.0/4294967296.0,1,-nbitq), 
to_sfixed(-114930278.0/4294967296.0,1,-nbitq), 
to_sfixed(176508736.0/4294967296.0,1,-nbitq), 
to_sfixed(-217012537.0/4294967296.0,1,-nbitq), 
to_sfixed(-343862937.0/4294967296.0,1,-nbitq), 
to_sfixed(-251612118.0/4294967296.0,1,-nbitq), 
to_sfixed(-156609373.0/4294967296.0,1,-nbitq), 
to_sfixed(191999443.0/4294967296.0,1,-nbitq), 
to_sfixed(12287011.0/4294967296.0,1,-nbitq), 
to_sfixed(-242659809.0/4294967296.0,1,-nbitq), 
to_sfixed(-309274562.0/4294967296.0,1,-nbitq), 
to_sfixed(-91538194.0/4294967296.0,1,-nbitq), 
to_sfixed(19490427.0/4294967296.0,1,-nbitq), 
to_sfixed(274192401.0/4294967296.0,1,-nbitq), 
to_sfixed(58793972.0/4294967296.0,1,-nbitq), 
to_sfixed(52394293.0/4294967296.0,1,-nbitq), 
to_sfixed(284011946.0/4294967296.0,1,-nbitq), 
to_sfixed(91877431.0/4294967296.0,1,-nbitq), 
to_sfixed(47911168.0/4294967296.0,1,-nbitq), 
to_sfixed(141878700.0/4294967296.0,1,-nbitq), 
to_sfixed(334363533.0/4294967296.0,1,-nbitq), 
to_sfixed(69319910.0/4294967296.0,1,-nbitq), 
to_sfixed(345045707.0/4294967296.0,1,-nbitq), 
to_sfixed(96247690.0/4294967296.0,1,-nbitq), 
to_sfixed(-45350060.0/4294967296.0,1,-nbitq), 
to_sfixed(84347049.0/4294967296.0,1,-nbitq), 
to_sfixed(-58159554.0/4294967296.0,1,-nbitq), 
to_sfixed(-108514349.0/4294967296.0,1,-nbitq), 
to_sfixed(-557826688.0/4294967296.0,1,-nbitq), 
to_sfixed(-138118214.0/4294967296.0,1,-nbitq), 
to_sfixed(416173208.0/4294967296.0,1,-nbitq), 
to_sfixed(141223854.0/4294967296.0,1,-nbitq), 
to_sfixed(268783839.0/4294967296.0,1,-nbitq), 
to_sfixed(-236432069.0/4294967296.0,1,-nbitq), 
to_sfixed(353815225.0/4294967296.0,1,-nbitq), 
to_sfixed(480129317.0/4294967296.0,1,-nbitq), 
to_sfixed(75862999.0/4294967296.0,1,-nbitq), 
to_sfixed(-257269618.0/4294967296.0,1,-nbitq), 
to_sfixed(23280553.0/4294967296.0,1,-nbitq), 
to_sfixed(104249280.0/4294967296.0,1,-nbitq), 
to_sfixed(163475458.0/4294967296.0,1,-nbitq), 
to_sfixed(141689413.0/4294967296.0,1,-nbitq), 
to_sfixed(-155509028.0/4294967296.0,1,-nbitq), 
to_sfixed(97009719.0/4294967296.0,1,-nbitq), 
to_sfixed(129476272.0/4294967296.0,1,-nbitq), 
to_sfixed(-217995526.0/4294967296.0,1,-nbitq), 
to_sfixed(278504177.0/4294967296.0,1,-nbitq), 
to_sfixed(-43571873.0/4294967296.0,1,-nbitq), 
to_sfixed(81482168.0/4294967296.0,1,-nbitq), 
to_sfixed(68424843.0/4294967296.0,1,-nbitq), 
to_sfixed(-30496944.0/4294967296.0,1,-nbitq), 
to_sfixed(167001485.0/4294967296.0,1,-nbitq), 
to_sfixed(379093663.0/4294967296.0,1,-nbitq), 
to_sfixed(147442045.0/4294967296.0,1,-nbitq), 
to_sfixed(294194471.0/4294967296.0,1,-nbitq), 
to_sfixed(-225075944.0/4294967296.0,1,-nbitq), 
to_sfixed(57418194.0/4294967296.0,1,-nbitq), 
to_sfixed(215190698.0/4294967296.0,1,-nbitq), 
to_sfixed(-359645896.0/4294967296.0,1,-nbitq), 
to_sfixed(49315484.0/4294967296.0,1,-nbitq), 
to_sfixed(-88895890.0/4294967296.0,1,-nbitq), 
to_sfixed(159091425.0/4294967296.0,1,-nbitq), 
to_sfixed(-35878347.0/4294967296.0,1,-nbitq), 
to_sfixed(-389589798.0/4294967296.0,1,-nbitq), 
to_sfixed(624065148.0/4294967296.0,1,-nbitq), 
to_sfixed(-23589193.0/4294967296.0,1,-nbitq), 
to_sfixed(407139223.0/4294967296.0,1,-nbitq), 
to_sfixed(-47869499.0/4294967296.0,1,-nbitq), 
to_sfixed(274373092.0/4294967296.0,1,-nbitq), 
to_sfixed(387622910.0/4294967296.0,1,-nbitq), 
to_sfixed(-163011812.0/4294967296.0,1,-nbitq), 
to_sfixed(308134471.0/4294967296.0,1,-nbitq), 
to_sfixed(346576186.0/4294967296.0,1,-nbitq), 
to_sfixed(-396524265.0/4294967296.0,1,-nbitq), 
to_sfixed(-429105389.0/4294967296.0,1,-nbitq), 
to_sfixed(234578729.0/4294967296.0,1,-nbitq), 
to_sfixed(-551175562.0/4294967296.0,1,-nbitq), 
to_sfixed(224573577.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-61401043.0/4294967296.0,1,-nbitq), 
to_sfixed(-512722727.0/4294967296.0,1,-nbitq), 
to_sfixed(189567008.0/4294967296.0,1,-nbitq), 
to_sfixed(-244436387.0/4294967296.0,1,-nbitq), 
to_sfixed(406824772.0/4294967296.0,1,-nbitq), 
to_sfixed(-144104737.0/4294967296.0,1,-nbitq), 
to_sfixed(-170227996.0/4294967296.0,1,-nbitq), 
to_sfixed(392637059.0/4294967296.0,1,-nbitq), 
to_sfixed(-54471531.0/4294967296.0,1,-nbitq), 
to_sfixed(176055424.0/4294967296.0,1,-nbitq), 
to_sfixed(71019177.0/4294967296.0,1,-nbitq), 
to_sfixed(-224656893.0/4294967296.0,1,-nbitq), 
to_sfixed(-223546094.0/4294967296.0,1,-nbitq), 
to_sfixed(-264680304.0/4294967296.0,1,-nbitq), 
to_sfixed(231967946.0/4294967296.0,1,-nbitq), 
to_sfixed(-207721298.0/4294967296.0,1,-nbitq), 
to_sfixed(-344337191.0/4294967296.0,1,-nbitq), 
to_sfixed(337295310.0/4294967296.0,1,-nbitq), 
to_sfixed(98529500.0/4294967296.0,1,-nbitq), 
to_sfixed(253326665.0/4294967296.0,1,-nbitq), 
to_sfixed(-40076196.0/4294967296.0,1,-nbitq), 
to_sfixed(44844094.0/4294967296.0,1,-nbitq), 
to_sfixed(-370472360.0/4294967296.0,1,-nbitq), 
to_sfixed(222887729.0/4294967296.0,1,-nbitq), 
to_sfixed(154478478.0/4294967296.0,1,-nbitq), 
to_sfixed(314784497.0/4294967296.0,1,-nbitq), 
to_sfixed(284846122.0/4294967296.0,1,-nbitq), 
to_sfixed(-26302826.0/4294967296.0,1,-nbitq), 
to_sfixed(-52576901.0/4294967296.0,1,-nbitq), 
to_sfixed(223430027.0/4294967296.0,1,-nbitq), 
to_sfixed(-223858323.0/4294967296.0,1,-nbitq), 
to_sfixed(-245208620.0/4294967296.0,1,-nbitq), 
to_sfixed(358742142.0/4294967296.0,1,-nbitq), 
to_sfixed(4045563.0/4294967296.0,1,-nbitq), 
to_sfixed(-124693983.0/4294967296.0,1,-nbitq), 
to_sfixed(399598491.0/4294967296.0,1,-nbitq), 
to_sfixed(48770459.0/4294967296.0,1,-nbitq), 
to_sfixed(557104311.0/4294967296.0,1,-nbitq), 
to_sfixed(-266023865.0/4294967296.0,1,-nbitq), 
to_sfixed(-222643404.0/4294967296.0,1,-nbitq), 
to_sfixed(-425804238.0/4294967296.0,1,-nbitq), 
to_sfixed(174927951.0/4294967296.0,1,-nbitq), 
to_sfixed(130791708.0/4294967296.0,1,-nbitq), 
to_sfixed(-32085595.0/4294967296.0,1,-nbitq), 
to_sfixed(-142291509.0/4294967296.0,1,-nbitq), 
to_sfixed(431579428.0/4294967296.0,1,-nbitq), 
to_sfixed(-402864372.0/4294967296.0,1,-nbitq), 
to_sfixed(-27838692.0/4294967296.0,1,-nbitq), 
to_sfixed(-96858615.0/4294967296.0,1,-nbitq), 
to_sfixed(391595379.0/4294967296.0,1,-nbitq), 
to_sfixed(-308833567.0/4294967296.0,1,-nbitq), 
to_sfixed(572118500.0/4294967296.0,1,-nbitq), 
to_sfixed(-391476173.0/4294967296.0,1,-nbitq), 
to_sfixed(309734321.0/4294967296.0,1,-nbitq), 
to_sfixed(-72076599.0/4294967296.0,1,-nbitq), 
to_sfixed(-390965801.0/4294967296.0,1,-nbitq), 
to_sfixed(124413846.0/4294967296.0,1,-nbitq), 
to_sfixed(-495611897.0/4294967296.0,1,-nbitq), 
to_sfixed(130578856.0/4294967296.0,1,-nbitq), 
to_sfixed(364699500.0/4294967296.0,1,-nbitq), 
to_sfixed(-63620999.0/4294967296.0,1,-nbitq), 
to_sfixed(622055081.0/4294967296.0,1,-nbitq), 
to_sfixed(163686548.0/4294967296.0,1,-nbitq), 
to_sfixed(-168280180.0/4294967296.0,1,-nbitq), 
to_sfixed(89959117.0/4294967296.0,1,-nbitq), 
to_sfixed(-77048774.0/4294967296.0,1,-nbitq), 
to_sfixed(654042873.0/4294967296.0,1,-nbitq), 
to_sfixed(-122797202.0/4294967296.0,1,-nbitq), 
to_sfixed(-63546869.0/4294967296.0,1,-nbitq), 
to_sfixed(483712277.0/4294967296.0,1,-nbitq), 
to_sfixed(-428070508.0/4294967296.0,1,-nbitq), 
to_sfixed(-222619439.0/4294967296.0,1,-nbitq), 
to_sfixed(-256776793.0/4294967296.0,1,-nbitq), 
to_sfixed(-159767160.0/4294967296.0,1,-nbitq), 
to_sfixed(207140440.0/4294967296.0,1,-nbitq), 
to_sfixed(-442654652.0/4294967296.0,1,-nbitq), 
to_sfixed(246238922.0/4294967296.0,1,-nbitq), 
to_sfixed(-142285424.0/4294967296.0,1,-nbitq), 
to_sfixed(160531702.0/4294967296.0,1,-nbitq), 
to_sfixed(365646846.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-205387502.0/4294967296.0,1,-nbitq), 
to_sfixed(-723043224.0/4294967296.0,1,-nbitq), 
to_sfixed(485140733.0/4294967296.0,1,-nbitq), 
to_sfixed(-379580829.0/4294967296.0,1,-nbitq), 
to_sfixed(-13556314.0/4294967296.0,1,-nbitq), 
to_sfixed(-142596448.0/4294967296.0,1,-nbitq), 
to_sfixed(128497803.0/4294967296.0,1,-nbitq), 
to_sfixed(56161675.0/4294967296.0,1,-nbitq), 
to_sfixed(246618664.0/4294967296.0,1,-nbitq), 
to_sfixed(-173249382.0/4294967296.0,1,-nbitq), 
to_sfixed(344648085.0/4294967296.0,1,-nbitq), 
to_sfixed(291817371.0/4294967296.0,1,-nbitq), 
to_sfixed(279594875.0/4294967296.0,1,-nbitq), 
to_sfixed(-5016773.0/4294967296.0,1,-nbitq), 
to_sfixed(159935739.0/4294967296.0,1,-nbitq), 
to_sfixed(178611381.0/4294967296.0,1,-nbitq), 
to_sfixed(-98257578.0/4294967296.0,1,-nbitq), 
to_sfixed(291819046.0/4294967296.0,1,-nbitq), 
to_sfixed(-364680270.0/4294967296.0,1,-nbitq), 
to_sfixed(145045063.0/4294967296.0,1,-nbitq), 
to_sfixed(288446916.0/4294967296.0,1,-nbitq), 
to_sfixed(-329240994.0/4294967296.0,1,-nbitq), 
to_sfixed(-510008724.0/4294967296.0,1,-nbitq), 
to_sfixed(467143039.0/4294967296.0,1,-nbitq), 
to_sfixed(112232500.0/4294967296.0,1,-nbitq), 
to_sfixed(-491566601.0/4294967296.0,1,-nbitq), 
to_sfixed(-158283456.0/4294967296.0,1,-nbitq), 
to_sfixed(-373571117.0/4294967296.0,1,-nbitq), 
to_sfixed(-444984327.0/4294967296.0,1,-nbitq), 
to_sfixed(92128940.0/4294967296.0,1,-nbitq), 
to_sfixed(149835186.0/4294967296.0,1,-nbitq), 
to_sfixed(-813144445.0/4294967296.0,1,-nbitq), 
to_sfixed(-60043764.0/4294967296.0,1,-nbitq), 
to_sfixed(238887671.0/4294967296.0,1,-nbitq), 
to_sfixed(-275215770.0/4294967296.0,1,-nbitq), 
to_sfixed(455318049.0/4294967296.0,1,-nbitq), 
to_sfixed(545985048.0/4294967296.0,1,-nbitq), 
to_sfixed(335289735.0/4294967296.0,1,-nbitq), 
to_sfixed(-136422290.0/4294967296.0,1,-nbitq), 
to_sfixed(436626008.0/4294967296.0,1,-nbitq), 
to_sfixed(-549772146.0/4294967296.0,1,-nbitq), 
to_sfixed(34965242.0/4294967296.0,1,-nbitq), 
to_sfixed(101729073.0/4294967296.0,1,-nbitq), 
to_sfixed(-261732240.0/4294967296.0,1,-nbitq), 
to_sfixed(-426313119.0/4294967296.0,1,-nbitq), 
to_sfixed(188952378.0/4294967296.0,1,-nbitq), 
to_sfixed(224423607.0/4294967296.0,1,-nbitq), 
to_sfixed(-429369121.0/4294967296.0,1,-nbitq), 
to_sfixed(51703087.0/4294967296.0,1,-nbitq), 
to_sfixed(-59564676.0/4294967296.0,1,-nbitq), 
to_sfixed(406781960.0/4294967296.0,1,-nbitq), 
to_sfixed(137094354.0/4294967296.0,1,-nbitq), 
to_sfixed(-51882106.0/4294967296.0,1,-nbitq), 
to_sfixed(372303624.0/4294967296.0,1,-nbitq), 
to_sfixed(1194374.0/4294967296.0,1,-nbitq), 
to_sfixed(87354549.0/4294967296.0,1,-nbitq), 
to_sfixed(251571798.0/4294967296.0,1,-nbitq), 
to_sfixed(196009671.0/4294967296.0,1,-nbitq), 
to_sfixed(-304956487.0/4294967296.0,1,-nbitq), 
to_sfixed(239323036.0/4294967296.0,1,-nbitq), 
to_sfixed(-284191903.0/4294967296.0,1,-nbitq), 
to_sfixed(32910060.0/4294967296.0,1,-nbitq), 
to_sfixed(363843073.0/4294967296.0,1,-nbitq), 
to_sfixed(-64553501.0/4294967296.0,1,-nbitq), 
to_sfixed(-235237005.0/4294967296.0,1,-nbitq), 
to_sfixed(-441788662.0/4294967296.0,1,-nbitq), 
to_sfixed(-102062250.0/4294967296.0,1,-nbitq), 
to_sfixed(369655083.0/4294967296.0,1,-nbitq), 
to_sfixed(386573824.0/4294967296.0,1,-nbitq), 
to_sfixed(158399685.0/4294967296.0,1,-nbitq), 
to_sfixed(260033271.0/4294967296.0,1,-nbitq), 
to_sfixed(-230848954.0/4294967296.0,1,-nbitq), 
to_sfixed(29304496.0/4294967296.0,1,-nbitq), 
to_sfixed(396648814.0/4294967296.0,1,-nbitq), 
to_sfixed(391689368.0/4294967296.0,1,-nbitq), 
to_sfixed(-224946420.0/4294967296.0,1,-nbitq), 
to_sfixed(-92932575.0/4294967296.0,1,-nbitq), 
to_sfixed(134637114.0/4294967296.0,1,-nbitq), 
to_sfixed(-307287555.0/4294967296.0,1,-nbitq), 
to_sfixed(381564619.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-278753277.0/4294967296.0,1,-nbitq), 
to_sfixed(-774485182.0/4294967296.0,1,-nbitq), 
to_sfixed(294457744.0/4294967296.0,1,-nbitq), 
to_sfixed(299820240.0/4294967296.0,1,-nbitq), 
to_sfixed(57975596.0/4294967296.0,1,-nbitq), 
to_sfixed(499063585.0/4294967296.0,1,-nbitq), 
to_sfixed(-83832804.0/4294967296.0,1,-nbitq), 
to_sfixed(19602884.0/4294967296.0,1,-nbitq), 
to_sfixed(-118017231.0/4294967296.0,1,-nbitq), 
to_sfixed(-331031382.0/4294967296.0,1,-nbitq), 
to_sfixed(361748440.0/4294967296.0,1,-nbitq), 
to_sfixed(-199008098.0/4294967296.0,1,-nbitq), 
to_sfixed(-156695592.0/4294967296.0,1,-nbitq), 
to_sfixed(-853056451.0/4294967296.0,1,-nbitq), 
to_sfixed(137496400.0/4294967296.0,1,-nbitq), 
to_sfixed(182579546.0/4294967296.0,1,-nbitq), 
to_sfixed(384093014.0/4294967296.0,1,-nbitq), 
to_sfixed(-83855443.0/4294967296.0,1,-nbitq), 
to_sfixed(-670143790.0/4294967296.0,1,-nbitq), 
to_sfixed(173378878.0/4294967296.0,1,-nbitq), 
to_sfixed(239477516.0/4294967296.0,1,-nbitq), 
to_sfixed(-501897799.0/4294967296.0,1,-nbitq), 
to_sfixed(-1030524686.0/4294967296.0,1,-nbitq), 
to_sfixed(308534512.0/4294967296.0,1,-nbitq), 
to_sfixed(-326989666.0/4294967296.0,1,-nbitq), 
to_sfixed(-500415626.0/4294967296.0,1,-nbitq), 
to_sfixed(640281981.0/4294967296.0,1,-nbitq), 
to_sfixed(435723710.0/4294967296.0,1,-nbitq), 
to_sfixed(-432172670.0/4294967296.0,1,-nbitq), 
to_sfixed(-219666284.0/4294967296.0,1,-nbitq), 
to_sfixed(-281883409.0/4294967296.0,1,-nbitq), 
to_sfixed(-187613711.0/4294967296.0,1,-nbitq), 
to_sfixed(-36478376.0/4294967296.0,1,-nbitq), 
to_sfixed(687035730.0/4294967296.0,1,-nbitq), 
to_sfixed(-344705296.0/4294967296.0,1,-nbitq), 
to_sfixed(-220998616.0/4294967296.0,1,-nbitq), 
to_sfixed(424318199.0/4294967296.0,1,-nbitq), 
to_sfixed(253746531.0/4294967296.0,1,-nbitq), 
to_sfixed(-50750737.0/4294967296.0,1,-nbitq), 
to_sfixed(-256886188.0/4294967296.0,1,-nbitq), 
to_sfixed(128417760.0/4294967296.0,1,-nbitq), 
to_sfixed(-501788161.0/4294967296.0,1,-nbitq), 
to_sfixed(-95718190.0/4294967296.0,1,-nbitq), 
to_sfixed(-576858474.0/4294967296.0,1,-nbitq), 
to_sfixed(-648605081.0/4294967296.0,1,-nbitq), 
to_sfixed(370700547.0/4294967296.0,1,-nbitq), 
to_sfixed(-87507792.0/4294967296.0,1,-nbitq), 
to_sfixed(-369880793.0/4294967296.0,1,-nbitq), 
to_sfixed(215570866.0/4294967296.0,1,-nbitq), 
to_sfixed(-205963345.0/4294967296.0,1,-nbitq), 
to_sfixed(425450756.0/4294967296.0,1,-nbitq), 
to_sfixed(391607336.0/4294967296.0,1,-nbitq), 
to_sfixed(272196965.0/4294967296.0,1,-nbitq), 
to_sfixed(-234327840.0/4294967296.0,1,-nbitq), 
to_sfixed(444814510.0/4294967296.0,1,-nbitq), 
to_sfixed(-336689807.0/4294967296.0,1,-nbitq), 
to_sfixed(28346373.0/4294967296.0,1,-nbitq), 
to_sfixed(155831273.0/4294967296.0,1,-nbitq), 
to_sfixed(87500120.0/4294967296.0,1,-nbitq), 
to_sfixed(-301869625.0/4294967296.0,1,-nbitq), 
to_sfixed(-5823319.0/4294967296.0,1,-nbitq), 
to_sfixed(290873713.0/4294967296.0,1,-nbitq), 
to_sfixed(449083510.0/4294967296.0,1,-nbitq), 
to_sfixed(321635370.0/4294967296.0,1,-nbitq), 
to_sfixed(-367052712.0/4294967296.0,1,-nbitq), 
to_sfixed(-208980420.0/4294967296.0,1,-nbitq), 
to_sfixed(-1004828610.0/4294967296.0,1,-nbitq), 
to_sfixed(-31462246.0/4294967296.0,1,-nbitq), 
to_sfixed(371356656.0/4294967296.0,1,-nbitq), 
to_sfixed(752086872.0/4294967296.0,1,-nbitq), 
to_sfixed(-152825048.0/4294967296.0,1,-nbitq), 
to_sfixed(-85814573.0/4294967296.0,1,-nbitq), 
to_sfixed(357252231.0/4294967296.0,1,-nbitq), 
to_sfixed(35330252.0/4294967296.0,1,-nbitq), 
to_sfixed(71862212.0/4294967296.0,1,-nbitq), 
to_sfixed(-124932079.0/4294967296.0,1,-nbitq), 
to_sfixed(-298047188.0/4294967296.0,1,-nbitq), 
to_sfixed(93061152.0/4294967296.0,1,-nbitq), 
to_sfixed(-393419452.0/4294967296.0,1,-nbitq), 
to_sfixed(-28278501.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-248195936.0/4294967296.0,1,-nbitq), 
to_sfixed(105727885.0/4294967296.0,1,-nbitq), 
to_sfixed(459771473.0/4294967296.0,1,-nbitq), 
to_sfixed(809123669.0/4294967296.0,1,-nbitq), 
to_sfixed(-133388038.0/4294967296.0,1,-nbitq), 
to_sfixed(947360404.0/4294967296.0,1,-nbitq), 
to_sfixed(178814141.0/4294967296.0,1,-nbitq), 
to_sfixed(284726069.0/4294967296.0,1,-nbitq), 
to_sfixed(223221609.0/4294967296.0,1,-nbitq), 
to_sfixed(19105495.0/4294967296.0,1,-nbitq), 
to_sfixed(1103944807.0/4294967296.0,1,-nbitq), 
to_sfixed(-512896710.0/4294967296.0,1,-nbitq), 
to_sfixed(-1021906088.0/4294967296.0,1,-nbitq), 
to_sfixed(-755652293.0/4294967296.0,1,-nbitq), 
to_sfixed(139869938.0/4294967296.0,1,-nbitq), 
to_sfixed(647124833.0/4294967296.0,1,-nbitq), 
to_sfixed(158736985.0/4294967296.0,1,-nbitq), 
to_sfixed(-104274310.0/4294967296.0,1,-nbitq), 
to_sfixed(-1700658485.0/4294967296.0,1,-nbitq), 
to_sfixed(1100921281.0/4294967296.0,1,-nbitq), 
to_sfixed(-335723608.0/4294967296.0,1,-nbitq), 
to_sfixed(-147196119.0/4294967296.0,1,-nbitq), 
to_sfixed(-535148196.0/4294967296.0,1,-nbitq), 
to_sfixed(727677968.0/4294967296.0,1,-nbitq), 
to_sfixed(144767600.0/4294967296.0,1,-nbitq), 
to_sfixed(-767310851.0/4294967296.0,1,-nbitq), 
to_sfixed(287761861.0/4294967296.0,1,-nbitq), 
to_sfixed(624522823.0/4294967296.0,1,-nbitq), 
to_sfixed(-44715217.0/4294967296.0,1,-nbitq), 
to_sfixed(-373439867.0/4294967296.0,1,-nbitq), 
to_sfixed(193086651.0/4294967296.0,1,-nbitq), 
to_sfixed(-1511813.0/4294967296.0,1,-nbitq), 
to_sfixed(644249538.0/4294967296.0,1,-nbitq), 
to_sfixed(428117211.0/4294967296.0,1,-nbitq), 
to_sfixed(297871262.0/4294967296.0,1,-nbitq), 
to_sfixed(-708183702.0/4294967296.0,1,-nbitq), 
to_sfixed(-104370194.0/4294967296.0,1,-nbitq), 
to_sfixed(-440165733.0/4294967296.0,1,-nbitq), 
to_sfixed(-147812194.0/4294967296.0,1,-nbitq), 
to_sfixed(-8008221.0/4294967296.0,1,-nbitq), 
to_sfixed(-509975173.0/4294967296.0,1,-nbitq), 
to_sfixed(-841667098.0/4294967296.0,1,-nbitq), 
to_sfixed(-194707577.0/4294967296.0,1,-nbitq), 
to_sfixed(-210997960.0/4294967296.0,1,-nbitq), 
to_sfixed(-274744002.0/4294967296.0,1,-nbitq), 
to_sfixed(-376860110.0/4294967296.0,1,-nbitq), 
to_sfixed(-141132614.0/4294967296.0,1,-nbitq), 
to_sfixed(-267494336.0/4294967296.0,1,-nbitq), 
to_sfixed(-178366814.0/4294967296.0,1,-nbitq), 
to_sfixed(-825865545.0/4294967296.0,1,-nbitq), 
to_sfixed(-115621899.0/4294967296.0,1,-nbitq), 
to_sfixed(441946959.0/4294967296.0,1,-nbitq), 
to_sfixed(696468451.0/4294967296.0,1,-nbitq), 
to_sfixed(-530725207.0/4294967296.0,1,-nbitq), 
to_sfixed(-224830918.0/4294967296.0,1,-nbitq), 
to_sfixed(615301507.0/4294967296.0,1,-nbitq), 
to_sfixed(262601101.0/4294967296.0,1,-nbitq), 
to_sfixed(-71209234.0/4294967296.0,1,-nbitq), 
to_sfixed(-84673789.0/4294967296.0,1,-nbitq), 
to_sfixed(-251359305.0/4294967296.0,1,-nbitq), 
to_sfixed(290922958.0/4294967296.0,1,-nbitq), 
to_sfixed(-191235287.0/4294967296.0,1,-nbitq), 
to_sfixed(446366049.0/4294967296.0,1,-nbitq), 
to_sfixed(-477994283.0/4294967296.0,1,-nbitq), 
to_sfixed(-516551424.0/4294967296.0,1,-nbitq), 
to_sfixed(69448239.0/4294967296.0,1,-nbitq), 
to_sfixed(-1359762030.0/4294967296.0,1,-nbitq), 
to_sfixed(-643374984.0/4294967296.0,1,-nbitq), 
to_sfixed(170067621.0/4294967296.0,1,-nbitq), 
to_sfixed(427650748.0/4294967296.0,1,-nbitq), 
to_sfixed(-361782644.0/4294967296.0,1,-nbitq), 
to_sfixed(-311935967.0/4294967296.0,1,-nbitq), 
to_sfixed(641774632.0/4294967296.0,1,-nbitq), 
to_sfixed(-342486325.0/4294967296.0,1,-nbitq), 
to_sfixed(-74154351.0/4294967296.0,1,-nbitq), 
to_sfixed(537600287.0/4294967296.0,1,-nbitq), 
to_sfixed(-981530599.0/4294967296.0,1,-nbitq), 
to_sfixed(67396543.0/4294967296.0,1,-nbitq), 
to_sfixed(-797759195.0/4294967296.0,1,-nbitq), 
to_sfixed(-172782989.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-367105503.0/4294967296.0,1,-nbitq), 
to_sfixed(-189708613.0/4294967296.0,1,-nbitq), 
to_sfixed(872870643.0/4294967296.0,1,-nbitq), 
to_sfixed(1113725647.0/4294967296.0,1,-nbitq), 
to_sfixed(-263818805.0/4294967296.0,1,-nbitq), 
to_sfixed(1110001694.0/4294967296.0,1,-nbitq), 
to_sfixed(-147826934.0/4294967296.0,1,-nbitq), 
to_sfixed(236158035.0/4294967296.0,1,-nbitq), 
to_sfixed(444774437.0/4294967296.0,1,-nbitq), 
to_sfixed(-214657311.0/4294967296.0,1,-nbitq), 
to_sfixed(252158399.0/4294967296.0,1,-nbitq), 
to_sfixed(-362718564.0/4294967296.0,1,-nbitq), 
to_sfixed(-1594217086.0/4294967296.0,1,-nbitq), 
to_sfixed(-677570299.0/4294967296.0,1,-nbitq), 
to_sfixed(-124357048.0/4294967296.0,1,-nbitq), 
to_sfixed(168165080.0/4294967296.0,1,-nbitq), 
to_sfixed(137842255.0/4294967296.0,1,-nbitq), 
to_sfixed(-106922508.0/4294967296.0,1,-nbitq), 
to_sfixed(-1798251812.0/4294967296.0,1,-nbitq), 
to_sfixed(225011916.0/4294967296.0,1,-nbitq), 
to_sfixed(-278614366.0/4294967296.0,1,-nbitq), 
to_sfixed(-471539877.0/4294967296.0,1,-nbitq), 
to_sfixed(-122904398.0/4294967296.0,1,-nbitq), 
to_sfixed(81987122.0/4294967296.0,1,-nbitq), 
to_sfixed(-17236447.0/4294967296.0,1,-nbitq), 
to_sfixed(-1016037025.0/4294967296.0,1,-nbitq), 
to_sfixed(155022409.0/4294967296.0,1,-nbitq), 
to_sfixed(703071330.0/4294967296.0,1,-nbitq), 
to_sfixed(374792816.0/4294967296.0,1,-nbitq), 
to_sfixed(-864848061.0/4294967296.0,1,-nbitq), 
to_sfixed(544867948.0/4294967296.0,1,-nbitq), 
to_sfixed(-167220637.0/4294967296.0,1,-nbitq), 
to_sfixed(543223972.0/4294967296.0,1,-nbitq), 
to_sfixed(675293375.0/4294967296.0,1,-nbitq), 
to_sfixed(-333732189.0/4294967296.0,1,-nbitq), 
to_sfixed(-1260290452.0/4294967296.0,1,-nbitq), 
to_sfixed(-229376264.0/4294967296.0,1,-nbitq), 
to_sfixed(325505409.0/4294967296.0,1,-nbitq), 
to_sfixed(510458153.0/4294967296.0,1,-nbitq), 
to_sfixed(239573891.0/4294967296.0,1,-nbitq), 
to_sfixed(74892578.0/4294967296.0,1,-nbitq), 
to_sfixed(-1002805890.0/4294967296.0,1,-nbitq), 
to_sfixed(542681667.0/4294967296.0,1,-nbitq), 
to_sfixed(-356020302.0/4294967296.0,1,-nbitq), 
to_sfixed(500641914.0/4294967296.0,1,-nbitq), 
to_sfixed(-824597963.0/4294967296.0,1,-nbitq), 
to_sfixed(-70166767.0/4294967296.0,1,-nbitq), 
to_sfixed(102586974.0/4294967296.0,1,-nbitq), 
to_sfixed(48689505.0/4294967296.0,1,-nbitq), 
to_sfixed(-220497564.0/4294967296.0,1,-nbitq), 
to_sfixed(-401008751.0/4294967296.0,1,-nbitq), 
to_sfixed(336090602.0/4294967296.0,1,-nbitq), 
to_sfixed(1033523697.0/4294967296.0,1,-nbitq), 
to_sfixed(-811238184.0/4294967296.0,1,-nbitq), 
to_sfixed(-1131046140.0/4294967296.0,1,-nbitq), 
to_sfixed(659894287.0/4294967296.0,1,-nbitq), 
to_sfixed(-131239643.0/4294967296.0,1,-nbitq), 
to_sfixed(12794397.0/4294967296.0,1,-nbitq), 
to_sfixed(-130518581.0/4294967296.0,1,-nbitq), 
to_sfixed(-237115731.0/4294967296.0,1,-nbitq), 
to_sfixed(393044636.0/4294967296.0,1,-nbitq), 
to_sfixed(176904362.0/4294967296.0,1,-nbitq), 
to_sfixed(322107851.0/4294967296.0,1,-nbitq), 
to_sfixed(-340584953.0/4294967296.0,1,-nbitq), 
to_sfixed(16132588.0/4294967296.0,1,-nbitq), 
to_sfixed(-275748269.0/4294967296.0,1,-nbitq), 
to_sfixed(-1406160309.0/4294967296.0,1,-nbitq), 
to_sfixed(-751818548.0/4294967296.0,1,-nbitq), 
to_sfixed(-123368490.0/4294967296.0,1,-nbitq), 
to_sfixed(335355772.0/4294967296.0,1,-nbitq), 
to_sfixed(-506696095.0/4294967296.0,1,-nbitq), 
to_sfixed(473017819.0/4294967296.0,1,-nbitq), 
to_sfixed(84936415.0/4294967296.0,1,-nbitq), 
to_sfixed(-96115786.0/4294967296.0,1,-nbitq), 
to_sfixed(-27324023.0/4294967296.0,1,-nbitq), 
to_sfixed(467810657.0/4294967296.0,1,-nbitq), 
to_sfixed(-1042878000.0/4294967296.0,1,-nbitq), 
to_sfixed(-120883245.0/4294967296.0,1,-nbitq), 
to_sfixed(-990421901.0/4294967296.0,1,-nbitq), 
to_sfixed(-96043781.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-306961180.0/4294967296.0,1,-nbitq), 
to_sfixed(95904709.0/4294967296.0,1,-nbitq), 
to_sfixed(771831665.0/4294967296.0,1,-nbitq), 
to_sfixed(1625124986.0/4294967296.0,1,-nbitq), 
to_sfixed(1010770447.0/4294967296.0,1,-nbitq), 
to_sfixed(1337617721.0/4294967296.0,1,-nbitq), 
to_sfixed(240635078.0/4294967296.0,1,-nbitq), 
to_sfixed(696169770.0/4294967296.0,1,-nbitq), 
to_sfixed(473651148.0/4294967296.0,1,-nbitq), 
to_sfixed(381732332.0/4294967296.0,1,-nbitq), 
to_sfixed(-223355151.0/4294967296.0,1,-nbitq), 
to_sfixed(-27736467.0/4294967296.0,1,-nbitq), 
to_sfixed(-1203946591.0/4294967296.0,1,-nbitq), 
to_sfixed(-822028681.0/4294967296.0,1,-nbitq), 
to_sfixed(-272515066.0/4294967296.0,1,-nbitq), 
to_sfixed(521736909.0/4294967296.0,1,-nbitq), 
to_sfixed(-394984266.0/4294967296.0,1,-nbitq), 
to_sfixed(247124495.0/4294967296.0,1,-nbitq), 
to_sfixed(-1370863279.0/4294967296.0,1,-nbitq), 
to_sfixed(486694009.0/4294967296.0,1,-nbitq), 
to_sfixed(-277542163.0/4294967296.0,1,-nbitq), 
to_sfixed(533745038.0/4294967296.0,1,-nbitq), 
to_sfixed(526939408.0/4294967296.0,1,-nbitq), 
to_sfixed(-28028427.0/4294967296.0,1,-nbitq), 
to_sfixed(-326417328.0/4294967296.0,1,-nbitq), 
to_sfixed(-1122269109.0/4294967296.0,1,-nbitq), 
to_sfixed(167372073.0/4294967296.0,1,-nbitq), 
to_sfixed(-27808192.0/4294967296.0,1,-nbitq), 
to_sfixed(686536273.0/4294967296.0,1,-nbitq), 
to_sfixed(82610837.0/4294967296.0,1,-nbitq), 
to_sfixed(787597736.0/4294967296.0,1,-nbitq), 
to_sfixed(-649099030.0/4294967296.0,1,-nbitq), 
to_sfixed(831529305.0/4294967296.0,1,-nbitq), 
to_sfixed(1144108932.0/4294967296.0,1,-nbitq), 
to_sfixed(-379665654.0/4294967296.0,1,-nbitq), 
to_sfixed(-1125538423.0/4294967296.0,1,-nbitq), 
to_sfixed(158275697.0/4294967296.0,1,-nbitq), 
to_sfixed(56509598.0/4294967296.0,1,-nbitq), 
to_sfixed(312948703.0/4294967296.0,1,-nbitq), 
to_sfixed(-98807079.0/4294967296.0,1,-nbitq), 
to_sfixed(242073407.0/4294967296.0,1,-nbitq), 
to_sfixed(-1091293825.0/4294967296.0,1,-nbitq), 
to_sfixed(-410702468.0/4294967296.0,1,-nbitq), 
to_sfixed(-706229083.0/4294967296.0,1,-nbitq), 
to_sfixed(339612380.0/4294967296.0,1,-nbitq), 
to_sfixed(-1729535726.0/4294967296.0,1,-nbitq), 
to_sfixed(-368053489.0/4294967296.0,1,-nbitq), 
to_sfixed(515905900.0/4294967296.0,1,-nbitq), 
to_sfixed(325657575.0/4294967296.0,1,-nbitq), 
to_sfixed(-298879026.0/4294967296.0,1,-nbitq), 
to_sfixed(-190965561.0/4294967296.0,1,-nbitq), 
to_sfixed(114211226.0/4294967296.0,1,-nbitq), 
to_sfixed(329321410.0/4294967296.0,1,-nbitq), 
to_sfixed(-296583003.0/4294967296.0,1,-nbitq), 
to_sfixed(406229877.0/4294967296.0,1,-nbitq), 
to_sfixed(582209311.0/4294967296.0,1,-nbitq), 
to_sfixed(-644778156.0/4294967296.0,1,-nbitq), 
to_sfixed(702914876.0/4294967296.0,1,-nbitq), 
to_sfixed(-339594986.0/4294967296.0,1,-nbitq), 
to_sfixed(89812748.0/4294967296.0,1,-nbitq), 
to_sfixed(229435355.0/4294967296.0,1,-nbitq), 
to_sfixed(488529691.0/4294967296.0,1,-nbitq), 
to_sfixed(117430628.0/4294967296.0,1,-nbitq), 
to_sfixed(215997168.0/4294967296.0,1,-nbitq), 
to_sfixed(-508314495.0/4294967296.0,1,-nbitq), 
to_sfixed(68989296.0/4294967296.0,1,-nbitq), 
to_sfixed(-1390608819.0/4294967296.0,1,-nbitq), 
to_sfixed(-709632301.0/4294967296.0,1,-nbitq), 
to_sfixed(34679925.0/4294967296.0,1,-nbitq), 
to_sfixed(550556324.0/4294967296.0,1,-nbitq), 
to_sfixed(355273078.0/4294967296.0,1,-nbitq), 
to_sfixed(266817896.0/4294967296.0,1,-nbitq), 
to_sfixed(404966193.0/4294967296.0,1,-nbitq), 
to_sfixed(-54873568.0/4294967296.0,1,-nbitq), 
to_sfixed(-100049042.0/4294967296.0,1,-nbitq), 
to_sfixed(170145744.0/4294967296.0,1,-nbitq), 
to_sfixed(-152922067.0/4294967296.0,1,-nbitq), 
to_sfixed(130717861.0/4294967296.0,1,-nbitq), 
to_sfixed(-920142490.0/4294967296.0,1,-nbitq), 
to_sfixed(249807677.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-479065120.0/4294967296.0,1,-nbitq), 
to_sfixed(545323317.0/4294967296.0,1,-nbitq), 
to_sfixed(752626425.0/4294967296.0,1,-nbitq), 
to_sfixed(1851479255.0/4294967296.0,1,-nbitq), 
to_sfixed(598601670.0/4294967296.0,1,-nbitq), 
to_sfixed(1256179706.0/4294967296.0,1,-nbitq), 
to_sfixed(-561663866.0/4294967296.0,1,-nbitq), 
to_sfixed(469579782.0/4294967296.0,1,-nbitq), 
to_sfixed(590641505.0/4294967296.0,1,-nbitq), 
to_sfixed(147064698.0/4294967296.0,1,-nbitq), 
to_sfixed(-300816962.0/4294967296.0,1,-nbitq), 
to_sfixed(769927193.0/4294967296.0,1,-nbitq), 
to_sfixed(-871847393.0/4294967296.0,1,-nbitq), 
to_sfixed(-963349332.0/4294967296.0,1,-nbitq), 
to_sfixed(194053766.0/4294967296.0,1,-nbitq), 
to_sfixed(171750050.0/4294967296.0,1,-nbitq), 
to_sfixed(-463984814.0/4294967296.0,1,-nbitq), 
to_sfixed(-136682671.0/4294967296.0,1,-nbitq), 
to_sfixed(-942842376.0/4294967296.0,1,-nbitq), 
to_sfixed(218231881.0/4294967296.0,1,-nbitq), 
to_sfixed(-376916307.0/4294967296.0,1,-nbitq), 
to_sfixed(410154340.0/4294967296.0,1,-nbitq), 
to_sfixed(67787793.0/4294967296.0,1,-nbitq), 
to_sfixed(209005747.0/4294967296.0,1,-nbitq), 
to_sfixed(-360812083.0/4294967296.0,1,-nbitq), 
to_sfixed(104289432.0/4294967296.0,1,-nbitq), 
to_sfixed(268930809.0/4294967296.0,1,-nbitq), 
to_sfixed(601313981.0/4294967296.0,1,-nbitq), 
to_sfixed(-156366829.0/4294967296.0,1,-nbitq), 
to_sfixed(837293.0/4294967296.0,1,-nbitq), 
to_sfixed(514354048.0/4294967296.0,1,-nbitq), 
to_sfixed(-799518070.0/4294967296.0,1,-nbitq), 
to_sfixed(810205212.0/4294967296.0,1,-nbitq), 
to_sfixed(559242951.0/4294967296.0,1,-nbitq), 
to_sfixed(-1148235795.0/4294967296.0,1,-nbitq), 
to_sfixed(-573700987.0/4294967296.0,1,-nbitq), 
to_sfixed(-141821544.0/4294967296.0,1,-nbitq), 
to_sfixed(-807606260.0/4294967296.0,1,-nbitq), 
to_sfixed(-142931950.0/4294967296.0,1,-nbitq), 
to_sfixed(-25655070.0/4294967296.0,1,-nbitq), 
to_sfixed(-466465626.0/4294967296.0,1,-nbitq), 
to_sfixed(-904867195.0/4294967296.0,1,-nbitq), 
to_sfixed(58745431.0/4294967296.0,1,-nbitq), 
to_sfixed(181208258.0/4294967296.0,1,-nbitq), 
to_sfixed(259340162.0/4294967296.0,1,-nbitq), 
to_sfixed(-1700416084.0/4294967296.0,1,-nbitq), 
to_sfixed(60337760.0/4294967296.0,1,-nbitq), 
to_sfixed(-15605683.0/4294967296.0,1,-nbitq), 
to_sfixed(207235836.0/4294967296.0,1,-nbitq), 
to_sfixed(-494357068.0/4294967296.0,1,-nbitq), 
to_sfixed(-623728803.0/4294967296.0,1,-nbitq), 
to_sfixed(278545985.0/4294967296.0,1,-nbitq), 
to_sfixed(-1003740938.0/4294967296.0,1,-nbitq), 
to_sfixed(-382793832.0/4294967296.0,1,-nbitq), 
to_sfixed(796328183.0/4294967296.0,1,-nbitq), 
to_sfixed(-369904352.0/4294967296.0,1,-nbitq), 
to_sfixed(-481127592.0/4294967296.0,1,-nbitq), 
to_sfixed(450125438.0/4294967296.0,1,-nbitq), 
to_sfixed(-230532475.0/4294967296.0,1,-nbitq), 
to_sfixed(3053516.0/4294967296.0,1,-nbitq), 
to_sfixed(-245486569.0/4294967296.0,1,-nbitq), 
to_sfixed(447873542.0/4294967296.0,1,-nbitq), 
to_sfixed(-14344964.0/4294967296.0,1,-nbitq), 
to_sfixed(26497115.0/4294967296.0,1,-nbitq), 
to_sfixed(-709105484.0/4294967296.0,1,-nbitq), 
to_sfixed(310801447.0/4294967296.0,1,-nbitq), 
to_sfixed(-1726851375.0/4294967296.0,1,-nbitq), 
to_sfixed(-1071971402.0/4294967296.0,1,-nbitq), 
to_sfixed(204088263.0/4294967296.0,1,-nbitq), 
to_sfixed(355341810.0/4294967296.0,1,-nbitq), 
to_sfixed(42002159.0/4294967296.0,1,-nbitq), 
to_sfixed(-14243433.0/4294967296.0,1,-nbitq), 
to_sfixed(407319436.0/4294967296.0,1,-nbitq), 
to_sfixed(221819455.0/4294967296.0,1,-nbitq), 
to_sfixed(467650462.0/4294967296.0,1,-nbitq), 
to_sfixed(-632189919.0/4294967296.0,1,-nbitq), 
to_sfixed(-141000240.0/4294967296.0,1,-nbitq), 
to_sfixed(-770737186.0/4294967296.0,1,-nbitq), 
to_sfixed(92473990.0/4294967296.0,1,-nbitq), 
to_sfixed(-322818721.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-195488782.0/4294967296.0,1,-nbitq), 
to_sfixed(352224344.0/4294967296.0,1,-nbitq), 
to_sfixed(859625343.0/4294967296.0,1,-nbitq), 
to_sfixed(1579562919.0/4294967296.0,1,-nbitq), 
to_sfixed(480079044.0/4294967296.0,1,-nbitq), 
to_sfixed(-395773891.0/4294967296.0,1,-nbitq), 
to_sfixed(-174043978.0/4294967296.0,1,-nbitq), 
to_sfixed(709136315.0/4294967296.0,1,-nbitq), 
to_sfixed(869164640.0/4294967296.0,1,-nbitq), 
to_sfixed(244067604.0/4294967296.0,1,-nbitq), 
to_sfixed(-94544826.0/4294967296.0,1,-nbitq), 
to_sfixed(690700169.0/4294967296.0,1,-nbitq), 
to_sfixed(-999741029.0/4294967296.0,1,-nbitq), 
to_sfixed(-1095468698.0/4294967296.0,1,-nbitq), 
to_sfixed(137642374.0/4294967296.0,1,-nbitq), 
to_sfixed(219548655.0/4294967296.0,1,-nbitq), 
to_sfixed(-418633496.0/4294967296.0,1,-nbitq), 
to_sfixed(260567250.0/4294967296.0,1,-nbitq), 
to_sfixed(3506785.0/4294967296.0,1,-nbitq), 
to_sfixed(-346817316.0/4294967296.0,1,-nbitq), 
to_sfixed(5921368.0/4294967296.0,1,-nbitq), 
to_sfixed(134670774.0/4294967296.0,1,-nbitq), 
to_sfixed(-448537712.0/4294967296.0,1,-nbitq), 
to_sfixed(-590860732.0/4294967296.0,1,-nbitq), 
to_sfixed(-49170013.0/4294967296.0,1,-nbitq), 
to_sfixed(-380101457.0/4294967296.0,1,-nbitq), 
to_sfixed(-238058040.0/4294967296.0,1,-nbitq), 
to_sfixed(1305645818.0/4294967296.0,1,-nbitq), 
to_sfixed(717627187.0/4294967296.0,1,-nbitq), 
to_sfixed(366965862.0/4294967296.0,1,-nbitq), 
to_sfixed(217726230.0/4294967296.0,1,-nbitq), 
to_sfixed(242991507.0/4294967296.0,1,-nbitq), 
to_sfixed(773988815.0/4294967296.0,1,-nbitq), 
to_sfixed(276644223.0/4294967296.0,1,-nbitq), 
to_sfixed(-280270686.0/4294967296.0,1,-nbitq), 
to_sfixed(-1272156604.0/4294967296.0,1,-nbitq), 
to_sfixed(-504965073.0/4294967296.0,1,-nbitq), 
to_sfixed(-416861010.0/4294967296.0,1,-nbitq), 
to_sfixed(161536099.0/4294967296.0,1,-nbitq), 
to_sfixed(-421134885.0/4294967296.0,1,-nbitq), 
to_sfixed(-376519712.0/4294967296.0,1,-nbitq), 
to_sfixed(-858011876.0/4294967296.0,1,-nbitq), 
to_sfixed(274453182.0/4294967296.0,1,-nbitq), 
to_sfixed(512199897.0/4294967296.0,1,-nbitq), 
to_sfixed(-362510405.0/4294967296.0,1,-nbitq), 
to_sfixed(-1987360915.0/4294967296.0,1,-nbitq), 
to_sfixed(222478818.0/4294967296.0,1,-nbitq), 
to_sfixed(340826610.0/4294967296.0,1,-nbitq), 
to_sfixed(-109201957.0/4294967296.0,1,-nbitq), 
to_sfixed(-795708440.0/4294967296.0,1,-nbitq), 
to_sfixed(-645039271.0/4294967296.0,1,-nbitq), 
to_sfixed(-45985397.0/4294967296.0,1,-nbitq), 
to_sfixed(-1005546016.0/4294967296.0,1,-nbitq), 
to_sfixed(76700191.0/4294967296.0,1,-nbitq), 
to_sfixed(443697701.0/4294967296.0,1,-nbitq), 
to_sfixed(-370135572.0/4294967296.0,1,-nbitq), 
to_sfixed(-443961805.0/4294967296.0,1,-nbitq), 
to_sfixed(206390273.0/4294967296.0,1,-nbitq), 
to_sfixed(349271294.0/4294967296.0,1,-nbitq), 
to_sfixed(117580999.0/4294967296.0,1,-nbitq), 
to_sfixed(266604382.0/4294967296.0,1,-nbitq), 
to_sfixed(1149363660.0/4294967296.0,1,-nbitq), 
to_sfixed(1106721713.0/4294967296.0,1,-nbitq), 
to_sfixed(397002494.0/4294967296.0,1,-nbitq), 
to_sfixed(-189422988.0/4294967296.0,1,-nbitq), 
to_sfixed(-25938921.0/4294967296.0,1,-nbitq), 
to_sfixed(-1090601880.0/4294967296.0,1,-nbitq), 
to_sfixed(-744401966.0/4294967296.0,1,-nbitq), 
to_sfixed(237436390.0/4294967296.0,1,-nbitq), 
to_sfixed(770002800.0/4294967296.0,1,-nbitq), 
to_sfixed(-1174710901.0/4294967296.0,1,-nbitq), 
to_sfixed(-219980812.0/4294967296.0,1,-nbitq), 
to_sfixed(509076803.0/4294967296.0,1,-nbitq), 
to_sfixed(54944156.0/4294967296.0,1,-nbitq), 
to_sfixed(286421076.0/4294967296.0,1,-nbitq), 
to_sfixed(531525400.0/4294967296.0,1,-nbitq), 
to_sfixed(-1071064813.0/4294967296.0,1,-nbitq), 
to_sfixed(-330668669.0/4294967296.0,1,-nbitq), 
to_sfixed(465694619.0/4294967296.0,1,-nbitq), 
to_sfixed(104591256.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-503867606.0/4294967296.0,1,-nbitq), 
to_sfixed(207343405.0/4294967296.0,1,-nbitq), 
to_sfixed(1343676260.0/4294967296.0,1,-nbitq), 
to_sfixed(1434619586.0/4294967296.0,1,-nbitq), 
to_sfixed(791449061.0/4294967296.0,1,-nbitq), 
to_sfixed(-720231801.0/4294967296.0,1,-nbitq), 
to_sfixed(-144044607.0/4294967296.0,1,-nbitq), 
to_sfixed(-1327098158.0/4294967296.0,1,-nbitq), 
to_sfixed(536528665.0/4294967296.0,1,-nbitq), 
to_sfixed(-70444591.0/4294967296.0,1,-nbitq), 
to_sfixed(-390099122.0/4294967296.0,1,-nbitq), 
to_sfixed(621987481.0/4294967296.0,1,-nbitq), 
to_sfixed(-1383024629.0/4294967296.0,1,-nbitq), 
to_sfixed(-598521020.0/4294967296.0,1,-nbitq), 
to_sfixed(322279684.0/4294967296.0,1,-nbitq), 
to_sfixed(-120651416.0/4294967296.0,1,-nbitq), 
to_sfixed(-316966715.0/4294967296.0,1,-nbitq), 
to_sfixed(-57716262.0/4294967296.0,1,-nbitq), 
to_sfixed(-59509222.0/4294967296.0,1,-nbitq), 
to_sfixed(-1156043489.0/4294967296.0,1,-nbitq), 
to_sfixed(-313181139.0/4294967296.0,1,-nbitq), 
to_sfixed(-141545765.0/4294967296.0,1,-nbitq), 
to_sfixed(108676276.0/4294967296.0,1,-nbitq), 
to_sfixed(-209712539.0/4294967296.0,1,-nbitq), 
to_sfixed(149899358.0/4294967296.0,1,-nbitq), 
to_sfixed(-257089422.0/4294967296.0,1,-nbitq), 
to_sfixed(-480225141.0/4294967296.0,1,-nbitq), 
to_sfixed(767256215.0/4294967296.0,1,-nbitq), 
to_sfixed(1318359601.0/4294967296.0,1,-nbitq), 
to_sfixed(-205095609.0/4294967296.0,1,-nbitq), 
to_sfixed(700884573.0/4294967296.0,1,-nbitq), 
to_sfixed(-133908022.0/4294967296.0,1,-nbitq), 
to_sfixed(901839202.0/4294967296.0,1,-nbitq), 
to_sfixed(-300206131.0/4294967296.0,1,-nbitq), 
to_sfixed(-404627060.0/4294967296.0,1,-nbitq), 
to_sfixed(-547220403.0/4294967296.0,1,-nbitq), 
to_sfixed(-917805438.0/4294967296.0,1,-nbitq), 
to_sfixed(83971035.0/4294967296.0,1,-nbitq), 
to_sfixed(-97646220.0/4294967296.0,1,-nbitq), 
to_sfixed(-341555686.0/4294967296.0,1,-nbitq), 
to_sfixed(-419313189.0/4294967296.0,1,-nbitq), 
to_sfixed(-688194177.0/4294967296.0,1,-nbitq), 
to_sfixed(1003526130.0/4294967296.0,1,-nbitq), 
to_sfixed(807185076.0/4294967296.0,1,-nbitq), 
to_sfixed(-225214195.0/4294967296.0,1,-nbitq), 
to_sfixed(-1814128119.0/4294967296.0,1,-nbitq), 
to_sfixed(-43164795.0/4294967296.0,1,-nbitq), 
to_sfixed(858471829.0/4294967296.0,1,-nbitq), 
to_sfixed(-591186930.0/4294967296.0,1,-nbitq), 
to_sfixed(-544536303.0/4294967296.0,1,-nbitq), 
to_sfixed(-313788153.0/4294967296.0,1,-nbitq), 
to_sfixed(-396981917.0/4294967296.0,1,-nbitq), 
to_sfixed(-1081061772.0/4294967296.0,1,-nbitq), 
to_sfixed(947936157.0/4294967296.0,1,-nbitq), 
to_sfixed(387867793.0/4294967296.0,1,-nbitq), 
to_sfixed(295202335.0/4294967296.0,1,-nbitq), 
to_sfixed(-800045938.0/4294967296.0,1,-nbitq), 
to_sfixed(82594596.0/4294967296.0,1,-nbitq), 
to_sfixed(-294205229.0/4294967296.0,1,-nbitq), 
to_sfixed(50156528.0/4294967296.0,1,-nbitq), 
to_sfixed(69920279.0/4294967296.0,1,-nbitq), 
to_sfixed(1712073295.0/4294967296.0,1,-nbitq), 
to_sfixed(1625896579.0/4294967296.0,1,-nbitq), 
to_sfixed(340877232.0/4294967296.0,1,-nbitq), 
to_sfixed(-144454866.0/4294967296.0,1,-nbitq), 
to_sfixed(168745276.0/4294967296.0,1,-nbitq), 
to_sfixed(1058278360.0/4294967296.0,1,-nbitq), 
to_sfixed(-459141110.0/4294967296.0,1,-nbitq), 
to_sfixed(122049644.0/4294967296.0,1,-nbitq), 
to_sfixed(523646972.0/4294967296.0,1,-nbitq), 
to_sfixed(-1233927187.0/4294967296.0,1,-nbitq), 
to_sfixed(122106868.0/4294967296.0,1,-nbitq), 
to_sfixed(365406975.0/4294967296.0,1,-nbitq), 
to_sfixed(-272008029.0/4294967296.0,1,-nbitq), 
to_sfixed(108690369.0/4294967296.0,1,-nbitq), 
to_sfixed(-56036046.0/4294967296.0,1,-nbitq), 
to_sfixed(-202560163.0/4294967296.0,1,-nbitq), 
to_sfixed(-13651686.0/4294967296.0,1,-nbitq), 
to_sfixed(391977199.0/4294967296.0,1,-nbitq), 
to_sfixed(204156294.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-72017086.0/4294967296.0,1,-nbitq), 
to_sfixed(457176451.0/4294967296.0,1,-nbitq), 
to_sfixed(-418179142.0/4294967296.0,1,-nbitq), 
to_sfixed(601989121.0/4294967296.0,1,-nbitq), 
to_sfixed(-622240578.0/4294967296.0,1,-nbitq), 
to_sfixed(-310266064.0/4294967296.0,1,-nbitq), 
to_sfixed(-131037157.0/4294967296.0,1,-nbitq), 
to_sfixed(-969184915.0/4294967296.0,1,-nbitq), 
to_sfixed(18588690.0/4294967296.0,1,-nbitq), 
to_sfixed(-61086019.0/4294967296.0,1,-nbitq), 
to_sfixed(435668874.0/4294967296.0,1,-nbitq), 
to_sfixed(1147367006.0/4294967296.0,1,-nbitq), 
to_sfixed(-1588959519.0/4294967296.0,1,-nbitq), 
to_sfixed(-849208467.0/4294967296.0,1,-nbitq), 
to_sfixed(244420649.0/4294967296.0,1,-nbitq), 
to_sfixed(-345436568.0/4294967296.0,1,-nbitq), 
to_sfixed(358345678.0/4294967296.0,1,-nbitq), 
to_sfixed(184981807.0/4294967296.0,1,-nbitq), 
to_sfixed(491446295.0/4294967296.0,1,-nbitq), 
to_sfixed(-200429264.0/4294967296.0,1,-nbitq), 
to_sfixed(304352226.0/4294967296.0,1,-nbitq), 
to_sfixed(93758383.0/4294967296.0,1,-nbitq), 
to_sfixed(633070877.0/4294967296.0,1,-nbitq), 
to_sfixed(25055103.0/4294967296.0,1,-nbitq), 
to_sfixed(-24463827.0/4294967296.0,1,-nbitq), 
to_sfixed(-529770841.0/4294967296.0,1,-nbitq), 
to_sfixed(-618429447.0/4294967296.0,1,-nbitq), 
to_sfixed(513012685.0/4294967296.0,1,-nbitq), 
to_sfixed(-484377778.0/4294967296.0,1,-nbitq), 
to_sfixed(-822120675.0/4294967296.0,1,-nbitq), 
to_sfixed(1404639791.0/4294967296.0,1,-nbitq), 
to_sfixed(388477047.0/4294967296.0,1,-nbitq), 
to_sfixed(604428264.0/4294967296.0,1,-nbitq), 
to_sfixed(-413357980.0/4294967296.0,1,-nbitq), 
to_sfixed(84711672.0/4294967296.0,1,-nbitq), 
to_sfixed(1880294383.0/4294967296.0,1,-nbitq), 
to_sfixed(-487326386.0/4294967296.0,1,-nbitq), 
to_sfixed(-226458614.0/4294967296.0,1,-nbitq), 
to_sfixed(-8003662.0/4294967296.0,1,-nbitq), 
to_sfixed(119363770.0/4294967296.0,1,-nbitq), 
to_sfixed(-685548033.0/4294967296.0,1,-nbitq), 
to_sfixed(-41091503.0/4294967296.0,1,-nbitq), 
to_sfixed(1339363587.0/4294967296.0,1,-nbitq), 
to_sfixed(24748968.0/4294967296.0,1,-nbitq), 
to_sfixed(22909478.0/4294967296.0,1,-nbitq), 
to_sfixed(-816263073.0/4294967296.0,1,-nbitq), 
to_sfixed(173150344.0/4294967296.0,1,-nbitq), 
to_sfixed(325833489.0/4294967296.0,1,-nbitq), 
to_sfixed(-227157755.0/4294967296.0,1,-nbitq), 
to_sfixed(-953169774.0/4294967296.0,1,-nbitq), 
to_sfixed(-240640877.0/4294967296.0,1,-nbitq), 
to_sfixed(-794676162.0/4294967296.0,1,-nbitq), 
to_sfixed(-1668105908.0/4294967296.0,1,-nbitq), 
to_sfixed(228115867.0/4294967296.0,1,-nbitq), 
to_sfixed(154060791.0/4294967296.0,1,-nbitq), 
to_sfixed(223020893.0/4294967296.0,1,-nbitq), 
to_sfixed(-497234366.0/4294967296.0,1,-nbitq), 
to_sfixed(629945426.0/4294967296.0,1,-nbitq), 
to_sfixed(116153051.0/4294967296.0,1,-nbitq), 
to_sfixed(228952833.0/4294967296.0,1,-nbitq), 
to_sfixed(-109268256.0/4294967296.0,1,-nbitq), 
to_sfixed(452974042.0/4294967296.0,1,-nbitq), 
to_sfixed(1934130198.0/4294967296.0,1,-nbitq), 
to_sfixed(-393284416.0/4294967296.0,1,-nbitq), 
to_sfixed(59462917.0/4294967296.0,1,-nbitq), 
to_sfixed(53584711.0/4294967296.0,1,-nbitq), 
to_sfixed(1472235000.0/4294967296.0,1,-nbitq), 
to_sfixed(487861353.0/4294967296.0,1,-nbitq), 
to_sfixed(-98149708.0/4294967296.0,1,-nbitq), 
to_sfixed(218756646.0/4294967296.0,1,-nbitq), 
to_sfixed(-807273903.0/4294967296.0,1,-nbitq), 
to_sfixed(30423525.0/4294967296.0,1,-nbitq), 
to_sfixed(833671167.0/4294967296.0,1,-nbitq), 
to_sfixed(248640906.0/4294967296.0,1,-nbitq), 
to_sfixed(126667113.0/4294967296.0,1,-nbitq), 
to_sfixed(-111975179.0/4294967296.0,1,-nbitq), 
to_sfixed(-38242780.0/4294967296.0,1,-nbitq), 
to_sfixed(189214723.0/4294967296.0,1,-nbitq), 
to_sfixed(-56127195.0/4294967296.0,1,-nbitq), 
to_sfixed(-140616564.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-600736050.0/4294967296.0,1,-nbitq), 
to_sfixed(-971433064.0/4294967296.0,1,-nbitq), 
to_sfixed(-1205430888.0/4294967296.0,1,-nbitq), 
to_sfixed(445658702.0/4294967296.0,1,-nbitq), 
to_sfixed(-1012190931.0/4294967296.0,1,-nbitq), 
to_sfixed(375808188.0/4294967296.0,1,-nbitq), 
to_sfixed(500070480.0/4294967296.0,1,-nbitq), 
to_sfixed(-1203715083.0/4294967296.0,1,-nbitq), 
to_sfixed(115843584.0/4294967296.0,1,-nbitq), 
to_sfixed(94649952.0/4294967296.0,1,-nbitq), 
to_sfixed(599213169.0/4294967296.0,1,-nbitq), 
to_sfixed(1002169215.0/4294967296.0,1,-nbitq), 
to_sfixed(-1635623866.0/4294967296.0,1,-nbitq), 
to_sfixed(-516741525.0/4294967296.0,1,-nbitq), 
to_sfixed(-35995845.0/4294967296.0,1,-nbitq), 
to_sfixed(-285646559.0/4294967296.0,1,-nbitq), 
to_sfixed(-108348390.0/4294967296.0,1,-nbitq), 
to_sfixed(-252686614.0/4294967296.0,1,-nbitq), 
to_sfixed(568458321.0/4294967296.0,1,-nbitq), 
to_sfixed(-482304621.0/4294967296.0,1,-nbitq), 
to_sfixed(11319813.0/4294967296.0,1,-nbitq), 
to_sfixed(14732185.0/4294967296.0,1,-nbitq), 
to_sfixed(1196240951.0/4294967296.0,1,-nbitq), 
to_sfixed(993246943.0/4294967296.0,1,-nbitq), 
to_sfixed(-156786750.0/4294967296.0,1,-nbitq), 
to_sfixed(1098567931.0/4294967296.0,1,-nbitq), 
to_sfixed(-279797957.0/4294967296.0,1,-nbitq), 
to_sfixed(-599328256.0/4294967296.0,1,-nbitq), 
to_sfixed(-1496745001.0/4294967296.0,1,-nbitq), 
to_sfixed(-700567111.0/4294967296.0,1,-nbitq), 
to_sfixed(790976054.0/4294967296.0,1,-nbitq), 
to_sfixed(-143332008.0/4294967296.0,1,-nbitq), 
to_sfixed(290746969.0/4294967296.0,1,-nbitq), 
to_sfixed(-714859085.0/4294967296.0,1,-nbitq), 
to_sfixed(-380870657.0/4294967296.0,1,-nbitq), 
to_sfixed(2641678267.0/4294967296.0,1,-nbitq), 
to_sfixed(-880954431.0/4294967296.0,1,-nbitq), 
to_sfixed(-43299581.0/4294967296.0,1,-nbitq), 
to_sfixed(-594155536.0/4294967296.0,1,-nbitq), 
to_sfixed(421322580.0/4294967296.0,1,-nbitq), 
to_sfixed(-171039019.0/4294967296.0,1,-nbitq), 
to_sfixed(45501499.0/4294967296.0,1,-nbitq), 
to_sfixed(784518360.0/4294967296.0,1,-nbitq), 
to_sfixed(-916180877.0/4294967296.0,1,-nbitq), 
to_sfixed(-8118212.0/4294967296.0,1,-nbitq), 
to_sfixed(106259186.0/4294967296.0,1,-nbitq), 
to_sfixed(-176875104.0/4294967296.0,1,-nbitq), 
to_sfixed(753662747.0/4294967296.0,1,-nbitq), 
to_sfixed(317884649.0/4294967296.0,1,-nbitq), 
to_sfixed(-608402412.0/4294967296.0,1,-nbitq), 
to_sfixed(503833198.0/4294967296.0,1,-nbitq), 
to_sfixed(-309169855.0/4294967296.0,1,-nbitq), 
to_sfixed(-1611284367.0/4294967296.0,1,-nbitq), 
to_sfixed(-114750311.0/4294967296.0,1,-nbitq), 
to_sfixed(-27000603.0/4294967296.0,1,-nbitq), 
to_sfixed(-782284060.0/4294967296.0,1,-nbitq), 
to_sfixed(-1025171599.0/4294967296.0,1,-nbitq), 
to_sfixed(709510761.0/4294967296.0,1,-nbitq), 
to_sfixed(-170018384.0/4294967296.0,1,-nbitq), 
to_sfixed(-196176218.0/4294967296.0,1,-nbitq), 
to_sfixed(-283997727.0/4294967296.0,1,-nbitq), 
to_sfixed(228176603.0/4294967296.0,1,-nbitq), 
to_sfixed(792585508.0/4294967296.0,1,-nbitq), 
to_sfixed(-368248454.0/4294967296.0,1,-nbitq), 
to_sfixed(587496187.0/4294967296.0,1,-nbitq), 
to_sfixed(-280695585.0/4294967296.0,1,-nbitq), 
to_sfixed(283372453.0/4294967296.0,1,-nbitq), 
to_sfixed(660306222.0/4294967296.0,1,-nbitq), 
to_sfixed(293416643.0/4294967296.0,1,-nbitq), 
to_sfixed(-521792616.0/4294967296.0,1,-nbitq), 
to_sfixed(-366969956.0/4294967296.0,1,-nbitq), 
to_sfixed(314431412.0/4294967296.0,1,-nbitq), 
to_sfixed(124286037.0/4294967296.0,1,-nbitq), 
to_sfixed(124293909.0/4294967296.0,1,-nbitq), 
to_sfixed(129370625.0/4294967296.0,1,-nbitq), 
to_sfixed(-540047796.0/4294967296.0,1,-nbitq), 
to_sfixed(304037107.0/4294967296.0,1,-nbitq), 
to_sfixed(538050326.0/4294967296.0,1,-nbitq), 
to_sfixed(-563212174.0/4294967296.0,1,-nbitq), 
to_sfixed(-213594001.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-160807326.0/4294967296.0,1,-nbitq), 
to_sfixed(-448850125.0/4294967296.0,1,-nbitq), 
to_sfixed(-543022086.0/4294967296.0,1,-nbitq), 
to_sfixed(217093580.0/4294967296.0,1,-nbitq), 
to_sfixed(-953912517.0/4294967296.0,1,-nbitq), 
to_sfixed(-481051224.0/4294967296.0,1,-nbitq), 
to_sfixed(193365962.0/4294967296.0,1,-nbitq), 
to_sfixed(-514512249.0/4294967296.0,1,-nbitq), 
to_sfixed(1240764993.0/4294967296.0,1,-nbitq), 
to_sfixed(-384820983.0/4294967296.0,1,-nbitq), 
to_sfixed(209636864.0/4294967296.0,1,-nbitq), 
to_sfixed(58432458.0/4294967296.0,1,-nbitq), 
to_sfixed(-936340276.0/4294967296.0,1,-nbitq), 
to_sfixed(185632647.0/4294967296.0,1,-nbitq), 
to_sfixed(-146083249.0/4294967296.0,1,-nbitq), 
to_sfixed(-46049269.0/4294967296.0,1,-nbitq), 
to_sfixed(318789827.0/4294967296.0,1,-nbitq), 
to_sfixed(111064697.0/4294967296.0,1,-nbitq), 
to_sfixed(-1349859981.0/4294967296.0,1,-nbitq), 
to_sfixed(-293862882.0/4294967296.0,1,-nbitq), 
to_sfixed(216209752.0/4294967296.0,1,-nbitq), 
to_sfixed(56322965.0/4294967296.0,1,-nbitq), 
to_sfixed(1205355500.0/4294967296.0,1,-nbitq), 
to_sfixed(629425561.0/4294967296.0,1,-nbitq), 
to_sfixed(148910631.0/4294967296.0,1,-nbitq), 
to_sfixed(480197289.0/4294967296.0,1,-nbitq), 
to_sfixed(-879892890.0/4294967296.0,1,-nbitq), 
to_sfixed(-1663959502.0/4294967296.0,1,-nbitq), 
to_sfixed(-480831691.0/4294967296.0,1,-nbitq), 
to_sfixed(-282700843.0/4294967296.0,1,-nbitq), 
to_sfixed(152182044.0/4294967296.0,1,-nbitq), 
to_sfixed(246279939.0/4294967296.0,1,-nbitq), 
to_sfixed(463124848.0/4294967296.0,1,-nbitq), 
to_sfixed(-842806089.0/4294967296.0,1,-nbitq), 
to_sfixed(-37376720.0/4294967296.0,1,-nbitq), 
to_sfixed(1360777037.0/4294967296.0,1,-nbitq), 
to_sfixed(-337264627.0/4294967296.0,1,-nbitq), 
to_sfixed(200813964.0/4294967296.0,1,-nbitq), 
to_sfixed(-604706564.0/4294967296.0,1,-nbitq), 
to_sfixed(454726493.0/4294967296.0,1,-nbitq), 
to_sfixed(335043855.0/4294967296.0,1,-nbitq), 
to_sfixed(-74882945.0/4294967296.0,1,-nbitq), 
to_sfixed(367792649.0/4294967296.0,1,-nbitq), 
to_sfixed(-559136653.0/4294967296.0,1,-nbitq), 
to_sfixed(-112482229.0/4294967296.0,1,-nbitq), 
to_sfixed(-545829037.0/4294967296.0,1,-nbitq), 
to_sfixed(299035597.0/4294967296.0,1,-nbitq), 
to_sfixed(70230228.0/4294967296.0,1,-nbitq), 
to_sfixed(546661669.0/4294967296.0,1,-nbitq), 
to_sfixed(-861859348.0/4294967296.0,1,-nbitq), 
to_sfixed(1337238452.0/4294967296.0,1,-nbitq), 
to_sfixed(-217954721.0/4294967296.0,1,-nbitq), 
to_sfixed(-594380311.0/4294967296.0,1,-nbitq), 
to_sfixed(290287508.0/4294967296.0,1,-nbitq), 
to_sfixed(666798069.0/4294967296.0,1,-nbitq), 
to_sfixed(-85198083.0/4294967296.0,1,-nbitq), 
to_sfixed(-815102245.0/4294967296.0,1,-nbitq), 
to_sfixed(-52823067.0/4294967296.0,1,-nbitq), 
to_sfixed(227557439.0/4294967296.0,1,-nbitq), 
to_sfixed(-192041591.0/4294967296.0,1,-nbitq), 
to_sfixed(-59166019.0/4294967296.0,1,-nbitq), 
to_sfixed(499403320.0/4294967296.0,1,-nbitq), 
to_sfixed(655563116.0/4294967296.0,1,-nbitq), 
to_sfixed(-569864257.0/4294967296.0,1,-nbitq), 
to_sfixed(-289986225.0/4294967296.0,1,-nbitq), 
to_sfixed(-416090122.0/4294967296.0,1,-nbitq), 
to_sfixed(-51535923.0/4294967296.0,1,-nbitq), 
to_sfixed(531923362.0/4294967296.0,1,-nbitq), 
to_sfixed(336989238.0/4294967296.0,1,-nbitq), 
to_sfixed(305374282.0/4294967296.0,1,-nbitq), 
to_sfixed(193027988.0/4294967296.0,1,-nbitq), 
to_sfixed(767164410.0/4294967296.0,1,-nbitq), 
to_sfixed(-115530873.0/4294967296.0,1,-nbitq), 
to_sfixed(-272258295.0/4294967296.0,1,-nbitq), 
to_sfixed(404474542.0/4294967296.0,1,-nbitq), 
to_sfixed(525140646.0/4294967296.0,1,-nbitq), 
to_sfixed(-257525302.0/4294967296.0,1,-nbitq), 
to_sfixed(174530518.0/4294967296.0,1,-nbitq), 
to_sfixed(-221736805.0/4294967296.0,1,-nbitq), 
to_sfixed(-267008424.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(314251379.0/4294967296.0,1,-nbitq), 
to_sfixed(-197937931.0/4294967296.0,1,-nbitq), 
to_sfixed(-188491268.0/4294967296.0,1,-nbitq), 
to_sfixed(316422798.0/4294967296.0,1,-nbitq), 
to_sfixed(-786898189.0/4294967296.0,1,-nbitq), 
to_sfixed(-680786839.0/4294967296.0,1,-nbitq), 
to_sfixed(480829327.0/4294967296.0,1,-nbitq), 
to_sfixed(32027800.0/4294967296.0,1,-nbitq), 
to_sfixed(1081594991.0/4294967296.0,1,-nbitq), 
to_sfixed(-267968698.0/4294967296.0,1,-nbitq), 
to_sfixed(551190506.0/4294967296.0,1,-nbitq), 
to_sfixed(816088532.0/4294967296.0,1,-nbitq), 
to_sfixed(-227621994.0/4294967296.0,1,-nbitq), 
to_sfixed(608209249.0/4294967296.0,1,-nbitq), 
to_sfixed(61680207.0/4294967296.0,1,-nbitq), 
to_sfixed(155808385.0/4294967296.0,1,-nbitq), 
to_sfixed(364667054.0/4294967296.0,1,-nbitq), 
to_sfixed(243018758.0/4294967296.0,1,-nbitq), 
to_sfixed(-538018309.0/4294967296.0,1,-nbitq), 
to_sfixed(-453341318.0/4294967296.0,1,-nbitq), 
to_sfixed(-245595393.0/4294967296.0,1,-nbitq), 
to_sfixed(-602528447.0/4294967296.0,1,-nbitq), 
to_sfixed(489573569.0/4294967296.0,1,-nbitq), 
to_sfixed(-384748172.0/4294967296.0,1,-nbitq), 
to_sfixed(-171950891.0/4294967296.0,1,-nbitq), 
to_sfixed(-367542318.0/4294967296.0,1,-nbitq), 
to_sfixed(-1092581033.0/4294967296.0,1,-nbitq), 
to_sfixed(-758809100.0/4294967296.0,1,-nbitq), 
to_sfixed(-253850974.0/4294967296.0,1,-nbitq), 
to_sfixed(-1445436212.0/4294967296.0,1,-nbitq), 
to_sfixed(-730791653.0/4294967296.0,1,-nbitq), 
to_sfixed(-507133044.0/4294967296.0,1,-nbitq), 
to_sfixed(-274924466.0/4294967296.0,1,-nbitq), 
to_sfixed(-154803228.0/4294967296.0,1,-nbitq), 
to_sfixed(873412203.0/4294967296.0,1,-nbitq), 
to_sfixed(289986627.0/4294967296.0,1,-nbitq), 
to_sfixed(-451910417.0/4294967296.0,1,-nbitq), 
to_sfixed(241981727.0/4294967296.0,1,-nbitq), 
to_sfixed(-256624225.0/4294967296.0,1,-nbitq), 
to_sfixed(-349242731.0/4294967296.0,1,-nbitq), 
to_sfixed(839011525.0/4294967296.0,1,-nbitq), 
to_sfixed(-100463355.0/4294967296.0,1,-nbitq), 
to_sfixed(191365158.0/4294967296.0,1,-nbitq), 
to_sfixed(512291984.0/4294967296.0,1,-nbitq), 
to_sfixed(-313416049.0/4294967296.0,1,-nbitq), 
to_sfixed(-64247514.0/4294967296.0,1,-nbitq), 
to_sfixed(-338001223.0/4294967296.0,1,-nbitq), 
to_sfixed(-307663038.0/4294967296.0,1,-nbitq), 
to_sfixed(277118977.0/4294967296.0,1,-nbitq), 
to_sfixed(-587727726.0/4294967296.0,1,-nbitq), 
to_sfixed(1147991801.0/4294967296.0,1,-nbitq), 
to_sfixed(-192510643.0/4294967296.0,1,-nbitq), 
to_sfixed(-433560234.0/4294967296.0,1,-nbitq), 
to_sfixed(-1179001742.0/4294967296.0,1,-nbitq), 
to_sfixed(396140763.0/4294967296.0,1,-nbitq), 
to_sfixed(-262924835.0/4294967296.0,1,-nbitq), 
to_sfixed(-1436414899.0/4294967296.0,1,-nbitq), 
to_sfixed(250882588.0/4294967296.0,1,-nbitq), 
to_sfixed(241062605.0/4294967296.0,1,-nbitq), 
to_sfixed(172547800.0/4294967296.0,1,-nbitq), 
to_sfixed(-152175848.0/4294967296.0,1,-nbitq), 
to_sfixed(-31270258.0/4294967296.0,1,-nbitq), 
to_sfixed(52761198.0/4294967296.0,1,-nbitq), 
to_sfixed(-206031529.0/4294967296.0,1,-nbitq), 
to_sfixed(-328363818.0/4294967296.0,1,-nbitq), 
to_sfixed(-348553545.0/4294967296.0,1,-nbitq), 
to_sfixed(-689209021.0/4294967296.0,1,-nbitq), 
to_sfixed(302905350.0/4294967296.0,1,-nbitq), 
to_sfixed(115498668.0/4294967296.0,1,-nbitq), 
to_sfixed(-315812118.0/4294967296.0,1,-nbitq), 
to_sfixed(-324161410.0/4294967296.0,1,-nbitq), 
to_sfixed(-276403168.0/4294967296.0,1,-nbitq), 
to_sfixed(-733298598.0/4294967296.0,1,-nbitq), 
to_sfixed(71383975.0/4294967296.0,1,-nbitq), 
to_sfixed(-225933788.0/4294967296.0,1,-nbitq), 
to_sfixed(1036720385.0/4294967296.0,1,-nbitq), 
to_sfixed(-452346797.0/4294967296.0,1,-nbitq), 
to_sfixed(625976456.0/4294967296.0,1,-nbitq), 
to_sfixed(180097503.0/4294967296.0,1,-nbitq), 
to_sfixed(320720330.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(35763382.0/4294967296.0,1,-nbitq), 
to_sfixed(-388769245.0/4294967296.0,1,-nbitq), 
to_sfixed(701895207.0/4294967296.0,1,-nbitq), 
to_sfixed(449749613.0/4294967296.0,1,-nbitq), 
to_sfixed(-2536364.0/4294967296.0,1,-nbitq), 
to_sfixed(97657664.0/4294967296.0,1,-nbitq), 
to_sfixed(753541711.0/4294967296.0,1,-nbitq), 
to_sfixed(129835308.0/4294967296.0,1,-nbitq), 
to_sfixed(933897078.0/4294967296.0,1,-nbitq), 
to_sfixed(142335016.0/4294967296.0,1,-nbitq), 
to_sfixed(585637958.0/4294967296.0,1,-nbitq), 
to_sfixed(970034002.0/4294967296.0,1,-nbitq), 
to_sfixed(143701806.0/4294967296.0,1,-nbitq), 
to_sfixed(988180134.0/4294967296.0,1,-nbitq), 
to_sfixed(279077946.0/4294967296.0,1,-nbitq), 
to_sfixed(882727103.0/4294967296.0,1,-nbitq), 
to_sfixed(99481720.0/4294967296.0,1,-nbitq), 
to_sfixed(-94587782.0/4294967296.0,1,-nbitq), 
to_sfixed(-572034442.0/4294967296.0,1,-nbitq), 
to_sfixed(-81172397.0/4294967296.0,1,-nbitq), 
to_sfixed(262953101.0/4294967296.0,1,-nbitq), 
to_sfixed(-316880920.0/4294967296.0,1,-nbitq), 
to_sfixed(-341064950.0/4294967296.0,1,-nbitq), 
to_sfixed(-1246728415.0/4294967296.0,1,-nbitq), 
to_sfixed(122528716.0/4294967296.0,1,-nbitq), 
to_sfixed(-4812399.0/4294967296.0,1,-nbitq), 
to_sfixed(-456015214.0/4294967296.0,1,-nbitq), 
to_sfixed(-419596907.0/4294967296.0,1,-nbitq), 
to_sfixed(-182249482.0/4294967296.0,1,-nbitq), 
to_sfixed(-1047454532.0/4294967296.0,1,-nbitq), 
to_sfixed(-886563820.0/4294967296.0,1,-nbitq), 
to_sfixed(-543885371.0/4294967296.0,1,-nbitq), 
to_sfixed(-712960166.0/4294967296.0,1,-nbitq), 
to_sfixed(905311197.0/4294967296.0,1,-nbitq), 
to_sfixed(88664461.0/4294967296.0,1,-nbitq), 
to_sfixed(153979266.0/4294967296.0,1,-nbitq), 
to_sfixed(-355550754.0/4294967296.0,1,-nbitq), 
to_sfixed(869604783.0/4294967296.0,1,-nbitq), 
to_sfixed(-243740365.0/4294967296.0,1,-nbitq), 
to_sfixed(-219354644.0/4294967296.0,1,-nbitq), 
to_sfixed(936416146.0/4294967296.0,1,-nbitq), 
to_sfixed(90965145.0/4294967296.0,1,-nbitq), 
to_sfixed(65172532.0/4294967296.0,1,-nbitq), 
to_sfixed(1505372105.0/4294967296.0,1,-nbitq), 
to_sfixed(179618100.0/4294967296.0,1,-nbitq), 
to_sfixed(354937300.0/4294967296.0,1,-nbitq), 
to_sfixed(-127594867.0/4294967296.0,1,-nbitq), 
to_sfixed(-532464579.0/4294967296.0,1,-nbitq), 
to_sfixed(382943731.0/4294967296.0,1,-nbitq), 
to_sfixed(693612589.0/4294967296.0,1,-nbitq), 
to_sfixed(559893240.0/4294967296.0,1,-nbitq), 
to_sfixed(721729299.0/4294967296.0,1,-nbitq), 
to_sfixed(151341421.0/4294967296.0,1,-nbitq), 
to_sfixed(-541884694.0/4294967296.0,1,-nbitq), 
to_sfixed(345741575.0/4294967296.0,1,-nbitq), 
to_sfixed(627183811.0/4294967296.0,1,-nbitq), 
to_sfixed(-736501194.0/4294967296.0,1,-nbitq), 
to_sfixed(665555166.0/4294967296.0,1,-nbitq), 
to_sfixed(252222855.0/4294967296.0,1,-nbitq), 
to_sfixed(155776767.0/4294967296.0,1,-nbitq), 
to_sfixed(-365399156.0/4294967296.0,1,-nbitq), 
to_sfixed(-195226303.0/4294967296.0,1,-nbitq), 
to_sfixed(-958906763.0/4294967296.0,1,-nbitq), 
to_sfixed(-776828459.0/4294967296.0,1,-nbitq), 
to_sfixed(-654285964.0/4294967296.0,1,-nbitq), 
to_sfixed(-199115236.0/4294967296.0,1,-nbitq), 
to_sfixed(-1419347110.0/4294967296.0,1,-nbitq), 
to_sfixed(-95156519.0/4294967296.0,1,-nbitq), 
to_sfixed(321345627.0/4294967296.0,1,-nbitq), 
to_sfixed(-653995541.0/4294967296.0,1,-nbitq), 
to_sfixed(584530094.0/4294967296.0,1,-nbitq), 
to_sfixed(-166854262.0/4294967296.0,1,-nbitq), 
to_sfixed(-433366126.0/4294967296.0,1,-nbitq), 
to_sfixed(-71162930.0/4294967296.0,1,-nbitq), 
to_sfixed(-31067535.0/4294967296.0,1,-nbitq), 
to_sfixed(941513827.0/4294967296.0,1,-nbitq), 
to_sfixed(52483287.0/4294967296.0,1,-nbitq), 
to_sfixed(481712196.0/4294967296.0,1,-nbitq), 
to_sfixed(908479191.0/4294967296.0,1,-nbitq), 
to_sfixed(-147289861.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(221980815.0/4294967296.0,1,-nbitq), 
to_sfixed(255611966.0/4294967296.0,1,-nbitq), 
to_sfixed(1401071873.0/4294967296.0,1,-nbitq), 
to_sfixed(-391220754.0/4294967296.0,1,-nbitq), 
to_sfixed(70978727.0/4294967296.0,1,-nbitq), 
to_sfixed(241245322.0/4294967296.0,1,-nbitq), 
to_sfixed(190955996.0/4294967296.0,1,-nbitq), 
to_sfixed(603411355.0/4294967296.0,1,-nbitq), 
to_sfixed(456915660.0/4294967296.0,1,-nbitq), 
to_sfixed(-98515132.0/4294967296.0,1,-nbitq), 
to_sfixed(20597104.0/4294967296.0,1,-nbitq), 
to_sfixed(480086594.0/4294967296.0,1,-nbitq), 
to_sfixed(-30087558.0/4294967296.0,1,-nbitq), 
to_sfixed(243644723.0/4294967296.0,1,-nbitq), 
to_sfixed(233063276.0/4294967296.0,1,-nbitq), 
to_sfixed(660458362.0/4294967296.0,1,-nbitq), 
to_sfixed(209812762.0/4294967296.0,1,-nbitq), 
to_sfixed(238967059.0/4294967296.0,1,-nbitq), 
to_sfixed(-263046876.0/4294967296.0,1,-nbitq), 
to_sfixed(-41652822.0/4294967296.0,1,-nbitq), 
to_sfixed(-311096799.0/4294967296.0,1,-nbitq), 
to_sfixed(125955004.0/4294967296.0,1,-nbitq), 
to_sfixed(-1213916233.0/4294967296.0,1,-nbitq), 
to_sfixed(-33762563.0/4294967296.0,1,-nbitq), 
to_sfixed(-184319820.0/4294967296.0,1,-nbitq), 
to_sfixed(1173376684.0/4294967296.0,1,-nbitq), 
to_sfixed(-1060207247.0/4294967296.0,1,-nbitq), 
to_sfixed(-97415638.0/4294967296.0,1,-nbitq), 
to_sfixed(887896986.0/4294967296.0,1,-nbitq), 
to_sfixed(-817014394.0/4294967296.0,1,-nbitq), 
to_sfixed(-805545711.0/4294967296.0,1,-nbitq), 
to_sfixed(-1028634821.0/4294967296.0,1,-nbitq), 
to_sfixed(-885504045.0/4294967296.0,1,-nbitq), 
to_sfixed(826868402.0/4294967296.0,1,-nbitq), 
to_sfixed(-469750115.0/4294967296.0,1,-nbitq), 
to_sfixed(439012877.0/4294967296.0,1,-nbitq), 
to_sfixed(716838377.0/4294967296.0,1,-nbitq), 
to_sfixed(765390914.0/4294967296.0,1,-nbitq), 
to_sfixed(-258009481.0/4294967296.0,1,-nbitq), 
to_sfixed(28092068.0/4294967296.0,1,-nbitq), 
to_sfixed(1025063766.0/4294967296.0,1,-nbitq), 
to_sfixed(488242142.0/4294967296.0,1,-nbitq), 
to_sfixed(176917848.0/4294967296.0,1,-nbitq), 
to_sfixed(1405971341.0/4294967296.0,1,-nbitq), 
to_sfixed(360352039.0/4294967296.0,1,-nbitq), 
to_sfixed(637095301.0/4294967296.0,1,-nbitq), 
to_sfixed(-269637352.0/4294967296.0,1,-nbitq), 
to_sfixed(-557387252.0/4294967296.0,1,-nbitq), 
to_sfixed(84228656.0/4294967296.0,1,-nbitq), 
to_sfixed(616486779.0/4294967296.0,1,-nbitq), 
to_sfixed(447415664.0/4294967296.0,1,-nbitq), 
to_sfixed(336683882.0/4294967296.0,1,-nbitq), 
to_sfixed(-1546841780.0/4294967296.0,1,-nbitq), 
to_sfixed(139926645.0/4294967296.0,1,-nbitq), 
to_sfixed(-408318555.0/4294967296.0,1,-nbitq), 
to_sfixed(-94269758.0/4294967296.0,1,-nbitq), 
to_sfixed(-177128453.0/4294967296.0,1,-nbitq), 
to_sfixed(853375628.0/4294967296.0,1,-nbitq), 
to_sfixed(-126427157.0/4294967296.0,1,-nbitq), 
to_sfixed(-341544890.0/4294967296.0,1,-nbitq), 
to_sfixed(91330049.0/4294967296.0,1,-nbitq), 
to_sfixed(-692395971.0/4294967296.0,1,-nbitq), 
to_sfixed(-993653670.0/4294967296.0,1,-nbitq), 
to_sfixed(-805059477.0/4294967296.0,1,-nbitq), 
to_sfixed(-578413075.0/4294967296.0,1,-nbitq), 
to_sfixed(-392083794.0/4294967296.0,1,-nbitq), 
to_sfixed(-1551133454.0/4294967296.0,1,-nbitq), 
to_sfixed(465668299.0/4294967296.0,1,-nbitq), 
to_sfixed(234764062.0/4294967296.0,1,-nbitq), 
to_sfixed(-504450408.0/4294967296.0,1,-nbitq), 
to_sfixed(766466670.0/4294967296.0,1,-nbitq), 
to_sfixed(-350108975.0/4294967296.0,1,-nbitq), 
to_sfixed(-384674687.0/4294967296.0,1,-nbitq), 
to_sfixed(331856504.0/4294967296.0,1,-nbitq), 
to_sfixed(3901127.0/4294967296.0,1,-nbitq), 
to_sfixed(382940136.0/4294967296.0,1,-nbitq), 
to_sfixed(-167879147.0/4294967296.0,1,-nbitq), 
to_sfixed(163966836.0/4294967296.0,1,-nbitq), 
to_sfixed(566679657.0/4294967296.0,1,-nbitq), 
to_sfixed(154841730.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-99300239.0/4294967296.0,1,-nbitq), 
to_sfixed(136500689.0/4294967296.0,1,-nbitq), 
to_sfixed(1397515527.0/4294967296.0,1,-nbitq), 
to_sfixed(-155775185.0/4294967296.0,1,-nbitq), 
to_sfixed(-359772934.0/4294967296.0,1,-nbitq), 
to_sfixed(-542567322.0/4294967296.0,1,-nbitq), 
to_sfixed(-260946704.0/4294967296.0,1,-nbitq), 
to_sfixed(22623334.0/4294967296.0,1,-nbitq), 
to_sfixed(1187589206.0/4294967296.0,1,-nbitq), 
to_sfixed(218475796.0/4294967296.0,1,-nbitq), 
to_sfixed(54841208.0/4294967296.0,1,-nbitq), 
to_sfixed(19664154.0/4294967296.0,1,-nbitq), 
to_sfixed(-358244126.0/4294967296.0,1,-nbitq), 
to_sfixed(1219172789.0/4294967296.0,1,-nbitq), 
to_sfixed(-236225399.0/4294967296.0,1,-nbitq), 
to_sfixed(694292832.0/4294967296.0,1,-nbitq), 
to_sfixed(196889518.0/4294967296.0,1,-nbitq), 
to_sfixed(-170159400.0/4294967296.0,1,-nbitq), 
to_sfixed(-45429361.0/4294967296.0,1,-nbitq), 
to_sfixed(-294999658.0/4294967296.0,1,-nbitq), 
to_sfixed(326397282.0/4294967296.0,1,-nbitq), 
to_sfixed(157931700.0/4294967296.0,1,-nbitq), 
to_sfixed(-1094611671.0/4294967296.0,1,-nbitq), 
to_sfixed(149117482.0/4294967296.0,1,-nbitq), 
to_sfixed(-304263463.0/4294967296.0,1,-nbitq), 
to_sfixed(585173778.0/4294967296.0,1,-nbitq), 
to_sfixed(-408559727.0/4294967296.0,1,-nbitq), 
to_sfixed(650043424.0/4294967296.0,1,-nbitq), 
to_sfixed(477315779.0/4294967296.0,1,-nbitq), 
to_sfixed(-113024183.0/4294967296.0,1,-nbitq), 
to_sfixed(-389086912.0/4294967296.0,1,-nbitq), 
to_sfixed(-488867158.0/4294967296.0,1,-nbitq), 
to_sfixed(-544146729.0/4294967296.0,1,-nbitq), 
to_sfixed(667062100.0/4294967296.0,1,-nbitq), 
to_sfixed(201149373.0/4294967296.0,1,-nbitq), 
to_sfixed(425353731.0/4294967296.0,1,-nbitq), 
to_sfixed(698188212.0/4294967296.0,1,-nbitq), 
to_sfixed(782692780.0/4294967296.0,1,-nbitq), 
to_sfixed(262716370.0/4294967296.0,1,-nbitq), 
to_sfixed(200637898.0/4294967296.0,1,-nbitq), 
to_sfixed(804285268.0/4294967296.0,1,-nbitq), 
to_sfixed(997296666.0/4294967296.0,1,-nbitq), 
to_sfixed(-361131083.0/4294967296.0,1,-nbitq), 
to_sfixed(1901352254.0/4294967296.0,1,-nbitq), 
to_sfixed(273908908.0/4294967296.0,1,-nbitq), 
to_sfixed(344052092.0/4294967296.0,1,-nbitq), 
to_sfixed(-52142867.0/4294967296.0,1,-nbitq), 
to_sfixed(14943296.0/4294967296.0,1,-nbitq), 
to_sfixed(-478751525.0/4294967296.0,1,-nbitq), 
to_sfixed(639290786.0/4294967296.0,1,-nbitq), 
to_sfixed(635240039.0/4294967296.0,1,-nbitq), 
to_sfixed(822412926.0/4294967296.0,1,-nbitq), 
to_sfixed(-2193065250.0/4294967296.0,1,-nbitq), 
to_sfixed(401287238.0/4294967296.0,1,-nbitq), 
to_sfixed(-1082245152.0/4294967296.0,1,-nbitq), 
to_sfixed(869910803.0/4294967296.0,1,-nbitq), 
to_sfixed(570571730.0/4294967296.0,1,-nbitq), 
to_sfixed(1320516101.0/4294967296.0,1,-nbitq), 
to_sfixed(-118472672.0/4294967296.0,1,-nbitq), 
to_sfixed(-124774335.0/4294967296.0,1,-nbitq), 
to_sfixed(-159497515.0/4294967296.0,1,-nbitq), 
to_sfixed(-938438903.0/4294967296.0,1,-nbitq), 
to_sfixed(-24677435.0/4294967296.0,1,-nbitq), 
to_sfixed(-167440565.0/4294967296.0,1,-nbitq), 
to_sfixed(-131813646.0/4294967296.0,1,-nbitq), 
to_sfixed(-314013632.0/4294967296.0,1,-nbitq), 
to_sfixed(-693673223.0/4294967296.0,1,-nbitq), 
to_sfixed(-459792994.0/4294967296.0,1,-nbitq), 
to_sfixed(204538091.0/4294967296.0,1,-nbitq), 
to_sfixed(-692377335.0/4294967296.0,1,-nbitq), 
to_sfixed(463179174.0/4294967296.0,1,-nbitq), 
to_sfixed(70538603.0/4294967296.0,1,-nbitq), 
to_sfixed(-644819153.0/4294967296.0,1,-nbitq), 
to_sfixed(-230681441.0/4294967296.0,1,-nbitq), 
to_sfixed(131848187.0/4294967296.0,1,-nbitq), 
to_sfixed(-244368390.0/4294967296.0,1,-nbitq), 
to_sfixed(-166127860.0/4294967296.0,1,-nbitq), 
to_sfixed(-324240681.0/4294967296.0,1,-nbitq), 
to_sfixed(311714308.0/4294967296.0,1,-nbitq), 
to_sfixed(317395066.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-120933990.0/4294967296.0,1,-nbitq), 
to_sfixed(-718563241.0/4294967296.0,1,-nbitq), 
to_sfixed(1792983171.0/4294967296.0,1,-nbitq), 
to_sfixed(87960903.0/4294967296.0,1,-nbitq), 
to_sfixed(-485717003.0/4294967296.0,1,-nbitq), 
to_sfixed(-700182005.0/4294967296.0,1,-nbitq), 
to_sfixed(-251374830.0/4294967296.0,1,-nbitq), 
to_sfixed(245251455.0/4294967296.0,1,-nbitq), 
to_sfixed(796356574.0/4294967296.0,1,-nbitq), 
to_sfixed(152006611.0/4294967296.0,1,-nbitq), 
to_sfixed(-185950194.0/4294967296.0,1,-nbitq), 
to_sfixed(569039356.0/4294967296.0,1,-nbitq), 
to_sfixed(-237272286.0/4294967296.0,1,-nbitq), 
to_sfixed(547652880.0/4294967296.0,1,-nbitq), 
to_sfixed(380349678.0/4294967296.0,1,-nbitq), 
to_sfixed(658761587.0/4294967296.0,1,-nbitq), 
to_sfixed(30028295.0/4294967296.0,1,-nbitq), 
to_sfixed(154582657.0/4294967296.0,1,-nbitq), 
to_sfixed(-379742044.0/4294967296.0,1,-nbitq), 
to_sfixed(-541206472.0/4294967296.0,1,-nbitq), 
to_sfixed(-280599538.0/4294967296.0,1,-nbitq), 
to_sfixed(974019808.0/4294967296.0,1,-nbitq), 
to_sfixed(-952934763.0/4294967296.0,1,-nbitq), 
to_sfixed(124617165.0/4294967296.0,1,-nbitq), 
to_sfixed(-359529635.0/4294967296.0,1,-nbitq), 
to_sfixed(-760998679.0/4294967296.0,1,-nbitq), 
to_sfixed(311006006.0/4294967296.0,1,-nbitq), 
to_sfixed(1025323065.0/4294967296.0,1,-nbitq), 
to_sfixed(-306036617.0/4294967296.0,1,-nbitq), 
to_sfixed(1140479483.0/4294967296.0,1,-nbitq), 
to_sfixed(454250053.0/4294967296.0,1,-nbitq), 
to_sfixed(-471113384.0/4294967296.0,1,-nbitq), 
to_sfixed(-792887520.0/4294967296.0,1,-nbitq), 
to_sfixed(397822825.0/4294967296.0,1,-nbitq), 
to_sfixed(344942569.0/4294967296.0,1,-nbitq), 
to_sfixed(440723438.0/4294967296.0,1,-nbitq), 
to_sfixed(692978929.0/4294967296.0,1,-nbitq), 
to_sfixed(422615137.0/4294967296.0,1,-nbitq), 
to_sfixed(525323534.0/4294967296.0,1,-nbitq), 
to_sfixed(46857529.0/4294967296.0,1,-nbitq), 
to_sfixed(526726082.0/4294967296.0,1,-nbitq), 
to_sfixed(313457528.0/4294967296.0,1,-nbitq), 
to_sfixed(-980707225.0/4294967296.0,1,-nbitq), 
to_sfixed(1169422380.0/4294967296.0,1,-nbitq), 
to_sfixed(-115561450.0/4294967296.0,1,-nbitq), 
to_sfixed(350171276.0/4294967296.0,1,-nbitq), 
to_sfixed(183903067.0/4294967296.0,1,-nbitq), 
to_sfixed(42100756.0/4294967296.0,1,-nbitq), 
to_sfixed(-1009048167.0/4294967296.0,1,-nbitq), 
to_sfixed(317850200.0/4294967296.0,1,-nbitq), 
to_sfixed(70840364.0/4294967296.0,1,-nbitq), 
to_sfixed(948111945.0/4294967296.0,1,-nbitq), 
to_sfixed(-761923670.0/4294967296.0,1,-nbitq), 
to_sfixed(853123983.0/4294967296.0,1,-nbitq), 
to_sfixed(-1224291625.0/4294967296.0,1,-nbitq), 
to_sfixed(1307914551.0/4294967296.0,1,-nbitq), 
to_sfixed(475951415.0/4294967296.0,1,-nbitq), 
to_sfixed(1091069529.0/4294967296.0,1,-nbitq), 
to_sfixed(-155039760.0/4294967296.0,1,-nbitq), 
to_sfixed(82337100.0/4294967296.0,1,-nbitq), 
to_sfixed(-184670150.0/4294967296.0,1,-nbitq), 
to_sfixed(-289126323.0/4294967296.0,1,-nbitq), 
to_sfixed(-603598334.0/4294967296.0,1,-nbitq), 
to_sfixed(-190250712.0/4294967296.0,1,-nbitq), 
to_sfixed(-79720211.0/4294967296.0,1,-nbitq), 
to_sfixed(-343033587.0/4294967296.0,1,-nbitq), 
to_sfixed(160691169.0/4294967296.0,1,-nbitq), 
to_sfixed(-68871851.0/4294967296.0,1,-nbitq), 
to_sfixed(-144510926.0/4294967296.0,1,-nbitq), 
to_sfixed(201731924.0/4294967296.0,1,-nbitq), 
to_sfixed(350403400.0/4294967296.0,1,-nbitq), 
to_sfixed(108134430.0/4294967296.0,1,-nbitq), 
to_sfixed(-367216163.0/4294967296.0,1,-nbitq), 
to_sfixed(384096449.0/4294967296.0,1,-nbitq), 
to_sfixed(-188560486.0/4294967296.0,1,-nbitq), 
to_sfixed(440703690.0/4294967296.0,1,-nbitq), 
to_sfixed(-265854688.0/4294967296.0,1,-nbitq), 
to_sfixed(-367249203.0/4294967296.0,1,-nbitq), 
to_sfixed(812787126.0/4294967296.0,1,-nbitq), 
to_sfixed(-69674492.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(214351220.0/4294967296.0,1,-nbitq), 
to_sfixed(-883850153.0/4294967296.0,1,-nbitq), 
to_sfixed(894794818.0/4294967296.0,1,-nbitq), 
to_sfixed(635023013.0/4294967296.0,1,-nbitq), 
to_sfixed(-637569489.0/4294967296.0,1,-nbitq), 
to_sfixed(-748060493.0/4294967296.0,1,-nbitq), 
to_sfixed(-473967133.0/4294967296.0,1,-nbitq), 
to_sfixed(-176477553.0/4294967296.0,1,-nbitq), 
to_sfixed(925499103.0/4294967296.0,1,-nbitq), 
to_sfixed(-289313714.0/4294967296.0,1,-nbitq), 
to_sfixed(-918124827.0/4294967296.0,1,-nbitq), 
to_sfixed(145094559.0/4294967296.0,1,-nbitq), 
to_sfixed(-1053181805.0/4294967296.0,1,-nbitq), 
to_sfixed(398473370.0/4294967296.0,1,-nbitq), 
to_sfixed(142755527.0/4294967296.0,1,-nbitq), 
to_sfixed(687589657.0/4294967296.0,1,-nbitq), 
to_sfixed(-194717934.0/4294967296.0,1,-nbitq), 
to_sfixed(-246047392.0/4294967296.0,1,-nbitq), 
to_sfixed(-693635383.0/4294967296.0,1,-nbitq), 
to_sfixed(-343908475.0/4294967296.0,1,-nbitq), 
to_sfixed(113893664.0/4294967296.0,1,-nbitq), 
to_sfixed(683471037.0/4294967296.0,1,-nbitq), 
to_sfixed(-660025708.0/4294967296.0,1,-nbitq), 
to_sfixed(312795986.0/4294967296.0,1,-nbitq), 
to_sfixed(263700946.0/4294967296.0,1,-nbitq), 
to_sfixed(-397132120.0/4294967296.0,1,-nbitq), 
to_sfixed(514498926.0/4294967296.0,1,-nbitq), 
to_sfixed(816639467.0/4294967296.0,1,-nbitq), 
to_sfixed(-13550489.0/4294967296.0,1,-nbitq), 
to_sfixed(1237649456.0/4294967296.0,1,-nbitq), 
to_sfixed(1017286694.0/4294967296.0,1,-nbitq), 
to_sfixed(-112779837.0/4294967296.0,1,-nbitq), 
to_sfixed(-1234779565.0/4294967296.0,1,-nbitq), 
to_sfixed(-122586135.0/4294967296.0,1,-nbitq), 
to_sfixed(60985509.0/4294967296.0,1,-nbitq), 
to_sfixed(-79283849.0/4294967296.0,1,-nbitq), 
to_sfixed(-208784645.0/4294967296.0,1,-nbitq), 
to_sfixed(452995577.0/4294967296.0,1,-nbitq), 
to_sfixed(37282657.0/4294967296.0,1,-nbitq), 
to_sfixed(-37105667.0/4294967296.0,1,-nbitq), 
to_sfixed(457964918.0/4294967296.0,1,-nbitq), 
to_sfixed(-500368012.0/4294967296.0,1,-nbitq), 
to_sfixed(-821990280.0/4294967296.0,1,-nbitq), 
to_sfixed(222760325.0/4294967296.0,1,-nbitq), 
to_sfixed(671191959.0/4294967296.0,1,-nbitq), 
to_sfixed(-28104877.0/4294967296.0,1,-nbitq), 
to_sfixed(189555995.0/4294967296.0,1,-nbitq), 
to_sfixed(-452632987.0/4294967296.0,1,-nbitq), 
to_sfixed(-1308333437.0/4294967296.0,1,-nbitq), 
to_sfixed(262412525.0/4294967296.0,1,-nbitq), 
to_sfixed(-308422735.0/4294967296.0,1,-nbitq), 
to_sfixed(234507065.0/4294967296.0,1,-nbitq), 
to_sfixed(-173844169.0/4294967296.0,1,-nbitq), 
to_sfixed(-101468693.0/4294967296.0,1,-nbitq), 
to_sfixed(-1765533018.0/4294967296.0,1,-nbitq), 
to_sfixed(401907536.0/4294967296.0,1,-nbitq), 
to_sfixed(136250031.0/4294967296.0,1,-nbitq), 
to_sfixed(349117765.0/4294967296.0,1,-nbitq), 
to_sfixed(76735572.0/4294967296.0,1,-nbitq), 
to_sfixed(112135256.0/4294967296.0,1,-nbitq), 
to_sfixed(-513334443.0/4294967296.0,1,-nbitq), 
to_sfixed(-212174501.0/4294967296.0,1,-nbitq), 
to_sfixed(89187050.0/4294967296.0,1,-nbitq), 
to_sfixed(-218453787.0/4294967296.0,1,-nbitq), 
to_sfixed(316809337.0/4294967296.0,1,-nbitq), 
to_sfixed(-193583659.0/4294967296.0,1,-nbitq), 
to_sfixed(504821790.0/4294967296.0,1,-nbitq), 
to_sfixed(-183363081.0/4294967296.0,1,-nbitq), 
to_sfixed(-245525399.0/4294967296.0,1,-nbitq), 
to_sfixed(276488431.0/4294967296.0,1,-nbitq), 
to_sfixed(182627600.0/4294967296.0,1,-nbitq), 
to_sfixed(570851944.0/4294967296.0,1,-nbitq), 
to_sfixed(-863490501.0/4294967296.0,1,-nbitq), 
to_sfixed(-140800724.0/4294967296.0,1,-nbitq), 
to_sfixed(33282531.0/4294967296.0,1,-nbitq), 
to_sfixed(424161506.0/4294967296.0,1,-nbitq), 
to_sfixed(98136584.0/4294967296.0,1,-nbitq), 
to_sfixed(-301172195.0/4294967296.0,1,-nbitq), 
to_sfixed(93570755.0/4294967296.0,1,-nbitq), 
to_sfixed(-324138815.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(129592619.0/4294967296.0,1,-nbitq), 
to_sfixed(-1603941268.0/4294967296.0,1,-nbitq), 
to_sfixed(750658095.0/4294967296.0,1,-nbitq), 
to_sfixed(674051529.0/4294967296.0,1,-nbitq), 
to_sfixed(-165391511.0/4294967296.0,1,-nbitq), 
to_sfixed(-472253465.0/4294967296.0,1,-nbitq), 
to_sfixed(-1112075.0/4294967296.0,1,-nbitq), 
to_sfixed(76772297.0/4294967296.0,1,-nbitq), 
to_sfixed(733217209.0/4294967296.0,1,-nbitq), 
to_sfixed(-302554470.0/4294967296.0,1,-nbitq), 
to_sfixed(-233261639.0/4294967296.0,1,-nbitq), 
to_sfixed(612175933.0/4294967296.0,1,-nbitq), 
to_sfixed(404686769.0/4294967296.0,1,-nbitq), 
to_sfixed(587404421.0/4294967296.0,1,-nbitq), 
to_sfixed(331263231.0/4294967296.0,1,-nbitq), 
to_sfixed(241868797.0/4294967296.0,1,-nbitq), 
to_sfixed(389223577.0/4294967296.0,1,-nbitq), 
to_sfixed(60800457.0/4294967296.0,1,-nbitq), 
to_sfixed(-1714555678.0/4294967296.0,1,-nbitq), 
to_sfixed(-564458956.0/4294967296.0,1,-nbitq), 
to_sfixed(93276384.0/4294967296.0,1,-nbitq), 
to_sfixed(1136652417.0/4294967296.0,1,-nbitq), 
to_sfixed(-668397734.0/4294967296.0,1,-nbitq), 
to_sfixed(1082040186.0/4294967296.0,1,-nbitq), 
to_sfixed(266938811.0/4294967296.0,1,-nbitq), 
to_sfixed(-415314547.0/4294967296.0,1,-nbitq), 
to_sfixed(509870219.0/4294967296.0,1,-nbitq), 
to_sfixed(556280566.0/4294967296.0,1,-nbitq), 
to_sfixed(637866597.0/4294967296.0,1,-nbitq), 
to_sfixed(892710984.0/4294967296.0,1,-nbitq), 
to_sfixed(1441693351.0/4294967296.0,1,-nbitq), 
to_sfixed(428584391.0/4294967296.0,1,-nbitq), 
to_sfixed(-1032212278.0/4294967296.0,1,-nbitq), 
to_sfixed(150660636.0/4294967296.0,1,-nbitq), 
to_sfixed(506142147.0/4294967296.0,1,-nbitq), 
to_sfixed(376407438.0/4294967296.0,1,-nbitq), 
to_sfixed(9878609.0/4294967296.0,1,-nbitq), 
to_sfixed(318106757.0/4294967296.0,1,-nbitq), 
to_sfixed(421329797.0/4294967296.0,1,-nbitq), 
to_sfixed(-126594085.0/4294967296.0,1,-nbitq), 
to_sfixed(279815184.0/4294967296.0,1,-nbitq), 
to_sfixed(-139890198.0/4294967296.0,1,-nbitq), 
to_sfixed(-414568129.0/4294967296.0,1,-nbitq), 
to_sfixed(-400902462.0/4294967296.0,1,-nbitq), 
to_sfixed(-43346057.0/4294967296.0,1,-nbitq), 
to_sfixed(23303717.0/4294967296.0,1,-nbitq), 
to_sfixed(-216558521.0/4294967296.0,1,-nbitq), 
to_sfixed(-310335589.0/4294967296.0,1,-nbitq), 
to_sfixed(-753868442.0/4294967296.0,1,-nbitq), 
to_sfixed(-228321594.0/4294967296.0,1,-nbitq), 
to_sfixed(532411248.0/4294967296.0,1,-nbitq), 
to_sfixed(801292234.0/4294967296.0,1,-nbitq), 
to_sfixed(333606743.0/4294967296.0,1,-nbitq), 
to_sfixed(-524215364.0/4294967296.0,1,-nbitq), 
to_sfixed(-1960275055.0/4294967296.0,1,-nbitq), 
to_sfixed(308249489.0/4294967296.0,1,-nbitq), 
to_sfixed(-99743402.0/4294967296.0,1,-nbitq), 
to_sfixed(247123330.0/4294967296.0,1,-nbitq), 
to_sfixed(90013519.0/4294967296.0,1,-nbitq), 
to_sfixed(-128476151.0/4294967296.0,1,-nbitq), 
to_sfixed(-478633153.0/4294967296.0,1,-nbitq), 
to_sfixed(-368122468.0/4294967296.0,1,-nbitq), 
to_sfixed(-180377654.0/4294967296.0,1,-nbitq), 
to_sfixed(648583495.0/4294967296.0,1,-nbitq), 
to_sfixed(-91227692.0/4294967296.0,1,-nbitq), 
to_sfixed(-77422474.0/4294967296.0,1,-nbitq), 
to_sfixed(549930428.0/4294967296.0,1,-nbitq), 
to_sfixed(-497883210.0/4294967296.0,1,-nbitq), 
to_sfixed(279479828.0/4294967296.0,1,-nbitq), 
to_sfixed(862963969.0/4294967296.0,1,-nbitq), 
to_sfixed(355170369.0/4294967296.0,1,-nbitq), 
to_sfixed(-22765918.0/4294967296.0,1,-nbitq), 
to_sfixed(-153073232.0/4294967296.0,1,-nbitq), 
to_sfixed(-208430682.0/4294967296.0,1,-nbitq), 
to_sfixed(-113681784.0/4294967296.0,1,-nbitq), 
to_sfixed(149624613.0/4294967296.0,1,-nbitq), 
to_sfixed(607564840.0/4294967296.0,1,-nbitq), 
to_sfixed(24807284.0/4294967296.0,1,-nbitq), 
to_sfixed(-28616404.0/4294967296.0,1,-nbitq), 
to_sfixed(59741314.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-401617883.0/4294967296.0,1,-nbitq), 
to_sfixed(-1244876179.0/4294967296.0,1,-nbitq), 
to_sfixed(1241994938.0/4294967296.0,1,-nbitq), 
to_sfixed(265138795.0/4294967296.0,1,-nbitq), 
to_sfixed(-465961599.0/4294967296.0,1,-nbitq), 
to_sfixed(-372876604.0/4294967296.0,1,-nbitq), 
to_sfixed(-66302275.0/4294967296.0,1,-nbitq), 
to_sfixed(985093933.0/4294967296.0,1,-nbitq), 
to_sfixed(335556773.0/4294967296.0,1,-nbitq), 
to_sfixed(-54305959.0/4294967296.0,1,-nbitq), 
to_sfixed(433824369.0/4294967296.0,1,-nbitq), 
to_sfixed(787380206.0/4294967296.0,1,-nbitq), 
to_sfixed(-31936141.0/4294967296.0,1,-nbitq), 
to_sfixed(1220333554.0/4294967296.0,1,-nbitq), 
to_sfixed(312377238.0/4294967296.0,1,-nbitq), 
to_sfixed(462826857.0/4294967296.0,1,-nbitq), 
to_sfixed(224724897.0/4294967296.0,1,-nbitq), 
to_sfixed(-105004186.0/4294967296.0,1,-nbitq), 
to_sfixed(-1280073323.0/4294967296.0,1,-nbitq), 
to_sfixed(-480596166.0/4294967296.0,1,-nbitq), 
to_sfixed(-144295723.0/4294967296.0,1,-nbitq), 
to_sfixed(777581745.0/4294967296.0,1,-nbitq), 
to_sfixed(-287608840.0/4294967296.0,1,-nbitq), 
to_sfixed(524271613.0/4294967296.0,1,-nbitq), 
to_sfixed(35658451.0/4294967296.0,1,-nbitq), 
to_sfixed(-303090534.0/4294967296.0,1,-nbitq), 
to_sfixed(240311297.0/4294967296.0,1,-nbitq), 
to_sfixed(374180368.0/4294967296.0,1,-nbitq), 
to_sfixed(389761946.0/4294967296.0,1,-nbitq), 
to_sfixed(970288812.0/4294967296.0,1,-nbitq), 
to_sfixed(692412791.0/4294967296.0,1,-nbitq), 
to_sfixed(129988625.0/4294967296.0,1,-nbitq), 
to_sfixed(-813799279.0/4294967296.0,1,-nbitq), 
to_sfixed(-174879609.0/4294967296.0,1,-nbitq), 
to_sfixed(-201909899.0/4294967296.0,1,-nbitq), 
to_sfixed(-149121149.0/4294967296.0,1,-nbitq), 
to_sfixed(-215460896.0/4294967296.0,1,-nbitq), 
to_sfixed(418674078.0/4294967296.0,1,-nbitq), 
to_sfixed(-107656034.0/4294967296.0,1,-nbitq), 
to_sfixed(-267828098.0/4294967296.0,1,-nbitq), 
to_sfixed(-103585541.0/4294967296.0,1,-nbitq), 
to_sfixed(-166075678.0/4294967296.0,1,-nbitq), 
to_sfixed(-466227814.0/4294967296.0,1,-nbitq), 
to_sfixed(-430736339.0/4294967296.0,1,-nbitq), 
to_sfixed(379077409.0/4294967296.0,1,-nbitq), 
to_sfixed(158740689.0/4294967296.0,1,-nbitq), 
to_sfixed(-209892182.0/4294967296.0,1,-nbitq), 
to_sfixed(74972298.0/4294967296.0,1,-nbitq), 
to_sfixed(-71844202.0/4294967296.0,1,-nbitq), 
to_sfixed(-691367874.0/4294967296.0,1,-nbitq), 
to_sfixed(474270608.0/4294967296.0,1,-nbitq), 
to_sfixed(973993935.0/4294967296.0,1,-nbitq), 
to_sfixed(527854037.0/4294967296.0,1,-nbitq), 
to_sfixed(-815650644.0/4294967296.0,1,-nbitq), 
to_sfixed(-1459033137.0/4294967296.0,1,-nbitq), 
to_sfixed(689063102.0/4294967296.0,1,-nbitq), 
to_sfixed(-213897141.0/4294967296.0,1,-nbitq), 
to_sfixed(464514410.0/4294967296.0,1,-nbitq), 
to_sfixed(-5883884.0/4294967296.0,1,-nbitq), 
to_sfixed(-32377383.0/4294967296.0,1,-nbitq), 
to_sfixed(135367606.0/4294967296.0,1,-nbitq), 
to_sfixed(-401488323.0/4294967296.0,1,-nbitq), 
to_sfixed(-545291523.0/4294967296.0,1,-nbitq), 
to_sfixed(580297528.0/4294967296.0,1,-nbitq), 
to_sfixed(202374334.0/4294967296.0,1,-nbitq), 
to_sfixed(-80179275.0/4294967296.0,1,-nbitq), 
to_sfixed(550122388.0/4294967296.0,1,-nbitq), 
to_sfixed(-88354362.0/4294967296.0,1,-nbitq), 
to_sfixed(-98125711.0/4294967296.0,1,-nbitq), 
to_sfixed(810796368.0/4294967296.0,1,-nbitq), 
to_sfixed(-420614353.0/4294967296.0,1,-nbitq), 
to_sfixed(134374815.0/4294967296.0,1,-nbitq), 
to_sfixed(-144060523.0/4294967296.0,1,-nbitq), 
to_sfixed(-151502799.0/4294967296.0,1,-nbitq), 
to_sfixed(328639240.0/4294967296.0,1,-nbitq), 
to_sfixed(23251093.0/4294967296.0,1,-nbitq), 
to_sfixed(1201885187.0/4294967296.0,1,-nbitq), 
to_sfixed(195053680.0/4294967296.0,1,-nbitq), 
to_sfixed(-339882660.0/4294967296.0,1,-nbitq), 
to_sfixed(-106020511.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-257187017.0/4294967296.0,1,-nbitq), 
to_sfixed(-1202782538.0/4294967296.0,1,-nbitq), 
to_sfixed(286367419.0/4294967296.0,1,-nbitq), 
to_sfixed(336154895.0/4294967296.0,1,-nbitq), 
to_sfixed(-345273560.0/4294967296.0,1,-nbitq), 
to_sfixed(-48655806.0/4294967296.0,1,-nbitq), 
to_sfixed(350553561.0/4294967296.0,1,-nbitq), 
to_sfixed(899971520.0/4294967296.0,1,-nbitq), 
to_sfixed(62661898.0/4294967296.0,1,-nbitq), 
to_sfixed(259960409.0/4294967296.0,1,-nbitq), 
to_sfixed(110339567.0/4294967296.0,1,-nbitq), 
to_sfixed(759078881.0/4294967296.0,1,-nbitq), 
to_sfixed(-181489447.0/4294967296.0,1,-nbitq), 
to_sfixed(215798814.0/4294967296.0,1,-nbitq), 
to_sfixed(-378205.0/4294967296.0,1,-nbitq), 
to_sfixed(-126324496.0/4294967296.0,1,-nbitq), 
to_sfixed(113947649.0/4294967296.0,1,-nbitq), 
to_sfixed(-370089830.0/4294967296.0,1,-nbitq), 
to_sfixed(-725856141.0/4294967296.0,1,-nbitq), 
to_sfixed(-422762771.0/4294967296.0,1,-nbitq), 
to_sfixed(142582553.0/4294967296.0,1,-nbitq), 
to_sfixed(432137782.0/4294967296.0,1,-nbitq), 
to_sfixed(-302686942.0/4294967296.0,1,-nbitq), 
to_sfixed(-613147549.0/4294967296.0,1,-nbitq), 
to_sfixed(-205724307.0/4294967296.0,1,-nbitq), 
to_sfixed(-315274942.0/4294967296.0,1,-nbitq), 
to_sfixed(-279672543.0/4294967296.0,1,-nbitq), 
to_sfixed(356191718.0/4294967296.0,1,-nbitq), 
to_sfixed(-19498843.0/4294967296.0,1,-nbitq), 
to_sfixed(923441447.0/4294967296.0,1,-nbitq), 
to_sfixed(-8472030.0/4294967296.0,1,-nbitq), 
to_sfixed(-360669437.0/4294967296.0,1,-nbitq), 
to_sfixed(-505071257.0/4294967296.0,1,-nbitq), 
to_sfixed(135656067.0/4294967296.0,1,-nbitq), 
to_sfixed(-68329614.0/4294967296.0,1,-nbitq), 
to_sfixed(352444580.0/4294967296.0,1,-nbitq), 
to_sfixed(-409965526.0/4294967296.0,1,-nbitq), 
to_sfixed(779164759.0/4294967296.0,1,-nbitq), 
to_sfixed(-192818284.0/4294967296.0,1,-nbitq), 
to_sfixed(-173289484.0/4294967296.0,1,-nbitq), 
to_sfixed(-62643787.0/4294967296.0,1,-nbitq), 
to_sfixed(3591919.0/4294967296.0,1,-nbitq), 
to_sfixed(-825295329.0/4294967296.0,1,-nbitq), 
to_sfixed(-627845678.0/4294967296.0,1,-nbitq), 
to_sfixed(750363228.0/4294967296.0,1,-nbitq), 
to_sfixed(-76724666.0/4294967296.0,1,-nbitq), 
to_sfixed(139345578.0/4294967296.0,1,-nbitq), 
to_sfixed(422342605.0/4294967296.0,1,-nbitq), 
to_sfixed(-190160972.0/4294967296.0,1,-nbitq), 
to_sfixed(-636562829.0/4294967296.0,1,-nbitq), 
to_sfixed(133240621.0/4294967296.0,1,-nbitq), 
to_sfixed(754705020.0/4294967296.0,1,-nbitq), 
to_sfixed(256677654.0/4294967296.0,1,-nbitq), 
to_sfixed(-726269817.0/4294967296.0,1,-nbitq), 
to_sfixed(-1280808778.0/4294967296.0,1,-nbitq), 
to_sfixed(405432660.0/4294967296.0,1,-nbitq), 
to_sfixed(374905361.0/4294967296.0,1,-nbitq), 
to_sfixed(249360272.0/4294967296.0,1,-nbitq), 
to_sfixed(-107621396.0/4294967296.0,1,-nbitq), 
to_sfixed(137500841.0/4294967296.0,1,-nbitq), 
to_sfixed(-201923275.0/4294967296.0,1,-nbitq), 
to_sfixed(-364778264.0/4294967296.0,1,-nbitq), 
to_sfixed(358324028.0/4294967296.0,1,-nbitq), 
to_sfixed(385065587.0/4294967296.0,1,-nbitq), 
to_sfixed(-48466758.0/4294967296.0,1,-nbitq), 
to_sfixed(237895989.0/4294967296.0,1,-nbitq), 
to_sfixed(797146853.0/4294967296.0,1,-nbitq), 
to_sfixed(345024936.0/4294967296.0,1,-nbitq), 
to_sfixed(-141870543.0/4294967296.0,1,-nbitq), 
to_sfixed(680397987.0/4294967296.0,1,-nbitq), 
to_sfixed(-412281698.0/4294967296.0,1,-nbitq), 
to_sfixed(324546412.0/4294967296.0,1,-nbitq), 
to_sfixed(384797881.0/4294967296.0,1,-nbitq), 
to_sfixed(399305958.0/4294967296.0,1,-nbitq), 
to_sfixed(-199904552.0/4294967296.0,1,-nbitq), 
to_sfixed(230090708.0/4294967296.0,1,-nbitq), 
to_sfixed(481763065.0/4294967296.0,1,-nbitq), 
to_sfixed(-283542719.0/4294967296.0,1,-nbitq), 
to_sfixed(-145982444.0/4294967296.0,1,-nbitq), 
to_sfixed(254764633.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(286064691.0/4294967296.0,1,-nbitq), 
to_sfixed(-105337703.0/4294967296.0,1,-nbitq), 
to_sfixed(932129495.0/4294967296.0,1,-nbitq), 
to_sfixed(-409364558.0/4294967296.0,1,-nbitq), 
to_sfixed(-161400705.0/4294967296.0,1,-nbitq), 
to_sfixed(-632396437.0/4294967296.0,1,-nbitq), 
to_sfixed(417517771.0/4294967296.0,1,-nbitq), 
to_sfixed(377667011.0/4294967296.0,1,-nbitq), 
to_sfixed(-408149415.0/4294967296.0,1,-nbitq), 
to_sfixed(156379342.0/4294967296.0,1,-nbitq), 
to_sfixed(357254133.0/4294967296.0,1,-nbitq), 
to_sfixed(-19187303.0/4294967296.0,1,-nbitq), 
to_sfixed(423895248.0/4294967296.0,1,-nbitq), 
to_sfixed(685231526.0/4294967296.0,1,-nbitq), 
to_sfixed(-209843475.0/4294967296.0,1,-nbitq), 
to_sfixed(450474290.0/4294967296.0,1,-nbitq), 
to_sfixed(199658713.0/4294967296.0,1,-nbitq), 
to_sfixed(-397710605.0/4294967296.0,1,-nbitq), 
to_sfixed(332855810.0/4294967296.0,1,-nbitq), 
to_sfixed(211603194.0/4294967296.0,1,-nbitq), 
to_sfixed(-318511305.0/4294967296.0,1,-nbitq), 
to_sfixed(716806.0/4294967296.0,1,-nbitq), 
to_sfixed(-331893712.0/4294967296.0,1,-nbitq), 
to_sfixed(605429129.0/4294967296.0,1,-nbitq), 
to_sfixed(-5001997.0/4294967296.0,1,-nbitq), 
to_sfixed(-650896664.0/4294967296.0,1,-nbitq), 
to_sfixed(-317185021.0/4294967296.0,1,-nbitq), 
to_sfixed(315591291.0/4294967296.0,1,-nbitq), 
to_sfixed(121050734.0/4294967296.0,1,-nbitq), 
to_sfixed(989254312.0/4294967296.0,1,-nbitq), 
to_sfixed(72482915.0/4294967296.0,1,-nbitq), 
to_sfixed(307562323.0/4294967296.0,1,-nbitq), 
to_sfixed(6793269.0/4294967296.0,1,-nbitq), 
to_sfixed(-454649008.0/4294967296.0,1,-nbitq), 
to_sfixed(-679575455.0/4294967296.0,1,-nbitq), 
to_sfixed(-170291634.0/4294967296.0,1,-nbitq), 
to_sfixed(124821757.0/4294967296.0,1,-nbitq), 
to_sfixed(-247851242.0/4294967296.0,1,-nbitq), 
to_sfixed(-214073747.0/4294967296.0,1,-nbitq), 
to_sfixed(483831227.0/4294967296.0,1,-nbitq), 
to_sfixed(134605787.0/4294967296.0,1,-nbitq), 
to_sfixed(-319699765.0/4294967296.0,1,-nbitq), 
to_sfixed(-35473694.0/4294967296.0,1,-nbitq), 
to_sfixed(-673601917.0/4294967296.0,1,-nbitq), 
to_sfixed(476227984.0/4294967296.0,1,-nbitq), 
to_sfixed(-687736213.0/4294967296.0,1,-nbitq), 
to_sfixed(-358059042.0/4294967296.0,1,-nbitq), 
to_sfixed(-10455716.0/4294967296.0,1,-nbitq), 
to_sfixed(-104894575.0/4294967296.0,1,-nbitq), 
to_sfixed(-459693863.0/4294967296.0,1,-nbitq), 
to_sfixed(-90306552.0/4294967296.0,1,-nbitq), 
to_sfixed(-199119595.0/4294967296.0,1,-nbitq), 
to_sfixed(79265695.0/4294967296.0,1,-nbitq), 
to_sfixed(125918955.0/4294967296.0,1,-nbitq), 
to_sfixed(-165305163.0/4294967296.0,1,-nbitq), 
to_sfixed(-210548474.0/4294967296.0,1,-nbitq), 
to_sfixed(-197952191.0/4294967296.0,1,-nbitq), 
to_sfixed(-24506584.0/4294967296.0,1,-nbitq), 
to_sfixed(-259315794.0/4294967296.0,1,-nbitq), 
to_sfixed(294574839.0/4294967296.0,1,-nbitq), 
to_sfixed(116322188.0/4294967296.0,1,-nbitq), 
to_sfixed(-328086878.0/4294967296.0,1,-nbitq), 
to_sfixed(3852545.0/4294967296.0,1,-nbitq), 
to_sfixed(405811045.0/4294967296.0,1,-nbitq), 
to_sfixed(-395386335.0/4294967296.0,1,-nbitq), 
to_sfixed(-199664638.0/4294967296.0,1,-nbitq), 
to_sfixed(252283061.0/4294967296.0,1,-nbitq), 
to_sfixed(-263382158.0/4294967296.0,1,-nbitq), 
to_sfixed(161596857.0/4294967296.0,1,-nbitq), 
to_sfixed(782850109.0/4294967296.0,1,-nbitq), 
to_sfixed(-498271965.0/4294967296.0,1,-nbitq), 
to_sfixed(-183259480.0/4294967296.0,1,-nbitq), 
to_sfixed(472088192.0/4294967296.0,1,-nbitq), 
to_sfixed(-33620968.0/4294967296.0,1,-nbitq), 
to_sfixed(46214097.0/4294967296.0,1,-nbitq), 
to_sfixed(-243737247.0/4294967296.0,1,-nbitq), 
to_sfixed(-186281234.0/4294967296.0,1,-nbitq), 
to_sfixed(252096191.0/4294967296.0,1,-nbitq), 
to_sfixed(98144006.0/4294967296.0,1,-nbitq), 
to_sfixed(-262067160.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-144526940.0/4294967296.0,1,-nbitq), 
to_sfixed(191423263.0/4294967296.0,1,-nbitq), 
to_sfixed(422260336.0/4294967296.0,1,-nbitq), 
to_sfixed(8906772.0/4294967296.0,1,-nbitq), 
to_sfixed(-56224919.0/4294967296.0,1,-nbitq), 
to_sfixed(-474112242.0/4294967296.0,1,-nbitq), 
to_sfixed(-166444569.0/4294967296.0,1,-nbitq), 
to_sfixed(170149007.0/4294967296.0,1,-nbitq), 
to_sfixed(-544874725.0/4294967296.0,1,-nbitq), 
to_sfixed(-26790618.0/4294967296.0,1,-nbitq), 
to_sfixed(201179294.0/4294967296.0,1,-nbitq), 
to_sfixed(148423487.0/4294967296.0,1,-nbitq), 
to_sfixed(257430299.0/4294967296.0,1,-nbitq), 
to_sfixed(434519731.0/4294967296.0,1,-nbitq), 
to_sfixed(-152083513.0/4294967296.0,1,-nbitq), 
to_sfixed(-312241856.0/4294967296.0,1,-nbitq), 
to_sfixed(72415049.0/4294967296.0,1,-nbitq), 
to_sfixed(-57799608.0/4294967296.0,1,-nbitq), 
to_sfixed(460118799.0/4294967296.0,1,-nbitq), 
to_sfixed(355411020.0/4294967296.0,1,-nbitq), 
to_sfixed(-78014140.0/4294967296.0,1,-nbitq), 
to_sfixed(-448265124.0/4294967296.0,1,-nbitq), 
to_sfixed(-178469948.0/4294967296.0,1,-nbitq), 
to_sfixed(154144481.0/4294967296.0,1,-nbitq), 
to_sfixed(-161864857.0/4294967296.0,1,-nbitq), 
to_sfixed(-382690053.0/4294967296.0,1,-nbitq), 
to_sfixed(435078322.0/4294967296.0,1,-nbitq), 
to_sfixed(-30876294.0/4294967296.0,1,-nbitq), 
to_sfixed(490770669.0/4294967296.0,1,-nbitq), 
to_sfixed(601790301.0/4294967296.0,1,-nbitq), 
to_sfixed(-143196862.0/4294967296.0,1,-nbitq), 
to_sfixed(49637500.0/4294967296.0,1,-nbitq), 
to_sfixed(357512721.0/4294967296.0,1,-nbitq), 
to_sfixed(82167432.0/4294967296.0,1,-nbitq), 
to_sfixed(-207492590.0/4294967296.0,1,-nbitq), 
to_sfixed(-210244057.0/4294967296.0,1,-nbitq), 
to_sfixed(-234599135.0/4294967296.0,1,-nbitq), 
to_sfixed(53751674.0/4294967296.0,1,-nbitq), 
to_sfixed(68425470.0/4294967296.0,1,-nbitq), 
to_sfixed(394746039.0/4294967296.0,1,-nbitq), 
to_sfixed(-75061276.0/4294967296.0,1,-nbitq), 
to_sfixed(-18734641.0/4294967296.0,1,-nbitq), 
to_sfixed(-420024685.0/4294967296.0,1,-nbitq), 
to_sfixed(-316185789.0/4294967296.0,1,-nbitq), 
to_sfixed(-211842111.0/4294967296.0,1,-nbitq), 
to_sfixed(-546905329.0/4294967296.0,1,-nbitq), 
to_sfixed(-148308886.0/4294967296.0,1,-nbitq), 
to_sfixed(-70054761.0/4294967296.0,1,-nbitq), 
to_sfixed(178749133.0/4294967296.0,1,-nbitq), 
to_sfixed(-162552887.0/4294967296.0,1,-nbitq), 
to_sfixed(-201397797.0/4294967296.0,1,-nbitq), 
to_sfixed(451551313.0/4294967296.0,1,-nbitq), 
to_sfixed(-85730003.0/4294967296.0,1,-nbitq), 
to_sfixed(-313576808.0/4294967296.0,1,-nbitq), 
to_sfixed(43961302.0/4294967296.0,1,-nbitq), 
to_sfixed(-402127043.0/4294967296.0,1,-nbitq), 
to_sfixed(-201356451.0/4294967296.0,1,-nbitq), 
to_sfixed(485143253.0/4294967296.0,1,-nbitq), 
to_sfixed(-69183941.0/4294967296.0,1,-nbitq), 
to_sfixed(-268612091.0/4294967296.0,1,-nbitq), 
to_sfixed(-181531219.0/4294967296.0,1,-nbitq), 
to_sfixed(310085478.0/4294967296.0,1,-nbitq), 
to_sfixed(389528853.0/4294967296.0,1,-nbitq), 
to_sfixed(290099727.0/4294967296.0,1,-nbitq), 
to_sfixed(272922328.0/4294967296.0,1,-nbitq), 
to_sfixed(53718378.0/4294967296.0,1,-nbitq), 
to_sfixed(690520711.0/4294967296.0,1,-nbitq), 
to_sfixed(-390366550.0/4294967296.0,1,-nbitq), 
to_sfixed(-287311319.0/4294967296.0,1,-nbitq), 
to_sfixed(337822061.0/4294967296.0,1,-nbitq), 
to_sfixed(-278026894.0/4294967296.0,1,-nbitq), 
to_sfixed(346991484.0/4294967296.0,1,-nbitq), 
to_sfixed(182221803.0/4294967296.0,1,-nbitq), 
to_sfixed(25966771.0/4294967296.0,1,-nbitq), 
to_sfixed(-90871580.0/4294967296.0,1,-nbitq), 
to_sfixed(-405249949.0/4294967296.0,1,-nbitq), 
to_sfixed(-567860353.0/4294967296.0,1,-nbitq), 
to_sfixed(157097121.0/4294967296.0,1,-nbitq), 
to_sfixed(-316028555.0/4294967296.0,1,-nbitq), 
to_sfixed(87122464.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-275521127.0/4294967296.0,1,-nbitq), 
to_sfixed(-513519474.0/4294967296.0,1,-nbitq), 
to_sfixed(508548698.0/4294967296.0,1,-nbitq), 
to_sfixed(185508371.0/4294967296.0,1,-nbitq), 
to_sfixed(168967397.0/4294967296.0,1,-nbitq), 
to_sfixed(-312587720.0/4294967296.0,1,-nbitq), 
to_sfixed(259200530.0/4294967296.0,1,-nbitq), 
to_sfixed(325801136.0/4294967296.0,1,-nbitq), 
to_sfixed(173821825.0/4294967296.0,1,-nbitq), 
to_sfixed(-257601610.0/4294967296.0,1,-nbitq), 
to_sfixed(220348396.0/4294967296.0,1,-nbitq), 
to_sfixed(63613506.0/4294967296.0,1,-nbitq), 
to_sfixed(-275013908.0/4294967296.0,1,-nbitq), 
to_sfixed(247543426.0/4294967296.0,1,-nbitq), 
to_sfixed(121766174.0/4294967296.0,1,-nbitq), 
to_sfixed(-33677190.0/4294967296.0,1,-nbitq), 
to_sfixed(-184373286.0/4294967296.0,1,-nbitq), 
to_sfixed(-412914817.0/4294967296.0,1,-nbitq), 
to_sfixed(120945553.0/4294967296.0,1,-nbitq), 
to_sfixed(-98240145.0/4294967296.0,1,-nbitq), 
to_sfixed(-375364727.0/4294967296.0,1,-nbitq), 
to_sfixed(119415631.0/4294967296.0,1,-nbitq), 
to_sfixed(214199513.0/4294967296.0,1,-nbitq), 
to_sfixed(185535143.0/4294967296.0,1,-nbitq), 
to_sfixed(226805392.0/4294967296.0,1,-nbitq), 
to_sfixed(-438409240.0/4294967296.0,1,-nbitq), 
to_sfixed(-204848763.0/4294967296.0,1,-nbitq), 
to_sfixed(-321458018.0/4294967296.0,1,-nbitq), 
to_sfixed(-154816758.0/4294967296.0,1,-nbitq), 
to_sfixed(-224557860.0/4294967296.0,1,-nbitq), 
to_sfixed(81941969.0/4294967296.0,1,-nbitq), 
to_sfixed(-160771965.0/4294967296.0,1,-nbitq), 
to_sfixed(-219206252.0/4294967296.0,1,-nbitq), 
to_sfixed(-321598113.0/4294967296.0,1,-nbitq), 
to_sfixed(-277828634.0/4294967296.0,1,-nbitq), 
to_sfixed(-483077843.0/4294967296.0,1,-nbitq), 
to_sfixed(268728054.0/4294967296.0,1,-nbitq), 
to_sfixed(-259739329.0/4294967296.0,1,-nbitq), 
to_sfixed(-225535785.0/4294967296.0,1,-nbitq), 
to_sfixed(-286188837.0/4294967296.0,1,-nbitq), 
to_sfixed(-418231629.0/4294967296.0,1,-nbitq), 
to_sfixed(105099703.0/4294967296.0,1,-nbitq), 
to_sfixed(10917872.0/4294967296.0,1,-nbitq), 
to_sfixed(-336823424.0/4294967296.0,1,-nbitq), 
to_sfixed(-172232784.0/4294967296.0,1,-nbitq), 
to_sfixed(-138894730.0/4294967296.0,1,-nbitq), 
to_sfixed(-186639605.0/4294967296.0,1,-nbitq), 
to_sfixed(-316987594.0/4294967296.0,1,-nbitq), 
to_sfixed(277128001.0/4294967296.0,1,-nbitq), 
to_sfixed(78787834.0/4294967296.0,1,-nbitq), 
to_sfixed(-219115538.0/4294967296.0,1,-nbitq), 
to_sfixed(-176273365.0/4294967296.0,1,-nbitq), 
to_sfixed(282743057.0/4294967296.0,1,-nbitq), 
to_sfixed(-155189790.0/4294967296.0,1,-nbitq), 
to_sfixed(-83362602.0/4294967296.0,1,-nbitq), 
to_sfixed(-154475975.0/4294967296.0,1,-nbitq), 
to_sfixed(233052282.0/4294967296.0,1,-nbitq), 
to_sfixed(-340883651.0/4294967296.0,1,-nbitq), 
to_sfixed(-133416039.0/4294967296.0,1,-nbitq), 
to_sfixed(-93321698.0/4294967296.0,1,-nbitq), 
to_sfixed(316522878.0/4294967296.0,1,-nbitq), 
to_sfixed(280385744.0/4294967296.0,1,-nbitq), 
to_sfixed(2366677.0/4294967296.0,1,-nbitq), 
to_sfixed(-298479912.0/4294967296.0,1,-nbitq), 
to_sfixed(262313305.0/4294967296.0,1,-nbitq), 
to_sfixed(-389562522.0/4294967296.0,1,-nbitq), 
to_sfixed(175654551.0/4294967296.0,1,-nbitq), 
to_sfixed(-168451309.0/4294967296.0,1,-nbitq), 
to_sfixed(170242963.0/4294967296.0,1,-nbitq), 
to_sfixed(226068441.0/4294967296.0,1,-nbitq), 
to_sfixed(-26064190.0/4294967296.0,1,-nbitq), 
to_sfixed(-312703012.0/4294967296.0,1,-nbitq), 
to_sfixed(-134118231.0/4294967296.0,1,-nbitq), 
to_sfixed(-250097062.0/4294967296.0,1,-nbitq), 
to_sfixed(27489034.0/4294967296.0,1,-nbitq), 
to_sfixed(167867527.0/4294967296.0,1,-nbitq), 
to_sfixed(41504294.0/4294967296.0,1,-nbitq), 
to_sfixed(4874714.0/4294967296.0,1,-nbitq), 
to_sfixed(-185251050.0/4294967296.0,1,-nbitq), 
to_sfixed(-155108874.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(109989815.0/4294967296.0,1,-nbitq), 
to_sfixed(110415942.0/4294967296.0,1,-nbitq), 
to_sfixed(-197651279.0/4294967296.0,1,-nbitq), 
to_sfixed(-95265948.0/4294967296.0,1,-nbitq), 
to_sfixed(260904056.0/4294967296.0,1,-nbitq), 
to_sfixed(231597592.0/4294967296.0,1,-nbitq), 
to_sfixed(-322325077.0/4294967296.0,1,-nbitq), 
to_sfixed(255611369.0/4294967296.0,1,-nbitq), 
to_sfixed(-346930612.0/4294967296.0,1,-nbitq), 
to_sfixed(-102123588.0/4294967296.0,1,-nbitq), 
to_sfixed(-401051629.0/4294967296.0,1,-nbitq), 
to_sfixed(15941594.0/4294967296.0,1,-nbitq), 
to_sfixed(79693080.0/4294967296.0,1,-nbitq), 
to_sfixed(-68159589.0/4294967296.0,1,-nbitq), 
to_sfixed(77939386.0/4294967296.0,1,-nbitq), 
to_sfixed(-88071159.0/4294967296.0,1,-nbitq), 
to_sfixed(-4953821.0/4294967296.0,1,-nbitq), 
to_sfixed(105241206.0/4294967296.0,1,-nbitq), 
to_sfixed(297492711.0/4294967296.0,1,-nbitq), 
to_sfixed(-356858335.0/4294967296.0,1,-nbitq), 
to_sfixed(-237955527.0/4294967296.0,1,-nbitq), 
to_sfixed(-28707995.0/4294967296.0,1,-nbitq), 
to_sfixed(374413629.0/4294967296.0,1,-nbitq), 
to_sfixed(-337196307.0/4294967296.0,1,-nbitq), 
to_sfixed(-314207361.0/4294967296.0,1,-nbitq), 
to_sfixed(-30948261.0/4294967296.0,1,-nbitq), 
to_sfixed(-330388660.0/4294967296.0,1,-nbitq), 
to_sfixed(-537171091.0/4294967296.0,1,-nbitq), 
to_sfixed(11174101.0/4294967296.0,1,-nbitq), 
to_sfixed(-18948659.0/4294967296.0,1,-nbitq), 
to_sfixed(-319078547.0/4294967296.0,1,-nbitq), 
to_sfixed(-245103652.0/4294967296.0,1,-nbitq), 
to_sfixed(-42566066.0/4294967296.0,1,-nbitq), 
to_sfixed(-142935768.0/4294967296.0,1,-nbitq), 
to_sfixed(67332955.0/4294967296.0,1,-nbitq), 
to_sfixed(21281806.0/4294967296.0,1,-nbitq), 
to_sfixed(-269142894.0/4294967296.0,1,-nbitq), 
to_sfixed(425914743.0/4294967296.0,1,-nbitq), 
to_sfixed(-85457013.0/4294967296.0,1,-nbitq), 
to_sfixed(339237432.0/4294967296.0,1,-nbitq), 
to_sfixed(41359062.0/4294967296.0,1,-nbitq), 
to_sfixed(-131500195.0/4294967296.0,1,-nbitq), 
to_sfixed(-342010827.0/4294967296.0,1,-nbitq), 
to_sfixed(-370030269.0/4294967296.0,1,-nbitq), 
to_sfixed(-75285188.0/4294967296.0,1,-nbitq), 
to_sfixed(360399949.0/4294967296.0,1,-nbitq), 
to_sfixed(-390247625.0/4294967296.0,1,-nbitq), 
to_sfixed(247188968.0/4294967296.0,1,-nbitq), 
to_sfixed(-187502352.0/4294967296.0,1,-nbitq), 
to_sfixed(336977518.0/4294967296.0,1,-nbitq), 
to_sfixed(76158371.0/4294967296.0,1,-nbitq), 
to_sfixed(312803335.0/4294967296.0,1,-nbitq), 
to_sfixed(-228074684.0/4294967296.0,1,-nbitq), 
to_sfixed(211532889.0/4294967296.0,1,-nbitq), 
to_sfixed(-244356472.0/4294967296.0,1,-nbitq), 
to_sfixed(-91282101.0/4294967296.0,1,-nbitq), 
to_sfixed(-246738666.0/4294967296.0,1,-nbitq), 
to_sfixed(-5189038.0/4294967296.0,1,-nbitq), 
to_sfixed(-81140897.0/4294967296.0,1,-nbitq), 
to_sfixed(-332502886.0/4294967296.0,1,-nbitq), 
to_sfixed(-7269825.0/4294967296.0,1,-nbitq), 
to_sfixed(382405638.0/4294967296.0,1,-nbitq), 
to_sfixed(-353293783.0/4294967296.0,1,-nbitq), 
to_sfixed(-83100239.0/4294967296.0,1,-nbitq), 
to_sfixed(-362798407.0/4294967296.0,1,-nbitq), 
to_sfixed(-321990547.0/4294967296.0,1,-nbitq), 
to_sfixed(184441609.0/4294967296.0,1,-nbitq), 
to_sfixed(-62126249.0/4294967296.0,1,-nbitq), 
to_sfixed(207423802.0/4294967296.0,1,-nbitq), 
to_sfixed(80616400.0/4294967296.0,1,-nbitq), 
to_sfixed(-89495144.0/4294967296.0,1,-nbitq), 
to_sfixed(-172346199.0/4294967296.0,1,-nbitq), 
to_sfixed(232587757.0/4294967296.0,1,-nbitq), 
to_sfixed(437808578.0/4294967296.0,1,-nbitq), 
to_sfixed(-128985958.0/4294967296.0,1,-nbitq), 
to_sfixed(-168978817.0/4294967296.0,1,-nbitq), 
to_sfixed(-222372021.0/4294967296.0,1,-nbitq), 
to_sfixed(251769205.0/4294967296.0,1,-nbitq), 
to_sfixed(-98766786.0/4294967296.0,1,-nbitq), 
to_sfixed(-310763439.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-275137881.0/4294967296.0,1,-nbitq), 
to_sfixed(-294885217.0/4294967296.0,1,-nbitq), 
to_sfixed(359364387.0/4294967296.0,1,-nbitq), 
to_sfixed(-252612530.0/4294967296.0,1,-nbitq), 
to_sfixed(-10154934.0/4294967296.0,1,-nbitq), 
to_sfixed(-90891465.0/4294967296.0,1,-nbitq), 
to_sfixed(-213045146.0/4294967296.0,1,-nbitq), 
to_sfixed(-354024157.0/4294967296.0,1,-nbitq), 
to_sfixed(161191921.0/4294967296.0,1,-nbitq), 
to_sfixed(316324162.0/4294967296.0,1,-nbitq), 
to_sfixed(367469424.0/4294967296.0,1,-nbitq), 
to_sfixed(-5196263.0/4294967296.0,1,-nbitq), 
to_sfixed(-35007451.0/4294967296.0,1,-nbitq), 
to_sfixed(-333198444.0/4294967296.0,1,-nbitq), 
to_sfixed(145389909.0/4294967296.0,1,-nbitq), 
to_sfixed(-3396591.0/4294967296.0,1,-nbitq), 
to_sfixed(-297331875.0/4294967296.0,1,-nbitq), 
to_sfixed(308214526.0/4294967296.0,1,-nbitq), 
to_sfixed(-39299063.0/4294967296.0,1,-nbitq), 
to_sfixed(-193501772.0/4294967296.0,1,-nbitq), 
to_sfixed(-18371800.0/4294967296.0,1,-nbitq), 
to_sfixed(163911557.0/4294967296.0,1,-nbitq), 
to_sfixed(320015749.0/4294967296.0,1,-nbitq), 
to_sfixed(-306357887.0/4294967296.0,1,-nbitq), 
to_sfixed(-310159291.0/4294967296.0,1,-nbitq), 
to_sfixed(-227860711.0/4294967296.0,1,-nbitq), 
to_sfixed(-232284553.0/4294967296.0,1,-nbitq), 
to_sfixed(31470100.0/4294967296.0,1,-nbitq), 
to_sfixed(-282365398.0/4294967296.0,1,-nbitq), 
to_sfixed(339949617.0/4294967296.0,1,-nbitq), 
to_sfixed(-624610909.0/4294967296.0,1,-nbitq), 
to_sfixed(126319146.0/4294967296.0,1,-nbitq), 
to_sfixed(231639568.0/4294967296.0,1,-nbitq), 
to_sfixed(237255773.0/4294967296.0,1,-nbitq), 
to_sfixed(12841947.0/4294967296.0,1,-nbitq), 
to_sfixed(-43865015.0/4294967296.0,1,-nbitq), 
to_sfixed(114095648.0/4294967296.0,1,-nbitq), 
to_sfixed(-311572313.0/4294967296.0,1,-nbitq), 
to_sfixed(368714113.0/4294967296.0,1,-nbitq), 
to_sfixed(81227501.0/4294967296.0,1,-nbitq), 
to_sfixed(-281907149.0/4294967296.0,1,-nbitq), 
to_sfixed(152141681.0/4294967296.0,1,-nbitq), 
to_sfixed(-327214596.0/4294967296.0,1,-nbitq), 
to_sfixed(186440087.0/4294967296.0,1,-nbitq), 
to_sfixed(-141902352.0/4294967296.0,1,-nbitq), 
to_sfixed(66269880.0/4294967296.0,1,-nbitq), 
to_sfixed(-275370229.0/4294967296.0,1,-nbitq), 
to_sfixed(-64779787.0/4294967296.0,1,-nbitq), 
to_sfixed(-56780460.0/4294967296.0,1,-nbitq), 
to_sfixed(177992727.0/4294967296.0,1,-nbitq), 
to_sfixed(36373824.0/4294967296.0,1,-nbitq), 
to_sfixed(449812526.0/4294967296.0,1,-nbitq), 
to_sfixed(89896422.0/4294967296.0,1,-nbitq), 
to_sfixed(-248480790.0/4294967296.0,1,-nbitq), 
to_sfixed(-18493831.0/4294967296.0,1,-nbitq), 
to_sfixed(112885876.0/4294967296.0,1,-nbitq), 
to_sfixed(68903337.0/4294967296.0,1,-nbitq), 
to_sfixed(-477069814.0/4294967296.0,1,-nbitq), 
to_sfixed(-171092942.0/4294967296.0,1,-nbitq), 
to_sfixed(-29194432.0/4294967296.0,1,-nbitq), 
to_sfixed(174865075.0/4294967296.0,1,-nbitq), 
to_sfixed(-122987697.0/4294967296.0,1,-nbitq), 
to_sfixed(-439917213.0/4294967296.0,1,-nbitq), 
to_sfixed(-12547841.0/4294967296.0,1,-nbitq), 
to_sfixed(-236492515.0/4294967296.0,1,-nbitq), 
to_sfixed(153820808.0/4294967296.0,1,-nbitq), 
to_sfixed(498101655.0/4294967296.0,1,-nbitq), 
to_sfixed(-7484341.0/4294967296.0,1,-nbitq), 
to_sfixed(366206024.0/4294967296.0,1,-nbitq), 
to_sfixed(533689393.0/4294967296.0,1,-nbitq), 
to_sfixed(-104100365.0/4294967296.0,1,-nbitq), 
to_sfixed(-82399808.0/4294967296.0,1,-nbitq), 
to_sfixed(-198425791.0/4294967296.0,1,-nbitq), 
to_sfixed(-293585757.0/4294967296.0,1,-nbitq), 
to_sfixed(306584889.0/4294967296.0,1,-nbitq), 
to_sfixed(-360945571.0/4294967296.0,1,-nbitq), 
to_sfixed(-316945591.0/4294967296.0,1,-nbitq), 
to_sfixed(-437303925.0/4294967296.0,1,-nbitq), 
to_sfixed(-275147486.0/4294967296.0,1,-nbitq), 
to_sfixed(63710037.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(39528595.0/4294967296.0,1,-nbitq), 
to_sfixed(-62117173.0/4294967296.0,1,-nbitq), 
to_sfixed(732554392.0/4294967296.0,1,-nbitq), 
to_sfixed(-280836078.0/4294967296.0,1,-nbitq), 
to_sfixed(-246448176.0/4294967296.0,1,-nbitq), 
to_sfixed(-181215561.0/4294967296.0,1,-nbitq), 
to_sfixed(331458601.0/4294967296.0,1,-nbitq), 
to_sfixed(-187010047.0/4294967296.0,1,-nbitq), 
to_sfixed(-271820716.0/4294967296.0,1,-nbitq), 
to_sfixed(-114041050.0/4294967296.0,1,-nbitq), 
to_sfixed(133026588.0/4294967296.0,1,-nbitq), 
to_sfixed(-285120645.0/4294967296.0,1,-nbitq), 
to_sfixed(-337929305.0/4294967296.0,1,-nbitq), 
to_sfixed(-263404650.0/4294967296.0,1,-nbitq), 
to_sfixed(67202704.0/4294967296.0,1,-nbitq), 
to_sfixed(370022136.0/4294967296.0,1,-nbitq), 
to_sfixed(67396700.0/4294967296.0,1,-nbitq), 
to_sfixed(-82432467.0/4294967296.0,1,-nbitq), 
to_sfixed(-714740504.0/4294967296.0,1,-nbitq), 
to_sfixed(423503016.0/4294967296.0,1,-nbitq), 
to_sfixed(-184385816.0/4294967296.0,1,-nbitq), 
to_sfixed(-96538143.0/4294967296.0,1,-nbitq), 
to_sfixed(-178438261.0/4294967296.0,1,-nbitq), 
to_sfixed(223101513.0/4294967296.0,1,-nbitq), 
to_sfixed(-95557356.0/4294967296.0,1,-nbitq), 
to_sfixed(147133541.0/4294967296.0,1,-nbitq), 
to_sfixed(95571593.0/4294967296.0,1,-nbitq), 
to_sfixed(-309299767.0/4294967296.0,1,-nbitq), 
to_sfixed(-224455048.0/4294967296.0,1,-nbitq), 
to_sfixed(448874225.0/4294967296.0,1,-nbitq), 
to_sfixed(55773905.0/4294967296.0,1,-nbitq), 
to_sfixed(-316122023.0/4294967296.0,1,-nbitq), 
to_sfixed(-95551228.0/4294967296.0,1,-nbitq), 
to_sfixed(-51712488.0/4294967296.0,1,-nbitq), 
to_sfixed(-279767991.0/4294967296.0,1,-nbitq), 
to_sfixed(-112790487.0/4294967296.0,1,-nbitq), 
to_sfixed(351455416.0/4294967296.0,1,-nbitq), 
to_sfixed(385270442.0/4294967296.0,1,-nbitq), 
to_sfixed(-218308636.0/4294967296.0,1,-nbitq), 
to_sfixed(-171308534.0/4294967296.0,1,-nbitq), 
to_sfixed(198474090.0/4294967296.0,1,-nbitq), 
to_sfixed(-114448129.0/4294967296.0,1,-nbitq), 
to_sfixed(-101499742.0/4294967296.0,1,-nbitq), 
to_sfixed(153217609.0/4294967296.0,1,-nbitq), 
to_sfixed(-420120827.0/4294967296.0,1,-nbitq), 
to_sfixed(-81872106.0/4294967296.0,1,-nbitq), 
to_sfixed(137130307.0/4294967296.0,1,-nbitq), 
to_sfixed(-21608897.0/4294967296.0,1,-nbitq), 
to_sfixed(-177630770.0/4294967296.0,1,-nbitq), 
to_sfixed(-297034572.0/4294967296.0,1,-nbitq), 
to_sfixed(-371580454.0/4294967296.0,1,-nbitq), 
to_sfixed(-293983686.0/4294967296.0,1,-nbitq), 
to_sfixed(-189068999.0/4294967296.0,1,-nbitq), 
to_sfixed(-198075168.0/4294967296.0,1,-nbitq), 
to_sfixed(-192269304.0/4294967296.0,1,-nbitq), 
to_sfixed(-104830286.0/4294967296.0,1,-nbitq), 
to_sfixed(-159404828.0/4294967296.0,1,-nbitq), 
to_sfixed(117168988.0/4294967296.0,1,-nbitq), 
to_sfixed(-176533282.0/4294967296.0,1,-nbitq), 
to_sfixed(-132722813.0/4294967296.0,1,-nbitq), 
to_sfixed(-27405730.0/4294967296.0,1,-nbitq), 
to_sfixed(383572308.0/4294967296.0,1,-nbitq), 
to_sfixed(-177406826.0/4294967296.0,1,-nbitq), 
to_sfixed(-297082497.0/4294967296.0,1,-nbitq), 
to_sfixed(-59870800.0/4294967296.0,1,-nbitq), 
to_sfixed(-181744948.0/4294967296.0,1,-nbitq), 
to_sfixed(532798266.0/4294967296.0,1,-nbitq), 
to_sfixed(-230245887.0/4294967296.0,1,-nbitq), 
to_sfixed(368128908.0/4294967296.0,1,-nbitq), 
to_sfixed(383620246.0/4294967296.0,1,-nbitq), 
to_sfixed(-117016811.0/4294967296.0,1,-nbitq), 
to_sfixed(326980599.0/4294967296.0,1,-nbitq), 
to_sfixed(193406716.0/4294967296.0,1,-nbitq), 
to_sfixed(274481812.0/4294967296.0,1,-nbitq), 
to_sfixed(340863890.0/4294967296.0,1,-nbitq), 
to_sfixed(185537909.0/4294967296.0,1,-nbitq), 
to_sfixed(-72736452.0/4294967296.0,1,-nbitq), 
to_sfixed(69519292.0/4294967296.0,1,-nbitq), 
to_sfixed(104776638.0/4294967296.0,1,-nbitq), 
to_sfixed(301995715.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-337185294.0/4294967296.0,1,-nbitq), 
to_sfixed(76121479.0/4294967296.0,1,-nbitq), 
to_sfixed(168270440.0/4294967296.0,1,-nbitq), 
to_sfixed(-147974925.0/4294967296.0,1,-nbitq), 
to_sfixed(291766827.0/4294967296.0,1,-nbitq), 
to_sfixed(325903345.0/4294967296.0,1,-nbitq), 
to_sfixed(-178966695.0/4294967296.0,1,-nbitq), 
to_sfixed(128769576.0/4294967296.0,1,-nbitq), 
to_sfixed(-407505669.0/4294967296.0,1,-nbitq), 
to_sfixed(-107534235.0/4294967296.0,1,-nbitq), 
to_sfixed(148222906.0/4294967296.0,1,-nbitq), 
to_sfixed(-389155145.0/4294967296.0,1,-nbitq), 
to_sfixed(-307220982.0/4294967296.0,1,-nbitq), 
to_sfixed(250167358.0/4294967296.0,1,-nbitq), 
to_sfixed(-388916971.0/4294967296.0,1,-nbitq), 
to_sfixed(479686792.0/4294967296.0,1,-nbitq), 
to_sfixed(-285303360.0/4294967296.0,1,-nbitq), 
to_sfixed(69896029.0/4294967296.0,1,-nbitq), 
to_sfixed(-533708077.0/4294967296.0,1,-nbitq), 
to_sfixed(443599810.0/4294967296.0,1,-nbitq), 
to_sfixed(-111497510.0/4294967296.0,1,-nbitq), 
to_sfixed(195478612.0/4294967296.0,1,-nbitq), 
to_sfixed(-603185145.0/4294967296.0,1,-nbitq), 
to_sfixed(471070436.0/4294967296.0,1,-nbitq), 
to_sfixed(402608997.0/4294967296.0,1,-nbitq), 
to_sfixed(24092239.0/4294967296.0,1,-nbitq), 
to_sfixed(105807231.0/4294967296.0,1,-nbitq), 
to_sfixed(187063751.0/4294967296.0,1,-nbitq), 
to_sfixed(-349888069.0/4294967296.0,1,-nbitq), 
to_sfixed(394114685.0/4294967296.0,1,-nbitq), 
to_sfixed(-319627333.0/4294967296.0,1,-nbitq), 
to_sfixed(-442560922.0/4294967296.0,1,-nbitq), 
to_sfixed(228584560.0/4294967296.0,1,-nbitq), 
to_sfixed(91114709.0/4294967296.0,1,-nbitq), 
to_sfixed(-236659581.0/4294967296.0,1,-nbitq), 
to_sfixed(-41410064.0/4294967296.0,1,-nbitq), 
to_sfixed(80561883.0/4294967296.0,1,-nbitq), 
to_sfixed(487021605.0/4294967296.0,1,-nbitq), 
to_sfixed(-291286901.0/4294967296.0,1,-nbitq), 
to_sfixed(22679296.0/4294967296.0,1,-nbitq), 
to_sfixed(-92910974.0/4294967296.0,1,-nbitq), 
to_sfixed(153610041.0/4294967296.0,1,-nbitq), 
to_sfixed(-480880544.0/4294967296.0,1,-nbitq), 
to_sfixed(207404422.0/4294967296.0,1,-nbitq), 
to_sfixed(-289262160.0/4294967296.0,1,-nbitq), 
to_sfixed(441248375.0/4294967296.0,1,-nbitq), 
to_sfixed(84068178.0/4294967296.0,1,-nbitq), 
to_sfixed(-170330573.0/4294967296.0,1,-nbitq), 
to_sfixed(102865524.0/4294967296.0,1,-nbitq), 
to_sfixed(146737959.0/4294967296.0,1,-nbitq), 
to_sfixed(39882446.0/4294967296.0,1,-nbitq), 
to_sfixed(-448819977.0/4294967296.0,1,-nbitq), 
to_sfixed(190128204.0/4294967296.0,1,-nbitq), 
to_sfixed(-87842713.0/4294967296.0,1,-nbitq), 
to_sfixed(467325566.0/4294967296.0,1,-nbitq), 
to_sfixed(-557585291.0/4294967296.0,1,-nbitq), 
to_sfixed(406059765.0/4294967296.0,1,-nbitq), 
to_sfixed(24628162.0/4294967296.0,1,-nbitq), 
to_sfixed(-154894965.0/4294967296.0,1,-nbitq), 
to_sfixed(328690092.0/4294967296.0,1,-nbitq), 
to_sfixed(-320189233.0/4294967296.0,1,-nbitq), 
to_sfixed(-305638520.0/4294967296.0,1,-nbitq), 
to_sfixed(-211027486.0/4294967296.0,1,-nbitq), 
to_sfixed(134368734.0/4294967296.0,1,-nbitq), 
to_sfixed(34982960.0/4294967296.0,1,-nbitq), 
to_sfixed(-102370199.0/4294967296.0,1,-nbitq), 
to_sfixed(204846081.0/4294967296.0,1,-nbitq), 
to_sfixed(661983835.0/4294967296.0,1,-nbitq), 
to_sfixed(-213688048.0/4294967296.0,1,-nbitq), 
to_sfixed(785535938.0/4294967296.0,1,-nbitq), 
to_sfixed(-451060529.0/4294967296.0,1,-nbitq), 
to_sfixed(233900069.0/4294967296.0,1,-nbitq), 
to_sfixed(191022339.0/4294967296.0,1,-nbitq), 
to_sfixed(346899510.0/4294967296.0,1,-nbitq), 
to_sfixed(-728283.0/4294967296.0,1,-nbitq), 
to_sfixed(583884630.0/4294967296.0,1,-nbitq), 
to_sfixed(-139762265.0/4294967296.0,1,-nbitq), 
to_sfixed(-123080995.0/4294967296.0,1,-nbitq), 
to_sfixed(253455408.0/4294967296.0,1,-nbitq), 
to_sfixed(332187967.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(436881232.0/4294967296.0,1,-nbitq), 
to_sfixed(-151623509.0/4294967296.0,1,-nbitq), 
to_sfixed(680038634.0/4294967296.0,1,-nbitq), 
to_sfixed(-89054357.0/4294967296.0,1,-nbitq), 
to_sfixed(8216913.0/4294967296.0,1,-nbitq), 
to_sfixed(510189967.0/4294967296.0,1,-nbitq), 
to_sfixed(-43519979.0/4294967296.0,1,-nbitq), 
to_sfixed(-289815516.0/4294967296.0,1,-nbitq), 
to_sfixed(-169453896.0/4294967296.0,1,-nbitq), 
to_sfixed(231468076.0/4294967296.0,1,-nbitq), 
to_sfixed(642417130.0/4294967296.0,1,-nbitq), 
to_sfixed(-607075166.0/4294967296.0,1,-nbitq), 
to_sfixed(33510637.0/4294967296.0,1,-nbitq), 
to_sfixed(-445573676.0/4294967296.0,1,-nbitq), 
to_sfixed(-188192638.0/4294967296.0,1,-nbitq), 
to_sfixed(574262875.0/4294967296.0,1,-nbitq), 
to_sfixed(-58004125.0/4294967296.0,1,-nbitq), 
to_sfixed(374530787.0/4294967296.0,1,-nbitq), 
to_sfixed(-895940281.0/4294967296.0,1,-nbitq), 
to_sfixed(362807767.0/4294967296.0,1,-nbitq), 
to_sfixed(-257406404.0/4294967296.0,1,-nbitq), 
to_sfixed(-526140237.0/4294967296.0,1,-nbitq), 
to_sfixed(-934441213.0/4294967296.0,1,-nbitq), 
to_sfixed(223881200.0/4294967296.0,1,-nbitq), 
to_sfixed(118179948.0/4294967296.0,1,-nbitq), 
to_sfixed(-589920559.0/4294967296.0,1,-nbitq), 
to_sfixed(506746787.0/4294967296.0,1,-nbitq), 
to_sfixed(354261646.0/4294967296.0,1,-nbitq), 
to_sfixed(-396873274.0/4294967296.0,1,-nbitq), 
to_sfixed(462268611.0/4294967296.0,1,-nbitq), 
to_sfixed(-92940057.0/4294967296.0,1,-nbitq), 
to_sfixed(15788353.0/4294967296.0,1,-nbitq), 
to_sfixed(76067349.0/4294967296.0,1,-nbitq), 
to_sfixed(557390533.0/4294967296.0,1,-nbitq), 
to_sfixed(-40410718.0/4294967296.0,1,-nbitq), 
to_sfixed(-157424311.0/4294967296.0,1,-nbitq), 
to_sfixed(180982503.0/4294967296.0,1,-nbitq), 
to_sfixed(230145659.0/4294967296.0,1,-nbitq), 
to_sfixed(316559118.0/4294967296.0,1,-nbitq), 
to_sfixed(433977520.0/4294967296.0,1,-nbitq), 
to_sfixed(-114556657.0/4294967296.0,1,-nbitq), 
to_sfixed(-611042621.0/4294967296.0,1,-nbitq), 
to_sfixed(-664370683.0/4294967296.0,1,-nbitq), 
to_sfixed(-869683612.0/4294967296.0,1,-nbitq), 
to_sfixed(-265941313.0/4294967296.0,1,-nbitq), 
to_sfixed(-155124960.0/4294967296.0,1,-nbitq), 
to_sfixed(-230994131.0/4294967296.0,1,-nbitq), 
to_sfixed(-275329883.0/4294967296.0,1,-nbitq), 
to_sfixed(75693681.0/4294967296.0,1,-nbitq), 
to_sfixed(-652770943.0/4294967296.0,1,-nbitq), 
to_sfixed(-139726953.0/4294967296.0,1,-nbitq), 
to_sfixed(-296297185.0/4294967296.0,1,-nbitq), 
to_sfixed(362182337.0/4294967296.0,1,-nbitq), 
to_sfixed(-304670069.0/4294967296.0,1,-nbitq), 
to_sfixed(98249023.0/4294967296.0,1,-nbitq), 
to_sfixed(-96148311.0/4294967296.0,1,-nbitq), 
to_sfixed(-90703937.0/4294967296.0,1,-nbitq), 
to_sfixed(503014123.0/4294967296.0,1,-nbitq), 
to_sfixed(-198897998.0/4294967296.0,1,-nbitq), 
to_sfixed(389216382.0/4294967296.0,1,-nbitq), 
to_sfixed(-85991775.0/4294967296.0,1,-nbitq), 
to_sfixed(-136064525.0/4294967296.0,1,-nbitq), 
to_sfixed(-314574164.0/4294967296.0,1,-nbitq), 
to_sfixed(-338190571.0/4294967296.0,1,-nbitq), 
to_sfixed(-261363682.0/4294967296.0,1,-nbitq), 
to_sfixed(-38436747.0/4294967296.0,1,-nbitq), 
to_sfixed(-355780818.0/4294967296.0,1,-nbitq), 
to_sfixed(-16540639.0/4294967296.0,1,-nbitq), 
to_sfixed(38137164.0/4294967296.0,1,-nbitq), 
to_sfixed(935159988.0/4294967296.0,1,-nbitq), 
to_sfixed(-92053874.0/4294967296.0,1,-nbitq), 
to_sfixed(310191495.0/4294967296.0,1,-nbitq), 
to_sfixed(570660931.0/4294967296.0,1,-nbitq), 
to_sfixed(149415044.0/4294967296.0,1,-nbitq), 
to_sfixed(413882867.0/4294967296.0,1,-nbitq), 
to_sfixed(223668451.0/4294967296.0,1,-nbitq), 
to_sfixed(-174213109.0/4294967296.0,1,-nbitq), 
to_sfixed(223304349.0/4294967296.0,1,-nbitq), 
to_sfixed(-250612116.0/4294967296.0,1,-nbitq), 
to_sfixed(250684409.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-117208057.0/4294967296.0,1,-nbitq), 
to_sfixed(-182451145.0/4294967296.0,1,-nbitq), 
to_sfixed(394642821.0/4294967296.0,1,-nbitq), 
to_sfixed(583332658.0/4294967296.0,1,-nbitq), 
to_sfixed(-579792881.0/4294967296.0,1,-nbitq), 
to_sfixed(1056829089.0/4294967296.0,1,-nbitq), 
to_sfixed(457021236.0/4294967296.0,1,-nbitq), 
to_sfixed(282016426.0/4294967296.0,1,-nbitq), 
to_sfixed(112136297.0/4294967296.0,1,-nbitq), 
to_sfixed(-202628685.0/4294967296.0,1,-nbitq), 
to_sfixed(1228347646.0/4294967296.0,1,-nbitq), 
to_sfixed(-263763085.0/4294967296.0,1,-nbitq), 
to_sfixed(-677811597.0/4294967296.0,1,-nbitq), 
to_sfixed(288147953.0/4294967296.0,1,-nbitq), 
to_sfixed(-232008155.0/4294967296.0,1,-nbitq), 
to_sfixed(531579604.0/4294967296.0,1,-nbitq), 
to_sfixed(140890391.0/4294967296.0,1,-nbitq), 
to_sfixed(-364645656.0/4294967296.0,1,-nbitq), 
to_sfixed(-1454690659.0/4294967296.0,1,-nbitq), 
to_sfixed(732348303.0/4294967296.0,1,-nbitq), 
to_sfixed(-246028203.0/4294967296.0,1,-nbitq), 
to_sfixed(-494912704.0/4294967296.0,1,-nbitq), 
to_sfixed(-433759109.0/4294967296.0,1,-nbitq), 
to_sfixed(392015704.0/4294967296.0,1,-nbitq), 
to_sfixed(185578282.0/4294967296.0,1,-nbitq), 
to_sfixed(-574893541.0/4294967296.0,1,-nbitq), 
to_sfixed(400658247.0/4294967296.0,1,-nbitq), 
to_sfixed(690630100.0/4294967296.0,1,-nbitq), 
to_sfixed(-13710070.0/4294967296.0,1,-nbitq), 
to_sfixed(-72939990.0/4294967296.0,1,-nbitq), 
to_sfixed(336366025.0/4294967296.0,1,-nbitq), 
to_sfixed(528003563.0/4294967296.0,1,-nbitq), 
to_sfixed(548486032.0/4294967296.0,1,-nbitq), 
to_sfixed(74314767.0/4294967296.0,1,-nbitq), 
to_sfixed(166292497.0/4294967296.0,1,-nbitq), 
to_sfixed(-452885015.0/4294967296.0,1,-nbitq), 
to_sfixed(-267964155.0/4294967296.0,1,-nbitq), 
to_sfixed(-661609030.0/4294967296.0,1,-nbitq), 
to_sfixed(357619111.0/4294967296.0,1,-nbitq), 
to_sfixed(88806767.0/4294967296.0,1,-nbitq), 
to_sfixed(84458361.0/4294967296.0,1,-nbitq), 
to_sfixed(-253873085.0/4294967296.0,1,-nbitq), 
to_sfixed(207712388.0/4294967296.0,1,-nbitq), 
to_sfixed(-1081167983.0/4294967296.0,1,-nbitq), 
to_sfixed(-413673726.0/4294967296.0,1,-nbitq), 
to_sfixed(-521795136.0/4294967296.0,1,-nbitq), 
to_sfixed(-326410210.0/4294967296.0,1,-nbitq), 
to_sfixed(557937501.0/4294967296.0,1,-nbitq), 
to_sfixed(-329320624.0/4294967296.0,1,-nbitq), 
to_sfixed(-424181325.0/4294967296.0,1,-nbitq), 
to_sfixed(-213531479.0/4294967296.0,1,-nbitq), 
to_sfixed(-1201244.0/4294967296.0,1,-nbitq), 
to_sfixed(962554797.0/4294967296.0,1,-nbitq), 
to_sfixed(-987743901.0/4294967296.0,1,-nbitq), 
to_sfixed(-901970796.0/4294967296.0,1,-nbitq), 
to_sfixed(946891886.0/4294967296.0,1,-nbitq), 
to_sfixed(300265126.0/4294967296.0,1,-nbitq), 
to_sfixed(30800483.0/4294967296.0,1,-nbitq), 
to_sfixed(153658474.0/4294967296.0,1,-nbitq), 
to_sfixed(323515545.0/4294967296.0,1,-nbitq), 
to_sfixed(87932087.0/4294967296.0,1,-nbitq), 
to_sfixed(-590995.0/4294967296.0,1,-nbitq), 
to_sfixed(471429473.0/4294967296.0,1,-nbitq), 
to_sfixed(-299185312.0/4294967296.0,1,-nbitq), 
to_sfixed(211087313.0/4294967296.0,1,-nbitq), 
to_sfixed(-207470108.0/4294967296.0,1,-nbitq), 
to_sfixed(-1002195002.0/4294967296.0,1,-nbitq), 
to_sfixed(-228411035.0/4294967296.0,1,-nbitq), 
to_sfixed(292198829.0/4294967296.0,1,-nbitq), 
to_sfixed(-71886831.0/4294967296.0,1,-nbitq), 
to_sfixed(-42651897.0/4294967296.0,1,-nbitq), 
to_sfixed(376248115.0/4294967296.0,1,-nbitq), 
to_sfixed(305598785.0/4294967296.0,1,-nbitq), 
to_sfixed(-223820312.0/4294967296.0,1,-nbitq), 
to_sfixed(61742232.0/4294967296.0,1,-nbitq), 
to_sfixed(-132744347.0/4294967296.0,1,-nbitq), 
to_sfixed(-962865292.0/4294967296.0,1,-nbitq), 
to_sfixed(-29601690.0/4294967296.0,1,-nbitq), 
to_sfixed(-1197715663.0/4294967296.0,1,-nbitq), 
to_sfixed(-97699639.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-422032400.0/4294967296.0,1,-nbitq), 
to_sfixed(109963417.0/4294967296.0,1,-nbitq), 
to_sfixed(914254407.0/4294967296.0,1,-nbitq), 
to_sfixed(1197705180.0/4294967296.0,1,-nbitq), 
to_sfixed(440520808.0/4294967296.0,1,-nbitq), 
to_sfixed(1733793599.0/4294967296.0,1,-nbitq), 
to_sfixed(210910456.0/4294967296.0,1,-nbitq), 
to_sfixed(655984209.0/4294967296.0,1,-nbitq), 
to_sfixed(982853087.0/4294967296.0,1,-nbitq), 
to_sfixed(-169775348.0/4294967296.0,1,-nbitq), 
to_sfixed(299838326.0/4294967296.0,1,-nbitq), 
to_sfixed(-821791800.0/4294967296.0,1,-nbitq), 
to_sfixed(-1650608781.0/4294967296.0,1,-nbitq), 
to_sfixed(-544947769.0/4294967296.0,1,-nbitq), 
to_sfixed(-59736327.0/4294967296.0,1,-nbitq), 
to_sfixed(562157654.0/4294967296.0,1,-nbitq), 
to_sfixed(-187590953.0/4294967296.0,1,-nbitq), 
to_sfixed(-260318680.0/4294967296.0,1,-nbitq), 
to_sfixed(-1344158982.0/4294967296.0,1,-nbitq), 
to_sfixed(774364756.0/4294967296.0,1,-nbitq), 
to_sfixed(-347001.0/4294967296.0,1,-nbitq), 
to_sfixed(-18095217.0/4294967296.0,1,-nbitq), 
to_sfixed(-25354437.0/4294967296.0,1,-nbitq), 
to_sfixed(20318602.0/4294967296.0,1,-nbitq), 
to_sfixed(-182399517.0/4294967296.0,1,-nbitq), 
to_sfixed(-850275541.0/4294967296.0,1,-nbitq), 
to_sfixed(781965223.0/4294967296.0,1,-nbitq), 
to_sfixed(502398679.0/4294967296.0,1,-nbitq), 
to_sfixed(58878426.0/4294967296.0,1,-nbitq), 
to_sfixed(-579200513.0/4294967296.0,1,-nbitq), 
to_sfixed(1054388486.0/4294967296.0,1,-nbitq), 
to_sfixed(-159681958.0/4294967296.0,1,-nbitq), 
to_sfixed(222642279.0/4294967296.0,1,-nbitq), 
to_sfixed(52527308.0/4294967296.0,1,-nbitq), 
to_sfixed(-128373488.0/4294967296.0,1,-nbitq), 
to_sfixed(-1932941128.0/4294967296.0,1,-nbitq), 
to_sfixed(-523807049.0/4294967296.0,1,-nbitq), 
to_sfixed(-186978184.0/4294967296.0,1,-nbitq), 
to_sfixed(92711443.0/4294967296.0,1,-nbitq), 
to_sfixed(376080884.0/4294967296.0,1,-nbitq), 
to_sfixed(325179606.0/4294967296.0,1,-nbitq), 
to_sfixed(-263783189.0/4294967296.0,1,-nbitq), 
to_sfixed(206778297.0/4294967296.0,1,-nbitq), 
to_sfixed(-848662036.0/4294967296.0,1,-nbitq), 
to_sfixed(300226376.0/4294967296.0,1,-nbitq), 
to_sfixed(-379098443.0/4294967296.0,1,-nbitq), 
to_sfixed(-206751898.0/4294967296.0,1,-nbitq), 
to_sfixed(462963823.0/4294967296.0,1,-nbitq), 
to_sfixed(-105361173.0/4294967296.0,1,-nbitq), 
to_sfixed(411053123.0/4294967296.0,1,-nbitq), 
to_sfixed(-802123966.0/4294967296.0,1,-nbitq), 
to_sfixed(-78246784.0/4294967296.0,1,-nbitq), 
to_sfixed(1197710141.0/4294967296.0,1,-nbitq), 
to_sfixed(-583640824.0/4294967296.0,1,-nbitq), 
to_sfixed(-1527324764.0/4294967296.0,1,-nbitq), 
to_sfixed(346557738.0/4294967296.0,1,-nbitq), 
to_sfixed(516854580.0/4294967296.0,1,-nbitq), 
to_sfixed(16702849.0/4294967296.0,1,-nbitq), 
to_sfixed(416027903.0/4294967296.0,1,-nbitq), 
to_sfixed(-226891787.0/4294967296.0,1,-nbitq), 
to_sfixed(169954752.0/4294967296.0,1,-nbitq), 
to_sfixed(641626171.0/4294967296.0,1,-nbitq), 
to_sfixed(1326516651.0/4294967296.0,1,-nbitq), 
to_sfixed(260075466.0/4294967296.0,1,-nbitq), 
to_sfixed(-435855468.0/4294967296.0,1,-nbitq), 
to_sfixed(-33260477.0/4294967296.0,1,-nbitq), 
to_sfixed(-1520125182.0/4294967296.0,1,-nbitq), 
to_sfixed(-21160226.0/4294967296.0,1,-nbitq), 
to_sfixed(-383251927.0/4294967296.0,1,-nbitq), 
to_sfixed(-110796352.0/4294967296.0,1,-nbitq), 
to_sfixed(-451344978.0/4294967296.0,1,-nbitq), 
to_sfixed(168157542.0/4294967296.0,1,-nbitq), 
to_sfixed(709453249.0/4294967296.0,1,-nbitq), 
to_sfixed(-225117579.0/4294967296.0,1,-nbitq), 
to_sfixed(-254568561.0/4294967296.0,1,-nbitq), 
to_sfixed(-406483588.0/4294967296.0,1,-nbitq), 
to_sfixed(-996949661.0/4294967296.0,1,-nbitq), 
to_sfixed(-225577752.0/4294967296.0,1,-nbitq), 
to_sfixed(-1099005302.0/4294967296.0,1,-nbitq), 
to_sfixed(401268351.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-357395598.0/4294967296.0,1,-nbitq), 
to_sfixed(401713178.0/4294967296.0,1,-nbitq), 
to_sfixed(521784531.0/4294967296.0,1,-nbitq), 
to_sfixed(937257312.0/4294967296.0,1,-nbitq), 
to_sfixed(458666652.0/4294967296.0,1,-nbitq), 
to_sfixed(1533710599.0/4294967296.0,1,-nbitq), 
to_sfixed(245424053.0/4294967296.0,1,-nbitq), 
to_sfixed(1202799573.0/4294967296.0,1,-nbitq), 
to_sfixed(740466284.0/4294967296.0,1,-nbitq), 
to_sfixed(-381788869.0/4294967296.0,1,-nbitq), 
to_sfixed(89605991.0/4294967296.0,1,-nbitq), 
to_sfixed(-634298301.0/4294967296.0,1,-nbitq), 
to_sfixed(-620730862.0/4294967296.0,1,-nbitq), 
to_sfixed(-738012950.0/4294967296.0,1,-nbitq), 
to_sfixed(221269818.0/4294967296.0,1,-nbitq), 
to_sfixed(504644918.0/4294967296.0,1,-nbitq), 
to_sfixed(-162103835.0/4294967296.0,1,-nbitq), 
to_sfixed(285664638.0/4294967296.0,1,-nbitq), 
to_sfixed(-753010703.0/4294967296.0,1,-nbitq), 
to_sfixed(-39389191.0/4294967296.0,1,-nbitq), 
to_sfixed(-134229972.0/4294967296.0,1,-nbitq), 
to_sfixed(251212017.0/4294967296.0,1,-nbitq), 
to_sfixed(-628712430.0/4294967296.0,1,-nbitq), 
to_sfixed(-133358459.0/4294967296.0,1,-nbitq), 
to_sfixed(-55734480.0/4294967296.0,1,-nbitq), 
to_sfixed(-1395947627.0/4294967296.0,1,-nbitq), 
to_sfixed(282809868.0/4294967296.0,1,-nbitq), 
to_sfixed(115722106.0/4294967296.0,1,-nbitq), 
to_sfixed(425250846.0/4294967296.0,1,-nbitq), 
to_sfixed(-94494121.0/4294967296.0,1,-nbitq), 
to_sfixed(462467445.0/4294967296.0,1,-nbitq), 
to_sfixed(-22373755.0/4294967296.0,1,-nbitq), 
to_sfixed(422107033.0/4294967296.0,1,-nbitq), 
to_sfixed(675919387.0/4294967296.0,1,-nbitq), 
to_sfixed(-364143905.0/4294967296.0,1,-nbitq), 
to_sfixed(-1774223858.0/4294967296.0,1,-nbitq), 
to_sfixed(-545467530.0/4294967296.0,1,-nbitq), 
to_sfixed(553114122.0/4294967296.0,1,-nbitq), 
to_sfixed(243519689.0/4294967296.0,1,-nbitq), 
to_sfixed(386412457.0/4294967296.0,1,-nbitq), 
to_sfixed(313144001.0/4294967296.0,1,-nbitq), 
to_sfixed(-664939492.0/4294967296.0,1,-nbitq), 
to_sfixed(-471143668.0/4294967296.0,1,-nbitq), 
to_sfixed(-669744036.0/4294967296.0,1,-nbitq), 
to_sfixed(6056425.0/4294967296.0,1,-nbitq), 
to_sfixed(-800164964.0/4294967296.0,1,-nbitq), 
to_sfixed(182719691.0/4294967296.0,1,-nbitq), 
to_sfixed(282360647.0/4294967296.0,1,-nbitq), 
to_sfixed(-36854214.0/4294967296.0,1,-nbitq), 
to_sfixed(492006297.0/4294967296.0,1,-nbitq), 
to_sfixed(-245285478.0/4294967296.0,1,-nbitq), 
to_sfixed(-808206666.0/4294967296.0,1,-nbitq), 
to_sfixed(913518422.0/4294967296.0,1,-nbitq), 
to_sfixed(32939587.0/4294967296.0,1,-nbitq), 
to_sfixed(-158697703.0/4294967296.0,1,-nbitq), 
to_sfixed(637996385.0/4294967296.0,1,-nbitq), 
to_sfixed(310824162.0/4294967296.0,1,-nbitq), 
to_sfixed(14682084.0/4294967296.0,1,-nbitq), 
to_sfixed(-54259055.0/4294967296.0,1,-nbitq), 
to_sfixed(172003705.0/4294967296.0,1,-nbitq), 
to_sfixed(3370781.0/4294967296.0,1,-nbitq), 
to_sfixed(104261970.0/4294967296.0,1,-nbitq), 
to_sfixed(1045317232.0/4294967296.0,1,-nbitq), 
to_sfixed(125339959.0/4294967296.0,1,-nbitq), 
to_sfixed(-219547407.0/4294967296.0,1,-nbitq), 
to_sfixed(7209391.0/4294967296.0,1,-nbitq), 
to_sfixed(-2112830209.0/4294967296.0,1,-nbitq), 
to_sfixed(-183927203.0/4294967296.0,1,-nbitq), 
to_sfixed(173064791.0/4294967296.0,1,-nbitq), 
to_sfixed(611745883.0/4294967296.0,1,-nbitq), 
to_sfixed(-103569886.0/4294967296.0,1,-nbitq), 
to_sfixed(-149056853.0/4294967296.0,1,-nbitq), 
to_sfixed(551654679.0/4294967296.0,1,-nbitq), 
to_sfixed(-165892545.0/4294967296.0,1,-nbitq), 
to_sfixed(41318650.0/4294967296.0,1,-nbitq), 
to_sfixed(-528251672.0/4294967296.0,1,-nbitq), 
to_sfixed(-852205337.0/4294967296.0,1,-nbitq), 
to_sfixed(41509802.0/4294967296.0,1,-nbitq), 
to_sfixed(-699066255.0/4294967296.0,1,-nbitq), 
to_sfixed(306345882.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-231273081.0/4294967296.0,1,-nbitq), 
to_sfixed(574390069.0/4294967296.0,1,-nbitq), 
to_sfixed(181872153.0/4294967296.0,1,-nbitq), 
to_sfixed(1706334860.0/4294967296.0,1,-nbitq), 
to_sfixed(728340849.0/4294967296.0,1,-nbitq), 
to_sfixed(1192296325.0/4294967296.0,1,-nbitq), 
to_sfixed(-651883111.0/4294967296.0,1,-nbitq), 
to_sfixed(1359132477.0/4294967296.0,1,-nbitq), 
to_sfixed(-85099455.0/4294967296.0,1,-nbitq), 
to_sfixed(-108162757.0/4294967296.0,1,-nbitq), 
to_sfixed(315303633.0/4294967296.0,1,-nbitq), 
to_sfixed(266748030.0/4294967296.0,1,-nbitq), 
to_sfixed(-946570221.0/4294967296.0,1,-nbitq), 
to_sfixed(-652908801.0/4294967296.0,1,-nbitq), 
to_sfixed(61954383.0/4294967296.0,1,-nbitq), 
to_sfixed(-195222835.0/4294967296.0,1,-nbitq), 
to_sfixed(-18441961.0/4294967296.0,1,-nbitq), 
to_sfixed(42797673.0/4294967296.0,1,-nbitq), 
to_sfixed(223422345.0/4294967296.0,1,-nbitq), 
to_sfixed(448366548.0/4294967296.0,1,-nbitq), 
to_sfixed(83451549.0/4294967296.0,1,-nbitq), 
to_sfixed(352382785.0/4294967296.0,1,-nbitq), 
to_sfixed(-224609091.0/4294967296.0,1,-nbitq), 
to_sfixed(506151470.0/4294967296.0,1,-nbitq), 
to_sfixed(272850918.0/4294967296.0,1,-nbitq), 
to_sfixed(-548214947.0/4294967296.0,1,-nbitq), 
to_sfixed(284709801.0/4294967296.0,1,-nbitq), 
to_sfixed(631032371.0/4294967296.0,1,-nbitq), 
to_sfixed(16284480.0/4294967296.0,1,-nbitq), 
to_sfixed(-73301681.0/4294967296.0,1,-nbitq), 
to_sfixed(202904745.0/4294967296.0,1,-nbitq), 
to_sfixed(463244754.0/4294967296.0,1,-nbitq), 
to_sfixed(1287063869.0/4294967296.0,1,-nbitq), 
to_sfixed(1006399234.0/4294967296.0,1,-nbitq), 
to_sfixed(-1095941354.0/4294967296.0,1,-nbitq), 
to_sfixed(-1047406378.0/4294967296.0,1,-nbitq), 
to_sfixed(-1467754965.0/4294967296.0,1,-nbitq), 
to_sfixed(-105451223.0/4294967296.0,1,-nbitq), 
to_sfixed(-489825816.0/4294967296.0,1,-nbitq), 
to_sfixed(112493745.0/4294967296.0,1,-nbitq), 
to_sfixed(-470314999.0/4294967296.0,1,-nbitq), 
to_sfixed(-658968202.0/4294967296.0,1,-nbitq), 
to_sfixed(668054807.0/4294967296.0,1,-nbitq), 
to_sfixed(-235009824.0/4294967296.0,1,-nbitq), 
to_sfixed(481065573.0/4294967296.0,1,-nbitq), 
to_sfixed(-672492403.0/4294967296.0,1,-nbitq), 
to_sfixed(47457199.0/4294967296.0,1,-nbitq), 
to_sfixed(623051458.0/4294967296.0,1,-nbitq), 
to_sfixed(441561779.0/4294967296.0,1,-nbitq), 
to_sfixed(438416358.0/4294967296.0,1,-nbitq), 
to_sfixed(-194557363.0/4294967296.0,1,-nbitq), 
to_sfixed(-25743403.0/4294967296.0,1,-nbitq), 
to_sfixed(59501148.0/4294967296.0,1,-nbitq), 
to_sfixed(-83882038.0/4294967296.0,1,-nbitq), 
to_sfixed(130903893.0/4294967296.0,1,-nbitq), 
to_sfixed(115973773.0/4294967296.0,1,-nbitq), 
to_sfixed(-239882928.0/4294967296.0,1,-nbitq), 
to_sfixed(-107963773.0/4294967296.0,1,-nbitq), 
to_sfixed(344806905.0/4294967296.0,1,-nbitq), 
to_sfixed(-247464321.0/4294967296.0,1,-nbitq), 
to_sfixed(365051745.0/4294967296.0,1,-nbitq), 
to_sfixed(275361732.0/4294967296.0,1,-nbitq), 
to_sfixed(228537438.0/4294967296.0,1,-nbitq), 
to_sfixed(-89039981.0/4294967296.0,1,-nbitq), 
to_sfixed(-592964265.0/4294967296.0,1,-nbitq), 
to_sfixed(18468384.0/4294967296.0,1,-nbitq), 
to_sfixed(-2237238137.0/4294967296.0,1,-nbitq), 
to_sfixed(-268128506.0/4294967296.0,1,-nbitq), 
to_sfixed(-248717543.0/4294967296.0,1,-nbitq), 
to_sfixed(-235960939.0/4294967296.0,1,-nbitq), 
to_sfixed(-943460841.0/4294967296.0,1,-nbitq), 
to_sfixed(-352496497.0/4294967296.0,1,-nbitq), 
to_sfixed(47752649.0/4294967296.0,1,-nbitq), 
to_sfixed(189882491.0/4294967296.0,1,-nbitq), 
to_sfixed(-76710122.0/4294967296.0,1,-nbitq), 
to_sfixed(-196347536.0/4294967296.0,1,-nbitq), 
to_sfixed(-601613594.0/4294967296.0,1,-nbitq), 
to_sfixed(-763214407.0/4294967296.0,1,-nbitq), 
to_sfixed(-144074693.0/4294967296.0,1,-nbitq), 
to_sfixed(39887289.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-785068126.0/4294967296.0,1,-nbitq), 
to_sfixed(-185928688.0/4294967296.0,1,-nbitq), 
to_sfixed(398886129.0/4294967296.0,1,-nbitq), 
to_sfixed(1713721649.0/4294967296.0,1,-nbitq), 
to_sfixed(617249032.0/4294967296.0,1,-nbitq), 
to_sfixed(-87383509.0/4294967296.0,1,-nbitq), 
to_sfixed(-84500335.0/4294967296.0,1,-nbitq), 
to_sfixed(1553005560.0/4294967296.0,1,-nbitq), 
to_sfixed(-906674046.0/4294967296.0,1,-nbitq), 
to_sfixed(370427160.0/4294967296.0,1,-nbitq), 
to_sfixed(326668637.0/4294967296.0,1,-nbitq), 
to_sfixed(1102497607.0/4294967296.0,1,-nbitq), 
to_sfixed(-790791752.0/4294967296.0,1,-nbitq), 
to_sfixed(-1204387018.0/4294967296.0,1,-nbitq), 
to_sfixed(-384894968.0/4294967296.0,1,-nbitq), 
to_sfixed(337818270.0/4294967296.0,1,-nbitq), 
to_sfixed(292911734.0/4294967296.0,1,-nbitq), 
to_sfixed(-33951232.0/4294967296.0,1,-nbitq), 
to_sfixed(399564586.0/4294967296.0,1,-nbitq), 
to_sfixed(495440878.0/4294967296.0,1,-nbitq), 
to_sfixed(314733859.0/4294967296.0,1,-nbitq), 
to_sfixed(118826304.0/4294967296.0,1,-nbitq), 
to_sfixed(396613925.0/4294967296.0,1,-nbitq), 
to_sfixed(517778404.0/4294967296.0,1,-nbitq), 
to_sfixed(-101144992.0/4294967296.0,1,-nbitq), 
to_sfixed(-895753696.0/4294967296.0,1,-nbitq), 
to_sfixed(202097878.0/4294967296.0,1,-nbitq), 
to_sfixed(506731593.0/4294967296.0,1,-nbitq), 
to_sfixed(768444826.0/4294967296.0,1,-nbitq), 
to_sfixed(805347347.0/4294967296.0,1,-nbitq), 
to_sfixed(741524595.0/4294967296.0,1,-nbitq), 
to_sfixed(1519390953.0/4294967296.0,1,-nbitq), 
to_sfixed(1040336985.0/4294967296.0,1,-nbitq), 
to_sfixed(1321549072.0/4294967296.0,1,-nbitq), 
to_sfixed(-963089920.0/4294967296.0,1,-nbitq), 
to_sfixed(-785778493.0/4294967296.0,1,-nbitq), 
to_sfixed(-2053562571.0/4294967296.0,1,-nbitq), 
to_sfixed(-488499313.0/4294967296.0,1,-nbitq), 
to_sfixed(-181422532.0/4294967296.0,1,-nbitq), 
to_sfixed(-176944567.0/4294967296.0,1,-nbitq), 
to_sfixed(-8527655.0/4294967296.0,1,-nbitq), 
to_sfixed(-488360957.0/4294967296.0,1,-nbitq), 
to_sfixed(731204562.0/4294967296.0,1,-nbitq), 
to_sfixed(592031857.0/4294967296.0,1,-nbitq), 
to_sfixed(-319582648.0/4294967296.0,1,-nbitq), 
to_sfixed(-709898175.0/4294967296.0,1,-nbitq), 
to_sfixed(268691335.0/4294967296.0,1,-nbitq), 
to_sfixed(761405673.0/4294967296.0,1,-nbitq), 
to_sfixed(132395716.0/4294967296.0,1,-nbitq), 
to_sfixed(493208230.0/4294967296.0,1,-nbitq), 
to_sfixed(-698317186.0/4294967296.0,1,-nbitq), 
to_sfixed(-187218569.0/4294967296.0,1,-nbitq), 
to_sfixed(-674951488.0/4294967296.0,1,-nbitq), 
to_sfixed(903038643.0/4294967296.0,1,-nbitq), 
to_sfixed(1061424708.0/4294967296.0,1,-nbitq), 
to_sfixed(179250333.0/4294967296.0,1,-nbitq), 
to_sfixed(-127870755.0/4294967296.0,1,-nbitq), 
to_sfixed(215714990.0/4294967296.0,1,-nbitq), 
to_sfixed(-239769963.0/4294967296.0,1,-nbitq), 
to_sfixed(-301321597.0/4294967296.0,1,-nbitq), 
to_sfixed(-5085443.0/4294967296.0,1,-nbitq), 
to_sfixed(185386770.0/4294967296.0,1,-nbitq), 
to_sfixed(688535780.0/4294967296.0,1,-nbitq), 
to_sfixed(276394267.0/4294967296.0,1,-nbitq), 
to_sfixed(-728957715.0/4294967296.0,1,-nbitq), 
to_sfixed(-119569509.0/4294967296.0,1,-nbitq), 
to_sfixed(-2145309845.0/4294967296.0,1,-nbitq), 
to_sfixed(-81455318.0/4294967296.0,1,-nbitq), 
to_sfixed(156017738.0/4294967296.0,1,-nbitq), 
to_sfixed(-75642556.0/4294967296.0,1,-nbitq), 
to_sfixed(401163368.0/4294967296.0,1,-nbitq), 
to_sfixed(-490036854.0/4294967296.0,1,-nbitq), 
to_sfixed(364822473.0/4294967296.0,1,-nbitq), 
to_sfixed(154395918.0/4294967296.0,1,-nbitq), 
to_sfixed(-183373011.0/4294967296.0,1,-nbitq), 
to_sfixed(170461149.0/4294967296.0,1,-nbitq), 
to_sfixed(-284807909.0/4294967296.0,1,-nbitq), 
to_sfixed(-165605544.0/4294967296.0,1,-nbitq), 
to_sfixed(334980939.0/4294967296.0,1,-nbitq), 
to_sfixed(-303847870.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-645832912.0/4294967296.0,1,-nbitq), 
to_sfixed(-336824658.0/4294967296.0,1,-nbitq), 
to_sfixed(1232004459.0/4294967296.0,1,-nbitq), 
to_sfixed(1136547626.0/4294967296.0,1,-nbitq), 
to_sfixed(913361816.0/4294967296.0,1,-nbitq), 
to_sfixed(-1371784636.0/4294967296.0,1,-nbitq), 
to_sfixed(-409593442.0/4294967296.0,1,-nbitq), 
to_sfixed(-713206546.0/4294967296.0,1,-nbitq), 
to_sfixed(-1109211468.0/4294967296.0,1,-nbitq), 
to_sfixed(-388533404.0/4294967296.0,1,-nbitq), 
to_sfixed(-141255051.0/4294967296.0,1,-nbitq), 
to_sfixed(1087750649.0/4294967296.0,1,-nbitq), 
to_sfixed(-989828008.0/4294967296.0,1,-nbitq), 
to_sfixed(-1622948475.0/4294967296.0,1,-nbitq), 
to_sfixed(-244635620.0/4294967296.0,1,-nbitq), 
to_sfixed(367138678.0/4294967296.0,1,-nbitq), 
to_sfixed(193161671.0/4294967296.0,1,-nbitq), 
to_sfixed(-169567742.0/4294967296.0,1,-nbitq), 
to_sfixed(696334466.0/4294967296.0,1,-nbitq), 
to_sfixed(4433991.0/4294967296.0,1,-nbitq), 
to_sfixed(152907178.0/4294967296.0,1,-nbitq), 
to_sfixed(-356570726.0/4294967296.0,1,-nbitq), 
to_sfixed(387231507.0/4294967296.0,1,-nbitq), 
to_sfixed(121216222.0/4294967296.0,1,-nbitq), 
to_sfixed(196946608.0/4294967296.0,1,-nbitq), 
to_sfixed(-382876127.0/4294967296.0,1,-nbitq), 
to_sfixed(247923006.0/4294967296.0,1,-nbitq), 
to_sfixed(1207636534.0/4294967296.0,1,-nbitq), 
to_sfixed(744144185.0/4294967296.0,1,-nbitq), 
to_sfixed(41687805.0/4294967296.0,1,-nbitq), 
to_sfixed(1430182789.0/4294967296.0,1,-nbitq), 
to_sfixed(1060033547.0/4294967296.0,1,-nbitq), 
to_sfixed(820042669.0/4294967296.0,1,-nbitq), 
to_sfixed(1052501544.0/4294967296.0,1,-nbitq), 
to_sfixed(-55267870.0/4294967296.0,1,-nbitq), 
to_sfixed(-103403649.0/4294967296.0,1,-nbitq), 
to_sfixed(-1916680909.0/4294967296.0,1,-nbitq), 
to_sfixed(-160917496.0/4294967296.0,1,-nbitq), 
to_sfixed(-145540590.0/4294967296.0,1,-nbitq), 
to_sfixed(-46967898.0/4294967296.0,1,-nbitq), 
to_sfixed(-483161985.0/4294967296.0,1,-nbitq), 
to_sfixed(-487348412.0/4294967296.0,1,-nbitq), 
to_sfixed(1391118540.0/4294967296.0,1,-nbitq), 
to_sfixed(747733041.0/4294967296.0,1,-nbitq), 
to_sfixed(-469407129.0/4294967296.0,1,-nbitq), 
to_sfixed(-1684330392.0/4294967296.0,1,-nbitq), 
to_sfixed(111568780.0/4294967296.0,1,-nbitq), 
to_sfixed(1061813351.0/4294967296.0,1,-nbitq), 
to_sfixed(-423675582.0/4294967296.0,1,-nbitq), 
to_sfixed(685881392.0/4294967296.0,1,-nbitq), 
to_sfixed(-379670917.0/4294967296.0,1,-nbitq), 
to_sfixed(1998872.0/4294967296.0,1,-nbitq), 
to_sfixed(-1235222302.0/4294967296.0,1,-nbitq), 
to_sfixed(758608338.0/4294967296.0,1,-nbitq), 
to_sfixed(-144161255.0/4294967296.0,1,-nbitq), 
to_sfixed(554908847.0/4294967296.0,1,-nbitq), 
to_sfixed(-59788980.0/4294967296.0,1,-nbitq), 
to_sfixed(-583283841.0/4294967296.0,1,-nbitq), 
to_sfixed(-218585536.0/4294967296.0,1,-nbitq), 
to_sfixed(-335952741.0/4294967296.0,1,-nbitq), 
to_sfixed(71188326.0/4294967296.0,1,-nbitq), 
to_sfixed(136923262.0/4294967296.0,1,-nbitq), 
to_sfixed(1517052932.0/4294967296.0,1,-nbitq), 
to_sfixed(79313373.0/4294967296.0,1,-nbitq), 
to_sfixed(-558835630.0/4294967296.0,1,-nbitq), 
to_sfixed(-409963725.0/4294967296.0,1,-nbitq), 
to_sfixed(-132120932.0/4294967296.0,1,-nbitq), 
to_sfixed(-597780522.0/4294967296.0,1,-nbitq), 
to_sfixed(-154387226.0/4294967296.0,1,-nbitq), 
to_sfixed(264502612.0/4294967296.0,1,-nbitq), 
to_sfixed(-400259563.0/4294967296.0,1,-nbitq), 
to_sfixed(-126301042.0/4294967296.0,1,-nbitq), 
to_sfixed(1066852166.0/4294967296.0,1,-nbitq), 
to_sfixed(-50297835.0/4294967296.0,1,-nbitq), 
to_sfixed(201812577.0/4294967296.0,1,-nbitq), 
to_sfixed(417240843.0/4294967296.0,1,-nbitq), 
to_sfixed(-961067674.0/4294967296.0,1,-nbitq), 
to_sfixed(-161049803.0/4294967296.0,1,-nbitq), 
to_sfixed(973753876.0/4294967296.0,1,-nbitq), 
to_sfixed(-23957581.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-702375114.0/4294967296.0,1,-nbitq), 
to_sfixed(235791303.0/4294967296.0,1,-nbitq), 
to_sfixed(-23299974.0/4294967296.0,1,-nbitq), 
to_sfixed(14041696.0/4294967296.0,1,-nbitq), 
to_sfixed(495986464.0/4294967296.0,1,-nbitq), 
to_sfixed(-941559268.0/4294967296.0,1,-nbitq), 
to_sfixed(207247805.0/4294967296.0,1,-nbitq), 
to_sfixed(-1149998113.0/4294967296.0,1,-nbitq), 
to_sfixed(-450323918.0/4294967296.0,1,-nbitq), 
to_sfixed(-38426096.0/4294967296.0,1,-nbitq), 
to_sfixed(105869908.0/4294967296.0,1,-nbitq), 
to_sfixed(793332889.0/4294967296.0,1,-nbitq), 
to_sfixed(-902919196.0/4294967296.0,1,-nbitq), 
to_sfixed(-1143003658.0/4294967296.0,1,-nbitq), 
to_sfixed(-404387860.0/4294967296.0,1,-nbitq), 
to_sfixed(482740753.0/4294967296.0,1,-nbitq), 
to_sfixed(59671903.0/4294967296.0,1,-nbitq), 
to_sfixed(74474909.0/4294967296.0,1,-nbitq), 
to_sfixed(1572012396.0/4294967296.0,1,-nbitq), 
to_sfixed(80944856.0/4294967296.0,1,-nbitq), 
to_sfixed(293922299.0/4294967296.0,1,-nbitq), 
to_sfixed(-485386583.0/4294967296.0,1,-nbitq), 
to_sfixed(464923748.0/4294967296.0,1,-nbitq), 
to_sfixed(408766511.0/4294967296.0,1,-nbitq), 
to_sfixed(-134463771.0/4294967296.0,1,-nbitq), 
to_sfixed(-322768981.0/4294967296.0,1,-nbitq), 
to_sfixed(-347077305.0/4294967296.0,1,-nbitq), 
to_sfixed(599591067.0/4294967296.0,1,-nbitq), 
to_sfixed(-841999247.0/4294967296.0,1,-nbitq), 
to_sfixed(-180032616.0/4294967296.0,1,-nbitq), 
to_sfixed(1600995726.0/4294967296.0,1,-nbitq), 
to_sfixed(1568748762.0/4294967296.0,1,-nbitq), 
to_sfixed(1135608141.0/4294967296.0,1,-nbitq), 
to_sfixed(497513338.0/4294967296.0,1,-nbitq), 
to_sfixed(-242730399.0/4294967296.0,1,-nbitq), 
to_sfixed(2051939235.0/4294967296.0,1,-nbitq), 
to_sfixed(-1647350940.0/4294967296.0,1,-nbitq), 
to_sfixed(-464349129.0/4294967296.0,1,-nbitq), 
to_sfixed(-565484372.0/4294967296.0,1,-nbitq), 
to_sfixed(-580084707.0/4294967296.0,1,-nbitq), 
to_sfixed(-892637293.0/4294967296.0,1,-nbitq), 
to_sfixed(-1125385393.0/4294967296.0,1,-nbitq), 
to_sfixed(699346641.0/4294967296.0,1,-nbitq), 
to_sfixed(12968834.0/4294967296.0,1,-nbitq), 
to_sfixed(-572086723.0/4294967296.0,1,-nbitq), 
to_sfixed(-939119211.0/4294967296.0,1,-nbitq), 
to_sfixed(-18001454.0/4294967296.0,1,-nbitq), 
to_sfixed(193643530.0/4294967296.0,1,-nbitq), 
to_sfixed(-628891284.0/4294967296.0,1,-nbitq), 
to_sfixed(-165801447.0/4294967296.0,1,-nbitq), 
to_sfixed(24326011.0/4294967296.0,1,-nbitq), 
to_sfixed(-956780414.0/4294967296.0,1,-nbitq), 
to_sfixed(-1783362893.0/4294967296.0,1,-nbitq), 
to_sfixed(553459941.0/4294967296.0,1,-nbitq), 
to_sfixed(875817810.0/4294967296.0,1,-nbitq), 
to_sfixed(596315373.0/4294967296.0,1,-nbitq), 
to_sfixed(-894331470.0/4294967296.0,1,-nbitq), 
to_sfixed(133936205.0/4294967296.0,1,-nbitq), 
to_sfixed(-86790991.0/4294967296.0,1,-nbitq), 
to_sfixed(-237310123.0/4294967296.0,1,-nbitq), 
to_sfixed(-287909357.0/4294967296.0,1,-nbitq), 
to_sfixed(1129919435.0/4294967296.0,1,-nbitq), 
to_sfixed(1145232740.0/4294967296.0,1,-nbitq), 
to_sfixed(-73354653.0/4294967296.0,1,-nbitq), 
to_sfixed(-264147742.0/4294967296.0,1,-nbitq), 
to_sfixed(-337965826.0/4294967296.0,1,-nbitq), 
to_sfixed(1085141657.0/4294967296.0,1,-nbitq), 
to_sfixed(1058530985.0/4294967296.0,1,-nbitq), 
to_sfixed(71441698.0/4294967296.0,1,-nbitq), 
to_sfixed(255569551.0/4294967296.0,1,-nbitq), 
to_sfixed(-505870940.0/4294967296.0,1,-nbitq), 
to_sfixed(-4000216.0/4294967296.0,1,-nbitq), 
to_sfixed(950745516.0/4294967296.0,1,-nbitq), 
to_sfixed(63668960.0/4294967296.0,1,-nbitq), 
to_sfixed(418541582.0/4294967296.0,1,-nbitq), 
to_sfixed(-577465434.0/4294967296.0,1,-nbitq), 
to_sfixed(-468374513.0/4294967296.0,1,-nbitq), 
to_sfixed(377169553.0/4294967296.0,1,-nbitq), 
to_sfixed(774329927.0/4294967296.0,1,-nbitq), 
to_sfixed(-23307292.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-259770601.0/4294967296.0,1,-nbitq), 
to_sfixed(-966648707.0/4294967296.0,1,-nbitq), 
to_sfixed(-591885070.0/4294967296.0,1,-nbitq), 
to_sfixed(-137311940.0/4294967296.0,1,-nbitq), 
to_sfixed(-1083664962.0/4294967296.0,1,-nbitq), 
to_sfixed(-305302387.0/4294967296.0,1,-nbitq), 
to_sfixed(-10708009.0/4294967296.0,1,-nbitq), 
to_sfixed(-820584914.0/4294967296.0,1,-nbitq), 
to_sfixed(-322492800.0/4294967296.0,1,-nbitq), 
to_sfixed(270629418.0/4294967296.0,1,-nbitq), 
to_sfixed(731380613.0/4294967296.0,1,-nbitq), 
to_sfixed(1161032400.0/4294967296.0,1,-nbitq), 
to_sfixed(-2040316065.0/4294967296.0,1,-nbitq), 
to_sfixed(-1655956325.0/4294967296.0,1,-nbitq), 
to_sfixed(-434020562.0/4294967296.0,1,-nbitq), 
to_sfixed(-235017976.0/4294967296.0,1,-nbitq), 
to_sfixed(77791598.0/4294967296.0,1,-nbitq), 
to_sfixed(-148911721.0/4294967296.0,1,-nbitq), 
to_sfixed(406945897.0/4294967296.0,1,-nbitq), 
to_sfixed(427942873.0/4294967296.0,1,-nbitq), 
to_sfixed(-373119701.0/4294967296.0,1,-nbitq), 
to_sfixed(-679805930.0/4294967296.0,1,-nbitq), 
to_sfixed(1074237571.0/4294967296.0,1,-nbitq), 
to_sfixed(932309357.0/4294967296.0,1,-nbitq), 
to_sfixed(82290264.0/4294967296.0,1,-nbitq), 
to_sfixed(702244919.0/4294967296.0,1,-nbitq), 
to_sfixed(-669625638.0/4294967296.0,1,-nbitq), 
to_sfixed(-947104716.0/4294967296.0,1,-nbitq), 
to_sfixed(-1715616891.0/4294967296.0,1,-nbitq), 
to_sfixed(-412594741.0/4294967296.0,1,-nbitq), 
to_sfixed(1372748892.0/4294967296.0,1,-nbitq), 
to_sfixed(559443245.0/4294967296.0,1,-nbitq), 
to_sfixed(1271562018.0/4294967296.0,1,-nbitq), 
to_sfixed(-613459904.0/4294967296.0,1,-nbitq), 
to_sfixed(653398385.0/4294967296.0,1,-nbitq), 
to_sfixed(2600327589.0/4294967296.0,1,-nbitq), 
to_sfixed(-1460290411.0/4294967296.0,1,-nbitq), 
to_sfixed(-522727164.0/4294967296.0,1,-nbitq), 
to_sfixed(-520809965.0/4294967296.0,1,-nbitq), 
to_sfixed(79417196.0/4294967296.0,1,-nbitq), 
to_sfixed(-84410834.0/4294967296.0,1,-nbitq), 
to_sfixed(-498806546.0/4294967296.0,1,-nbitq), 
to_sfixed(-422304840.0/4294967296.0,1,-nbitq), 
to_sfixed(-172830117.0/4294967296.0,1,-nbitq), 
to_sfixed(-966687627.0/4294967296.0,1,-nbitq), 
to_sfixed(-693483468.0/4294967296.0,1,-nbitq), 
to_sfixed(202427292.0/4294967296.0,1,-nbitq), 
to_sfixed(-402757995.0/4294967296.0,1,-nbitq), 
to_sfixed(-301175680.0/4294967296.0,1,-nbitq), 
to_sfixed(-850590200.0/4294967296.0,1,-nbitq), 
to_sfixed(669434098.0/4294967296.0,1,-nbitq), 
to_sfixed(-266498498.0/4294967296.0,1,-nbitq), 
to_sfixed(-2527114604.0/4294967296.0,1,-nbitq), 
to_sfixed(-317516683.0/4294967296.0,1,-nbitq), 
to_sfixed(-346613159.0/4294967296.0,1,-nbitq), 
to_sfixed(-76793843.0/4294967296.0,1,-nbitq), 
to_sfixed(-620468768.0/4294967296.0,1,-nbitq), 
to_sfixed(475342412.0/4294967296.0,1,-nbitq), 
to_sfixed(-201755734.0/4294967296.0,1,-nbitq), 
to_sfixed(111497719.0/4294967296.0,1,-nbitq), 
to_sfixed(425815993.0/4294967296.0,1,-nbitq), 
to_sfixed(1068985538.0/4294967296.0,1,-nbitq), 
to_sfixed(901951466.0/4294967296.0,1,-nbitq), 
to_sfixed(154999714.0/4294967296.0,1,-nbitq), 
to_sfixed(329272802.0/4294967296.0,1,-nbitq), 
to_sfixed(-112773102.0/4294967296.0,1,-nbitq), 
to_sfixed(191512293.0/4294967296.0,1,-nbitq), 
to_sfixed(609354558.0/4294967296.0,1,-nbitq), 
to_sfixed(310030755.0/4294967296.0,1,-nbitq), 
to_sfixed(-370138895.0/4294967296.0,1,-nbitq), 
to_sfixed(-1083770621.0/4294967296.0,1,-nbitq), 
to_sfixed(-91498127.0/4294967296.0,1,-nbitq), 
to_sfixed(258254653.0/4294967296.0,1,-nbitq), 
to_sfixed(-273083962.0/4294967296.0,1,-nbitq), 
to_sfixed(-231252123.0/4294967296.0,1,-nbitq), 
to_sfixed(-493717936.0/4294967296.0,1,-nbitq), 
to_sfixed(-1052815897.0/4294967296.0,1,-nbitq), 
to_sfixed(-85953191.0/4294967296.0,1,-nbitq), 
to_sfixed(308954005.0/4294967296.0,1,-nbitq), 
to_sfixed(-393952752.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-384344417.0/4294967296.0,1,-nbitq), 
to_sfixed(-543650086.0/4294967296.0,1,-nbitq), 
to_sfixed(-776120474.0/4294967296.0,1,-nbitq), 
to_sfixed(457431919.0/4294967296.0,1,-nbitq), 
to_sfixed(-2430780868.0/4294967296.0,1,-nbitq), 
to_sfixed(-460520394.0/4294967296.0,1,-nbitq), 
to_sfixed(655403780.0/4294967296.0,1,-nbitq), 
to_sfixed(-425501174.0/4294967296.0,1,-nbitq), 
to_sfixed(-79226314.0/4294967296.0,1,-nbitq), 
to_sfixed(49616577.0/4294967296.0,1,-nbitq), 
to_sfixed(163738712.0/4294967296.0,1,-nbitq), 
to_sfixed(361234024.0/4294967296.0,1,-nbitq), 
to_sfixed(-2382552102.0/4294967296.0,1,-nbitq), 
to_sfixed(-1260771553.0/4294967296.0,1,-nbitq), 
to_sfixed(-28192954.0/4294967296.0,1,-nbitq), 
to_sfixed(-213137908.0/4294967296.0,1,-nbitq), 
to_sfixed(-366549425.0/4294967296.0,1,-nbitq), 
to_sfixed(98684638.0/4294967296.0,1,-nbitq), 
to_sfixed(-1755246268.0/4294967296.0,1,-nbitq), 
to_sfixed(473667903.0/4294967296.0,1,-nbitq), 
to_sfixed(-361478986.0/4294967296.0,1,-nbitq), 
to_sfixed(-1036556344.0/4294967296.0,1,-nbitq), 
to_sfixed(821691672.0/4294967296.0,1,-nbitq), 
to_sfixed(101317041.0/4294967296.0,1,-nbitq), 
to_sfixed(-260307058.0/4294967296.0,1,-nbitq), 
to_sfixed(1237571980.0/4294967296.0,1,-nbitq), 
to_sfixed(-1022233793.0/4294967296.0,1,-nbitq), 
to_sfixed(-1378681501.0/4294967296.0,1,-nbitq), 
to_sfixed(-635840333.0/4294967296.0,1,-nbitq), 
to_sfixed(-601625324.0/4294967296.0,1,-nbitq), 
to_sfixed(47869500.0/4294967296.0,1,-nbitq), 
to_sfixed(300001161.0/4294967296.0,1,-nbitq), 
to_sfixed(1066845724.0/4294967296.0,1,-nbitq), 
to_sfixed(-1455322702.0/4294967296.0,1,-nbitq), 
to_sfixed(982671961.0/4294967296.0,1,-nbitq), 
to_sfixed(1216663537.0/4294967296.0,1,-nbitq), 
to_sfixed(-513168914.0/4294967296.0,1,-nbitq), 
to_sfixed(15873097.0/4294967296.0,1,-nbitq), 
to_sfixed(-79520185.0/4294967296.0,1,-nbitq), 
to_sfixed(-324624153.0/4294967296.0,1,-nbitq), 
to_sfixed(241638465.0/4294967296.0,1,-nbitq), 
to_sfixed(-90288148.0/4294967296.0,1,-nbitq), 
to_sfixed(-1083107997.0/4294967296.0,1,-nbitq), 
to_sfixed(-171459402.0/4294967296.0,1,-nbitq), 
to_sfixed(167808714.0/4294967296.0,1,-nbitq), 
to_sfixed(-345362296.0/4294967296.0,1,-nbitq), 
to_sfixed(-347698406.0/4294967296.0,1,-nbitq), 
to_sfixed(-1020388025.0/4294967296.0,1,-nbitq), 
to_sfixed(54761849.0/4294967296.0,1,-nbitq), 
to_sfixed(-220678400.0/4294967296.0,1,-nbitq), 
to_sfixed(723460542.0/4294967296.0,1,-nbitq), 
to_sfixed(-271794800.0/4294967296.0,1,-nbitq), 
to_sfixed(-2607780603.0/4294967296.0,1,-nbitq), 
to_sfixed(-49761245.0/4294967296.0,1,-nbitq), 
to_sfixed(556580891.0/4294967296.0,1,-nbitq), 
to_sfixed(-85982899.0/4294967296.0,1,-nbitq), 
to_sfixed(-1198976289.0/4294967296.0,1,-nbitq), 
to_sfixed(198980909.0/4294967296.0,1,-nbitq), 
to_sfixed(-257761976.0/4294967296.0,1,-nbitq), 
to_sfixed(-205723025.0/4294967296.0,1,-nbitq), 
to_sfixed(-259044939.0/4294967296.0,1,-nbitq), 
to_sfixed(1447615138.0/4294967296.0,1,-nbitq), 
to_sfixed(511772143.0/4294967296.0,1,-nbitq), 
to_sfixed(-288172116.0/4294967296.0,1,-nbitq), 
to_sfixed(272571964.0/4294967296.0,1,-nbitq), 
to_sfixed(2482856.0/4294967296.0,1,-nbitq), 
to_sfixed(-59425439.0/4294967296.0,1,-nbitq), 
to_sfixed(1559032787.0/4294967296.0,1,-nbitq), 
to_sfixed(303292885.0/4294967296.0,1,-nbitq), 
to_sfixed(-651369290.0/4294967296.0,1,-nbitq), 
to_sfixed(241882668.0/4294967296.0,1,-nbitq), 
to_sfixed(537607660.0/4294967296.0,1,-nbitq), 
to_sfixed(-590205179.0/4294967296.0,1,-nbitq), 
to_sfixed(358625215.0/4294967296.0,1,-nbitq), 
to_sfixed(266430879.0/4294967296.0,1,-nbitq), 
to_sfixed(35260277.0/4294967296.0,1,-nbitq), 
to_sfixed(-750001598.0/4294967296.0,1,-nbitq), 
to_sfixed(-24863287.0/4294967296.0,1,-nbitq), 
to_sfixed(-445560554.0/4294967296.0,1,-nbitq), 
to_sfixed(-360997994.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-90411022.0/4294967296.0,1,-nbitq), 
to_sfixed(-74131625.0/4294967296.0,1,-nbitq), 
to_sfixed(12370298.0/4294967296.0,1,-nbitq), 
to_sfixed(348705925.0/4294967296.0,1,-nbitq), 
to_sfixed(-1987312652.0/4294967296.0,1,-nbitq), 
to_sfixed(89932472.0/4294967296.0,1,-nbitq), 
to_sfixed(340776817.0/4294967296.0,1,-nbitq), 
to_sfixed(-385858732.0/4294967296.0,1,-nbitq), 
to_sfixed(816859926.0/4294967296.0,1,-nbitq), 
to_sfixed(358664379.0/4294967296.0,1,-nbitq), 
to_sfixed(303969268.0/4294967296.0,1,-nbitq), 
to_sfixed(372582143.0/4294967296.0,1,-nbitq), 
to_sfixed(-458784959.0/4294967296.0,1,-nbitq), 
to_sfixed(-706148464.0/4294967296.0,1,-nbitq), 
to_sfixed(254221000.0/4294967296.0,1,-nbitq), 
to_sfixed(-458378215.0/4294967296.0,1,-nbitq), 
to_sfixed(250799340.0/4294967296.0,1,-nbitq), 
to_sfixed(-394665810.0/4294967296.0,1,-nbitq), 
to_sfixed(-827366924.0/4294967296.0,1,-nbitq), 
to_sfixed(929238160.0/4294967296.0,1,-nbitq), 
to_sfixed(195920696.0/4294967296.0,1,-nbitq), 
to_sfixed(-247471322.0/4294967296.0,1,-nbitq), 
to_sfixed(354121174.0/4294967296.0,1,-nbitq), 
to_sfixed(-357414.0/4294967296.0,1,-nbitq), 
to_sfixed(377028949.0/4294967296.0,1,-nbitq), 
to_sfixed(460207441.0/4294967296.0,1,-nbitq), 
to_sfixed(-532487320.0/4294967296.0,1,-nbitq), 
to_sfixed(-811351523.0/4294967296.0,1,-nbitq), 
to_sfixed(235437511.0/4294967296.0,1,-nbitq), 
to_sfixed(-598506266.0/4294967296.0,1,-nbitq), 
to_sfixed(-766682352.0/4294967296.0,1,-nbitq), 
to_sfixed(-272143026.0/4294967296.0,1,-nbitq), 
to_sfixed(754434335.0/4294967296.0,1,-nbitq), 
to_sfixed(-237648376.0/4294967296.0,1,-nbitq), 
to_sfixed(1081749495.0/4294967296.0,1,-nbitq), 
to_sfixed(208314764.0/4294967296.0,1,-nbitq), 
to_sfixed(170299856.0/4294967296.0,1,-nbitq), 
to_sfixed(441862465.0/4294967296.0,1,-nbitq), 
to_sfixed(333403093.0/4294967296.0,1,-nbitq), 
to_sfixed(-13647983.0/4294967296.0,1,-nbitq), 
to_sfixed(931687002.0/4294967296.0,1,-nbitq), 
to_sfixed(432445579.0/4294967296.0,1,-nbitq), 
to_sfixed(-1289120675.0/4294967296.0,1,-nbitq), 
to_sfixed(244662556.0/4294967296.0,1,-nbitq), 
to_sfixed(10315499.0/4294967296.0,1,-nbitq), 
to_sfixed(-518974861.0/4294967296.0,1,-nbitq), 
to_sfixed(346058217.0/4294967296.0,1,-nbitq), 
to_sfixed(-407267590.0/4294967296.0,1,-nbitq), 
to_sfixed(73830623.0/4294967296.0,1,-nbitq), 
to_sfixed(130133334.0/4294967296.0,1,-nbitq), 
to_sfixed(722851030.0/4294967296.0,1,-nbitq), 
to_sfixed(-42928708.0/4294967296.0,1,-nbitq), 
to_sfixed(-1476463917.0/4294967296.0,1,-nbitq), 
to_sfixed(-456356000.0/4294967296.0,1,-nbitq), 
to_sfixed(130829833.0/4294967296.0,1,-nbitq), 
to_sfixed(-4736087.0/4294967296.0,1,-nbitq), 
to_sfixed(-1180216292.0/4294967296.0,1,-nbitq), 
to_sfixed(925941288.0/4294967296.0,1,-nbitq), 
to_sfixed(-354847740.0/4294967296.0,1,-nbitq), 
to_sfixed(72339318.0/4294967296.0,1,-nbitq), 
to_sfixed(94363392.0/4294967296.0,1,-nbitq), 
to_sfixed(1262052462.0/4294967296.0,1,-nbitq), 
to_sfixed(-1287547862.0/4294967296.0,1,-nbitq), 
to_sfixed(-424289334.0/4294967296.0,1,-nbitq), 
to_sfixed(-213160103.0/4294967296.0,1,-nbitq), 
to_sfixed(-391664601.0/4294967296.0,1,-nbitq), 
to_sfixed(-1031827274.0/4294967296.0,1,-nbitq), 
to_sfixed(1251372399.0/4294967296.0,1,-nbitq), 
to_sfixed(-100476107.0/4294967296.0,1,-nbitq), 
to_sfixed(-702653300.0/4294967296.0,1,-nbitq), 
to_sfixed(1030899077.0/4294967296.0,1,-nbitq), 
to_sfixed(339487339.0/4294967296.0,1,-nbitq), 
to_sfixed(-1060273744.0/4294967296.0,1,-nbitq), 
to_sfixed(177684383.0/4294967296.0,1,-nbitq), 
to_sfixed(-94060519.0/4294967296.0,1,-nbitq), 
to_sfixed(338750612.0/4294967296.0,1,-nbitq), 
to_sfixed(55283843.0/4294967296.0,1,-nbitq), 
to_sfixed(547511858.0/4294967296.0,1,-nbitq), 
to_sfixed(-583009610.0/4294967296.0,1,-nbitq), 
to_sfixed(-10238717.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-162357116.0/4294967296.0,1,-nbitq), 
to_sfixed(-86594561.0/4294967296.0,1,-nbitq), 
to_sfixed(595989942.0/4294967296.0,1,-nbitq), 
to_sfixed(-357040097.0/4294967296.0,1,-nbitq), 
to_sfixed(-1172310028.0/4294967296.0,1,-nbitq), 
to_sfixed(1100106097.0/4294967296.0,1,-nbitq), 
to_sfixed(144610995.0/4294967296.0,1,-nbitq), 
to_sfixed(579282585.0/4294967296.0,1,-nbitq), 
to_sfixed(647954981.0/4294967296.0,1,-nbitq), 
to_sfixed(65133680.0/4294967296.0,1,-nbitq), 
to_sfixed(-7610806.0/4294967296.0,1,-nbitq), 
to_sfixed(516471572.0/4294967296.0,1,-nbitq), 
to_sfixed(721749669.0/4294967296.0,1,-nbitq), 
to_sfixed(16853663.0/4294967296.0,1,-nbitq), 
to_sfixed(243036616.0/4294967296.0,1,-nbitq), 
to_sfixed(-226703748.0/4294967296.0,1,-nbitq), 
to_sfixed(33322413.0/4294967296.0,1,-nbitq), 
to_sfixed(247849663.0/4294967296.0,1,-nbitq), 
to_sfixed(-894443946.0/4294967296.0,1,-nbitq), 
to_sfixed(967280480.0/4294967296.0,1,-nbitq), 
to_sfixed(-50177888.0/4294967296.0,1,-nbitq), 
to_sfixed(60132245.0/4294967296.0,1,-nbitq), 
to_sfixed(258758236.0/4294967296.0,1,-nbitq), 
to_sfixed(-1146793520.0/4294967296.0,1,-nbitq), 
to_sfixed(372278538.0/4294967296.0,1,-nbitq), 
to_sfixed(664774431.0/4294967296.0,1,-nbitq), 
to_sfixed(-707803132.0/4294967296.0,1,-nbitq), 
to_sfixed(-607980062.0/4294967296.0,1,-nbitq), 
to_sfixed(-522509894.0/4294967296.0,1,-nbitq), 
to_sfixed(-288971253.0/4294967296.0,1,-nbitq), 
to_sfixed(-1091687550.0/4294967296.0,1,-nbitq), 
to_sfixed(-718613394.0/4294967296.0,1,-nbitq), 
to_sfixed(545480639.0/4294967296.0,1,-nbitq), 
to_sfixed(161786829.0/4294967296.0,1,-nbitq), 
to_sfixed(242033572.0/4294967296.0,1,-nbitq), 
to_sfixed(198307806.0/4294967296.0,1,-nbitq), 
to_sfixed(671119084.0/4294967296.0,1,-nbitq), 
to_sfixed(278103447.0/4294967296.0,1,-nbitq), 
to_sfixed(45940039.0/4294967296.0,1,-nbitq), 
to_sfixed(68186003.0/4294967296.0,1,-nbitq), 
to_sfixed(1117192752.0/4294967296.0,1,-nbitq), 
to_sfixed(725418016.0/4294967296.0,1,-nbitq), 
to_sfixed(-1489652129.0/4294967296.0,1,-nbitq), 
to_sfixed(1402565996.0/4294967296.0,1,-nbitq), 
to_sfixed(454498827.0/4294967296.0,1,-nbitq), 
to_sfixed(-69471618.0/4294967296.0,1,-nbitq), 
to_sfixed(-104183571.0/4294967296.0,1,-nbitq), 
to_sfixed(-639723729.0/4294967296.0,1,-nbitq), 
to_sfixed(112791682.0/4294967296.0,1,-nbitq), 
to_sfixed(575241408.0/4294967296.0,1,-nbitq), 
to_sfixed(224228503.0/4294967296.0,1,-nbitq), 
to_sfixed(74833466.0/4294967296.0,1,-nbitq), 
to_sfixed(-429689524.0/4294967296.0,1,-nbitq), 
to_sfixed(-782027147.0/4294967296.0,1,-nbitq), 
to_sfixed(-905371749.0/4294967296.0,1,-nbitq), 
to_sfixed(-40033020.0/4294967296.0,1,-nbitq), 
to_sfixed(-530242717.0/4294967296.0,1,-nbitq), 
to_sfixed(1331178786.0/4294967296.0,1,-nbitq), 
to_sfixed(75804036.0/4294967296.0,1,-nbitq), 
to_sfixed(155206279.0/4294967296.0,1,-nbitq), 
to_sfixed(272010249.0/4294967296.0,1,-nbitq), 
to_sfixed(636884622.0/4294967296.0,1,-nbitq), 
to_sfixed(-1173986334.0/4294967296.0,1,-nbitq), 
to_sfixed(-478784821.0/4294967296.0,1,-nbitq), 
to_sfixed(-791445711.0/4294967296.0,1,-nbitq), 
to_sfixed(154722469.0/4294967296.0,1,-nbitq), 
to_sfixed(-2107835357.0/4294967296.0,1,-nbitq), 
to_sfixed(205212552.0/4294967296.0,1,-nbitq), 
to_sfixed(148025524.0/4294967296.0,1,-nbitq), 
to_sfixed(-45412121.0/4294967296.0,1,-nbitq), 
to_sfixed(958175257.0/4294967296.0,1,-nbitq), 
to_sfixed(-522804284.0/4294967296.0,1,-nbitq), 
to_sfixed(-1443245702.0/4294967296.0,1,-nbitq), 
to_sfixed(232842981.0/4294967296.0,1,-nbitq), 
to_sfixed(-222737841.0/4294967296.0,1,-nbitq), 
to_sfixed(1067289617.0/4294967296.0,1,-nbitq), 
to_sfixed(-185638038.0/4294967296.0,1,-nbitq), 
to_sfixed(820781391.0/4294967296.0,1,-nbitq), 
to_sfixed(-555703196.0/4294967296.0,1,-nbitq), 
to_sfixed(-203510165.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(197522370.0/4294967296.0,1,-nbitq), 
to_sfixed(392932284.0/4294967296.0,1,-nbitq), 
to_sfixed(1154156791.0/4294967296.0,1,-nbitq), 
to_sfixed(-929388759.0/4294967296.0,1,-nbitq), 
to_sfixed(-751647829.0/4294967296.0,1,-nbitq), 
to_sfixed(475286277.0/4294967296.0,1,-nbitq), 
to_sfixed(242564160.0/4294967296.0,1,-nbitq), 
to_sfixed(1064775830.0/4294967296.0,1,-nbitq), 
to_sfixed(90055847.0/4294967296.0,1,-nbitq), 
to_sfixed(-187455712.0/4294967296.0,1,-nbitq), 
to_sfixed(505383171.0/4294967296.0,1,-nbitq), 
to_sfixed(1031023398.0/4294967296.0,1,-nbitq), 
to_sfixed(493971054.0/4294967296.0,1,-nbitq), 
to_sfixed(598311802.0/4294967296.0,1,-nbitq), 
to_sfixed(-307980899.0/4294967296.0,1,-nbitq), 
to_sfixed(-248787277.0/4294967296.0,1,-nbitq), 
to_sfixed(-303148992.0/4294967296.0,1,-nbitq), 
to_sfixed(-216587942.0/4294967296.0,1,-nbitq), 
to_sfixed(-964074671.0/4294967296.0,1,-nbitq), 
to_sfixed(41832196.0/4294967296.0,1,-nbitq), 
to_sfixed(-299036942.0/4294967296.0,1,-nbitq), 
to_sfixed(-376892031.0/4294967296.0,1,-nbitq), 
to_sfixed(-745441074.0/4294967296.0,1,-nbitq), 
to_sfixed(48013033.0/4294967296.0,1,-nbitq), 
to_sfixed(27784011.0/4294967296.0,1,-nbitq), 
to_sfixed(575759440.0/4294967296.0,1,-nbitq), 
to_sfixed(-522489707.0/4294967296.0,1,-nbitq), 
to_sfixed(508623241.0/4294967296.0,1,-nbitq), 
to_sfixed(685415268.0/4294967296.0,1,-nbitq), 
to_sfixed(110472355.0/4294967296.0,1,-nbitq), 
to_sfixed(-1064531607.0/4294967296.0,1,-nbitq), 
to_sfixed(-378189832.0/4294967296.0,1,-nbitq), 
to_sfixed(1053943703.0/4294967296.0,1,-nbitq), 
to_sfixed(1354457132.0/4294967296.0,1,-nbitq), 
to_sfixed(443513983.0/4294967296.0,1,-nbitq), 
to_sfixed(179643572.0/4294967296.0,1,-nbitq), 
to_sfixed(860923088.0/4294967296.0,1,-nbitq), 
to_sfixed(257966899.0/4294967296.0,1,-nbitq), 
to_sfixed(29251385.0/4294967296.0,1,-nbitq), 
to_sfixed(240399917.0/4294967296.0,1,-nbitq), 
to_sfixed(595710723.0/4294967296.0,1,-nbitq), 
to_sfixed(1066132255.0/4294967296.0,1,-nbitq), 
to_sfixed(-1188363347.0/4294967296.0,1,-nbitq), 
to_sfixed(2225594628.0/4294967296.0,1,-nbitq), 
to_sfixed(140503111.0/4294967296.0,1,-nbitq), 
to_sfixed(-229884212.0/4294967296.0,1,-nbitq), 
to_sfixed(-205760683.0/4294967296.0,1,-nbitq), 
to_sfixed(-620543194.0/4294967296.0,1,-nbitq), 
to_sfixed(-572060184.0/4294967296.0,1,-nbitq), 
to_sfixed(111977775.0/4294967296.0,1,-nbitq), 
to_sfixed(319365186.0/4294967296.0,1,-nbitq), 
to_sfixed(-25139067.0/4294967296.0,1,-nbitq), 
to_sfixed(-517765994.0/4294967296.0,1,-nbitq), 
to_sfixed(13153425.0/4294967296.0,1,-nbitq), 
to_sfixed(-1240658640.0/4294967296.0,1,-nbitq), 
to_sfixed(-293387340.0/4294967296.0,1,-nbitq), 
to_sfixed(-640915564.0/4294967296.0,1,-nbitq), 
to_sfixed(1568592626.0/4294967296.0,1,-nbitq), 
to_sfixed(122605290.0/4294967296.0,1,-nbitq), 
to_sfixed(-78720567.0/4294967296.0,1,-nbitq), 
to_sfixed(207520055.0/4294967296.0,1,-nbitq), 
to_sfixed(-327090667.0/4294967296.0,1,-nbitq), 
to_sfixed(207382781.0/4294967296.0,1,-nbitq), 
to_sfixed(-760942915.0/4294967296.0,1,-nbitq), 
to_sfixed(-460882541.0/4294967296.0,1,-nbitq), 
to_sfixed(-1545262.0/4294967296.0,1,-nbitq), 
to_sfixed(-2752393896.0/4294967296.0,1,-nbitq), 
to_sfixed(40164661.0/4294967296.0,1,-nbitq), 
to_sfixed(221917193.0/4294967296.0,1,-nbitq), 
to_sfixed(-247524186.0/4294967296.0,1,-nbitq), 
to_sfixed(1220187303.0/4294967296.0,1,-nbitq), 
to_sfixed(-282364341.0/4294967296.0,1,-nbitq), 
to_sfixed(-445670774.0/4294967296.0,1,-nbitq), 
to_sfixed(128892801.0/4294967296.0,1,-nbitq), 
to_sfixed(270443706.0/4294967296.0,1,-nbitq), 
to_sfixed(795684411.0/4294967296.0,1,-nbitq), 
to_sfixed(-625375042.0/4294967296.0,1,-nbitq), 
to_sfixed(-194504539.0/4294967296.0,1,-nbitq), 
to_sfixed(135002239.0/4294967296.0,1,-nbitq), 
to_sfixed(-278371659.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-252243054.0/4294967296.0,1,-nbitq), 
to_sfixed(329274303.0/4294967296.0,1,-nbitq), 
to_sfixed(1288669276.0/4294967296.0,1,-nbitq), 
to_sfixed(-139232069.0/4294967296.0,1,-nbitq), 
to_sfixed(-968690107.0/4294967296.0,1,-nbitq), 
to_sfixed(604335373.0/4294967296.0,1,-nbitq), 
to_sfixed(-383541244.0/4294967296.0,1,-nbitq), 
to_sfixed(308365526.0/4294967296.0,1,-nbitq), 
to_sfixed(349119538.0/4294967296.0,1,-nbitq), 
to_sfixed(176017926.0/4294967296.0,1,-nbitq), 
to_sfixed(576761799.0/4294967296.0,1,-nbitq), 
to_sfixed(803127462.0/4294967296.0,1,-nbitq), 
to_sfixed(-351204470.0/4294967296.0,1,-nbitq), 
to_sfixed(605887365.0/4294967296.0,1,-nbitq), 
to_sfixed(346730395.0/4294967296.0,1,-nbitq), 
to_sfixed(291317957.0/4294967296.0,1,-nbitq), 
to_sfixed(-271880276.0/4294967296.0,1,-nbitq), 
to_sfixed(-234084974.0/4294967296.0,1,-nbitq), 
to_sfixed(-505060319.0/4294967296.0,1,-nbitq), 
to_sfixed(-268922182.0/4294967296.0,1,-nbitq), 
to_sfixed(335158593.0/4294967296.0,1,-nbitq), 
to_sfixed(87204009.0/4294967296.0,1,-nbitq), 
to_sfixed(-1093647063.0/4294967296.0,1,-nbitq), 
to_sfixed(-573941691.0/4294967296.0,1,-nbitq), 
to_sfixed(-14438383.0/4294967296.0,1,-nbitq), 
to_sfixed(-296517684.0/4294967296.0,1,-nbitq), 
to_sfixed(15350689.0/4294967296.0,1,-nbitq), 
to_sfixed(534065685.0/4294967296.0,1,-nbitq), 
to_sfixed(358363349.0/4294967296.0,1,-nbitq), 
to_sfixed(485388402.0/4294967296.0,1,-nbitq), 
to_sfixed(-573545028.0/4294967296.0,1,-nbitq), 
to_sfixed(162073123.0/4294967296.0,1,-nbitq), 
to_sfixed(513245445.0/4294967296.0,1,-nbitq), 
to_sfixed(730988545.0/4294967296.0,1,-nbitq), 
to_sfixed(151640016.0/4294967296.0,1,-nbitq), 
to_sfixed(-337459729.0/4294967296.0,1,-nbitq), 
to_sfixed(1213575020.0/4294967296.0,1,-nbitq), 
to_sfixed(650590518.0/4294967296.0,1,-nbitq), 
to_sfixed(-180849941.0/4294967296.0,1,-nbitq), 
to_sfixed(308539643.0/4294967296.0,1,-nbitq), 
to_sfixed(396803916.0/4294967296.0,1,-nbitq), 
to_sfixed(956514686.0/4294967296.0,1,-nbitq), 
to_sfixed(-1096977135.0/4294967296.0,1,-nbitq), 
to_sfixed(897984218.0/4294967296.0,1,-nbitq), 
to_sfixed(592580017.0/4294967296.0,1,-nbitq), 
to_sfixed(-854996271.0/4294967296.0,1,-nbitq), 
to_sfixed(-161828582.0/4294967296.0,1,-nbitq), 
to_sfixed(-179782904.0/4294967296.0,1,-nbitq), 
to_sfixed(-519097776.0/4294967296.0,1,-nbitq), 
to_sfixed(1098691627.0/4294967296.0,1,-nbitq), 
to_sfixed(930338030.0/4294967296.0,1,-nbitq), 
to_sfixed(605001883.0/4294967296.0,1,-nbitq), 
to_sfixed(75669573.0/4294967296.0,1,-nbitq), 
to_sfixed(274423918.0/4294967296.0,1,-nbitq), 
to_sfixed(-2081514966.0/4294967296.0,1,-nbitq), 
to_sfixed(773270170.0/4294967296.0,1,-nbitq), 
to_sfixed(182556580.0/4294967296.0,1,-nbitq), 
to_sfixed(1554963831.0/4294967296.0,1,-nbitq), 
to_sfixed(-198329879.0/4294967296.0,1,-nbitq), 
to_sfixed(-28499087.0/4294967296.0,1,-nbitq), 
to_sfixed(299273444.0/4294967296.0,1,-nbitq), 
to_sfixed(-976627007.0/4294967296.0,1,-nbitq), 
to_sfixed(-30581692.0/4294967296.0,1,-nbitq), 
to_sfixed(-1273774692.0/4294967296.0,1,-nbitq), 
to_sfixed(-560345891.0/4294967296.0,1,-nbitq), 
to_sfixed(-188108964.0/4294967296.0,1,-nbitq), 
to_sfixed(-1572965175.0/4294967296.0,1,-nbitq), 
to_sfixed(-34753012.0/4294967296.0,1,-nbitq), 
to_sfixed(-148010052.0/4294967296.0,1,-nbitq), 
to_sfixed(-87797368.0/4294967296.0,1,-nbitq), 
to_sfixed(800774669.0/4294967296.0,1,-nbitq), 
to_sfixed(-362328244.0/4294967296.0,1,-nbitq), 
to_sfixed(-270152892.0/4294967296.0,1,-nbitq), 
to_sfixed(-190322706.0/4294967296.0,1,-nbitq), 
to_sfixed(-206662086.0/4294967296.0,1,-nbitq), 
to_sfixed(1179854931.0/4294967296.0,1,-nbitq), 
to_sfixed(-981682656.0/4294967296.0,1,-nbitq), 
to_sfixed(-249325887.0/4294967296.0,1,-nbitq), 
to_sfixed(45957871.0/4294967296.0,1,-nbitq), 
to_sfixed(102490541.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(297728312.0/4294967296.0,1,-nbitq), 
to_sfixed(-1122090237.0/4294967296.0,1,-nbitq), 
to_sfixed(1548023261.0/4294967296.0,1,-nbitq), 
to_sfixed(843821749.0/4294967296.0,1,-nbitq), 
to_sfixed(-656830164.0/4294967296.0,1,-nbitq), 
to_sfixed(-121485233.0/4294967296.0,1,-nbitq), 
to_sfixed(-106357808.0/4294967296.0,1,-nbitq), 
to_sfixed(226969038.0/4294967296.0,1,-nbitq), 
to_sfixed(840865719.0/4294967296.0,1,-nbitq), 
to_sfixed(-27357922.0/4294967296.0,1,-nbitq), 
to_sfixed(-862166255.0/4294967296.0,1,-nbitq), 
to_sfixed(894226627.0/4294967296.0,1,-nbitq), 
to_sfixed(-22282068.0/4294967296.0,1,-nbitq), 
to_sfixed(-636817839.0/4294967296.0,1,-nbitq), 
to_sfixed(381640032.0/4294967296.0,1,-nbitq), 
to_sfixed(885129081.0/4294967296.0,1,-nbitq), 
to_sfixed(388630656.0/4294967296.0,1,-nbitq), 
to_sfixed(41391601.0/4294967296.0,1,-nbitq), 
to_sfixed(-996674344.0/4294967296.0,1,-nbitq), 
to_sfixed(-329997710.0/4294967296.0,1,-nbitq), 
to_sfixed(-12805348.0/4294967296.0,1,-nbitq), 
to_sfixed(207387623.0/4294967296.0,1,-nbitq), 
to_sfixed(-1323995891.0/4294967296.0,1,-nbitq), 
to_sfixed(-596740572.0/4294967296.0,1,-nbitq), 
to_sfixed(208685310.0/4294967296.0,1,-nbitq), 
to_sfixed(-727852097.0/4294967296.0,1,-nbitq), 
to_sfixed(571756590.0/4294967296.0,1,-nbitq), 
to_sfixed(822656360.0/4294967296.0,1,-nbitq), 
to_sfixed(-141974110.0/4294967296.0,1,-nbitq), 
to_sfixed(1715949450.0/4294967296.0,1,-nbitq), 
to_sfixed(14506763.0/4294967296.0,1,-nbitq), 
to_sfixed(-156906718.0/4294967296.0,1,-nbitq), 
to_sfixed(320330011.0/4294967296.0,1,-nbitq), 
to_sfixed(400821299.0/4294967296.0,1,-nbitq), 
to_sfixed(500303825.0/4294967296.0,1,-nbitq), 
to_sfixed(744428348.0/4294967296.0,1,-nbitq), 
to_sfixed(991374815.0/4294967296.0,1,-nbitq), 
to_sfixed(1027820509.0/4294967296.0,1,-nbitq), 
to_sfixed(-201706776.0/4294967296.0,1,-nbitq), 
to_sfixed(513320577.0/4294967296.0,1,-nbitq), 
to_sfixed(-29440262.0/4294967296.0,1,-nbitq), 
to_sfixed(-102283016.0/4294967296.0,1,-nbitq), 
to_sfixed(-836788449.0/4294967296.0,1,-nbitq), 
to_sfixed(312021100.0/4294967296.0,1,-nbitq), 
to_sfixed(259128312.0/4294967296.0,1,-nbitq), 
to_sfixed(-637609570.0/4294967296.0,1,-nbitq), 
to_sfixed(191228470.0/4294967296.0,1,-nbitq), 
to_sfixed(-366837972.0/4294967296.0,1,-nbitq), 
to_sfixed(-1134683055.0/4294967296.0,1,-nbitq), 
to_sfixed(876818543.0/4294967296.0,1,-nbitq), 
to_sfixed(439640088.0/4294967296.0,1,-nbitq), 
to_sfixed(448872512.0/4294967296.0,1,-nbitq), 
to_sfixed(74737299.0/4294967296.0,1,-nbitq), 
to_sfixed(195760295.0/4294967296.0,1,-nbitq), 
to_sfixed(-2167963907.0/4294967296.0,1,-nbitq), 
to_sfixed(1098932762.0/4294967296.0,1,-nbitq), 
to_sfixed(179508667.0/4294967296.0,1,-nbitq), 
to_sfixed(1568098112.0/4294967296.0,1,-nbitq), 
to_sfixed(403561691.0/4294967296.0,1,-nbitq), 
to_sfixed(-64128156.0/4294967296.0,1,-nbitq), 
to_sfixed(-73258585.0/4294967296.0,1,-nbitq), 
to_sfixed(100780163.0/4294967296.0,1,-nbitq), 
to_sfixed(-585057269.0/4294967296.0,1,-nbitq), 
to_sfixed(-996398544.0/4294967296.0,1,-nbitq), 
to_sfixed(423410327.0/4294967296.0,1,-nbitq), 
to_sfixed(146654811.0/4294967296.0,1,-nbitq), 
to_sfixed(314307212.0/4294967296.0,1,-nbitq), 
to_sfixed(-305483787.0/4294967296.0,1,-nbitq), 
to_sfixed(-233093698.0/4294967296.0,1,-nbitq), 
to_sfixed(610318895.0/4294967296.0,1,-nbitq), 
to_sfixed(556018908.0/4294967296.0,1,-nbitq), 
to_sfixed(-432481824.0/4294967296.0,1,-nbitq), 
to_sfixed(106275046.0/4294967296.0,1,-nbitq), 
to_sfixed(-154768884.0/4294967296.0,1,-nbitq), 
to_sfixed(4119735.0/4294967296.0,1,-nbitq), 
to_sfixed(802085855.0/4294967296.0,1,-nbitq), 
to_sfixed(-149360515.0/4294967296.0,1,-nbitq), 
to_sfixed(-286597837.0/4294967296.0,1,-nbitq), 
to_sfixed(705003007.0/4294967296.0,1,-nbitq), 
to_sfixed(-104028622.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-325495221.0/4294967296.0,1,-nbitq), 
to_sfixed(-1120484642.0/4294967296.0,1,-nbitq), 
to_sfixed(741305293.0/4294967296.0,1,-nbitq), 
to_sfixed(1045163924.0/4294967296.0,1,-nbitq), 
to_sfixed(-866617473.0/4294967296.0,1,-nbitq), 
to_sfixed(-120564944.0/4294967296.0,1,-nbitq), 
to_sfixed(-270370989.0/4294967296.0,1,-nbitq), 
to_sfixed(779621047.0/4294967296.0,1,-nbitq), 
to_sfixed(672443142.0/4294967296.0,1,-nbitq), 
to_sfixed(136372431.0/4294967296.0,1,-nbitq), 
to_sfixed(-348213799.0/4294967296.0,1,-nbitq), 
to_sfixed(336162102.0/4294967296.0,1,-nbitq), 
to_sfixed(180684601.0/4294967296.0,1,-nbitq), 
to_sfixed(626580573.0/4294967296.0,1,-nbitq), 
to_sfixed(-66988164.0/4294967296.0,1,-nbitq), 
to_sfixed(598221124.0/4294967296.0,1,-nbitq), 
to_sfixed(-335297654.0/4294967296.0,1,-nbitq), 
to_sfixed(56488604.0/4294967296.0,1,-nbitq), 
to_sfixed(-642496810.0/4294967296.0,1,-nbitq), 
to_sfixed(-699258641.0/4294967296.0,1,-nbitq), 
to_sfixed(-80506069.0/4294967296.0,1,-nbitq), 
to_sfixed(450413511.0/4294967296.0,1,-nbitq), 
to_sfixed(-1033105474.0/4294967296.0,1,-nbitq), 
to_sfixed(561496772.0/4294967296.0,1,-nbitq), 
to_sfixed(42086430.0/4294967296.0,1,-nbitq), 
to_sfixed(-544959585.0/4294967296.0,1,-nbitq), 
to_sfixed(389011962.0/4294967296.0,1,-nbitq), 
to_sfixed(156131389.0/4294967296.0,1,-nbitq), 
to_sfixed(-32501474.0/4294967296.0,1,-nbitq), 
to_sfixed(1570168543.0/4294967296.0,1,-nbitq), 
to_sfixed(850264897.0/4294967296.0,1,-nbitq), 
to_sfixed(349878718.0/4294967296.0,1,-nbitq), 
to_sfixed(-64561640.0/4294967296.0,1,-nbitq), 
to_sfixed(-268358801.0/4294967296.0,1,-nbitq), 
to_sfixed(441792115.0/4294967296.0,1,-nbitq), 
to_sfixed(210086692.0/4294967296.0,1,-nbitq), 
to_sfixed(476417391.0/4294967296.0,1,-nbitq), 
to_sfixed(620210765.0/4294967296.0,1,-nbitq), 
to_sfixed(-208859646.0/4294967296.0,1,-nbitq), 
to_sfixed(564845212.0/4294967296.0,1,-nbitq), 
to_sfixed(-235640188.0/4294967296.0,1,-nbitq), 
to_sfixed(-216894797.0/4294967296.0,1,-nbitq), 
to_sfixed(-1095535137.0/4294967296.0,1,-nbitq), 
to_sfixed(66420085.0/4294967296.0,1,-nbitq), 
to_sfixed(444301921.0/4294967296.0,1,-nbitq), 
to_sfixed(-1090074913.0/4294967296.0,1,-nbitq), 
to_sfixed(-197809259.0/4294967296.0,1,-nbitq), 
to_sfixed(-3772786.0/4294967296.0,1,-nbitq), 
to_sfixed(-1124585978.0/4294967296.0,1,-nbitq), 
to_sfixed(467818147.0/4294967296.0,1,-nbitq), 
to_sfixed(-21156061.0/4294967296.0,1,-nbitq), 
to_sfixed(257392920.0/4294967296.0,1,-nbitq), 
to_sfixed(328789274.0/4294967296.0,1,-nbitq), 
to_sfixed(-311380547.0/4294967296.0,1,-nbitq), 
to_sfixed(-1619289410.0/4294967296.0,1,-nbitq), 
to_sfixed(833536084.0/4294967296.0,1,-nbitq), 
to_sfixed(574050164.0/4294967296.0,1,-nbitq), 
to_sfixed(894736871.0/4294967296.0,1,-nbitq), 
to_sfixed(-70097248.0/4294967296.0,1,-nbitq), 
to_sfixed(133721289.0/4294967296.0,1,-nbitq), 
to_sfixed(-221859528.0/4294967296.0,1,-nbitq), 
to_sfixed(-640799950.0/4294967296.0,1,-nbitq), 
to_sfixed(-251635669.0/4294967296.0,1,-nbitq), 
to_sfixed(256428862.0/4294967296.0,1,-nbitq), 
to_sfixed(-145209858.0/4294967296.0,1,-nbitq), 
to_sfixed(170339856.0/4294967296.0,1,-nbitq), 
to_sfixed(866353704.0/4294967296.0,1,-nbitq), 
to_sfixed(-527449599.0/4294967296.0,1,-nbitq), 
to_sfixed(366106005.0/4294967296.0,1,-nbitq), 
to_sfixed(731833588.0/4294967296.0,1,-nbitq), 
to_sfixed(214574262.0/4294967296.0,1,-nbitq), 
to_sfixed(190731404.0/4294967296.0,1,-nbitq), 
to_sfixed(-39208092.0/4294967296.0,1,-nbitq), 
to_sfixed(252260859.0/4294967296.0,1,-nbitq), 
to_sfixed(107427600.0/4294967296.0,1,-nbitq), 
to_sfixed(552792582.0/4294967296.0,1,-nbitq), 
to_sfixed(-58446981.0/4294967296.0,1,-nbitq), 
to_sfixed(-44763560.0/4294967296.0,1,-nbitq), 
to_sfixed(323825295.0/4294967296.0,1,-nbitq), 
to_sfixed(256197047.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-37767630.0/4294967296.0,1,-nbitq), 
to_sfixed(-1158500116.0/4294967296.0,1,-nbitq), 
to_sfixed(465916173.0/4294967296.0,1,-nbitq), 
to_sfixed(1341558841.0/4294967296.0,1,-nbitq), 
to_sfixed(-415664121.0/4294967296.0,1,-nbitq), 
to_sfixed(-119235688.0/4294967296.0,1,-nbitq), 
to_sfixed(159204935.0/4294967296.0,1,-nbitq), 
to_sfixed(42830874.0/4294967296.0,1,-nbitq), 
to_sfixed(307151404.0/4294967296.0,1,-nbitq), 
to_sfixed(389206183.0/4294967296.0,1,-nbitq), 
to_sfixed(-126567584.0/4294967296.0,1,-nbitq), 
to_sfixed(653305961.0/4294967296.0,1,-nbitq), 
to_sfixed(334603435.0/4294967296.0,1,-nbitq), 
to_sfixed(143024427.0/4294967296.0,1,-nbitq), 
to_sfixed(-27516168.0/4294967296.0,1,-nbitq), 
to_sfixed(256159304.0/4294967296.0,1,-nbitq), 
to_sfixed(63372399.0/4294967296.0,1,-nbitq), 
to_sfixed(-231325599.0/4294967296.0,1,-nbitq), 
to_sfixed(-1017539264.0/4294967296.0,1,-nbitq), 
to_sfixed(-114257012.0/4294967296.0,1,-nbitq), 
to_sfixed(9771287.0/4294967296.0,1,-nbitq), 
to_sfixed(229852280.0/4294967296.0,1,-nbitq), 
to_sfixed(-870162940.0/4294967296.0,1,-nbitq), 
to_sfixed(-124017468.0/4294967296.0,1,-nbitq), 
to_sfixed(-79861845.0/4294967296.0,1,-nbitq), 
to_sfixed(-556532307.0/4294967296.0,1,-nbitq), 
to_sfixed(214296845.0/4294967296.0,1,-nbitq), 
to_sfixed(-186743742.0/4294967296.0,1,-nbitq), 
to_sfixed(-167656582.0/4294967296.0,1,-nbitq), 
to_sfixed(1175876604.0/4294967296.0,1,-nbitq), 
to_sfixed(1406984470.0/4294967296.0,1,-nbitq), 
to_sfixed(467821189.0/4294967296.0,1,-nbitq), 
to_sfixed(-361843815.0/4294967296.0,1,-nbitq), 
to_sfixed(17520767.0/4294967296.0,1,-nbitq), 
to_sfixed(-158327340.0/4294967296.0,1,-nbitq), 
to_sfixed(239143444.0/4294967296.0,1,-nbitq), 
to_sfixed(181177563.0/4294967296.0,1,-nbitq), 
to_sfixed(314209873.0/4294967296.0,1,-nbitq), 
to_sfixed(204111727.0/4294967296.0,1,-nbitq), 
to_sfixed(295472810.0/4294967296.0,1,-nbitq), 
to_sfixed(185510961.0/4294967296.0,1,-nbitq), 
to_sfixed(235120079.0/4294967296.0,1,-nbitq), 
to_sfixed(-834418307.0/4294967296.0,1,-nbitq), 
to_sfixed(-872108097.0/4294967296.0,1,-nbitq), 
to_sfixed(84462453.0/4294967296.0,1,-nbitq), 
to_sfixed(-383421872.0/4294967296.0,1,-nbitq), 
to_sfixed(-152178708.0/4294967296.0,1,-nbitq), 
to_sfixed(229536355.0/4294967296.0,1,-nbitq), 
to_sfixed(-419303834.0/4294967296.0,1,-nbitq), 
to_sfixed(-537026208.0/4294967296.0,1,-nbitq), 
to_sfixed(477281885.0/4294967296.0,1,-nbitq), 
to_sfixed(738595125.0/4294967296.0,1,-nbitq), 
to_sfixed(1128878110.0/4294967296.0,1,-nbitq), 
to_sfixed(-465290741.0/4294967296.0,1,-nbitq), 
to_sfixed(-2023875220.0/4294967296.0,1,-nbitq), 
to_sfixed(896359519.0/4294967296.0,1,-nbitq), 
to_sfixed(434955892.0/4294967296.0,1,-nbitq), 
to_sfixed(688013622.0/4294967296.0,1,-nbitq), 
to_sfixed(131844030.0/4294967296.0,1,-nbitq), 
to_sfixed(399577649.0/4294967296.0,1,-nbitq), 
to_sfixed(258261792.0/4294967296.0,1,-nbitq), 
to_sfixed(-841101466.0/4294967296.0,1,-nbitq), 
to_sfixed(-54833648.0/4294967296.0,1,-nbitq), 
to_sfixed(302990274.0/4294967296.0,1,-nbitq), 
to_sfixed(219288986.0/4294967296.0,1,-nbitq), 
to_sfixed(115325302.0/4294967296.0,1,-nbitq), 
to_sfixed(957475689.0/4294967296.0,1,-nbitq), 
to_sfixed(-259758562.0/4294967296.0,1,-nbitq), 
to_sfixed(-109348492.0/4294967296.0,1,-nbitq), 
to_sfixed(854639141.0/4294967296.0,1,-nbitq), 
to_sfixed(716346935.0/4294967296.0,1,-nbitq), 
to_sfixed(517930934.0/4294967296.0,1,-nbitq), 
to_sfixed(-114230486.0/4294967296.0,1,-nbitq), 
to_sfixed(-136885421.0/4294967296.0,1,-nbitq), 
to_sfixed(76220898.0/4294967296.0,1,-nbitq), 
to_sfixed(53884811.0/4294967296.0,1,-nbitq), 
to_sfixed(12290113.0/4294967296.0,1,-nbitq), 
to_sfixed(-357707281.0/4294967296.0,1,-nbitq), 
to_sfixed(584578370.0/4294967296.0,1,-nbitq), 
to_sfixed(146397943.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(196633563.0/4294967296.0,1,-nbitq), 
to_sfixed(-1879884518.0/4294967296.0,1,-nbitq), 
to_sfixed(955188235.0/4294967296.0,1,-nbitq), 
to_sfixed(957751717.0/4294967296.0,1,-nbitq), 
to_sfixed(-928325681.0/4294967296.0,1,-nbitq), 
to_sfixed(-498533793.0/4294967296.0,1,-nbitq), 
to_sfixed(-241266441.0/4294967296.0,1,-nbitq), 
to_sfixed(1083651420.0/4294967296.0,1,-nbitq), 
to_sfixed(99143463.0/4294967296.0,1,-nbitq), 
to_sfixed(-217036482.0/4294967296.0,1,-nbitq), 
to_sfixed(335782864.0/4294967296.0,1,-nbitq), 
to_sfixed(513339597.0/4294967296.0,1,-nbitq), 
to_sfixed(147927712.0/4294967296.0,1,-nbitq), 
to_sfixed(1089990414.0/4294967296.0,1,-nbitq), 
to_sfixed(-26990706.0/4294967296.0,1,-nbitq), 
to_sfixed(432460765.0/4294967296.0,1,-nbitq), 
to_sfixed(322172498.0/4294967296.0,1,-nbitq), 
to_sfixed(-393502889.0/4294967296.0,1,-nbitq), 
to_sfixed(-1868803856.0/4294967296.0,1,-nbitq), 
to_sfixed(-352485628.0/4294967296.0,1,-nbitq), 
to_sfixed(312804588.0/4294967296.0,1,-nbitq), 
to_sfixed(376495113.0/4294967296.0,1,-nbitq), 
to_sfixed(-82818386.0/4294967296.0,1,-nbitq), 
to_sfixed(713205938.0/4294967296.0,1,-nbitq), 
to_sfixed(348540480.0/4294967296.0,1,-nbitq), 
to_sfixed(-147389597.0/4294967296.0,1,-nbitq), 
to_sfixed(44121949.0/4294967296.0,1,-nbitq), 
to_sfixed(-119083220.0/4294967296.0,1,-nbitq), 
to_sfixed(83221445.0/4294967296.0,1,-nbitq), 
to_sfixed(1571672099.0/4294967296.0,1,-nbitq), 
to_sfixed(327733074.0/4294967296.0,1,-nbitq), 
to_sfixed(691535295.0/4294967296.0,1,-nbitq), 
to_sfixed(-1147454352.0/4294967296.0,1,-nbitq), 
to_sfixed(539774999.0/4294967296.0,1,-nbitq), 
to_sfixed(-399275332.0/4294967296.0,1,-nbitq), 
to_sfixed(-399390587.0/4294967296.0,1,-nbitq), 
to_sfixed(-201017436.0/4294967296.0,1,-nbitq), 
to_sfixed(817460273.0/4294967296.0,1,-nbitq), 
to_sfixed(-221698117.0/4294967296.0,1,-nbitq), 
to_sfixed(-32387247.0/4294967296.0,1,-nbitq), 
to_sfixed(6862580.0/4294967296.0,1,-nbitq), 
to_sfixed(56628707.0/4294967296.0,1,-nbitq), 
to_sfixed(-1102524517.0/4294967296.0,1,-nbitq), 
to_sfixed(-922743151.0/4294967296.0,1,-nbitq), 
to_sfixed(309289486.0/4294967296.0,1,-nbitq), 
to_sfixed(-814097430.0/4294967296.0,1,-nbitq), 
to_sfixed(205225011.0/4294967296.0,1,-nbitq), 
to_sfixed(721521545.0/4294967296.0,1,-nbitq), 
to_sfixed(-95263316.0/4294967296.0,1,-nbitq), 
to_sfixed(-1201501931.0/4294967296.0,1,-nbitq), 
to_sfixed(8366469.0/4294967296.0,1,-nbitq), 
to_sfixed(876664242.0/4294967296.0,1,-nbitq), 
to_sfixed(873322566.0/4294967296.0,1,-nbitq), 
to_sfixed(-766706875.0/4294967296.0,1,-nbitq), 
to_sfixed(-1887373026.0/4294967296.0,1,-nbitq), 
to_sfixed(311746685.0/4294967296.0,1,-nbitq), 
to_sfixed(296688189.0/4294967296.0,1,-nbitq), 
to_sfixed(226209826.0/4294967296.0,1,-nbitq), 
to_sfixed(-84998520.0/4294967296.0,1,-nbitq), 
to_sfixed(14639835.0/4294967296.0,1,-nbitq), 
to_sfixed(261195588.0/4294967296.0,1,-nbitq), 
to_sfixed(-414616955.0/4294967296.0,1,-nbitq), 
to_sfixed(90158373.0/4294967296.0,1,-nbitq), 
to_sfixed(946953532.0/4294967296.0,1,-nbitq), 
to_sfixed(402227098.0/4294967296.0,1,-nbitq), 
to_sfixed(-175036395.0/4294967296.0,1,-nbitq), 
to_sfixed(516171701.0/4294967296.0,1,-nbitq), 
to_sfixed(-58690505.0/4294967296.0,1,-nbitq), 
to_sfixed(-3398474.0/4294967296.0,1,-nbitq), 
to_sfixed(885258928.0/4294967296.0,1,-nbitq), 
to_sfixed(-86171055.0/4294967296.0,1,-nbitq), 
to_sfixed(124309319.0/4294967296.0,1,-nbitq), 
to_sfixed(-602300926.0/4294967296.0,1,-nbitq), 
to_sfixed(-115268490.0/4294967296.0,1,-nbitq), 
to_sfixed(-48352554.0/4294967296.0,1,-nbitq), 
to_sfixed(255940463.0/4294967296.0,1,-nbitq), 
to_sfixed(1400228431.0/4294967296.0,1,-nbitq), 
to_sfixed(250152471.0/4294967296.0,1,-nbitq), 
to_sfixed(-177708941.0/4294967296.0,1,-nbitq), 
to_sfixed(84822916.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-150146195.0/4294967296.0,1,-nbitq), 
to_sfixed(-1399070609.0/4294967296.0,1,-nbitq), 
to_sfixed(124963622.0/4294967296.0,1,-nbitq), 
to_sfixed(314431375.0/4294967296.0,1,-nbitq), 
to_sfixed(-607174258.0/4294967296.0,1,-nbitq), 
to_sfixed(-240013773.0/4294967296.0,1,-nbitq), 
to_sfixed(-114230025.0/4294967296.0,1,-nbitq), 
to_sfixed(717705852.0/4294967296.0,1,-nbitq), 
to_sfixed(68010263.0/4294967296.0,1,-nbitq), 
to_sfixed(312275898.0/4294967296.0,1,-nbitq), 
to_sfixed(-78177593.0/4294967296.0,1,-nbitq), 
to_sfixed(799893079.0/4294967296.0,1,-nbitq), 
to_sfixed(112745755.0/4294967296.0,1,-nbitq), 
to_sfixed(443370487.0/4294967296.0,1,-nbitq), 
to_sfixed(-134572780.0/4294967296.0,1,-nbitq), 
to_sfixed(1075787.0/4294967296.0,1,-nbitq), 
to_sfixed(67098886.0/4294967296.0,1,-nbitq), 
to_sfixed(-87598957.0/4294967296.0,1,-nbitq), 
to_sfixed(-743625647.0/4294967296.0,1,-nbitq), 
to_sfixed(231009254.0/4294967296.0,1,-nbitq), 
to_sfixed(53917945.0/4294967296.0,1,-nbitq), 
to_sfixed(476446702.0/4294967296.0,1,-nbitq), 
to_sfixed(-476721765.0/4294967296.0,1,-nbitq), 
to_sfixed(-556739656.0/4294967296.0,1,-nbitq), 
to_sfixed(-242967493.0/4294967296.0,1,-nbitq), 
to_sfixed(-626736957.0/4294967296.0,1,-nbitq), 
to_sfixed(-579920129.0/4294967296.0,1,-nbitq), 
to_sfixed(60966570.0/4294967296.0,1,-nbitq), 
to_sfixed(-634093119.0/4294967296.0,1,-nbitq), 
to_sfixed(1420035150.0/4294967296.0,1,-nbitq), 
to_sfixed(150090440.0/4294967296.0,1,-nbitq), 
to_sfixed(396280097.0/4294967296.0,1,-nbitq), 
to_sfixed(-940234699.0/4294967296.0,1,-nbitq), 
to_sfixed(383585707.0/4294967296.0,1,-nbitq), 
to_sfixed(-493714310.0/4294967296.0,1,-nbitq), 
to_sfixed(105345701.0/4294967296.0,1,-nbitq), 
to_sfixed(79284554.0/4294967296.0,1,-nbitq), 
to_sfixed(373698910.0/4294967296.0,1,-nbitq), 
to_sfixed(244928697.0/4294967296.0,1,-nbitq), 
to_sfixed(-269559973.0/4294967296.0,1,-nbitq), 
to_sfixed(228363158.0/4294967296.0,1,-nbitq), 
to_sfixed(-142441377.0/4294967296.0,1,-nbitq), 
to_sfixed(-1129972874.0/4294967296.0,1,-nbitq), 
to_sfixed(-1016206088.0/4294967296.0,1,-nbitq), 
to_sfixed(609784413.0/4294967296.0,1,-nbitq), 
to_sfixed(4335509.0/4294967296.0,1,-nbitq), 
to_sfixed(151552980.0/4294967296.0,1,-nbitq), 
to_sfixed(107461523.0/4294967296.0,1,-nbitq), 
to_sfixed(167181229.0/4294967296.0,1,-nbitq), 
to_sfixed(-648171653.0/4294967296.0,1,-nbitq), 
to_sfixed(528748192.0/4294967296.0,1,-nbitq), 
to_sfixed(837370268.0/4294967296.0,1,-nbitq), 
to_sfixed(72341610.0/4294967296.0,1,-nbitq), 
to_sfixed(-739682762.0/4294967296.0,1,-nbitq), 
to_sfixed(-1727618914.0/4294967296.0,1,-nbitq), 
to_sfixed(208949327.0/4294967296.0,1,-nbitq), 
to_sfixed(-37513043.0/4294967296.0,1,-nbitq), 
to_sfixed(395153287.0/4294967296.0,1,-nbitq), 
to_sfixed(-66009696.0/4294967296.0,1,-nbitq), 
to_sfixed(-184854068.0/4294967296.0,1,-nbitq), 
to_sfixed(184329184.0/4294967296.0,1,-nbitq), 
to_sfixed(-5125864.0/4294967296.0,1,-nbitq), 
to_sfixed(56962051.0/4294967296.0,1,-nbitq), 
to_sfixed(649240950.0/4294967296.0,1,-nbitq), 
to_sfixed(404718202.0/4294967296.0,1,-nbitq), 
to_sfixed(-70576022.0/4294967296.0,1,-nbitq), 
to_sfixed(121921836.0/4294967296.0,1,-nbitq), 
to_sfixed(-318491036.0/4294967296.0,1,-nbitq), 
to_sfixed(21541753.0/4294967296.0,1,-nbitq), 
to_sfixed(1025812032.0/4294967296.0,1,-nbitq), 
to_sfixed(-128501974.0/4294967296.0,1,-nbitq), 
to_sfixed(-14629854.0/4294967296.0,1,-nbitq), 
to_sfixed(-14227858.0/4294967296.0,1,-nbitq), 
to_sfixed(-62831339.0/4294967296.0,1,-nbitq), 
to_sfixed(277683258.0/4294967296.0,1,-nbitq), 
to_sfixed(57425931.0/4294967296.0,1,-nbitq), 
to_sfixed(35234634.0/4294967296.0,1,-nbitq), 
to_sfixed(-67995508.0/4294967296.0,1,-nbitq), 
to_sfixed(68974744.0/4294967296.0,1,-nbitq), 
to_sfixed(307202847.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(397246071.0/4294967296.0,1,-nbitq), 
to_sfixed(-25451785.0/4294967296.0,1,-nbitq), 
to_sfixed(453173440.0/4294967296.0,1,-nbitq), 
to_sfixed(-143701199.0/4294967296.0,1,-nbitq), 
to_sfixed(-184801298.0/4294967296.0,1,-nbitq), 
to_sfixed(-708249537.0/4294967296.0,1,-nbitq), 
to_sfixed(276204488.0/4294967296.0,1,-nbitq), 
to_sfixed(800828342.0/4294967296.0,1,-nbitq), 
to_sfixed(-219184136.0/4294967296.0,1,-nbitq), 
to_sfixed(24290473.0/4294967296.0,1,-nbitq), 
to_sfixed(327755807.0/4294967296.0,1,-nbitq), 
to_sfixed(183699117.0/4294967296.0,1,-nbitq), 
to_sfixed(-56973520.0/4294967296.0,1,-nbitq), 
to_sfixed(732644374.0/4294967296.0,1,-nbitq), 
to_sfixed(361826934.0/4294967296.0,1,-nbitq), 
to_sfixed(83993755.0/4294967296.0,1,-nbitq), 
to_sfixed(18607893.0/4294967296.0,1,-nbitq), 
to_sfixed(-229605568.0/4294967296.0,1,-nbitq), 
to_sfixed(-9969500.0/4294967296.0,1,-nbitq), 
to_sfixed(-146857595.0/4294967296.0,1,-nbitq), 
to_sfixed(-346979643.0/4294967296.0,1,-nbitq), 
to_sfixed(260422325.0/4294967296.0,1,-nbitq), 
to_sfixed(1012837.0/4294967296.0,1,-nbitq), 
to_sfixed(399632448.0/4294967296.0,1,-nbitq), 
to_sfixed(-243205599.0/4294967296.0,1,-nbitq), 
to_sfixed(-571850064.0/4294967296.0,1,-nbitq), 
to_sfixed(355383191.0/4294967296.0,1,-nbitq), 
to_sfixed(127924843.0/4294967296.0,1,-nbitq), 
to_sfixed(301214262.0/4294967296.0,1,-nbitq), 
to_sfixed(1041085792.0/4294967296.0,1,-nbitq), 
to_sfixed(67497309.0/4294967296.0,1,-nbitq), 
to_sfixed(56552818.0/4294967296.0,1,-nbitq), 
to_sfixed(-285106780.0/4294967296.0,1,-nbitq), 
to_sfixed(-124720835.0/4294967296.0,1,-nbitq), 
to_sfixed(-461060250.0/4294967296.0,1,-nbitq), 
to_sfixed(-525761909.0/4294967296.0,1,-nbitq), 
to_sfixed(145962905.0/4294967296.0,1,-nbitq), 
to_sfixed(-97632898.0/4294967296.0,1,-nbitq), 
to_sfixed(-76311922.0/4294967296.0,1,-nbitq), 
to_sfixed(421908496.0/4294967296.0,1,-nbitq), 
to_sfixed(46444326.0/4294967296.0,1,-nbitq), 
to_sfixed(-239315848.0/4294967296.0,1,-nbitq), 
to_sfixed(-246045830.0/4294967296.0,1,-nbitq), 
to_sfixed(-1044535999.0/4294967296.0,1,-nbitq), 
to_sfixed(135661363.0/4294967296.0,1,-nbitq), 
to_sfixed(-641361924.0/4294967296.0,1,-nbitq), 
to_sfixed(-328107576.0/4294967296.0,1,-nbitq), 
to_sfixed(-199048145.0/4294967296.0,1,-nbitq), 
to_sfixed(76042774.0/4294967296.0,1,-nbitq), 
to_sfixed(-421253523.0/4294967296.0,1,-nbitq), 
to_sfixed(294984023.0/4294967296.0,1,-nbitq), 
to_sfixed(114369867.0/4294967296.0,1,-nbitq), 
to_sfixed(363206614.0/4294967296.0,1,-nbitq), 
to_sfixed(35052379.0/4294967296.0,1,-nbitq), 
to_sfixed(-670818525.0/4294967296.0,1,-nbitq), 
to_sfixed(60580800.0/4294967296.0,1,-nbitq), 
to_sfixed(-39147868.0/4294967296.0,1,-nbitq), 
to_sfixed(295099859.0/4294967296.0,1,-nbitq), 
to_sfixed(-231557789.0/4294967296.0,1,-nbitq), 
to_sfixed(-52468362.0/4294967296.0,1,-nbitq), 
to_sfixed(207855393.0/4294967296.0,1,-nbitq), 
to_sfixed(-264643415.0/4294967296.0,1,-nbitq), 
to_sfixed(476748812.0/4294967296.0,1,-nbitq), 
to_sfixed(-41380671.0/4294967296.0,1,-nbitq), 
to_sfixed(93453902.0/4294967296.0,1,-nbitq), 
to_sfixed(-224934754.0/4294967296.0,1,-nbitq), 
to_sfixed(170408370.0/4294967296.0,1,-nbitq), 
to_sfixed(122677211.0/4294967296.0,1,-nbitq), 
to_sfixed(-14682801.0/4294967296.0,1,-nbitq), 
to_sfixed(124150704.0/4294967296.0,1,-nbitq), 
to_sfixed(-487061963.0/4294967296.0,1,-nbitq), 
to_sfixed(205659552.0/4294967296.0,1,-nbitq), 
to_sfixed(396570216.0/4294967296.0,1,-nbitq), 
to_sfixed(440831774.0/4294967296.0,1,-nbitq), 
to_sfixed(127041457.0/4294967296.0,1,-nbitq), 
to_sfixed(-70664917.0/4294967296.0,1,-nbitq), 
to_sfixed(-337062356.0/4294967296.0,1,-nbitq), 
to_sfixed(-178599722.0/4294967296.0,1,-nbitq), 
to_sfixed(172721475.0/4294967296.0,1,-nbitq), 
to_sfixed(-31796081.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-31707908.0/4294967296.0,1,-nbitq), 
to_sfixed(-39501649.0/4294967296.0,1,-nbitq), 
to_sfixed(664475112.0/4294967296.0,1,-nbitq), 
to_sfixed(-218692294.0/4294967296.0,1,-nbitq), 
to_sfixed(-331872035.0/4294967296.0,1,-nbitq), 
to_sfixed(-740923740.0/4294967296.0,1,-nbitq), 
to_sfixed(254469101.0/4294967296.0,1,-nbitq), 
to_sfixed(14530363.0/4294967296.0,1,-nbitq), 
to_sfixed(-322378542.0/4294967296.0,1,-nbitq), 
to_sfixed(382099141.0/4294967296.0,1,-nbitq), 
to_sfixed(487917095.0/4294967296.0,1,-nbitq), 
to_sfixed(61501950.0/4294967296.0,1,-nbitq), 
to_sfixed(-240032049.0/4294967296.0,1,-nbitq), 
to_sfixed(527160181.0/4294967296.0,1,-nbitq), 
to_sfixed(171814171.0/4294967296.0,1,-nbitq), 
to_sfixed(410381220.0/4294967296.0,1,-nbitq), 
to_sfixed(-229217546.0/4294967296.0,1,-nbitq), 
to_sfixed(-29690929.0/4294967296.0,1,-nbitq), 
to_sfixed(-191251109.0/4294967296.0,1,-nbitq), 
to_sfixed(-306208124.0/4294967296.0,1,-nbitq), 
to_sfixed(-29792271.0/4294967296.0,1,-nbitq), 
to_sfixed(-26363871.0/4294967296.0,1,-nbitq), 
to_sfixed(-538504450.0/4294967296.0,1,-nbitq), 
to_sfixed(419440359.0/4294967296.0,1,-nbitq), 
to_sfixed(379031307.0/4294967296.0,1,-nbitq), 
to_sfixed(-633792527.0/4294967296.0,1,-nbitq), 
to_sfixed(53555541.0/4294967296.0,1,-nbitq), 
to_sfixed(-239397386.0/4294967296.0,1,-nbitq), 
to_sfixed(355658602.0/4294967296.0,1,-nbitq), 
to_sfixed(-14625325.0/4294967296.0,1,-nbitq), 
to_sfixed(-552497522.0/4294967296.0,1,-nbitq), 
to_sfixed(-295882183.0/4294967296.0,1,-nbitq), 
to_sfixed(65238746.0/4294967296.0,1,-nbitq), 
to_sfixed(243796725.0/4294967296.0,1,-nbitq), 
to_sfixed(-307566034.0/4294967296.0,1,-nbitq), 
to_sfixed(-190009769.0/4294967296.0,1,-nbitq), 
to_sfixed(121129468.0/4294967296.0,1,-nbitq), 
to_sfixed(-132298187.0/4294967296.0,1,-nbitq), 
to_sfixed(141702626.0/4294967296.0,1,-nbitq), 
to_sfixed(432573844.0/4294967296.0,1,-nbitq), 
to_sfixed(-75333067.0/4294967296.0,1,-nbitq), 
to_sfixed(172818064.0/4294967296.0,1,-nbitq), 
to_sfixed(-320640395.0/4294967296.0,1,-nbitq), 
to_sfixed(-595222757.0/4294967296.0,1,-nbitq), 
to_sfixed(-76231241.0/4294967296.0,1,-nbitq), 
to_sfixed(-371813128.0/4294967296.0,1,-nbitq), 
to_sfixed(-212306484.0/4294967296.0,1,-nbitq), 
to_sfixed(261836814.0/4294967296.0,1,-nbitq), 
to_sfixed(-414172727.0/4294967296.0,1,-nbitq), 
to_sfixed(212378999.0/4294967296.0,1,-nbitq), 
to_sfixed(253467673.0/4294967296.0,1,-nbitq), 
to_sfixed(60352862.0/4294967296.0,1,-nbitq), 
to_sfixed(8148112.0/4294967296.0,1,-nbitq), 
to_sfixed(26528127.0/4294967296.0,1,-nbitq), 
to_sfixed(-382819836.0/4294967296.0,1,-nbitq), 
to_sfixed(101037595.0/4294967296.0,1,-nbitq), 
to_sfixed(484785218.0/4294967296.0,1,-nbitq), 
to_sfixed(280421895.0/4294967296.0,1,-nbitq), 
to_sfixed(-263936342.0/4294967296.0,1,-nbitq), 
to_sfixed(-197544711.0/4294967296.0,1,-nbitq), 
to_sfixed(166613834.0/4294967296.0,1,-nbitq), 
to_sfixed(329731873.0/4294967296.0,1,-nbitq), 
to_sfixed(-141648125.0/4294967296.0,1,-nbitq), 
to_sfixed(-138859965.0/4294967296.0,1,-nbitq), 
to_sfixed(56315023.0/4294967296.0,1,-nbitq), 
to_sfixed(-331961266.0/4294967296.0,1,-nbitq), 
to_sfixed(257834889.0/4294967296.0,1,-nbitq), 
to_sfixed(1315596.0/4294967296.0,1,-nbitq), 
to_sfixed(325354785.0/4294967296.0,1,-nbitq), 
to_sfixed(82460227.0/4294967296.0,1,-nbitq), 
to_sfixed(126806765.0/4294967296.0,1,-nbitq), 
to_sfixed(181823622.0/4294967296.0,1,-nbitq), 
to_sfixed(419130444.0/4294967296.0,1,-nbitq), 
to_sfixed(144399253.0/4294967296.0,1,-nbitq), 
to_sfixed(325788846.0/4294967296.0,1,-nbitq), 
to_sfixed(75396721.0/4294967296.0,1,-nbitq), 
to_sfixed(49844030.0/4294967296.0,1,-nbitq), 
to_sfixed(-284128107.0/4294967296.0,1,-nbitq), 
to_sfixed(-235910439.0/4294967296.0,1,-nbitq), 
to_sfixed(-374650898.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-358098391.0/4294967296.0,1,-nbitq), 
to_sfixed(94645196.0/4294967296.0,1,-nbitq), 
to_sfixed(523335069.0/4294967296.0,1,-nbitq), 
to_sfixed(-623391489.0/4294967296.0,1,-nbitq), 
to_sfixed(113174163.0/4294967296.0,1,-nbitq), 
to_sfixed(70762644.0/4294967296.0,1,-nbitq), 
to_sfixed(235593170.0/4294967296.0,1,-nbitq), 
to_sfixed(-5695914.0/4294967296.0,1,-nbitq), 
to_sfixed(-369587236.0/4294967296.0,1,-nbitq), 
to_sfixed(439131393.0/4294967296.0,1,-nbitq), 
to_sfixed(480979763.0/4294967296.0,1,-nbitq), 
to_sfixed(192453435.0/4294967296.0,1,-nbitq), 
to_sfixed(312521421.0/4294967296.0,1,-nbitq), 
to_sfixed(353370167.0/4294967296.0,1,-nbitq), 
to_sfixed(229162689.0/4294967296.0,1,-nbitq), 
to_sfixed(137895133.0/4294967296.0,1,-nbitq), 
to_sfixed(153239840.0/4294967296.0,1,-nbitq), 
to_sfixed(248952773.0/4294967296.0,1,-nbitq), 
to_sfixed(370123400.0/4294967296.0,1,-nbitq), 
to_sfixed(86361484.0/4294967296.0,1,-nbitq), 
to_sfixed(283012640.0/4294967296.0,1,-nbitq), 
to_sfixed(173999532.0/4294967296.0,1,-nbitq), 
to_sfixed(284245813.0/4294967296.0,1,-nbitq), 
to_sfixed(132896419.0/4294967296.0,1,-nbitq), 
to_sfixed(410785058.0/4294967296.0,1,-nbitq), 
to_sfixed(253115524.0/4294967296.0,1,-nbitq), 
to_sfixed(-160238142.0/4294967296.0,1,-nbitq), 
to_sfixed(33301624.0/4294967296.0,1,-nbitq), 
to_sfixed(232329341.0/4294967296.0,1,-nbitq), 
to_sfixed(3882946.0/4294967296.0,1,-nbitq), 
to_sfixed(-212136780.0/4294967296.0,1,-nbitq), 
to_sfixed(52346663.0/4294967296.0,1,-nbitq), 
to_sfixed(-20962514.0/4294967296.0,1,-nbitq), 
to_sfixed(257315794.0/4294967296.0,1,-nbitq), 
to_sfixed(-357812795.0/4294967296.0,1,-nbitq), 
to_sfixed(-4308407.0/4294967296.0,1,-nbitq), 
to_sfixed(188610904.0/4294967296.0,1,-nbitq), 
to_sfixed(-436902727.0/4294967296.0,1,-nbitq), 
to_sfixed(-4052455.0/4294967296.0,1,-nbitq), 
to_sfixed(-228442157.0/4294967296.0,1,-nbitq), 
to_sfixed(-54251209.0/4294967296.0,1,-nbitq), 
to_sfixed(-386410190.0/4294967296.0,1,-nbitq), 
to_sfixed(-14012533.0/4294967296.0,1,-nbitq), 
to_sfixed(-426665829.0/4294967296.0,1,-nbitq), 
to_sfixed(263801158.0/4294967296.0,1,-nbitq), 
to_sfixed(-370745895.0/4294967296.0,1,-nbitq), 
to_sfixed(293086780.0/4294967296.0,1,-nbitq), 
to_sfixed(-401331944.0/4294967296.0,1,-nbitq), 
to_sfixed(334591528.0/4294967296.0,1,-nbitq), 
to_sfixed(325049591.0/4294967296.0,1,-nbitq), 
to_sfixed(45965588.0/4294967296.0,1,-nbitq), 
to_sfixed(-43288581.0/4294967296.0,1,-nbitq), 
to_sfixed(115486908.0/4294967296.0,1,-nbitq), 
to_sfixed(-136963866.0/4294967296.0,1,-nbitq), 
to_sfixed(-221594316.0/4294967296.0,1,-nbitq), 
to_sfixed(-383967638.0/4294967296.0,1,-nbitq), 
to_sfixed(499320394.0/4294967296.0,1,-nbitq), 
to_sfixed(-46916369.0/4294967296.0,1,-nbitq), 
to_sfixed(166541354.0/4294967296.0,1,-nbitq), 
to_sfixed(409654566.0/4294967296.0,1,-nbitq), 
to_sfixed(50637668.0/4294967296.0,1,-nbitq), 
to_sfixed(281826102.0/4294967296.0,1,-nbitq), 
to_sfixed(92696998.0/4294967296.0,1,-nbitq), 
to_sfixed(76304248.0/4294967296.0,1,-nbitq), 
to_sfixed(155747730.0/4294967296.0,1,-nbitq), 
to_sfixed(84020300.0/4294967296.0,1,-nbitq), 
to_sfixed(562884517.0/4294967296.0,1,-nbitq), 
to_sfixed(295678076.0/4294967296.0,1,-nbitq), 
to_sfixed(-207833102.0/4294967296.0,1,-nbitq), 
to_sfixed(-232315176.0/4294967296.0,1,-nbitq), 
to_sfixed(198220456.0/4294967296.0,1,-nbitq), 
to_sfixed(44175707.0/4294967296.0,1,-nbitq), 
to_sfixed(273480346.0/4294967296.0,1,-nbitq), 
to_sfixed(221274994.0/4294967296.0,1,-nbitq), 
to_sfixed(-185021537.0/4294967296.0,1,-nbitq), 
to_sfixed(36524181.0/4294967296.0,1,-nbitq), 
to_sfixed(88531125.0/4294967296.0,1,-nbitq), 
to_sfixed(149129308.0/4294967296.0,1,-nbitq), 
to_sfixed(18050039.0/4294967296.0,1,-nbitq), 
to_sfixed(-314987364.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-274837755.0/4294967296.0,1,-nbitq), 
to_sfixed(-137686086.0/4294967296.0,1,-nbitq), 
to_sfixed(-283581255.0/4294967296.0,1,-nbitq), 
to_sfixed(-368045311.0/4294967296.0,1,-nbitq), 
to_sfixed(184977542.0/4294967296.0,1,-nbitq), 
to_sfixed(309395882.0/4294967296.0,1,-nbitq), 
to_sfixed(230658496.0/4294967296.0,1,-nbitq), 
to_sfixed(-376227499.0/4294967296.0,1,-nbitq), 
to_sfixed(-267465745.0/4294967296.0,1,-nbitq), 
to_sfixed(12164826.0/4294967296.0,1,-nbitq), 
to_sfixed(-287037921.0/4294967296.0,1,-nbitq), 
to_sfixed(412495778.0/4294967296.0,1,-nbitq), 
to_sfixed(-298057413.0/4294967296.0,1,-nbitq), 
to_sfixed(78692174.0/4294967296.0,1,-nbitq), 
to_sfixed(-291464285.0/4294967296.0,1,-nbitq), 
to_sfixed(-198918461.0/4294967296.0,1,-nbitq), 
to_sfixed(184167875.0/4294967296.0,1,-nbitq), 
to_sfixed(-300213136.0/4294967296.0,1,-nbitq), 
to_sfixed(95088637.0/4294967296.0,1,-nbitq), 
to_sfixed(-37512491.0/4294967296.0,1,-nbitq), 
to_sfixed(241967178.0/4294967296.0,1,-nbitq), 
to_sfixed(42361933.0/4294967296.0,1,-nbitq), 
to_sfixed(179444559.0/4294967296.0,1,-nbitq), 
to_sfixed(460211737.0/4294967296.0,1,-nbitq), 
to_sfixed(47775295.0/4294967296.0,1,-nbitq), 
to_sfixed(151485760.0/4294967296.0,1,-nbitq), 
to_sfixed(-127711072.0/4294967296.0,1,-nbitq), 
to_sfixed(114564433.0/4294967296.0,1,-nbitq), 
to_sfixed(3086548.0/4294967296.0,1,-nbitq), 
to_sfixed(104134666.0/4294967296.0,1,-nbitq), 
to_sfixed(-18976260.0/4294967296.0,1,-nbitq), 
to_sfixed(279062499.0/4294967296.0,1,-nbitq), 
to_sfixed(421033374.0/4294967296.0,1,-nbitq), 
to_sfixed(-166236752.0/4294967296.0,1,-nbitq), 
to_sfixed(301543722.0/4294967296.0,1,-nbitq), 
to_sfixed(-190668951.0/4294967296.0,1,-nbitq), 
to_sfixed(268825109.0/4294967296.0,1,-nbitq), 
to_sfixed(408194559.0/4294967296.0,1,-nbitq), 
to_sfixed(-39648983.0/4294967296.0,1,-nbitq), 
to_sfixed(-111887431.0/4294967296.0,1,-nbitq), 
to_sfixed(-2502971.0/4294967296.0,1,-nbitq), 
to_sfixed(-80905442.0/4294967296.0,1,-nbitq), 
to_sfixed(1405545.0/4294967296.0,1,-nbitq), 
to_sfixed(-216669667.0/4294967296.0,1,-nbitq), 
to_sfixed(-88417303.0/4294967296.0,1,-nbitq), 
to_sfixed(447530065.0/4294967296.0,1,-nbitq), 
to_sfixed(262137198.0/4294967296.0,1,-nbitq), 
to_sfixed(-167381130.0/4294967296.0,1,-nbitq), 
to_sfixed(305998576.0/4294967296.0,1,-nbitq), 
to_sfixed(227025369.0/4294967296.0,1,-nbitq), 
to_sfixed(-250683493.0/4294967296.0,1,-nbitq), 
to_sfixed(17143619.0/4294967296.0,1,-nbitq), 
to_sfixed(-535063150.0/4294967296.0,1,-nbitq), 
to_sfixed(-130909055.0/4294967296.0,1,-nbitq), 
to_sfixed(-121776097.0/4294967296.0,1,-nbitq), 
to_sfixed(323808965.0/4294967296.0,1,-nbitq), 
to_sfixed(396181385.0/4294967296.0,1,-nbitq), 
to_sfixed(-85124330.0/4294967296.0,1,-nbitq), 
to_sfixed(399232694.0/4294967296.0,1,-nbitq), 
to_sfixed(286846930.0/4294967296.0,1,-nbitq), 
to_sfixed(-364813089.0/4294967296.0,1,-nbitq), 
to_sfixed(471938775.0/4294967296.0,1,-nbitq), 
to_sfixed(-255699844.0/4294967296.0,1,-nbitq), 
to_sfixed(89562399.0/4294967296.0,1,-nbitq), 
to_sfixed(208701119.0/4294967296.0,1,-nbitq), 
to_sfixed(8705556.0/4294967296.0,1,-nbitq), 
to_sfixed(317283260.0/4294967296.0,1,-nbitq), 
to_sfixed(-393593272.0/4294967296.0,1,-nbitq), 
to_sfixed(-289287158.0/4294967296.0,1,-nbitq), 
to_sfixed(331289706.0/4294967296.0,1,-nbitq), 
to_sfixed(4098067.0/4294967296.0,1,-nbitq), 
to_sfixed(-236256593.0/4294967296.0,1,-nbitq), 
to_sfixed(-59065994.0/4294967296.0,1,-nbitq), 
to_sfixed(443979372.0/4294967296.0,1,-nbitq), 
to_sfixed(270644932.0/4294967296.0,1,-nbitq), 
to_sfixed(-328562205.0/4294967296.0,1,-nbitq), 
to_sfixed(-184537509.0/4294967296.0,1,-nbitq), 
to_sfixed(-235819784.0/4294967296.0,1,-nbitq), 
to_sfixed(-225106060.0/4294967296.0,1,-nbitq), 
to_sfixed(-100113762.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-433821936.0/4294967296.0,1,-nbitq), 
to_sfixed(-40374104.0/4294967296.0,1,-nbitq), 
to_sfixed(-235246696.0/4294967296.0,1,-nbitq), 
to_sfixed(228031490.0/4294967296.0,1,-nbitq), 
to_sfixed(467204414.0/4294967296.0,1,-nbitq), 
to_sfixed(217391500.0/4294967296.0,1,-nbitq), 
to_sfixed(-64491084.0/4294967296.0,1,-nbitq), 
to_sfixed(173666884.0/4294967296.0,1,-nbitq), 
to_sfixed(-193269822.0/4294967296.0,1,-nbitq), 
to_sfixed(-322134776.0/4294967296.0,1,-nbitq), 
to_sfixed(-216737087.0/4294967296.0,1,-nbitq), 
to_sfixed(50062675.0/4294967296.0,1,-nbitq), 
to_sfixed(-80467022.0/4294967296.0,1,-nbitq), 
to_sfixed(-41831937.0/4294967296.0,1,-nbitq), 
to_sfixed(-213462866.0/4294967296.0,1,-nbitq), 
to_sfixed(282349595.0/4294967296.0,1,-nbitq), 
to_sfixed(82200792.0/4294967296.0,1,-nbitq), 
to_sfixed(-376686968.0/4294967296.0,1,-nbitq), 
to_sfixed(-98514849.0/4294967296.0,1,-nbitq), 
to_sfixed(306055771.0/4294967296.0,1,-nbitq), 
to_sfixed(-271287777.0/4294967296.0,1,-nbitq), 
to_sfixed(120907424.0/4294967296.0,1,-nbitq), 
to_sfixed(156255373.0/4294967296.0,1,-nbitq), 
to_sfixed(309677930.0/4294967296.0,1,-nbitq), 
to_sfixed(49129793.0/4294967296.0,1,-nbitq), 
to_sfixed(458699268.0/4294967296.0,1,-nbitq), 
to_sfixed(288540738.0/4294967296.0,1,-nbitq), 
to_sfixed(-421286664.0/4294967296.0,1,-nbitq), 
to_sfixed(467966912.0/4294967296.0,1,-nbitq), 
to_sfixed(46217274.0/4294967296.0,1,-nbitq), 
to_sfixed(-531347390.0/4294967296.0,1,-nbitq), 
to_sfixed(-221743018.0/4294967296.0,1,-nbitq), 
to_sfixed(-98340546.0/4294967296.0,1,-nbitq), 
to_sfixed(-92524941.0/4294967296.0,1,-nbitq), 
to_sfixed(350627946.0/4294967296.0,1,-nbitq), 
to_sfixed(-138182773.0/4294967296.0,1,-nbitq), 
to_sfixed(258897954.0/4294967296.0,1,-nbitq), 
to_sfixed(465110927.0/4294967296.0,1,-nbitq), 
to_sfixed(-99670595.0/4294967296.0,1,-nbitq), 
to_sfixed(309441399.0/4294967296.0,1,-nbitq), 
to_sfixed(157799614.0/4294967296.0,1,-nbitq), 
to_sfixed(153917865.0/4294967296.0,1,-nbitq), 
to_sfixed(79854937.0/4294967296.0,1,-nbitq), 
to_sfixed(78013001.0/4294967296.0,1,-nbitq), 
to_sfixed(190580167.0/4294967296.0,1,-nbitq), 
to_sfixed(312392436.0/4294967296.0,1,-nbitq), 
to_sfixed(-106628918.0/4294967296.0,1,-nbitq), 
to_sfixed(-106407109.0/4294967296.0,1,-nbitq), 
to_sfixed(-91786145.0/4294967296.0,1,-nbitq), 
to_sfixed(114867982.0/4294967296.0,1,-nbitq), 
to_sfixed(402036734.0/4294967296.0,1,-nbitq), 
to_sfixed(-85229469.0/4294967296.0,1,-nbitq), 
to_sfixed(-252807451.0/4294967296.0,1,-nbitq), 
to_sfixed(-162911303.0/4294967296.0,1,-nbitq), 
to_sfixed(320103019.0/4294967296.0,1,-nbitq), 
to_sfixed(-232383552.0/4294967296.0,1,-nbitq), 
to_sfixed(112160279.0/4294967296.0,1,-nbitq), 
to_sfixed(114545579.0/4294967296.0,1,-nbitq), 
to_sfixed(381216426.0/4294967296.0,1,-nbitq), 
to_sfixed(351538578.0/4294967296.0,1,-nbitq), 
to_sfixed(333164493.0/4294967296.0,1,-nbitq), 
to_sfixed(81504881.0/4294967296.0,1,-nbitq), 
to_sfixed(-26646207.0/4294967296.0,1,-nbitq), 
to_sfixed(432936606.0/4294967296.0,1,-nbitq), 
to_sfixed(12285063.0/4294967296.0,1,-nbitq), 
to_sfixed(-327324056.0/4294967296.0,1,-nbitq), 
to_sfixed(263400825.0/4294967296.0,1,-nbitq), 
to_sfixed(-53912811.0/4294967296.0,1,-nbitq), 
to_sfixed(60915719.0/4294967296.0,1,-nbitq), 
to_sfixed(26390830.0/4294967296.0,1,-nbitq), 
to_sfixed(31249405.0/4294967296.0,1,-nbitq), 
to_sfixed(33110109.0/4294967296.0,1,-nbitq), 
to_sfixed(-480823426.0/4294967296.0,1,-nbitq), 
to_sfixed(-307259679.0/4294967296.0,1,-nbitq), 
to_sfixed(240639989.0/4294967296.0,1,-nbitq), 
to_sfixed(-118402714.0/4294967296.0,1,-nbitq), 
to_sfixed(-268748963.0/4294967296.0,1,-nbitq), 
to_sfixed(-410970668.0/4294967296.0,1,-nbitq), 
to_sfixed(146667930.0/4294967296.0,1,-nbitq), 
to_sfixed(115904415.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-3518145.0/4294967296.0,1,-nbitq), 
to_sfixed(124388105.0/4294967296.0,1,-nbitq), 
to_sfixed(-33926235.0/4294967296.0,1,-nbitq), 
to_sfixed(-257140789.0/4294967296.0,1,-nbitq), 
to_sfixed(316854306.0/4294967296.0,1,-nbitq), 
to_sfixed(-136862829.0/4294967296.0,1,-nbitq), 
to_sfixed(141676157.0/4294967296.0,1,-nbitq), 
to_sfixed(251411309.0/4294967296.0,1,-nbitq), 
to_sfixed(151906180.0/4294967296.0,1,-nbitq), 
to_sfixed(431013906.0/4294967296.0,1,-nbitq), 
to_sfixed(-361459978.0/4294967296.0,1,-nbitq), 
to_sfixed(-185867826.0/4294967296.0,1,-nbitq), 
to_sfixed(-78718184.0/4294967296.0,1,-nbitq), 
to_sfixed(23497433.0/4294967296.0,1,-nbitq), 
to_sfixed(90437950.0/4294967296.0,1,-nbitq), 
to_sfixed(36360948.0/4294967296.0,1,-nbitq), 
to_sfixed(-308375301.0/4294967296.0,1,-nbitq), 
to_sfixed(-342800676.0/4294967296.0,1,-nbitq), 
to_sfixed(-268748116.0/4294967296.0,1,-nbitq), 
to_sfixed(-69636235.0/4294967296.0,1,-nbitq), 
to_sfixed(306256024.0/4294967296.0,1,-nbitq), 
to_sfixed(53005021.0/4294967296.0,1,-nbitq), 
to_sfixed(-226250993.0/4294967296.0,1,-nbitq), 
to_sfixed(-110592220.0/4294967296.0,1,-nbitq), 
to_sfixed(198760494.0/4294967296.0,1,-nbitq), 
to_sfixed(-108212020.0/4294967296.0,1,-nbitq), 
to_sfixed(-140898114.0/4294967296.0,1,-nbitq), 
to_sfixed(-639900193.0/4294967296.0,1,-nbitq), 
to_sfixed(389796170.0/4294967296.0,1,-nbitq), 
to_sfixed(8864384.0/4294967296.0,1,-nbitq), 
to_sfixed(-105716109.0/4294967296.0,1,-nbitq), 
to_sfixed(102596571.0/4294967296.0,1,-nbitq), 
to_sfixed(-280346235.0/4294967296.0,1,-nbitq), 
to_sfixed(-386318619.0/4294967296.0,1,-nbitq), 
to_sfixed(534455513.0/4294967296.0,1,-nbitq), 
to_sfixed(456705243.0/4294967296.0,1,-nbitq), 
to_sfixed(371597297.0/4294967296.0,1,-nbitq), 
to_sfixed(208004059.0/4294967296.0,1,-nbitq), 
to_sfixed(-240118759.0/4294967296.0,1,-nbitq), 
to_sfixed(-246473994.0/4294967296.0,1,-nbitq), 
to_sfixed(-519847905.0/4294967296.0,1,-nbitq), 
to_sfixed(461258160.0/4294967296.0,1,-nbitq), 
to_sfixed(-306785664.0/4294967296.0,1,-nbitq), 
to_sfixed(92715396.0/4294967296.0,1,-nbitq), 
to_sfixed(-48030048.0/4294967296.0,1,-nbitq), 
to_sfixed(45429499.0/4294967296.0,1,-nbitq), 
to_sfixed(-339153567.0/4294967296.0,1,-nbitq), 
to_sfixed(182620552.0/4294967296.0,1,-nbitq), 
to_sfixed(61188073.0/4294967296.0,1,-nbitq), 
to_sfixed(98268744.0/4294967296.0,1,-nbitq), 
to_sfixed(-59928227.0/4294967296.0,1,-nbitq), 
to_sfixed(126191798.0/4294967296.0,1,-nbitq), 
to_sfixed(-368875566.0/4294967296.0,1,-nbitq), 
to_sfixed(-315851403.0/4294967296.0,1,-nbitq), 
to_sfixed(409254710.0/4294967296.0,1,-nbitq), 
to_sfixed(150723951.0/4294967296.0,1,-nbitq), 
to_sfixed(-337459917.0/4294967296.0,1,-nbitq), 
to_sfixed(192758789.0/4294967296.0,1,-nbitq), 
to_sfixed(203739649.0/4294967296.0,1,-nbitq), 
to_sfixed(-210681634.0/4294967296.0,1,-nbitq), 
to_sfixed(274354941.0/4294967296.0,1,-nbitq), 
to_sfixed(-28909915.0/4294967296.0,1,-nbitq), 
to_sfixed(-484837032.0/4294967296.0,1,-nbitq), 
to_sfixed(278093736.0/4294967296.0,1,-nbitq), 
to_sfixed(113718949.0/4294967296.0,1,-nbitq), 
to_sfixed(-132237832.0/4294967296.0,1,-nbitq), 
to_sfixed(380823002.0/4294967296.0,1,-nbitq), 
to_sfixed(-84808840.0/4294967296.0,1,-nbitq), 
to_sfixed(-275853199.0/4294967296.0,1,-nbitq), 
to_sfixed(203100451.0/4294967296.0,1,-nbitq), 
to_sfixed(383775197.0/4294967296.0,1,-nbitq), 
to_sfixed(-263143826.0/4294967296.0,1,-nbitq), 
to_sfixed(-553060167.0/4294967296.0,1,-nbitq), 
to_sfixed(322108335.0/4294967296.0,1,-nbitq), 
to_sfixed(-10284173.0/4294967296.0,1,-nbitq), 
to_sfixed(-408217884.0/4294967296.0,1,-nbitq), 
to_sfixed(134207611.0/4294967296.0,1,-nbitq), 
to_sfixed(-434260319.0/4294967296.0,1,-nbitq), 
to_sfixed(-223139772.0/4294967296.0,1,-nbitq), 
to_sfixed(-245925376.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(352558092.0/4294967296.0,1,-nbitq), 
to_sfixed(58058456.0/4294967296.0,1,-nbitq), 
to_sfixed(245943730.0/4294967296.0,1,-nbitq), 
to_sfixed(-141586543.0/4294967296.0,1,-nbitq), 
to_sfixed(147023413.0/4294967296.0,1,-nbitq), 
to_sfixed(-260741468.0/4294967296.0,1,-nbitq), 
to_sfixed(-300532737.0/4294967296.0,1,-nbitq), 
to_sfixed(377210791.0/4294967296.0,1,-nbitq), 
to_sfixed(132837217.0/4294967296.0,1,-nbitq), 
to_sfixed(-206743185.0/4294967296.0,1,-nbitq), 
to_sfixed(-323528706.0/4294967296.0,1,-nbitq), 
to_sfixed(-481598893.0/4294967296.0,1,-nbitq), 
to_sfixed(141473293.0/4294967296.0,1,-nbitq), 
to_sfixed(88160597.0/4294967296.0,1,-nbitq), 
to_sfixed(225003134.0/4294967296.0,1,-nbitq), 
to_sfixed(16749661.0/4294967296.0,1,-nbitq), 
to_sfixed(-7421713.0/4294967296.0,1,-nbitq), 
to_sfixed(-224340887.0/4294967296.0,1,-nbitq), 
to_sfixed(-41701073.0/4294967296.0,1,-nbitq), 
to_sfixed(-67571783.0/4294967296.0,1,-nbitq), 
to_sfixed(-418073674.0/4294967296.0,1,-nbitq), 
to_sfixed(12040659.0/4294967296.0,1,-nbitq), 
to_sfixed(-427667148.0/4294967296.0,1,-nbitq), 
to_sfixed(75749922.0/4294967296.0,1,-nbitq), 
to_sfixed(233728092.0/4294967296.0,1,-nbitq), 
to_sfixed(-168208539.0/4294967296.0,1,-nbitq), 
to_sfixed(-164112136.0/4294967296.0,1,-nbitq), 
to_sfixed(-441802238.0/4294967296.0,1,-nbitq), 
to_sfixed(318154558.0/4294967296.0,1,-nbitq), 
to_sfixed(574592903.0/4294967296.0,1,-nbitq), 
to_sfixed(174179797.0/4294967296.0,1,-nbitq), 
to_sfixed(-167711152.0/4294967296.0,1,-nbitq), 
to_sfixed(467478383.0/4294967296.0,1,-nbitq), 
to_sfixed(-233936058.0/4294967296.0,1,-nbitq), 
to_sfixed(331813943.0/4294967296.0,1,-nbitq), 
to_sfixed(-394313610.0/4294967296.0,1,-nbitq), 
to_sfixed(-34446170.0/4294967296.0,1,-nbitq), 
to_sfixed(374594783.0/4294967296.0,1,-nbitq), 
to_sfixed(225755696.0/4294967296.0,1,-nbitq), 
to_sfixed(159033686.0/4294967296.0,1,-nbitq), 
to_sfixed(-449466538.0/4294967296.0,1,-nbitq), 
to_sfixed(50432711.0/4294967296.0,1,-nbitq), 
to_sfixed(-154922051.0/4294967296.0,1,-nbitq), 
to_sfixed(391600185.0/4294967296.0,1,-nbitq), 
to_sfixed(192220416.0/4294967296.0,1,-nbitq), 
to_sfixed(257442659.0/4294967296.0,1,-nbitq), 
to_sfixed(-94671383.0/4294967296.0,1,-nbitq), 
to_sfixed(63408893.0/4294967296.0,1,-nbitq), 
to_sfixed(12702650.0/4294967296.0,1,-nbitq), 
to_sfixed(180253584.0/4294967296.0,1,-nbitq), 
to_sfixed(283921413.0/4294967296.0,1,-nbitq), 
to_sfixed(-486480807.0/4294967296.0,1,-nbitq), 
to_sfixed(-158621230.0/4294967296.0,1,-nbitq), 
to_sfixed(177772210.0/4294967296.0,1,-nbitq), 
to_sfixed(439317394.0/4294967296.0,1,-nbitq), 
to_sfixed(214763809.0/4294967296.0,1,-nbitq), 
to_sfixed(-224262742.0/4294967296.0,1,-nbitq), 
to_sfixed(-26270802.0/4294967296.0,1,-nbitq), 
to_sfixed(42398505.0/4294967296.0,1,-nbitq), 
to_sfixed(272542964.0/4294967296.0,1,-nbitq), 
to_sfixed(-221027587.0/4294967296.0,1,-nbitq), 
to_sfixed(-87562340.0/4294967296.0,1,-nbitq), 
to_sfixed(-365180322.0/4294967296.0,1,-nbitq), 
to_sfixed(282029028.0/4294967296.0,1,-nbitq), 
to_sfixed(-152679728.0/4294967296.0,1,-nbitq), 
to_sfixed(-197146059.0/4294967296.0,1,-nbitq), 
to_sfixed(279268946.0/4294967296.0,1,-nbitq), 
to_sfixed(269325473.0/4294967296.0,1,-nbitq), 
to_sfixed(16956798.0/4294967296.0,1,-nbitq), 
to_sfixed(389872166.0/4294967296.0,1,-nbitq), 
to_sfixed(-202597915.0/4294967296.0,1,-nbitq), 
to_sfixed(282872297.0/4294967296.0,1,-nbitq), 
to_sfixed(129590329.0/4294967296.0,1,-nbitq), 
to_sfixed(262879257.0/4294967296.0,1,-nbitq), 
to_sfixed(-57320193.0/4294967296.0,1,-nbitq), 
to_sfixed(317296219.0/4294967296.0,1,-nbitq), 
to_sfixed(-137440347.0/4294967296.0,1,-nbitq), 
to_sfixed(-213332506.0/4294967296.0,1,-nbitq), 
to_sfixed(-5043646.0/4294967296.0,1,-nbitq), 
to_sfixed(313766884.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(441092362.0/4294967296.0,1,-nbitq), 
to_sfixed(-573771979.0/4294967296.0,1,-nbitq), 
to_sfixed(702445971.0/4294967296.0,1,-nbitq), 
to_sfixed(27384434.0/4294967296.0,1,-nbitq), 
to_sfixed(-424225167.0/4294967296.0,1,-nbitq), 
to_sfixed(-344904559.0/4294967296.0,1,-nbitq), 
to_sfixed(46933536.0/4294967296.0,1,-nbitq), 
to_sfixed(161319012.0/4294967296.0,1,-nbitq), 
to_sfixed(-271858510.0/4294967296.0,1,-nbitq), 
to_sfixed(-361897387.0/4294967296.0,1,-nbitq), 
to_sfixed(-171574642.0/4294967296.0,1,-nbitq), 
to_sfixed(-359827667.0/4294967296.0,1,-nbitq), 
to_sfixed(-276924329.0/4294967296.0,1,-nbitq), 
to_sfixed(-88312583.0/4294967296.0,1,-nbitq), 
to_sfixed(-7999351.0/4294967296.0,1,-nbitq), 
to_sfixed(-26120207.0/4294967296.0,1,-nbitq), 
to_sfixed(71358925.0/4294967296.0,1,-nbitq), 
to_sfixed(24459860.0/4294967296.0,1,-nbitq), 
to_sfixed(-473083294.0/4294967296.0,1,-nbitq), 
to_sfixed(133872080.0/4294967296.0,1,-nbitq), 
to_sfixed(38493466.0/4294967296.0,1,-nbitq), 
to_sfixed(-195376586.0/4294967296.0,1,-nbitq), 
to_sfixed(-1286967057.0/4294967296.0,1,-nbitq), 
to_sfixed(570963501.0/4294967296.0,1,-nbitq), 
to_sfixed(89760439.0/4294967296.0,1,-nbitq), 
to_sfixed(-260918202.0/4294967296.0,1,-nbitq), 
to_sfixed(-47291349.0/4294967296.0,1,-nbitq), 
to_sfixed(-196216341.0/4294967296.0,1,-nbitq), 
to_sfixed(-348297778.0/4294967296.0,1,-nbitq), 
to_sfixed(-16291245.0/4294967296.0,1,-nbitq), 
to_sfixed(-360592443.0/4294967296.0,1,-nbitq), 
to_sfixed(-251788332.0/4294967296.0,1,-nbitq), 
to_sfixed(125563396.0/4294967296.0,1,-nbitq), 
to_sfixed(486524784.0/4294967296.0,1,-nbitq), 
to_sfixed(55141890.0/4294967296.0,1,-nbitq), 
to_sfixed(-507983766.0/4294967296.0,1,-nbitq), 
to_sfixed(91356053.0/4294967296.0,1,-nbitq), 
to_sfixed(468626593.0/4294967296.0,1,-nbitq), 
to_sfixed(200469064.0/4294967296.0,1,-nbitq), 
to_sfixed(68031470.0/4294967296.0,1,-nbitq), 
to_sfixed(-435698020.0/4294967296.0,1,-nbitq), 
to_sfixed(-166502222.0/4294967296.0,1,-nbitq), 
to_sfixed(-207380377.0/4294967296.0,1,-nbitq), 
to_sfixed(245295913.0/4294967296.0,1,-nbitq), 
to_sfixed(-232824411.0/4294967296.0,1,-nbitq), 
to_sfixed(64358430.0/4294967296.0,1,-nbitq), 
to_sfixed(293812762.0/4294967296.0,1,-nbitq), 
to_sfixed(23111948.0/4294967296.0,1,-nbitq), 
to_sfixed(-294019785.0/4294967296.0,1,-nbitq), 
to_sfixed(-184508681.0/4294967296.0,1,-nbitq), 
to_sfixed(-26672416.0/4294967296.0,1,-nbitq), 
to_sfixed(-485544412.0/4294967296.0,1,-nbitq), 
to_sfixed(391477227.0/4294967296.0,1,-nbitq), 
to_sfixed(-56592801.0/4294967296.0,1,-nbitq), 
to_sfixed(471869937.0/4294967296.0,1,-nbitq), 
to_sfixed(-228022711.0/4294967296.0,1,-nbitq), 
to_sfixed(-338089625.0/4294967296.0,1,-nbitq), 
to_sfixed(-294146350.0/4294967296.0,1,-nbitq), 
to_sfixed(-353383765.0/4294967296.0,1,-nbitq), 
to_sfixed(-211218310.0/4294967296.0,1,-nbitq), 
to_sfixed(-413627559.0/4294967296.0,1,-nbitq), 
to_sfixed(381595640.0/4294967296.0,1,-nbitq), 
to_sfixed(-337650598.0/4294967296.0,1,-nbitq), 
to_sfixed(155777280.0/4294967296.0,1,-nbitq), 
to_sfixed(-117782214.0/4294967296.0,1,-nbitq), 
to_sfixed(-431935490.0/4294967296.0,1,-nbitq), 
to_sfixed(49674791.0/4294967296.0,1,-nbitq), 
to_sfixed(645525891.0/4294967296.0,1,-nbitq), 
to_sfixed(75851942.0/4294967296.0,1,-nbitq), 
to_sfixed(251969918.0/4294967296.0,1,-nbitq), 
to_sfixed(-462270614.0/4294967296.0,1,-nbitq), 
to_sfixed(88271938.0/4294967296.0,1,-nbitq), 
to_sfixed(444073033.0/4294967296.0,1,-nbitq), 
to_sfixed(300157977.0/4294967296.0,1,-nbitq), 
to_sfixed(335050243.0/4294967296.0,1,-nbitq), 
to_sfixed(409741676.0/4294967296.0,1,-nbitq), 
to_sfixed(-326696870.0/4294967296.0,1,-nbitq), 
to_sfixed(-254471608.0/4294967296.0,1,-nbitq), 
to_sfixed(511884129.0/4294967296.0,1,-nbitq), 
to_sfixed(161319171.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-95709764.0/4294967296.0,1,-nbitq), 
to_sfixed(-173822321.0/4294967296.0,1,-nbitq), 
to_sfixed(778806228.0/4294967296.0,1,-nbitq), 
to_sfixed(-101444639.0/4294967296.0,1,-nbitq), 
to_sfixed(-394001356.0/4294967296.0,1,-nbitq), 
to_sfixed(212179215.0/4294967296.0,1,-nbitq), 
to_sfixed(-302927615.0/4294967296.0,1,-nbitq), 
to_sfixed(-307421435.0/4294967296.0,1,-nbitq), 
to_sfixed(2143856.0/4294967296.0,1,-nbitq), 
to_sfixed(426228398.0/4294967296.0,1,-nbitq), 
to_sfixed(249954211.0/4294967296.0,1,-nbitq), 
to_sfixed(-658550655.0/4294967296.0,1,-nbitq), 
to_sfixed(246460725.0/4294967296.0,1,-nbitq), 
to_sfixed(665582906.0/4294967296.0,1,-nbitq), 
to_sfixed(96052366.0/4294967296.0,1,-nbitq), 
to_sfixed(663007946.0/4294967296.0,1,-nbitq), 
to_sfixed(131094892.0/4294967296.0,1,-nbitq), 
to_sfixed(-396532073.0/4294967296.0,1,-nbitq), 
to_sfixed(-577541726.0/4294967296.0,1,-nbitq), 
to_sfixed(503830875.0/4294967296.0,1,-nbitq), 
to_sfixed(149502218.0/4294967296.0,1,-nbitq), 
to_sfixed(-395316994.0/4294967296.0,1,-nbitq), 
to_sfixed(-1496153995.0/4294967296.0,1,-nbitq), 
to_sfixed(107985611.0/4294967296.0,1,-nbitq), 
to_sfixed(-165052143.0/4294967296.0,1,-nbitq), 
to_sfixed(-928993211.0/4294967296.0,1,-nbitq), 
to_sfixed(756865650.0/4294967296.0,1,-nbitq), 
to_sfixed(352797733.0/4294967296.0,1,-nbitq), 
to_sfixed(434162743.0/4294967296.0,1,-nbitq), 
to_sfixed(357672785.0/4294967296.0,1,-nbitq), 
to_sfixed(-206475989.0/4294967296.0,1,-nbitq), 
to_sfixed(-118167106.0/4294967296.0,1,-nbitq), 
to_sfixed(515529974.0/4294967296.0,1,-nbitq), 
to_sfixed(409062257.0/4294967296.0,1,-nbitq), 
to_sfixed(-9367080.0/4294967296.0,1,-nbitq), 
to_sfixed(278680628.0/4294967296.0,1,-nbitq), 
to_sfixed(-385635389.0/4294967296.0,1,-nbitq), 
to_sfixed(-84546984.0/4294967296.0,1,-nbitq), 
to_sfixed(-393755228.0/4294967296.0,1,-nbitq), 
to_sfixed(-49996993.0/4294967296.0,1,-nbitq), 
to_sfixed(-383529752.0/4294967296.0,1,-nbitq), 
to_sfixed(-265195467.0/4294967296.0,1,-nbitq), 
to_sfixed(-657478703.0/4294967296.0,1,-nbitq), 
to_sfixed(-1363761456.0/4294967296.0,1,-nbitq), 
to_sfixed(-598196739.0/4294967296.0,1,-nbitq), 
to_sfixed(25888237.0/4294967296.0,1,-nbitq), 
to_sfixed(248728730.0/4294967296.0,1,-nbitq), 
to_sfixed(-121141276.0/4294967296.0,1,-nbitq), 
to_sfixed(155987522.0/4294967296.0,1,-nbitq), 
to_sfixed(-166318128.0/4294967296.0,1,-nbitq), 
to_sfixed(-27613871.0/4294967296.0,1,-nbitq), 
to_sfixed(-228968689.0/4294967296.0,1,-nbitq), 
to_sfixed(728575870.0/4294967296.0,1,-nbitq), 
to_sfixed(-556692837.0/4294967296.0,1,-nbitq), 
to_sfixed(-161686116.0/4294967296.0,1,-nbitq), 
to_sfixed(66320266.0/4294967296.0,1,-nbitq), 
to_sfixed(254064372.0/4294967296.0,1,-nbitq), 
to_sfixed(676602404.0/4294967296.0,1,-nbitq), 
to_sfixed(-208456384.0/4294967296.0,1,-nbitq), 
to_sfixed(12803153.0/4294967296.0,1,-nbitq), 
to_sfixed(-329411994.0/4294967296.0,1,-nbitq), 
to_sfixed(56876141.0/4294967296.0,1,-nbitq), 
to_sfixed(773599184.0/4294967296.0,1,-nbitq), 
to_sfixed(-550559141.0/4294967296.0,1,-nbitq), 
to_sfixed(-197294785.0/4294967296.0,1,-nbitq), 
to_sfixed(-281565637.0/4294967296.0,1,-nbitq), 
to_sfixed(467578127.0/4294967296.0,1,-nbitq), 
to_sfixed(38800313.0/4294967296.0,1,-nbitq), 
to_sfixed(-321762452.0/4294967296.0,1,-nbitq), 
to_sfixed(-294160390.0/4294967296.0,1,-nbitq), 
to_sfixed(141661440.0/4294967296.0,1,-nbitq), 
to_sfixed(-93578078.0/4294967296.0,1,-nbitq), 
to_sfixed(763813232.0/4294967296.0,1,-nbitq), 
to_sfixed(-295854134.0/4294967296.0,1,-nbitq), 
to_sfixed(317539316.0/4294967296.0,1,-nbitq), 
to_sfixed(170648794.0/4294967296.0,1,-nbitq), 
to_sfixed(-837677013.0/4294967296.0,1,-nbitq), 
to_sfixed(80223628.0/4294967296.0,1,-nbitq), 
to_sfixed(689039208.0/4294967296.0,1,-nbitq), 
to_sfixed(33566462.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-46519846.0/4294967296.0,1,-nbitq), 
to_sfixed(429598521.0/4294967296.0,1,-nbitq), 
to_sfixed(296906626.0/4294967296.0,1,-nbitq), 
to_sfixed(-236529367.0/4294967296.0,1,-nbitq), 
to_sfixed(-389071257.0/4294967296.0,1,-nbitq), 
to_sfixed(528538866.0/4294967296.0,1,-nbitq), 
to_sfixed(424604256.0/4294967296.0,1,-nbitq), 
to_sfixed(221646929.0/4294967296.0,1,-nbitq), 
to_sfixed(113317681.0/4294967296.0,1,-nbitq), 
to_sfixed(-324518611.0/4294967296.0,1,-nbitq), 
to_sfixed(551768638.0/4294967296.0,1,-nbitq), 
to_sfixed(-547935310.0/4294967296.0,1,-nbitq), 
to_sfixed(-685383753.0/4294967296.0,1,-nbitq), 
to_sfixed(877905129.0/4294967296.0,1,-nbitq), 
to_sfixed(41012575.0/4294967296.0,1,-nbitq), 
to_sfixed(515908516.0/4294967296.0,1,-nbitq), 
to_sfixed(370571377.0/4294967296.0,1,-nbitq), 
to_sfixed(-246644136.0/4294967296.0,1,-nbitq), 
to_sfixed(-518005912.0/4294967296.0,1,-nbitq), 
to_sfixed(941210147.0/4294967296.0,1,-nbitq), 
to_sfixed(-290340595.0/4294967296.0,1,-nbitq), 
to_sfixed(-8582541.0/4294967296.0,1,-nbitq), 
to_sfixed(-688169379.0/4294967296.0,1,-nbitq), 
to_sfixed(506987208.0/4294967296.0,1,-nbitq), 
to_sfixed(98047285.0/4294967296.0,1,-nbitq), 
to_sfixed(-645738333.0/4294967296.0,1,-nbitq), 
to_sfixed(322287251.0/4294967296.0,1,-nbitq), 
to_sfixed(737494754.0/4294967296.0,1,-nbitq), 
to_sfixed(726580033.0/4294967296.0,1,-nbitq), 
to_sfixed(-234254705.0/4294967296.0,1,-nbitq), 
to_sfixed(80527531.0/4294967296.0,1,-nbitq), 
to_sfixed(-69156850.0/4294967296.0,1,-nbitq), 
to_sfixed(300613767.0/4294967296.0,1,-nbitq), 
to_sfixed(-618059315.0/4294967296.0,1,-nbitq), 
to_sfixed(330964668.0/4294967296.0,1,-nbitq), 
to_sfixed(-519305040.0/4294967296.0,1,-nbitq), 
to_sfixed(-768982024.0/4294967296.0,1,-nbitq), 
to_sfixed(-380136657.0/4294967296.0,1,-nbitq), 
to_sfixed(-227618066.0/4294967296.0,1,-nbitq), 
to_sfixed(476583105.0/4294967296.0,1,-nbitq), 
to_sfixed(-281703000.0/4294967296.0,1,-nbitq), 
to_sfixed(-535777371.0/4294967296.0,1,-nbitq), 
to_sfixed(-344044996.0/4294967296.0,1,-nbitq), 
to_sfixed(-1234324468.0/4294967296.0,1,-nbitq), 
to_sfixed(-497104743.0/4294967296.0,1,-nbitq), 
to_sfixed(352812254.0/4294967296.0,1,-nbitq), 
to_sfixed(171058330.0/4294967296.0,1,-nbitq), 
to_sfixed(251483343.0/4294967296.0,1,-nbitq), 
to_sfixed(-24522945.0/4294967296.0,1,-nbitq), 
to_sfixed(-201470028.0/4294967296.0,1,-nbitq), 
to_sfixed(-377997272.0/4294967296.0,1,-nbitq), 
to_sfixed(-916246810.0/4294967296.0,1,-nbitq), 
to_sfixed(771732908.0/4294967296.0,1,-nbitq), 
to_sfixed(-495964465.0/4294967296.0,1,-nbitq), 
to_sfixed(-901645470.0/4294967296.0,1,-nbitq), 
to_sfixed(50948202.0/4294967296.0,1,-nbitq), 
to_sfixed(51361390.0/4294967296.0,1,-nbitq), 
to_sfixed(-353707476.0/4294967296.0,1,-nbitq), 
to_sfixed(416466037.0/4294967296.0,1,-nbitq), 
to_sfixed(428586179.0/4294967296.0,1,-nbitq), 
to_sfixed(331700202.0/4294967296.0,1,-nbitq), 
to_sfixed(168093509.0/4294967296.0,1,-nbitq), 
to_sfixed(388305118.0/4294967296.0,1,-nbitq), 
to_sfixed(141716786.0/4294967296.0,1,-nbitq), 
to_sfixed(-447131428.0/4294967296.0,1,-nbitq), 
to_sfixed(-104832186.0/4294967296.0,1,-nbitq), 
to_sfixed(-776586784.0/4294967296.0,1,-nbitq), 
to_sfixed(130084242.0/4294967296.0,1,-nbitq), 
to_sfixed(390581501.0/4294967296.0,1,-nbitq), 
to_sfixed(-967283782.0/4294967296.0,1,-nbitq), 
to_sfixed(303954854.0/4294967296.0,1,-nbitq), 
to_sfixed(-88718042.0/4294967296.0,1,-nbitq), 
to_sfixed(558407532.0/4294967296.0,1,-nbitq), 
to_sfixed(-149089819.0/4294967296.0,1,-nbitq), 
to_sfixed(387764674.0/4294967296.0,1,-nbitq), 
to_sfixed(-510367109.0/4294967296.0,1,-nbitq), 
to_sfixed(-1506269212.0/4294967296.0,1,-nbitq), 
to_sfixed(166324056.0/4294967296.0,1,-nbitq), 
to_sfixed(-591378694.0/4294967296.0,1,-nbitq), 
to_sfixed(2064135.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-51427278.0/4294967296.0,1,-nbitq), 
to_sfixed(348152328.0/4294967296.0,1,-nbitq), 
to_sfixed(-591529812.0/4294967296.0,1,-nbitq), 
to_sfixed(806176082.0/4294967296.0,1,-nbitq), 
to_sfixed(587971998.0/4294967296.0,1,-nbitq), 
to_sfixed(1190576972.0/4294967296.0,1,-nbitq), 
to_sfixed(503099609.0/4294967296.0,1,-nbitq), 
to_sfixed(1094827874.0/4294967296.0,1,-nbitq), 
to_sfixed(841131570.0/4294967296.0,1,-nbitq), 
to_sfixed(-336315741.0/4294967296.0,1,-nbitq), 
to_sfixed(211657090.0/4294967296.0,1,-nbitq), 
to_sfixed(-1489081990.0/4294967296.0,1,-nbitq), 
to_sfixed(-1034800534.0/4294967296.0,1,-nbitq), 
to_sfixed(-63626446.0/4294967296.0,1,-nbitq), 
to_sfixed(-134128176.0/4294967296.0,1,-nbitq), 
to_sfixed(516386715.0/4294967296.0,1,-nbitq), 
to_sfixed(-361768285.0/4294967296.0,1,-nbitq), 
to_sfixed(-34746150.0/4294967296.0,1,-nbitq), 
to_sfixed(-592559288.0/4294967296.0,1,-nbitq), 
to_sfixed(1000295643.0/4294967296.0,1,-nbitq), 
to_sfixed(-6832185.0/4294967296.0,1,-nbitq), 
to_sfixed(277517195.0/4294967296.0,1,-nbitq), 
to_sfixed(294131140.0/4294967296.0,1,-nbitq), 
to_sfixed(114429342.0/4294967296.0,1,-nbitq), 
to_sfixed(-246949739.0/4294967296.0,1,-nbitq), 
to_sfixed(-1288865188.0/4294967296.0,1,-nbitq), 
to_sfixed(396060793.0/4294967296.0,1,-nbitq), 
to_sfixed(891541029.0/4294967296.0,1,-nbitq), 
to_sfixed(562947732.0/4294967296.0,1,-nbitq), 
to_sfixed(302971286.0/4294967296.0,1,-nbitq), 
to_sfixed(46690445.0/4294967296.0,1,-nbitq), 
to_sfixed(204621307.0/4294967296.0,1,-nbitq), 
to_sfixed(758407650.0/4294967296.0,1,-nbitq), 
to_sfixed(309069629.0/4294967296.0,1,-nbitq), 
to_sfixed(-441543725.0/4294967296.0,1,-nbitq), 
to_sfixed(-1816063066.0/4294967296.0,1,-nbitq), 
to_sfixed(-936401746.0/4294967296.0,1,-nbitq), 
to_sfixed(434230336.0/4294967296.0,1,-nbitq), 
to_sfixed(493738239.0/4294967296.0,1,-nbitq), 
to_sfixed(171683499.0/4294967296.0,1,-nbitq), 
to_sfixed(-79903245.0/4294967296.0,1,-nbitq), 
to_sfixed(-154448928.0/4294967296.0,1,-nbitq), 
to_sfixed(216114368.0/4294967296.0,1,-nbitq), 
to_sfixed(-75177497.0/4294967296.0,1,-nbitq), 
to_sfixed(-105736480.0/4294967296.0,1,-nbitq), 
to_sfixed(-326877761.0/4294967296.0,1,-nbitq), 
to_sfixed(268613582.0/4294967296.0,1,-nbitq), 
to_sfixed(917200960.0/4294967296.0,1,-nbitq), 
to_sfixed(199701133.0/4294967296.0,1,-nbitq), 
to_sfixed(372869030.0/4294967296.0,1,-nbitq), 
to_sfixed(-598489851.0/4294967296.0,1,-nbitq), 
to_sfixed(-696286725.0/4294967296.0,1,-nbitq), 
to_sfixed(1204632249.0/4294967296.0,1,-nbitq), 
to_sfixed(758096533.0/4294967296.0,1,-nbitq), 
to_sfixed(-306860825.0/4294967296.0,1,-nbitq), 
to_sfixed(116120694.0/4294967296.0,1,-nbitq), 
to_sfixed(-155955345.0/4294967296.0,1,-nbitq), 
to_sfixed(-682166236.0/4294967296.0,1,-nbitq), 
to_sfixed(-355897943.0/4294967296.0,1,-nbitq), 
to_sfixed(233709680.0/4294967296.0,1,-nbitq), 
to_sfixed(-135632571.0/4294967296.0,1,-nbitq), 
to_sfixed(675806601.0/4294967296.0,1,-nbitq), 
to_sfixed(1818894692.0/4294967296.0,1,-nbitq), 
to_sfixed(629326077.0/4294967296.0,1,-nbitq), 
to_sfixed(166398491.0/4294967296.0,1,-nbitq), 
to_sfixed(-90332722.0/4294967296.0,1,-nbitq), 
to_sfixed(-783942878.0/4294967296.0,1,-nbitq), 
to_sfixed(139277213.0/4294967296.0,1,-nbitq), 
to_sfixed(358237836.0/4294967296.0,1,-nbitq), 
to_sfixed(-123025508.0/4294967296.0,1,-nbitq), 
to_sfixed(-426731403.0/4294967296.0,1,-nbitq), 
to_sfixed(-397228332.0/4294967296.0,1,-nbitq), 
to_sfixed(472912523.0/4294967296.0,1,-nbitq), 
to_sfixed(79568964.0/4294967296.0,1,-nbitq), 
to_sfixed(-187911498.0/4294967296.0,1,-nbitq), 
to_sfixed(256117345.0/4294967296.0,1,-nbitq), 
to_sfixed(-1332082252.0/4294967296.0,1,-nbitq), 
to_sfixed(211100588.0/4294967296.0,1,-nbitq), 
to_sfixed(-297097085.0/4294967296.0,1,-nbitq), 
to_sfixed(-113866212.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-424216705.0/4294967296.0,1,-nbitq), 
to_sfixed(-65433967.0/4294967296.0,1,-nbitq), 
to_sfixed(-554498274.0/4294967296.0,1,-nbitq), 
to_sfixed(1413283138.0/4294967296.0,1,-nbitq), 
to_sfixed(39224263.0/4294967296.0,1,-nbitq), 
to_sfixed(1835041144.0/4294967296.0,1,-nbitq), 
to_sfixed(499139340.0/4294967296.0,1,-nbitq), 
to_sfixed(1707105230.0/4294967296.0,1,-nbitq), 
to_sfixed(-24718621.0/4294967296.0,1,-nbitq), 
to_sfixed(-367091954.0/4294967296.0,1,-nbitq), 
to_sfixed(-81836976.0/4294967296.0,1,-nbitq), 
to_sfixed(-2342447366.0/4294967296.0,1,-nbitq), 
to_sfixed(-180423479.0/4294967296.0,1,-nbitq), 
to_sfixed(98893731.0/4294967296.0,1,-nbitq), 
to_sfixed(181933076.0/4294967296.0,1,-nbitq), 
to_sfixed(510042291.0/4294967296.0,1,-nbitq), 
to_sfixed(192445355.0/4294967296.0,1,-nbitq), 
to_sfixed(-170927709.0/4294967296.0,1,-nbitq), 
to_sfixed(-293618789.0/4294967296.0,1,-nbitq), 
to_sfixed(675975330.0/4294967296.0,1,-nbitq), 
to_sfixed(-81035570.0/4294967296.0,1,-nbitq), 
to_sfixed(213566056.0/4294967296.0,1,-nbitq), 
to_sfixed(30402546.0/4294967296.0,1,-nbitq), 
to_sfixed(464217609.0/4294967296.0,1,-nbitq), 
to_sfixed(-139565533.0/4294967296.0,1,-nbitq), 
to_sfixed(-1511551943.0/4294967296.0,1,-nbitq), 
to_sfixed(396965041.0/4294967296.0,1,-nbitq), 
to_sfixed(-173704570.0/4294967296.0,1,-nbitq), 
to_sfixed(474371044.0/4294967296.0,1,-nbitq), 
to_sfixed(369478028.0/4294967296.0,1,-nbitq), 
to_sfixed(168118096.0/4294967296.0,1,-nbitq), 
to_sfixed(814981823.0/4294967296.0,1,-nbitq), 
to_sfixed(537238811.0/4294967296.0,1,-nbitq), 
to_sfixed(-115754810.0/4294967296.0,1,-nbitq), 
to_sfixed(-752403025.0/4294967296.0,1,-nbitq), 
to_sfixed(-2406874076.0/4294967296.0,1,-nbitq), 
to_sfixed(-1379119076.0/4294967296.0,1,-nbitq), 
to_sfixed(-314149139.0/4294967296.0,1,-nbitq), 
to_sfixed(-292447601.0/4294967296.0,1,-nbitq), 
to_sfixed(150384456.0/4294967296.0,1,-nbitq), 
to_sfixed(-27172929.0/4294967296.0,1,-nbitq), 
to_sfixed(123686589.0/4294967296.0,1,-nbitq), 
to_sfixed(-271434173.0/4294967296.0,1,-nbitq), 
to_sfixed(-1056912370.0/4294967296.0,1,-nbitq), 
to_sfixed(-256452534.0/4294967296.0,1,-nbitq), 
to_sfixed(-141834063.0/4294967296.0,1,-nbitq), 
to_sfixed(-43136626.0/4294967296.0,1,-nbitq), 
to_sfixed(883042326.0/4294967296.0,1,-nbitq), 
to_sfixed(547732566.0/4294967296.0,1,-nbitq), 
to_sfixed(230937420.0/4294967296.0,1,-nbitq), 
to_sfixed(-187338247.0/4294967296.0,1,-nbitq), 
to_sfixed(-851999303.0/4294967296.0,1,-nbitq), 
to_sfixed(1090634914.0/4294967296.0,1,-nbitq), 
to_sfixed(709437648.0/4294967296.0,1,-nbitq), 
to_sfixed(-197011931.0/4294967296.0,1,-nbitq), 
to_sfixed(-476692369.0/4294967296.0,1,-nbitq), 
to_sfixed(175314261.0/4294967296.0,1,-nbitq), 
to_sfixed(-229257846.0/4294967296.0,1,-nbitq), 
to_sfixed(-198545720.0/4294967296.0,1,-nbitq), 
to_sfixed(421484503.0/4294967296.0,1,-nbitq), 
to_sfixed(308810213.0/4294967296.0,1,-nbitq), 
to_sfixed(247539659.0/4294967296.0,1,-nbitq), 
to_sfixed(1780014649.0/4294967296.0,1,-nbitq), 
to_sfixed(481683100.0/4294967296.0,1,-nbitq), 
to_sfixed(-113310610.0/4294967296.0,1,-nbitq), 
to_sfixed(324579075.0/4294967296.0,1,-nbitq), 
to_sfixed(-1426988936.0/4294967296.0,1,-nbitq), 
to_sfixed(542100185.0/4294967296.0,1,-nbitq), 
to_sfixed(-145550092.0/4294967296.0,1,-nbitq), 
to_sfixed(412713350.0/4294967296.0,1,-nbitq), 
to_sfixed(393074452.0/4294967296.0,1,-nbitq), 
to_sfixed(-574055557.0/4294967296.0,1,-nbitq), 
to_sfixed(803083764.0/4294967296.0,1,-nbitq), 
to_sfixed(-156929930.0/4294967296.0,1,-nbitq), 
to_sfixed(66528099.0/4294967296.0,1,-nbitq), 
to_sfixed(387228448.0/4294967296.0,1,-nbitq), 
to_sfixed(-1031340117.0/4294967296.0,1,-nbitq), 
to_sfixed(314706332.0/4294967296.0,1,-nbitq), 
to_sfixed(-217450079.0/4294967296.0,1,-nbitq), 
to_sfixed(400961373.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-1051991741.0/4294967296.0,1,-nbitq), 
to_sfixed(143194827.0/4294967296.0,1,-nbitq), 
to_sfixed(246604677.0/4294967296.0,1,-nbitq), 
to_sfixed(1639695116.0/4294967296.0,1,-nbitq), 
to_sfixed(399645669.0/4294967296.0,1,-nbitq), 
to_sfixed(1680506721.0/4294967296.0,1,-nbitq), 
to_sfixed(-125013586.0/4294967296.0,1,-nbitq), 
to_sfixed(1650327099.0/4294967296.0,1,-nbitq), 
to_sfixed(-516881872.0/4294967296.0,1,-nbitq), 
to_sfixed(-182242316.0/4294967296.0,1,-nbitq), 
to_sfixed(-153238406.0/4294967296.0,1,-nbitq), 
to_sfixed(-2065038431.0/4294967296.0,1,-nbitq), 
to_sfixed(-198812350.0/4294967296.0,1,-nbitq), 
to_sfixed(124919070.0/4294967296.0,1,-nbitq), 
to_sfixed(-152946740.0/4294967296.0,1,-nbitq), 
to_sfixed(526883660.0/4294967296.0,1,-nbitq), 
to_sfixed(-295048923.0/4294967296.0,1,-nbitq), 
to_sfixed(-185691242.0/4294967296.0,1,-nbitq), 
to_sfixed(857769573.0/4294967296.0,1,-nbitq), 
to_sfixed(908258691.0/4294967296.0,1,-nbitq), 
to_sfixed(193533425.0/4294967296.0,1,-nbitq), 
to_sfixed(197752872.0/4294967296.0,1,-nbitq), 
to_sfixed(-209000955.0/4294967296.0,1,-nbitq), 
to_sfixed(133156286.0/4294967296.0,1,-nbitq), 
to_sfixed(-17915938.0/4294967296.0,1,-nbitq), 
to_sfixed(-989339550.0/4294967296.0,1,-nbitq), 
to_sfixed(159608370.0/4294967296.0,1,-nbitq), 
to_sfixed(-138646896.0/4294967296.0,1,-nbitq), 
to_sfixed(-167599948.0/4294967296.0,1,-nbitq), 
to_sfixed(885203258.0/4294967296.0,1,-nbitq), 
to_sfixed(493708027.0/4294967296.0,1,-nbitq), 
to_sfixed(737501798.0/4294967296.0,1,-nbitq), 
to_sfixed(505329220.0/4294967296.0,1,-nbitq), 
to_sfixed(893885306.0/4294967296.0,1,-nbitq), 
to_sfixed(-364297566.0/4294967296.0,1,-nbitq), 
to_sfixed(-1007945625.0/4294967296.0,1,-nbitq), 
to_sfixed(-1614676438.0/4294967296.0,1,-nbitq), 
to_sfixed(-925413312.0/4294967296.0,1,-nbitq), 
to_sfixed(179097587.0/4294967296.0,1,-nbitq), 
to_sfixed(252711949.0/4294967296.0,1,-nbitq), 
to_sfixed(-439549545.0/4294967296.0,1,-nbitq), 
to_sfixed(400859436.0/4294967296.0,1,-nbitq), 
to_sfixed(318997542.0/4294967296.0,1,-nbitq), 
to_sfixed(-714463240.0/4294967296.0,1,-nbitq), 
to_sfixed(-345600843.0/4294967296.0,1,-nbitq), 
to_sfixed(-41792847.0/4294967296.0,1,-nbitq), 
to_sfixed(52970311.0/4294967296.0,1,-nbitq), 
to_sfixed(1067500863.0/4294967296.0,1,-nbitq), 
to_sfixed(740971812.0/4294967296.0,1,-nbitq), 
to_sfixed(-13230061.0/4294967296.0,1,-nbitq), 
to_sfixed(-680613386.0/4294967296.0,1,-nbitq), 
to_sfixed(-792274663.0/4294967296.0,1,-nbitq), 
to_sfixed(828623282.0/4294967296.0,1,-nbitq), 
to_sfixed(264630275.0/4294967296.0,1,-nbitq), 
to_sfixed(591028939.0/4294967296.0,1,-nbitq), 
to_sfixed(-260733504.0/4294967296.0,1,-nbitq), 
to_sfixed(-11275185.0/4294967296.0,1,-nbitq), 
to_sfixed(45351006.0/4294967296.0,1,-nbitq), 
to_sfixed(364188541.0/4294967296.0,1,-nbitq), 
to_sfixed(400965400.0/4294967296.0,1,-nbitq), 
to_sfixed(-7015168.0/4294967296.0,1,-nbitq), 
to_sfixed(-183555908.0/4294967296.0,1,-nbitq), 
to_sfixed(1772312835.0/4294967296.0,1,-nbitq), 
to_sfixed(79237481.0/4294967296.0,1,-nbitq), 
to_sfixed(-82093029.0/4294967296.0,1,-nbitq), 
to_sfixed(-63613377.0/4294967296.0,1,-nbitq), 
to_sfixed(-1680704794.0/4294967296.0,1,-nbitq), 
to_sfixed(-355154586.0/4294967296.0,1,-nbitq), 
to_sfixed(402259626.0/4294967296.0,1,-nbitq), 
to_sfixed(-125884889.0/4294967296.0,1,-nbitq), 
to_sfixed(384768465.0/4294967296.0,1,-nbitq), 
to_sfixed(-218322951.0/4294967296.0,1,-nbitq), 
to_sfixed(610479201.0/4294967296.0,1,-nbitq), 
to_sfixed(252293998.0/4294967296.0,1,-nbitq), 
to_sfixed(-228374044.0/4294967296.0,1,-nbitq), 
to_sfixed(65560253.0/4294967296.0,1,-nbitq), 
to_sfixed(-775365734.0/4294967296.0,1,-nbitq), 
to_sfixed(-284208102.0/4294967296.0,1,-nbitq), 
to_sfixed(-257581004.0/4294967296.0,1,-nbitq), 
to_sfixed(407056445.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-616852873.0/4294967296.0,1,-nbitq), 
to_sfixed(-902001625.0/4294967296.0,1,-nbitq), 
to_sfixed(740921476.0/4294967296.0,1,-nbitq), 
to_sfixed(921433480.0/4294967296.0,1,-nbitq), 
to_sfixed(295723020.0/4294967296.0,1,-nbitq), 
to_sfixed(419648518.0/4294967296.0,1,-nbitq), 
to_sfixed(21851450.0/4294967296.0,1,-nbitq), 
to_sfixed(1700782049.0/4294967296.0,1,-nbitq), 
to_sfixed(-885379811.0/4294967296.0,1,-nbitq), 
to_sfixed(-116574852.0/4294967296.0,1,-nbitq), 
to_sfixed(-666973532.0/4294967296.0,1,-nbitq), 
to_sfixed(-543552201.0/4294967296.0,1,-nbitq), 
to_sfixed(-712665023.0/4294967296.0,1,-nbitq), 
to_sfixed(-1160046272.0/4294967296.0,1,-nbitq), 
to_sfixed(285198366.0/4294967296.0,1,-nbitq), 
to_sfixed(850031859.0/4294967296.0,1,-nbitq), 
to_sfixed(-199422321.0/4294967296.0,1,-nbitq), 
to_sfixed(-323267293.0/4294967296.0,1,-nbitq), 
to_sfixed(1716093965.0/4294967296.0,1,-nbitq), 
to_sfixed(741055405.0/4294967296.0,1,-nbitq), 
to_sfixed(-223346432.0/4294967296.0,1,-nbitq), 
to_sfixed(154255528.0/4294967296.0,1,-nbitq), 
to_sfixed(-116759018.0/4294967296.0,1,-nbitq), 
to_sfixed(725205436.0/4294967296.0,1,-nbitq), 
to_sfixed(347932763.0/4294967296.0,1,-nbitq), 
to_sfixed(-984849495.0/4294967296.0,1,-nbitq), 
to_sfixed(-619742394.0/4294967296.0,1,-nbitq), 
to_sfixed(578578476.0/4294967296.0,1,-nbitq), 
to_sfixed(240148441.0/4294967296.0,1,-nbitq), 
to_sfixed(1106517537.0/4294967296.0,1,-nbitq), 
to_sfixed(572020994.0/4294967296.0,1,-nbitq), 
to_sfixed(1093541902.0/4294967296.0,1,-nbitq), 
to_sfixed(289357078.0/4294967296.0,1,-nbitq), 
to_sfixed(1863899564.0/4294967296.0,1,-nbitq), 
to_sfixed(-431870372.0/4294967296.0,1,-nbitq), 
to_sfixed(21415350.0/4294967296.0,1,-nbitq), 
to_sfixed(-1638421563.0/4294967296.0,1,-nbitq), 
to_sfixed(17347037.0/4294967296.0,1,-nbitq), 
to_sfixed(30408338.0/4294967296.0,1,-nbitq), 
to_sfixed(128975734.0/4294967296.0,1,-nbitq), 
to_sfixed(204712616.0/4294967296.0,1,-nbitq), 
to_sfixed(-41346531.0/4294967296.0,1,-nbitq), 
to_sfixed(795217023.0/4294967296.0,1,-nbitq), 
to_sfixed(-416607131.0/4294967296.0,1,-nbitq), 
to_sfixed(-19828968.0/4294967296.0,1,-nbitq), 
to_sfixed(-782416421.0/4294967296.0,1,-nbitq), 
to_sfixed(-277150305.0/4294967296.0,1,-nbitq), 
to_sfixed(1340962024.0/4294967296.0,1,-nbitq), 
to_sfixed(30243052.0/4294967296.0,1,-nbitq), 
to_sfixed(598164098.0/4294967296.0,1,-nbitq), 
to_sfixed(-831966427.0/4294967296.0,1,-nbitq), 
to_sfixed(256847355.0/4294967296.0,1,-nbitq), 
to_sfixed(688535943.0/4294967296.0,1,-nbitq), 
to_sfixed(286342235.0/4294967296.0,1,-nbitq), 
to_sfixed(724539392.0/4294967296.0,1,-nbitq), 
to_sfixed(-497868573.0/4294967296.0,1,-nbitq), 
to_sfixed(2121040.0/4294967296.0,1,-nbitq), 
to_sfixed(-627073297.0/4294967296.0,1,-nbitq), 
to_sfixed(442393502.0/4294967296.0,1,-nbitq), 
to_sfixed(-223420196.0/4294967296.0,1,-nbitq), 
to_sfixed(-269674545.0/4294967296.0,1,-nbitq), 
to_sfixed(-949070565.0/4294967296.0,1,-nbitq), 
to_sfixed(1603837771.0/4294967296.0,1,-nbitq), 
to_sfixed(145463083.0/4294967296.0,1,-nbitq), 
to_sfixed(-135446856.0/4294967296.0,1,-nbitq), 
to_sfixed(-247054043.0/4294967296.0,1,-nbitq), 
to_sfixed(-1575709059.0/4294967296.0,1,-nbitq), 
to_sfixed(-932654345.0/4294967296.0,1,-nbitq), 
to_sfixed(191460747.0/4294967296.0,1,-nbitq), 
to_sfixed(207152997.0/4294967296.0,1,-nbitq), 
to_sfixed(663817914.0/4294967296.0,1,-nbitq), 
to_sfixed(149698258.0/4294967296.0,1,-nbitq), 
to_sfixed(387463828.0/4294967296.0,1,-nbitq), 
to_sfixed(-245855174.0/4294967296.0,1,-nbitq), 
to_sfixed(399239262.0/4294967296.0,1,-nbitq), 
to_sfixed(-47029996.0/4294967296.0,1,-nbitq), 
to_sfixed(-1035935171.0/4294967296.0,1,-nbitq), 
to_sfixed(228118616.0/4294967296.0,1,-nbitq), 
to_sfixed(-101840862.0/4294967296.0,1,-nbitq), 
to_sfixed(-172866101.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-710710486.0/4294967296.0,1,-nbitq), 
to_sfixed(-455550977.0/4294967296.0,1,-nbitq), 
to_sfixed(770942336.0/4294967296.0,1,-nbitq), 
to_sfixed(896977536.0/4294967296.0,1,-nbitq), 
to_sfixed(578449525.0/4294967296.0,1,-nbitq), 
to_sfixed(-1085317814.0/4294967296.0,1,-nbitq), 
to_sfixed(241979937.0/4294967296.0,1,-nbitq), 
to_sfixed(-959410354.0/4294967296.0,1,-nbitq), 
to_sfixed(-1497930157.0/4294967296.0,1,-nbitq), 
to_sfixed(-127732194.0/4294967296.0,1,-nbitq), 
to_sfixed(-586077025.0/4294967296.0,1,-nbitq), 
to_sfixed(198862399.0/4294967296.0,1,-nbitq), 
to_sfixed(-791908886.0/4294967296.0,1,-nbitq), 
to_sfixed(-1190658402.0/4294967296.0,1,-nbitq), 
to_sfixed(-218629703.0/4294967296.0,1,-nbitq), 
to_sfixed(711885309.0/4294967296.0,1,-nbitq), 
to_sfixed(310065119.0/4294967296.0,1,-nbitq), 
to_sfixed(254055443.0/4294967296.0,1,-nbitq), 
to_sfixed(1981207053.0/4294967296.0,1,-nbitq), 
to_sfixed(641224252.0/4294967296.0,1,-nbitq), 
to_sfixed(182429888.0/4294967296.0,1,-nbitq), 
to_sfixed(124630543.0/4294967296.0,1,-nbitq), 
to_sfixed(420359888.0/4294967296.0,1,-nbitq), 
to_sfixed(219881459.0/4294967296.0,1,-nbitq), 
to_sfixed(320985086.0/4294967296.0,1,-nbitq), 
to_sfixed(225029057.0/4294967296.0,1,-nbitq), 
to_sfixed(238924954.0/4294967296.0,1,-nbitq), 
to_sfixed(920401406.0/4294967296.0,1,-nbitq), 
to_sfixed(1073377432.0/4294967296.0,1,-nbitq), 
to_sfixed(1094539962.0/4294967296.0,1,-nbitq), 
to_sfixed(-83279919.0/4294967296.0,1,-nbitq), 
to_sfixed(733314836.0/4294967296.0,1,-nbitq), 
to_sfixed(625288874.0/4294967296.0,1,-nbitq), 
to_sfixed(1375433526.0/4294967296.0,1,-nbitq), 
to_sfixed(-431233171.0/4294967296.0,1,-nbitq), 
to_sfixed(264633251.0/4294967296.0,1,-nbitq), 
to_sfixed(-958529137.0/4294967296.0,1,-nbitq), 
to_sfixed(32601647.0/4294967296.0,1,-nbitq), 
to_sfixed(114988828.0/4294967296.0,1,-nbitq), 
to_sfixed(9549225.0/4294967296.0,1,-nbitq), 
to_sfixed(257721635.0/4294967296.0,1,-nbitq), 
to_sfixed(-331364134.0/4294967296.0,1,-nbitq), 
to_sfixed(649281335.0/4294967296.0,1,-nbitq), 
to_sfixed(-133193989.0/4294967296.0,1,-nbitq), 
to_sfixed(-443800620.0/4294967296.0,1,-nbitq), 
to_sfixed(-598470912.0/4294967296.0,1,-nbitq), 
to_sfixed(295594115.0/4294967296.0,1,-nbitq), 
to_sfixed(791215384.0/4294967296.0,1,-nbitq), 
to_sfixed(44610480.0/4294967296.0,1,-nbitq), 
to_sfixed(507347822.0/4294967296.0,1,-nbitq), 
to_sfixed(-1271555930.0/4294967296.0,1,-nbitq), 
to_sfixed(268659674.0/4294967296.0,1,-nbitq), 
to_sfixed(-156297672.0/4294967296.0,1,-nbitq), 
to_sfixed(351259146.0/4294967296.0,1,-nbitq), 
to_sfixed(1365145855.0/4294967296.0,1,-nbitq), 
to_sfixed(386096681.0/4294967296.0,1,-nbitq), 
to_sfixed(137271320.0/4294967296.0,1,-nbitq), 
to_sfixed(-1003600796.0/4294967296.0,1,-nbitq), 
to_sfixed(-286545480.0/4294967296.0,1,-nbitq), 
to_sfixed(378700938.0/4294967296.0,1,-nbitq), 
to_sfixed(-431268423.0/4294967296.0,1,-nbitq), 
to_sfixed(-1814014295.0/4294967296.0,1,-nbitq), 
to_sfixed(-54406711.0/4294967296.0,1,-nbitq), 
to_sfixed(-276198817.0/4294967296.0,1,-nbitq), 
to_sfixed(-792156354.0/4294967296.0,1,-nbitq), 
to_sfixed(93941240.0/4294967296.0,1,-nbitq), 
to_sfixed(-143565724.0/4294967296.0,1,-nbitq), 
to_sfixed(-331192230.0/4294967296.0,1,-nbitq), 
to_sfixed(70405452.0/4294967296.0,1,-nbitq), 
to_sfixed(-224597692.0/4294967296.0,1,-nbitq), 
to_sfixed(208675429.0/4294967296.0,1,-nbitq), 
to_sfixed(-708163801.0/4294967296.0,1,-nbitq), 
to_sfixed(803276284.0/4294967296.0,1,-nbitq), 
to_sfixed(276771564.0/4294967296.0,1,-nbitq), 
to_sfixed(267326430.0/4294967296.0,1,-nbitq), 
to_sfixed(-739650880.0/4294967296.0,1,-nbitq), 
to_sfixed(-343201743.0/4294967296.0,1,-nbitq), 
to_sfixed(590429743.0/4294967296.0,1,-nbitq), 
to_sfixed(269548526.0/4294967296.0,1,-nbitq), 
to_sfixed(-31733957.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-750685939.0/4294967296.0,1,-nbitq), 
to_sfixed(-481721678.0/4294967296.0,1,-nbitq), 
to_sfixed(-734957860.0/4294967296.0,1,-nbitq), 
to_sfixed(324381217.0/4294967296.0,1,-nbitq), 
to_sfixed(1319145284.0/4294967296.0,1,-nbitq), 
to_sfixed(-626803716.0/4294967296.0,1,-nbitq), 
to_sfixed(226927119.0/4294967296.0,1,-nbitq), 
to_sfixed(-1885051089.0/4294967296.0,1,-nbitq), 
to_sfixed(-1185229510.0/4294967296.0,1,-nbitq), 
to_sfixed(-295668305.0/4294967296.0,1,-nbitq), 
to_sfixed(-698750810.0/4294967296.0,1,-nbitq), 
to_sfixed(548657723.0/4294967296.0,1,-nbitq), 
to_sfixed(-561484060.0/4294967296.0,1,-nbitq), 
to_sfixed(-713987632.0/4294967296.0,1,-nbitq), 
to_sfixed(-162298290.0/4294967296.0,1,-nbitq), 
to_sfixed(1660196142.0/4294967296.0,1,-nbitq), 
to_sfixed(-366868504.0/4294967296.0,1,-nbitq), 
to_sfixed(252952129.0/4294967296.0,1,-nbitq), 
to_sfixed(1765620301.0/4294967296.0,1,-nbitq), 
to_sfixed(653074790.0/4294967296.0,1,-nbitq), 
to_sfixed(232512215.0/4294967296.0,1,-nbitq), 
to_sfixed(-224736535.0/4294967296.0,1,-nbitq), 
to_sfixed(446407862.0/4294967296.0,1,-nbitq), 
to_sfixed(462405790.0/4294967296.0,1,-nbitq), 
to_sfixed(99906407.0/4294967296.0,1,-nbitq), 
to_sfixed(-191096497.0/4294967296.0,1,-nbitq), 
to_sfixed(-97607042.0/4294967296.0,1,-nbitq), 
to_sfixed(780010883.0/4294967296.0,1,-nbitq), 
to_sfixed(-742134643.0/4294967296.0,1,-nbitq), 
to_sfixed(1521926372.0/4294967296.0,1,-nbitq), 
to_sfixed(1005680965.0/4294967296.0,1,-nbitq), 
to_sfixed(873572960.0/4294967296.0,1,-nbitq), 
to_sfixed(583109496.0/4294967296.0,1,-nbitq), 
to_sfixed(763226206.0/4294967296.0,1,-nbitq), 
to_sfixed(-264269129.0/4294967296.0,1,-nbitq), 
to_sfixed(1840804433.0/4294967296.0,1,-nbitq), 
to_sfixed(-1482511197.0/4294967296.0,1,-nbitq), 
to_sfixed(-203509421.0/4294967296.0,1,-nbitq), 
to_sfixed(-122426063.0/4294967296.0,1,-nbitq), 
to_sfixed(-318122778.0/4294967296.0,1,-nbitq), 
to_sfixed(-169651609.0/4294967296.0,1,-nbitq), 
to_sfixed(-291126333.0/4294967296.0,1,-nbitq), 
to_sfixed(-219961368.0/4294967296.0,1,-nbitq), 
to_sfixed(1062755836.0/4294967296.0,1,-nbitq), 
to_sfixed(-662171617.0/4294967296.0,1,-nbitq), 
to_sfixed(130203385.0/4294967296.0,1,-nbitq), 
to_sfixed(-161122651.0/4294967296.0,1,-nbitq), 
to_sfixed(34509851.0/4294967296.0,1,-nbitq), 
to_sfixed(11573671.0/4294967296.0,1,-nbitq), 
to_sfixed(4261342.0/4294967296.0,1,-nbitq), 
to_sfixed(-683172692.0/4294967296.0,1,-nbitq), 
to_sfixed(-356756777.0/4294967296.0,1,-nbitq), 
to_sfixed(-796941938.0/4294967296.0,1,-nbitq), 
to_sfixed(229177345.0/4294967296.0,1,-nbitq), 
to_sfixed(2370731464.0/4294967296.0,1,-nbitq), 
to_sfixed(92795511.0/4294967296.0,1,-nbitq), 
to_sfixed(-408929346.0/4294967296.0,1,-nbitq), 
to_sfixed(-575264921.0/4294967296.0,1,-nbitq), 
to_sfixed(-204288345.0/4294967296.0,1,-nbitq), 
to_sfixed(-319793226.0/4294967296.0,1,-nbitq), 
to_sfixed(-434617880.0/4294967296.0,1,-nbitq), 
to_sfixed(-1226314462.0/4294967296.0,1,-nbitq), 
to_sfixed(194023816.0/4294967296.0,1,-nbitq), 
to_sfixed(-120315100.0/4294967296.0,1,-nbitq), 
to_sfixed(-81980739.0/4294967296.0,1,-nbitq), 
to_sfixed(72442639.0/4294967296.0,1,-nbitq), 
to_sfixed(1662233038.0/4294967296.0,1,-nbitq), 
to_sfixed(-148628507.0/4294967296.0,1,-nbitq), 
to_sfixed(-342871586.0/4294967296.0,1,-nbitq), 
to_sfixed(-313199994.0/4294967296.0,1,-nbitq), 
to_sfixed(274544270.0/4294967296.0,1,-nbitq), 
to_sfixed(-471129532.0/4294967296.0,1,-nbitq), 
to_sfixed(530624546.0/4294967296.0,1,-nbitq), 
to_sfixed(365829551.0/4294967296.0,1,-nbitq), 
to_sfixed(52121146.0/4294967296.0,1,-nbitq), 
to_sfixed(12021390.0/4294967296.0,1,-nbitq), 
to_sfixed(-70895460.0/4294967296.0,1,-nbitq), 
to_sfixed(527498728.0/4294967296.0,1,-nbitq), 
to_sfixed(1315002944.0/4294967296.0,1,-nbitq), 
to_sfixed(-169108811.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-403277922.0/4294967296.0,1,-nbitq), 
to_sfixed(-214076099.0/4294967296.0,1,-nbitq), 
to_sfixed(-1098141149.0/4294967296.0,1,-nbitq), 
to_sfixed(882035929.0/4294967296.0,1,-nbitq), 
to_sfixed(534154248.0/4294967296.0,1,-nbitq), 
to_sfixed(125292759.0/4294967296.0,1,-nbitq), 
to_sfixed(714083064.0/4294967296.0,1,-nbitq), 
to_sfixed(-972505504.0/4294967296.0,1,-nbitq), 
to_sfixed(-1760063036.0/4294967296.0,1,-nbitq), 
to_sfixed(-361207627.0/4294967296.0,1,-nbitq), 
to_sfixed(-501177016.0/4294967296.0,1,-nbitq), 
to_sfixed(1004794018.0/4294967296.0,1,-nbitq), 
to_sfixed(-1156743371.0/4294967296.0,1,-nbitq), 
to_sfixed(-1914166035.0/4294967296.0,1,-nbitq), 
to_sfixed(179528173.0/4294967296.0,1,-nbitq), 
to_sfixed(1312040098.0/4294967296.0,1,-nbitq), 
to_sfixed(146277424.0/4294967296.0,1,-nbitq), 
to_sfixed(-376751850.0/4294967296.0,1,-nbitq), 
to_sfixed(-162367985.0/4294967296.0,1,-nbitq), 
to_sfixed(43976307.0/4294967296.0,1,-nbitq), 
to_sfixed(184945797.0/4294967296.0,1,-nbitq), 
to_sfixed(-510278007.0/4294967296.0,1,-nbitq), 
to_sfixed(1439764192.0/4294967296.0,1,-nbitq), 
to_sfixed(650178070.0/4294967296.0,1,-nbitq), 
to_sfixed(-288948237.0/4294967296.0,1,-nbitq), 
to_sfixed(403735504.0/4294967296.0,1,-nbitq), 
to_sfixed(-155073963.0/4294967296.0,1,-nbitq), 
to_sfixed(-605194139.0/4294967296.0,1,-nbitq), 
to_sfixed(-1132037704.0/4294967296.0,1,-nbitq), 
to_sfixed(808952447.0/4294967296.0,1,-nbitq), 
to_sfixed(1076869081.0/4294967296.0,1,-nbitq), 
to_sfixed(-135328774.0/4294967296.0,1,-nbitq), 
to_sfixed(666252149.0/4294967296.0,1,-nbitq), 
to_sfixed(401683239.0/4294967296.0,1,-nbitq), 
to_sfixed(703031420.0/4294967296.0,1,-nbitq), 
to_sfixed(2167261619.0/4294967296.0,1,-nbitq), 
to_sfixed(-575910703.0/4294967296.0,1,-nbitq), 
to_sfixed(-802618281.0/4294967296.0,1,-nbitq), 
to_sfixed(-94290608.0/4294967296.0,1,-nbitq), 
to_sfixed(163038770.0/4294967296.0,1,-nbitq), 
to_sfixed(218919219.0/4294967296.0,1,-nbitq), 
to_sfixed(-1130062760.0/4294967296.0,1,-nbitq), 
to_sfixed(-1511714061.0/4294967296.0,1,-nbitq), 
to_sfixed(1112420223.0/4294967296.0,1,-nbitq), 
to_sfixed(-889450167.0/4294967296.0,1,-nbitq), 
to_sfixed(-72845448.0/4294967296.0,1,-nbitq), 
to_sfixed(-271866568.0/4294967296.0,1,-nbitq), 
to_sfixed(14336213.0/4294967296.0,1,-nbitq), 
to_sfixed(-371733559.0/4294967296.0,1,-nbitq), 
to_sfixed(-176029814.0/4294967296.0,1,-nbitq), 
to_sfixed(-876165811.0/4294967296.0,1,-nbitq), 
to_sfixed(105833549.0/4294967296.0,1,-nbitq), 
to_sfixed(-1528903672.0/4294967296.0,1,-nbitq), 
to_sfixed(-107503970.0/4294967296.0,1,-nbitq), 
to_sfixed(2100789390.0/4294967296.0,1,-nbitq), 
to_sfixed(307606224.0/4294967296.0,1,-nbitq), 
to_sfixed(-198203276.0/4294967296.0,1,-nbitq), 
to_sfixed(-68086907.0/4294967296.0,1,-nbitq), 
to_sfixed(-209580850.0/4294967296.0,1,-nbitq), 
to_sfixed(-164006645.0/4294967296.0,1,-nbitq), 
to_sfixed(147591840.0/4294967296.0,1,-nbitq), 
to_sfixed(-737564869.0/4294967296.0,1,-nbitq), 
to_sfixed(-158327882.0/4294967296.0,1,-nbitq), 
to_sfixed(299456372.0/4294967296.0,1,-nbitq), 
to_sfixed(-129261855.0/4294967296.0,1,-nbitq), 
to_sfixed(-341618451.0/4294967296.0,1,-nbitq), 
to_sfixed(481458808.0/4294967296.0,1,-nbitq), 
to_sfixed(434536149.0/4294967296.0,1,-nbitq), 
to_sfixed(-110708175.0/4294967296.0,1,-nbitq), 
to_sfixed(-574462937.0/4294967296.0,1,-nbitq), 
to_sfixed(185087848.0/4294967296.0,1,-nbitq), 
to_sfixed(18283814.0/4294967296.0,1,-nbitq), 
to_sfixed(607016252.0/4294967296.0,1,-nbitq), 
to_sfixed(242368198.0/4294967296.0,1,-nbitq), 
to_sfixed(413088276.0/4294967296.0,1,-nbitq), 
to_sfixed(-224399834.0/4294967296.0,1,-nbitq), 
to_sfixed(-729552104.0/4294967296.0,1,-nbitq), 
to_sfixed(-118229455.0/4294967296.0,1,-nbitq), 
to_sfixed(516418775.0/4294967296.0,1,-nbitq), 
to_sfixed(214189132.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(103813209.0/4294967296.0,1,-nbitq), 
to_sfixed(290494440.0/4294967296.0,1,-nbitq), 
to_sfixed(314661470.0/4294967296.0,1,-nbitq), 
to_sfixed(380639991.0/4294967296.0,1,-nbitq), 
to_sfixed(-1784142384.0/4294967296.0,1,-nbitq), 
to_sfixed(-62564324.0/4294967296.0,1,-nbitq), 
to_sfixed(314284656.0/4294967296.0,1,-nbitq), 
to_sfixed(-284919811.0/4294967296.0,1,-nbitq), 
to_sfixed(-637769608.0/4294967296.0,1,-nbitq), 
to_sfixed(-382884393.0/4294967296.0,1,-nbitq), 
to_sfixed(-939852986.0/4294967296.0,1,-nbitq), 
to_sfixed(713962389.0/4294967296.0,1,-nbitq), 
to_sfixed(-1066739750.0/4294967296.0,1,-nbitq), 
to_sfixed(-2538482147.0/4294967296.0,1,-nbitq), 
to_sfixed(-145879152.0/4294967296.0,1,-nbitq), 
to_sfixed(406520375.0/4294967296.0,1,-nbitq), 
to_sfixed(102285004.0/4294967296.0,1,-nbitq), 
to_sfixed(340219934.0/4294967296.0,1,-nbitq), 
to_sfixed(-1321231076.0/4294967296.0,1,-nbitq), 
to_sfixed(-130907302.0/4294967296.0,1,-nbitq), 
to_sfixed(314348879.0/4294967296.0,1,-nbitq), 
to_sfixed(-975962975.0/4294967296.0,1,-nbitq), 
to_sfixed(484555195.0/4294967296.0,1,-nbitq), 
to_sfixed(-1050520460.0/4294967296.0,1,-nbitq), 
to_sfixed(137651685.0/4294967296.0,1,-nbitq), 
to_sfixed(1190957751.0/4294967296.0,1,-nbitq), 
to_sfixed(-632155617.0/4294967296.0,1,-nbitq), 
to_sfixed(-1099561312.0/4294967296.0,1,-nbitq), 
to_sfixed(-33156996.0/4294967296.0,1,-nbitq), 
to_sfixed(21416493.0/4294967296.0,1,-nbitq), 
to_sfixed(883072672.0/4294967296.0,1,-nbitq), 
to_sfixed(-101479362.0/4294967296.0,1,-nbitq), 
to_sfixed(541084131.0/4294967296.0,1,-nbitq), 
to_sfixed(-410846384.0/4294967296.0,1,-nbitq), 
to_sfixed(1125883730.0/4294967296.0,1,-nbitq), 
to_sfixed(599069860.0/4294967296.0,1,-nbitq), 
to_sfixed(580978003.0/4294967296.0,1,-nbitq), 
to_sfixed(-1034044965.0/4294967296.0,1,-nbitq), 
to_sfixed(254377700.0/4294967296.0,1,-nbitq), 
to_sfixed(-290126681.0/4294967296.0,1,-nbitq), 
to_sfixed(81431073.0/4294967296.0,1,-nbitq), 
to_sfixed(-255079892.0/4294967296.0,1,-nbitq), 
to_sfixed(-2280206727.0/4294967296.0,1,-nbitq), 
to_sfixed(305031402.0/4294967296.0,1,-nbitq), 
to_sfixed(-157098878.0/4294967296.0,1,-nbitq), 
to_sfixed(-912862935.0/4294967296.0,1,-nbitq), 
to_sfixed(-89675318.0/4294967296.0,1,-nbitq), 
to_sfixed(-194515760.0/4294967296.0,1,-nbitq), 
to_sfixed(-108660536.0/4294967296.0,1,-nbitq), 
to_sfixed(-299445499.0/4294967296.0,1,-nbitq), 
to_sfixed(-662354425.0/4294967296.0,1,-nbitq), 
to_sfixed(-737941447.0/4294967296.0,1,-nbitq), 
to_sfixed(-1084727141.0/4294967296.0,1,-nbitq), 
to_sfixed(-649263943.0/4294967296.0,1,-nbitq), 
to_sfixed(228817702.0/4294967296.0,1,-nbitq), 
to_sfixed(135854234.0/4294967296.0,1,-nbitq), 
to_sfixed(-628351447.0/4294967296.0,1,-nbitq), 
to_sfixed(-69097006.0/4294967296.0,1,-nbitq), 
to_sfixed(-110119395.0/4294967296.0,1,-nbitq), 
to_sfixed(369473216.0/4294967296.0,1,-nbitq), 
to_sfixed(-451787805.0/4294967296.0,1,-nbitq), 
to_sfixed(660408020.0/4294967296.0,1,-nbitq), 
to_sfixed(114837093.0/4294967296.0,1,-nbitq), 
to_sfixed(-40128429.0/4294967296.0,1,-nbitq), 
to_sfixed(14498338.0/4294967296.0,1,-nbitq), 
to_sfixed(-166031754.0/4294967296.0,1,-nbitq), 
to_sfixed(519535196.0/4294967296.0,1,-nbitq), 
to_sfixed(1520574456.0/4294967296.0,1,-nbitq), 
to_sfixed(299591293.0/4294967296.0,1,-nbitq), 
to_sfixed(-379073130.0/4294967296.0,1,-nbitq), 
to_sfixed(1083155135.0/4294967296.0,1,-nbitq), 
to_sfixed(-92789682.0/4294967296.0,1,-nbitq), 
to_sfixed(-770783577.0/4294967296.0,1,-nbitq), 
to_sfixed(-240424730.0/4294967296.0,1,-nbitq), 
to_sfixed(49337631.0/4294967296.0,1,-nbitq), 
to_sfixed(223529259.0/4294967296.0,1,-nbitq), 
to_sfixed(-59690547.0/4294967296.0,1,-nbitq), 
to_sfixed(-442169492.0/4294967296.0,1,-nbitq), 
to_sfixed(128890680.0/4294967296.0,1,-nbitq), 
to_sfixed(-205785892.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(146008191.0/4294967296.0,1,-nbitq), 
to_sfixed(883229755.0/4294967296.0,1,-nbitq), 
to_sfixed(449539365.0/4294967296.0,1,-nbitq), 
to_sfixed(-215436508.0/4294967296.0,1,-nbitq), 
to_sfixed(-2521999204.0/4294967296.0,1,-nbitq), 
to_sfixed(62016159.0/4294967296.0,1,-nbitq), 
to_sfixed(282151312.0/4294967296.0,1,-nbitq), 
to_sfixed(327273379.0/4294967296.0,1,-nbitq), 
to_sfixed(-168225996.0/4294967296.0,1,-nbitq), 
to_sfixed(225028567.0/4294967296.0,1,-nbitq), 
to_sfixed(-41028167.0/4294967296.0,1,-nbitq), 
to_sfixed(823515345.0/4294967296.0,1,-nbitq), 
to_sfixed(-1073310875.0/4294967296.0,1,-nbitq), 
to_sfixed(-2848152386.0/4294967296.0,1,-nbitq), 
to_sfixed(-372724326.0/4294967296.0,1,-nbitq), 
to_sfixed(-120546412.0/4294967296.0,1,-nbitq), 
to_sfixed(373758732.0/4294967296.0,1,-nbitq), 
to_sfixed(319449576.0/4294967296.0,1,-nbitq), 
to_sfixed(-1172928501.0/4294967296.0,1,-nbitq), 
to_sfixed(2272274.0/4294967296.0,1,-nbitq), 
to_sfixed(208240746.0/4294967296.0,1,-nbitq), 
to_sfixed(-139378585.0/4294967296.0,1,-nbitq), 
to_sfixed(1109670755.0/4294967296.0,1,-nbitq), 
to_sfixed(-1853573567.0/4294967296.0,1,-nbitq), 
to_sfixed(-105918182.0/4294967296.0,1,-nbitq), 
to_sfixed(893774887.0/4294967296.0,1,-nbitq), 
to_sfixed(-777172699.0/4294967296.0,1,-nbitq), 
to_sfixed(-559378125.0/4294967296.0,1,-nbitq), 
to_sfixed(191182702.0/4294967296.0,1,-nbitq), 
to_sfixed(32951745.0/4294967296.0,1,-nbitq), 
to_sfixed(-1496297115.0/4294967296.0,1,-nbitq), 
to_sfixed(-11270909.0/4294967296.0,1,-nbitq), 
to_sfixed(1241458431.0/4294967296.0,1,-nbitq), 
to_sfixed(-602539917.0/4294967296.0,1,-nbitq), 
to_sfixed(1605088397.0/4294967296.0,1,-nbitq), 
to_sfixed(-243260758.0/4294967296.0,1,-nbitq), 
to_sfixed(-195946753.0/4294967296.0,1,-nbitq), 
to_sfixed(-669238634.0/4294967296.0,1,-nbitq), 
to_sfixed(690807575.0/4294967296.0,1,-nbitq), 
to_sfixed(75447587.0/4294967296.0,1,-nbitq), 
to_sfixed(1078544135.0/4294967296.0,1,-nbitq), 
to_sfixed(-266187354.0/4294967296.0,1,-nbitq), 
to_sfixed(-2222620923.0/4294967296.0,1,-nbitq), 
to_sfixed(770877583.0/4294967296.0,1,-nbitq), 
to_sfixed(-214359797.0/4294967296.0,1,-nbitq), 
to_sfixed(-605294161.0/4294967296.0,1,-nbitq), 
to_sfixed(-369437532.0/4294967296.0,1,-nbitq), 
to_sfixed(-7557354.0/4294967296.0,1,-nbitq), 
to_sfixed(60419970.0/4294967296.0,1,-nbitq), 
to_sfixed(574625752.0/4294967296.0,1,-nbitq), 
to_sfixed(-437663148.0/4294967296.0,1,-nbitq), 
to_sfixed(-187497542.0/4294967296.0,1,-nbitq), 
to_sfixed(-769391086.0/4294967296.0,1,-nbitq), 
to_sfixed(-994590045.0/4294967296.0,1,-nbitq), 
to_sfixed(-1175883845.0/4294967296.0,1,-nbitq), 
to_sfixed(137196642.0/4294967296.0,1,-nbitq), 
to_sfixed(-647721156.0/4294967296.0,1,-nbitq), 
to_sfixed(769281739.0/4294967296.0,1,-nbitq), 
to_sfixed(182544030.0/4294967296.0,1,-nbitq), 
to_sfixed(268343825.0/4294967296.0,1,-nbitq), 
to_sfixed(212856389.0/4294967296.0,1,-nbitq), 
to_sfixed(969354144.0/4294967296.0,1,-nbitq), 
to_sfixed(-623372192.0/4294967296.0,1,-nbitq), 
to_sfixed(-207494325.0/4294967296.0,1,-nbitq), 
to_sfixed(-81326191.0/4294967296.0,1,-nbitq), 
to_sfixed(-109124930.0/4294967296.0,1,-nbitq), 
to_sfixed(87122185.0/4294967296.0,1,-nbitq), 
to_sfixed(1387789663.0/4294967296.0,1,-nbitq), 
to_sfixed(193317727.0/4294967296.0,1,-nbitq), 
to_sfixed(386538525.0/4294967296.0,1,-nbitq), 
to_sfixed(2339147163.0/4294967296.0,1,-nbitq), 
to_sfixed(412055112.0/4294967296.0,1,-nbitq), 
to_sfixed(-1291014391.0/4294967296.0,1,-nbitq), 
to_sfixed(-148929209.0/4294967296.0,1,-nbitq), 
to_sfixed(-100044001.0/4294967296.0,1,-nbitq), 
to_sfixed(-379667974.0/4294967296.0,1,-nbitq), 
to_sfixed(-161945635.0/4294967296.0,1,-nbitq), 
to_sfixed(1051258.0/4294967296.0,1,-nbitq), 
to_sfixed(-8072719.0/4294967296.0,1,-nbitq), 
to_sfixed(-157233945.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(290945641.0/4294967296.0,1,-nbitq), 
to_sfixed(648225503.0/4294967296.0,1,-nbitq), 
to_sfixed(587170810.0/4294967296.0,1,-nbitq), 
to_sfixed(535964139.0/4294967296.0,1,-nbitq), 
to_sfixed(-2260879572.0/4294967296.0,1,-nbitq), 
to_sfixed(831266992.0/4294967296.0,1,-nbitq), 
to_sfixed(118994294.0/4294967296.0,1,-nbitq), 
to_sfixed(644893168.0/4294967296.0,1,-nbitq), 
to_sfixed(-48321643.0/4294967296.0,1,-nbitq), 
to_sfixed(80278358.0/4294967296.0,1,-nbitq), 
to_sfixed(237441555.0/4294967296.0,1,-nbitq), 
to_sfixed(1182963622.0/4294967296.0,1,-nbitq), 
to_sfixed(87415117.0/4294967296.0,1,-nbitq), 
to_sfixed(-1230921956.0/4294967296.0,1,-nbitq), 
to_sfixed(284162728.0/4294967296.0,1,-nbitq), 
to_sfixed(43787848.0/4294967296.0,1,-nbitq), 
to_sfixed(-391373808.0/4294967296.0,1,-nbitq), 
to_sfixed(179097690.0/4294967296.0,1,-nbitq), 
to_sfixed(-1264280939.0/4294967296.0,1,-nbitq), 
to_sfixed(763235481.0/4294967296.0,1,-nbitq), 
to_sfixed(70928121.0/4294967296.0,1,-nbitq), 
to_sfixed(-433994465.0/4294967296.0,1,-nbitq), 
to_sfixed(50960731.0/4294967296.0,1,-nbitq), 
to_sfixed(-923166472.0/4294967296.0,1,-nbitq), 
to_sfixed(342292372.0/4294967296.0,1,-nbitq), 
to_sfixed(822714042.0/4294967296.0,1,-nbitq), 
to_sfixed(-749890500.0/4294967296.0,1,-nbitq), 
to_sfixed(112767631.0/4294967296.0,1,-nbitq), 
to_sfixed(-145569854.0/4294967296.0,1,-nbitq), 
to_sfixed(413005905.0/4294967296.0,1,-nbitq), 
to_sfixed(-1023604749.0/4294967296.0,1,-nbitq), 
to_sfixed(-1148394236.0/4294967296.0,1,-nbitq), 
to_sfixed(1055765942.0/4294967296.0,1,-nbitq), 
to_sfixed(46122953.0/4294967296.0,1,-nbitq), 
to_sfixed(1259164112.0/4294967296.0,1,-nbitq), 
to_sfixed(187316362.0/4294967296.0,1,-nbitq), 
to_sfixed(-269880905.0/4294967296.0,1,-nbitq), 
to_sfixed(-32264165.0/4294967296.0,1,-nbitq), 
to_sfixed(84804876.0/4294967296.0,1,-nbitq), 
to_sfixed(20137529.0/4294967296.0,1,-nbitq), 
to_sfixed(451633496.0/4294967296.0,1,-nbitq), 
to_sfixed(1262773399.0/4294967296.0,1,-nbitq), 
to_sfixed(-1624835350.0/4294967296.0,1,-nbitq), 
to_sfixed(1506955488.0/4294967296.0,1,-nbitq), 
to_sfixed(46194723.0/4294967296.0,1,-nbitq), 
to_sfixed(-967994542.0/4294967296.0,1,-nbitq), 
to_sfixed(178366815.0/4294967296.0,1,-nbitq), 
to_sfixed(-204734736.0/4294967296.0,1,-nbitq), 
to_sfixed(-210334921.0/4294967296.0,1,-nbitq), 
to_sfixed(-67070872.0/4294967296.0,1,-nbitq), 
to_sfixed(-59124246.0/4294967296.0,1,-nbitq), 
to_sfixed(647888999.0/4294967296.0,1,-nbitq), 
to_sfixed(-285251953.0/4294967296.0,1,-nbitq), 
to_sfixed(-718418680.0/4294967296.0,1,-nbitq), 
to_sfixed(-923730084.0/4294967296.0,1,-nbitq), 
to_sfixed(52857220.0/4294967296.0,1,-nbitq), 
to_sfixed(-869106389.0/4294967296.0,1,-nbitq), 
to_sfixed(160575063.0/4294967296.0,1,-nbitq), 
to_sfixed(166388838.0/4294967296.0,1,-nbitq), 
to_sfixed(338030256.0/4294967296.0,1,-nbitq), 
to_sfixed(273141195.0/4294967296.0,1,-nbitq), 
to_sfixed(1221890410.0/4294967296.0,1,-nbitq), 
to_sfixed(-1001658072.0/4294967296.0,1,-nbitq), 
to_sfixed(-247948720.0/4294967296.0,1,-nbitq), 
to_sfixed(-416504092.0/4294967296.0,1,-nbitq), 
to_sfixed(273949763.0/4294967296.0,1,-nbitq), 
to_sfixed(-1896604093.0/4294967296.0,1,-nbitq), 
to_sfixed(-849472421.0/4294967296.0,1,-nbitq), 
to_sfixed(191042847.0/4294967296.0,1,-nbitq), 
to_sfixed(128305898.0/4294967296.0,1,-nbitq), 
to_sfixed(1681672431.0/4294967296.0,1,-nbitq), 
to_sfixed(-178438416.0/4294967296.0,1,-nbitq), 
to_sfixed(-1037604562.0/4294967296.0,1,-nbitq), 
to_sfixed(329749516.0/4294967296.0,1,-nbitq), 
to_sfixed(287549936.0/4294967296.0,1,-nbitq), 
to_sfixed(-126502906.0/4294967296.0,1,-nbitq), 
to_sfixed(540221379.0/4294967296.0,1,-nbitq), 
to_sfixed(263217277.0/4294967296.0,1,-nbitq), 
to_sfixed(-501940334.0/4294967296.0,1,-nbitq), 
to_sfixed(24102514.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(134247336.0/4294967296.0,1,-nbitq), 
to_sfixed(1207036127.0/4294967296.0,1,-nbitq), 
to_sfixed(755632005.0/4294967296.0,1,-nbitq), 
to_sfixed(1222465967.0/4294967296.0,1,-nbitq), 
to_sfixed(-2236047266.0/4294967296.0,1,-nbitq), 
to_sfixed(582697222.0/4294967296.0,1,-nbitq), 
to_sfixed(-351681804.0/4294967296.0,1,-nbitq), 
to_sfixed(717269131.0/4294967296.0,1,-nbitq), 
to_sfixed(-189786377.0/4294967296.0,1,-nbitq), 
to_sfixed(198580547.0/4294967296.0,1,-nbitq), 
to_sfixed(172488631.0/4294967296.0,1,-nbitq), 
to_sfixed(1014979151.0/4294967296.0,1,-nbitq), 
to_sfixed(-197392440.0/4294967296.0,1,-nbitq), 
to_sfixed(-1413561074.0/4294967296.0,1,-nbitq), 
to_sfixed(243714320.0/4294967296.0,1,-nbitq), 
to_sfixed(-460168919.0/4294967296.0,1,-nbitq), 
to_sfixed(-89681233.0/4294967296.0,1,-nbitq), 
to_sfixed(-145876504.0/4294967296.0,1,-nbitq), 
to_sfixed(-1679945179.0/4294967296.0,1,-nbitq), 
to_sfixed(168655063.0/4294967296.0,1,-nbitq), 
to_sfixed(70516542.0/4294967296.0,1,-nbitq), 
to_sfixed(-575917700.0/4294967296.0,1,-nbitq), 
to_sfixed(-732196695.0/4294967296.0,1,-nbitq), 
to_sfixed(-992319148.0/4294967296.0,1,-nbitq), 
to_sfixed(-166232806.0/4294967296.0,1,-nbitq), 
to_sfixed(377289151.0/4294967296.0,1,-nbitq), 
to_sfixed(-736849701.0/4294967296.0,1,-nbitq), 
to_sfixed(253536989.0/4294967296.0,1,-nbitq), 
to_sfixed(-487501519.0/4294967296.0,1,-nbitq), 
to_sfixed(960577637.0/4294967296.0,1,-nbitq), 
to_sfixed(-878789469.0/4294967296.0,1,-nbitq), 
to_sfixed(-81696517.0/4294967296.0,1,-nbitq), 
to_sfixed(928819248.0/4294967296.0,1,-nbitq), 
to_sfixed(574388634.0/4294967296.0,1,-nbitq), 
to_sfixed(-1035922.0/4294967296.0,1,-nbitq), 
to_sfixed(-685204360.0/4294967296.0,1,-nbitq), 
to_sfixed(-212593153.0/4294967296.0,1,-nbitq), 
to_sfixed(-94848564.0/4294967296.0,1,-nbitq), 
to_sfixed(161560253.0/4294967296.0,1,-nbitq), 
to_sfixed(-280873798.0/4294967296.0,1,-nbitq), 
to_sfixed(-86882316.0/4294967296.0,1,-nbitq), 
to_sfixed(1482705134.0/4294967296.0,1,-nbitq), 
to_sfixed(-1656268045.0/4294967296.0,1,-nbitq), 
to_sfixed(657085779.0/4294967296.0,1,-nbitq), 
to_sfixed(259090819.0/4294967296.0,1,-nbitq), 
to_sfixed(-316885048.0/4294967296.0,1,-nbitq), 
to_sfixed(-306853263.0/4294967296.0,1,-nbitq), 
to_sfixed(266688290.0/4294967296.0,1,-nbitq), 
to_sfixed(-391693283.0/4294967296.0,1,-nbitq), 
to_sfixed(256796762.0/4294967296.0,1,-nbitq), 
to_sfixed(499947775.0/4294967296.0,1,-nbitq), 
to_sfixed(711456953.0/4294967296.0,1,-nbitq), 
to_sfixed(413036131.0/4294967296.0,1,-nbitq), 
to_sfixed(159425382.0/4294967296.0,1,-nbitq), 
to_sfixed(-1340954841.0/4294967296.0,1,-nbitq), 
to_sfixed(303718084.0/4294967296.0,1,-nbitq), 
to_sfixed(-327687656.0/4294967296.0,1,-nbitq), 
to_sfixed(1256063681.0/4294967296.0,1,-nbitq), 
to_sfixed(73396451.0/4294967296.0,1,-nbitq), 
to_sfixed(23023322.0/4294967296.0,1,-nbitq), 
to_sfixed(382750983.0/4294967296.0,1,-nbitq), 
to_sfixed(430033168.0/4294967296.0,1,-nbitq), 
to_sfixed(268297076.0/4294967296.0,1,-nbitq), 
to_sfixed(-46919508.0/4294967296.0,1,-nbitq), 
to_sfixed(-751436375.0/4294967296.0,1,-nbitq), 
to_sfixed(274230699.0/4294967296.0,1,-nbitq), 
to_sfixed(-2761049464.0/4294967296.0,1,-nbitq), 
to_sfixed(-680111043.0/4294967296.0,1,-nbitq), 
to_sfixed(-65448959.0/4294967296.0,1,-nbitq), 
to_sfixed(430873461.0/4294967296.0,1,-nbitq), 
to_sfixed(809648473.0/4294967296.0,1,-nbitq), 
to_sfixed(-426106598.0/4294967296.0,1,-nbitq), 
to_sfixed(-354534154.0/4294967296.0,1,-nbitq), 
to_sfixed(359480465.0/4294967296.0,1,-nbitq), 
to_sfixed(-329781140.0/4294967296.0,1,-nbitq), 
to_sfixed(1171474319.0/4294967296.0,1,-nbitq), 
to_sfixed(-56690677.0/4294967296.0,1,-nbitq), 
to_sfixed(-289676935.0/4294967296.0,1,-nbitq), 
to_sfixed(182086131.0/4294967296.0,1,-nbitq), 
to_sfixed(9682434.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(124251791.0/4294967296.0,1,-nbitq), 
to_sfixed(126688169.0/4294967296.0,1,-nbitq), 
to_sfixed(1158844911.0/4294967296.0,1,-nbitq), 
to_sfixed(1062958705.0/4294967296.0,1,-nbitq), 
to_sfixed(-1616116603.0/4294967296.0,1,-nbitq), 
to_sfixed(159124156.0/4294967296.0,1,-nbitq), 
to_sfixed(-53724409.0/4294967296.0,1,-nbitq), 
to_sfixed(412528919.0/4294967296.0,1,-nbitq), 
to_sfixed(-409862879.0/4294967296.0,1,-nbitq), 
to_sfixed(-419413730.0/4294967296.0,1,-nbitq), 
to_sfixed(83234603.0/4294967296.0,1,-nbitq), 
to_sfixed(250490917.0/4294967296.0,1,-nbitq), 
to_sfixed(444687633.0/4294967296.0,1,-nbitq), 
to_sfixed(31689324.0/4294967296.0,1,-nbitq), 
to_sfixed(454631443.0/4294967296.0,1,-nbitq), 
to_sfixed(-137462055.0/4294967296.0,1,-nbitq), 
to_sfixed(-133516466.0/4294967296.0,1,-nbitq), 
to_sfixed(223291098.0/4294967296.0,1,-nbitq), 
to_sfixed(-1625522143.0/4294967296.0,1,-nbitq), 
to_sfixed(34922285.0/4294967296.0,1,-nbitq), 
to_sfixed(-429566525.0/4294967296.0,1,-nbitq), 
to_sfixed(-281483305.0/4294967296.0,1,-nbitq), 
to_sfixed(-612926447.0/4294967296.0,1,-nbitq), 
to_sfixed(-427171160.0/4294967296.0,1,-nbitq), 
to_sfixed(-148399147.0/4294967296.0,1,-nbitq), 
to_sfixed(106296832.0/4294967296.0,1,-nbitq), 
to_sfixed(-502233762.0/4294967296.0,1,-nbitq), 
to_sfixed(145368422.0/4294967296.0,1,-nbitq), 
to_sfixed(-131807911.0/4294967296.0,1,-nbitq), 
to_sfixed(2017768549.0/4294967296.0,1,-nbitq), 
to_sfixed(-778280816.0/4294967296.0,1,-nbitq), 
to_sfixed(840731862.0/4294967296.0,1,-nbitq), 
to_sfixed(730379934.0/4294967296.0,1,-nbitq), 
to_sfixed(481190401.0/4294967296.0,1,-nbitq), 
to_sfixed(374803838.0/4294967296.0,1,-nbitq), 
to_sfixed(-636376052.0/4294967296.0,1,-nbitq), 
to_sfixed(-257236722.0/4294967296.0,1,-nbitq), 
to_sfixed(-53512648.0/4294967296.0,1,-nbitq), 
to_sfixed(-15756170.0/4294967296.0,1,-nbitq), 
to_sfixed(-146408081.0/4294967296.0,1,-nbitq), 
to_sfixed(-710189869.0/4294967296.0,1,-nbitq), 
to_sfixed(1387715985.0/4294967296.0,1,-nbitq), 
to_sfixed(-1425424113.0/4294967296.0,1,-nbitq), 
to_sfixed(-37789695.0/4294967296.0,1,-nbitq), 
to_sfixed(-138177577.0/4294967296.0,1,-nbitq), 
to_sfixed(-1080218017.0/4294967296.0,1,-nbitq), 
to_sfixed(162158099.0/4294967296.0,1,-nbitq), 
to_sfixed(360783536.0/4294967296.0,1,-nbitq), 
to_sfixed(-735122994.0/4294967296.0,1,-nbitq), 
to_sfixed(352015101.0/4294967296.0,1,-nbitq), 
to_sfixed(312762281.0/4294967296.0,1,-nbitq), 
to_sfixed(61522080.0/4294967296.0,1,-nbitq), 
to_sfixed(301946327.0/4294967296.0,1,-nbitq), 
to_sfixed(565336501.0/4294967296.0,1,-nbitq), 
to_sfixed(-2037069265.0/4294967296.0,1,-nbitq), 
to_sfixed(1240008172.0/4294967296.0,1,-nbitq), 
to_sfixed(-741666707.0/4294967296.0,1,-nbitq), 
to_sfixed(1212460574.0/4294967296.0,1,-nbitq), 
to_sfixed(116520525.0/4294967296.0,1,-nbitq), 
to_sfixed(60886041.0/4294967296.0,1,-nbitq), 
to_sfixed(516354345.0/4294967296.0,1,-nbitq), 
to_sfixed(-62906339.0/4294967296.0,1,-nbitq), 
to_sfixed(421700149.0/4294967296.0,1,-nbitq), 
to_sfixed(-642129758.0/4294967296.0,1,-nbitq), 
to_sfixed(88899643.0/4294967296.0,1,-nbitq), 
to_sfixed(321154857.0/4294967296.0,1,-nbitq), 
to_sfixed(-1262703661.0/4294967296.0,1,-nbitq), 
to_sfixed(-478524813.0/4294967296.0,1,-nbitq), 
to_sfixed(-368250733.0/4294967296.0,1,-nbitq), 
to_sfixed(278050887.0/4294967296.0,1,-nbitq), 
to_sfixed(980084109.0/4294967296.0,1,-nbitq), 
to_sfixed(-682816801.0/4294967296.0,1,-nbitq), 
to_sfixed(-1245094542.0/4294967296.0,1,-nbitq), 
to_sfixed(-62329966.0/4294967296.0,1,-nbitq), 
to_sfixed(227654215.0/4294967296.0,1,-nbitq), 
to_sfixed(1371368027.0/4294967296.0,1,-nbitq), 
to_sfixed(-88559750.0/4294967296.0,1,-nbitq), 
to_sfixed(91632772.0/4294967296.0,1,-nbitq), 
to_sfixed(301934551.0/4294967296.0,1,-nbitq), 
to_sfixed(-217172958.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-409727312.0/4294967296.0,1,-nbitq), 
to_sfixed(-159317673.0/4294967296.0,1,-nbitq), 
to_sfixed(472213568.0/4294967296.0,1,-nbitq), 
to_sfixed(1964395349.0/4294967296.0,1,-nbitq), 
to_sfixed(-928597226.0/4294967296.0,1,-nbitq), 
to_sfixed(837747884.0/4294967296.0,1,-nbitq), 
to_sfixed(-93148420.0/4294967296.0,1,-nbitq), 
to_sfixed(113857156.0/4294967296.0,1,-nbitq), 
to_sfixed(355416445.0/4294967296.0,1,-nbitq), 
to_sfixed(236096047.0/4294967296.0,1,-nbitq), 
to_sfixed(-600255986.0/4294967296.0,1,-nbitq), 
to_sfixed(1403001985.0/4294967296.0,1,-nbitq), 
to_sfixed(505825316.0/4294967296.0,1,-nbitq), 
to_sfixed(-273350466.0/4294967296.0,1,-nbitq), 
to_sfixed(262836737.0/4294967296.0,1,-nbitq), 
to_sfixed(661067368.0/4294967296.0,1,-nbitq), 
to_sfixed(-96882042.0/4294967296.0,1,-nbitq), 
to_sfixed(843356.0/4294967296.0,1,-nbitq), 
to_sfixed(-1470620024.0/4294967296.0,1,-nbitq), 
to_sfixed(-154999862.0/4294967296.0,1,-nbitq), 
to_sfixed(315288538.0/4294967296.0,1,-nbitq), 
to_sfixed(-26712192.0/4294967296.0,1,-nbitq), 
to_sfixed(-701186675.0/4294967296.0,1,-nbitq), 
to_sfixed(-169286452.0/4294967296.0,1,-nbitq), 
to_sfixed(-361797771.0/4294967296.0,1,-nbitq), 
to_sfixed(-222969943.0/4294967296.0,1,-nbitq), 
to_sfixed(27043822.0/4294967296.0,1,-nbitq), 
to_sfixed(357346418.0/4294967296.0,1,-nbitq), 
to_sfixed(-729902419.0/4294967296.0,1,-nbitq), 
to_sfixed(1718896173.0/4294967296.0,1,-nbitq), 
to_sfixed(-36997226.0/4294967296.0,1,-nbitq), 
to_sfixed(330620112.0/4294967296.0,1,-nbitq), 
to_sfixed(849852758.0/4294967296.0,1,-nbitq), 
to_sfixed(131340838.0/4294967296.0,1,-nbitq), 
to_sfixed(-159035509.0/4294967296.0,1,-nbitq), 
to_sfixed(336533532.0/4294967296.0,1,-nbitq), 
to_sfixed(-471226801.0/4294967296.0,1,-nbitq), 
to_sfixed(-39396174.0/4294967296.0,1,-nbitq), 
to_sfixed(-22929801.0/4294967296.0,1,-nbitq), 
to_sfixed(582308340.0/4294967296.0,1,-nbitq), 
to_sfixed(-890411464.0/4294967296.0,1,-nbitq), 
to_sfixed(674642215.0/4294967296.0,1,-nbitq), 
to_sfixed(-1416165302.0/4294967296.0,1,-nbitq), 
to_sfixed(-13267168.0/4294967296.0,1,-nbitq), 
to_sfixed(354261528.0/4294967296.0,1,-nbitq), 
to_sfixed(-2173229620.0/4294967296.0,1,-nbitq), 
to_sfixed(-110830781.0/4294967296.0,1,-nbitq), 
to_sfixed(40172851.0/4294967296.0,1,-nbitq), 
to_sfixed(-107310036.0/4294967296.0,1,-nbitq), 
to_sfixed(486217361.0/4294967296.0,1,-nbitq), 
to_sfixed(851682457.0/4294967296.0,1,-nbitq), 
to_sfixed(866847040.0/4294967296.0,1,-nbitq), 
to_sfixed(1026390765.0/4294967296.0,1,-nbitq), 
to_sfixed(653883439.0/4294967296.0,1,-nbitq), 
to_sfixed(-1779280492.0/4294967296.0,1,-nbitq), 
to_sfixed(1531806738.0/4294967296.0,1,-nbitq), 
to_sfixed(-26676937.0/4294967296.0,1,-nbitq), 
to_sfixed(1346219380.0/4294967296.0,1,-nbitq), 
to_sfixed(-85775066.0/4294967296.0,1,-nbitq), 
to_sfixed(-28127293.0/4294967296.0,1,-nbitq), 
to_sfixed(512732867.0/4294967296.0,1,-nbitq), 
to_sfixed(240888222.0/4294967296.0,1,-nbitq), 
to_sfixed(313319043.0/4294967296.0,1,-nbitq), 
to_sfixed(-417606877.0/4294967296.0,1,-nbitq), 
to_sfixed(81295510.0/4294967296.0,1,-nbitq), 
to_sfixed(99192634.0/4294967296.0,1,-nbitq), 
to_sfixed(-626016801.0/4294967296.0,1,-nbitq), 
to_sfixed(-775656320.0/4294967296.0,1,-nbitq), 
to_sfixed(-46159563.0/4294967296.0,1,-nbitq), 
to_sfixed(773816227.0/4294967296.0,1,-nbitq), 
to_sfixed(721876061.0/4294967296.0,1,-nbitq), 
to_sfixed(-608174326.0/4294967296.0,1,-nbitq), 
to_sfixed(-180574734.0/4294967296.0,1,-nbitq), 
to_sfixed(-143911750.0/4294967296.0,1,-nbitq), 
to_sfixed(166364663.0/4294967296.0,1,-nbitq), 
to_sfixed(600817423.0/4294967296.0,1,-nbitq), 
to_sfixed(91182712.0/4294967296.0,1,-nbitq), 
to_sfixed(134635855.0/4294967296.0,1,-nbitq), 
to_sfixed(63377518.0/4294967296.0,1,-nbitq), 
to_sfixed(298274285.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-293144087.0/4294967296.0,1,-nbitq), 
to_sfixed(-817902699.0/4294967296.0,1,-nbitq), 
to_sfixed(596274864.0/4294967296.0,1,-nbitq), 
to_sfixed(1974518023.0/4294967296.0,1,-nbitq), 
to_sfixed(-943835575.0/4294967296.0,1,-nbitq), 
to_sfixed(11179351.0/4294967296.0,1,-nbitq), 
to_sfixed(191733057.0/4294967296.0,1,-nbitq), 
to_sfixed(266960333.0/4294967296.0,1,-nbitq), 
to_sfixed(803669963.0/4294967296.0,1,-nbitq), 
to_sfixed(254670347.0/4294967296.0,1,-nbitq), 
to_sfixed(-420564855.0/4294967296.0,1,-nbitq), 
to_sfixed(562343414.0/4294967296.0,1,-nbitq), 
to_sfixed(851061597.0/4294967296.0,1,-nbitq), 
to_sfixed(-543323954.0/4294967296.0,1,-nbitq), 
to_sfixed(-20512398.0/4294967296.0,1,-nbitq), 
to_sfixed(794939056.0/4294967296.0,1,-nbitq), 
to_sfixed(-318903614.0/4294967296.0,1,-nbitq), 
to_sfixed(196705906.0/4294967296.0,1,-nbitq), 
to_sfixed(-743372426.0/4294967296.0,1,-nbitq), 
to_sfixed(-562228796.0/4294967296.0,1,-nbitq), 
to_sfixed(-183048068.0/4294967296.0,1,-nbitq), 
to_sfixed(242287777.0/4294967296.0,1,-nbitq), 
to_sfixed(-1410751387.0/4294967296.0,1,-nbitq), 
to_sfixed(-107031321.0/4294967296.0,1,-nbitq), 
to_sfixed(244964127.0/4294967296.0,1,-nbitq), 
to_sfixed(-427989118.0/4294967296.0,1,-nbitq), 
to_sfixed(-48649767.0/4294967296.0,1,-nbitq), 
to_sfixed(280301862.0/4294967296.0,1,-nbitq), 
to_sfixed(-668284627.0/4294967296.0,1,-nbitq), 
to_sfixed(2303932280.0/4294967296.0,1,-nbitq), 
to_sfixed(324098926.0/4294967296.0,1,-nbitq), 
to_sfixed(216825598.0/4294967296.0,1,-nbitq), 
to_sfixed(306901825.0/4294967296.0,1,-nbitq), 
to_sfixed(87677180.0/4294967296.0,1,-nbitq), 
to_sfixed(-13525473.0/4294967296.0,1,-nbitq), 
to_sfixed(-170094936.0/4294967296.0,1,-nbitq), 
to_sfixed(-131797617.0/4294967296.0,1,-nbitq), 
to_sfixed(239689041.0/4294967296.0,1,-nbitq), 
to_sfixed(6831839.0/4294967296.0,1,-nbitq), 
to_sfixed(-154424833.0/4294967296.0,1,-nbitq), 
to_sfixed(-722634810.0/4294967296.0,1,-nbitq), 
to_sfixed(49366872.0/4294967296.0,1,-nbitq), 
to_sfixed(-1695897386.0/4294967296.0,1,-nbitq), 
to_sfixed(127494193.0/4294967296.0,1,-nbitq), 
to_sfixed(103140177.0/4294967296.0,1,-nbitq), 
to_sfixed(-1721111226.0/4294967296.0,1,-nbitq), 
to_sfixed(-109286103.0/4294967296.0,1,-nbitq), 
to_sfixed(-123488823.0/4294967296.0,1,-nbitq), 
to_sfixed(144231260.0/4294967296.0,1,-nbitq), 
to_sfixed(267226445.0/4294967296.0,1,-nbitq), 
to_sfixed(219115290.0/4294967296.0,1,-nbitq), 
to_sfixed(-11042574.0/4294967296.0,1,-nbitq), 
to_sfixed(1877963752.0/4294967296.0,1,-nbitq), 
to_sfixed(266774184.0/4294967296.0,1,-nbitq), 
to_sfixed(-1658663345.0/4294967296.0,1,-nbitq), 
to_sfixed(1654908736.0/4294967296.0,1,-nbitq), 
to_sfixed(105805942.0/4294967296.0,1,-nbitq), 
to_sfixed(652625196.0/4294967296.0,1,-nbitq), 
to_sfixed(110923764.0/4294967296.0,1,-nbitq), 
to_sfixed(-70278135.0/4294967296.0,1,-nbitq), 
to_sfixed(535702329.0/4294967296.0,1,-nbitq), 
to_sfixed(-408898702.0/4294967296.0,1,-nbitq), 
to_sfixed(121816733.0/4294967296.0,1,-nbitq), 
to_sfixed(-28812570.0/4294967296.0,1,-nbitq), 
to_sfixed(85437797.0/4294967296.0,1,-nbitq), 
to_sfixed(341298573.0/4294967296.0,1,-nbitq), 
to_sfixed(840535930.0/4294967296.0,1,-nbitq), 
to_sfixed(-123028758.0/4294967296.0,1,-nbitq), 
to_sfixed(-116326413.0/4294967296.0,1,-nbitq), 
to_sfixed(814977460.0/4294967296.0,1,-nbitq), 
to_sfixed(627307030.0/4294967296.0,1,-nbitq), 
to_sfixed(505545700.0/4294967296.0,1,-nbitq), 
to_sfixed(-546040759.0/4294967296.0,1,-nbitq), 
to_sfixed(-217852590.0/4294967296.0,1,-nbitq), 
to_sfixed(145805719.0/4294967296.0,1,-nbitq), 
to_sfixed(213822252.0/4294967296.0,1,-nbitq), 
to_sfixed(500833477.0/4294967296.0,1,-nbitq), 
to_sfixed(-544022356.0/4294967296.0,1,-nbitq), 
to_sfixed(313183648.0/4294967296.0,1,-nbitq), 
to_sfixed(-263933765.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-33647934.0/4294967296.0,1,-nbitq), 
to_sfixed(-103233397.0/4294967296.0,1,-nbitq), 
to_sfixed(-786023471.0/4294967296.0,1,-nbitq), 
to_sfixed(1729029879.0/4294967296.0,1,-nbitq), 
to_sfixed(-489660782.0/4294967296.0,1,-nbitq), 
to_sfixed(-609311358.0/4294967296.0,1,-nbitq), 
to_sfixed(-232944897.0/4294967296.0,1,-nbitq), 
to_sfixed(669018292.0/4294967296.0,1,-nbitq), 
to_sfixed(-529293043.0/4294967296.0,1,-nbitq), 
to_sfixed(-243990047.0/4294967296.0,1,-nbitq), 
to_sfixed(-261602094.0/4294967296.0,1,-nbitq), 
to_sfixed(438351827.0/4294967296.0,1,-nbitq), 
to_sfixed(248782494.0/4294967296.0,1,-nbitq), 
to_sfixed(-831762700.0/4294967296.0,1,-nbitq), 
to_sfixed(118968356.0/4294967296.0,1,-nbitq), 
to_sfixed(195741090.0/4294967296.0,1,-nbitq), 
to_sfixed(-50341674.0/4294967296.0,1,-nbitq), 
to_sfixed(-344228745.0/4294967296.0,1,-nbitq), 
to_sfixed(-986925057.0/4294967296.0,1,-nbitq), 
to_sfixed(-289292674.0/4294967296.0,1,-nbitq), 
to_sfixed(-300472679.0/4294967296.0,1,-nbitq), 
to_sfixed(-519911636.0/4294967296.0,1,-nbitq), 
to_sfixed(-1099504017.0/4294967296.0,1,-nbitq), 
to_sfixed(-348482923.0/4294967296.0,1,-nbitq), 
to_sfixed(-51306371.0/4294967296.0,1,-nbitq), 
to_sfixed(-457165007.0/4294967296.0,1,-nbitq), 
to_sfixed(-268405019.0/4294967296.0,1,-nbitq), 
to_sfixed(-184942685.0/4294967296.0,1,-nbitq), 
to_sfixed(-288874958.0/4294967296.0,1,-nbitq), 
to_sfixed(1230366996.0/4294967296.0,1,-nbitq), 
to_sfixed(1706796406.0/4294967296.0,1,-nbitq), 
to_sfixed(848110009.0/4294967296.0,1,-nbitq), 
to_sfixed(359589214.0/4294967296.0,1,-nbitq), 
to_sfixed(249556798.0/4294967296.0,1,-nbitq), 
to_sfixed(-232678657.0/4294967296.0,1,-nbitq), 
to_sfixed(94019473.0/4294967296.0,1,-nbitq), 
to_sfixed(67794923.0/4294967296.0,1,-nbitq), 
to_sfixed(-67550799.0/4294967296.0,1,-nbitq), 
to_sfixed(307110231.0/4294967296.0,1,-nbitq), 
to_sfixed(82917523.0/4294967296.0,1,-nbitq), 
to_sfixed(-173721601.0/4294967296.0,1,-nbitq), 
to_sfixed(-451462425.0/4294967296.0,1,-nbitq), 
to_sfixed(-1534053186.0/4294967296.0,1,-nbitq), 
to_sfixed(-609673300.0/4294967296.0,1,-nbitq), 
to_sfixed(-195980666.0/4294967296.0,1,-nbitq), 
to_sfixed(-775215041.0/4294967296.0,1,-nbitq), 
to_sfixed(-225969611.0/4294967296.0,1,-nbitq), 
to_sfixed(-58091906.0/4294967296.0,1,-nbitq), 
to_sfixed(-645109545.0/4294967296.0,1,-nbitq), 
to_sfixed(-651136978.0/4294967296.0,1,-nbitq), 
to_sfixed(749124304.0/4294967296.0,1,-nbitq), 
to_sfixed(292603689.0/4294967296.0,1,-nbitq), 
to_sfixed(2015864002.0/4294967296.0,1,-nbitq), 
to_sfixed(-502763887.0/4294967296.0,1,-nbitq), 
to_sfixed(-1068318653.0/4294967296.0,1,-nbitq), 
to_sfixed(604816820.0/4294967296.0,1,-nbitq), 
to_sfixed(153463634.0/4294967296.0,1,-nbitq), 
to_sfixed(1124687467.0/4294967296.0,1,-nbitq), 
to_sfixed(369719120.0/4294967296.0,1,-nbitq), 
to_sfixed(-148682215.0/4294967296.0,1,-nbitq), 
to_sfixed(378156403.0/4294967296.0,1,-nbitq), 
to_sfixed(-282765477.0/4294967296.0,1,-nbitq), 
to_sfixed(796989108.0/4294967296.0,1,-nbitq), 
to_sfixed(404009845.0/4294967296.0,1,-nbitq), 
to_sfixed(234371325.0/4294967296.0,1,-nbitq), 
to_sfixed(407992205.0/4294967296.0,1,-nbitq), 
to_sfixed(1406801691.0/4294967296.0,1,-nbitq), 
to_sfixed(209267871.0/4294967296.0,1,-nbitq), 
to_sfixed(214238199.0/4294967296.0,1,-nbitq), 
to_sfixed(773694219.0/4294967296.0,1,-nbitq), 
to_sfixed(544521350.0/4294967296.0,1,-nbitq), 
to_sfixed(-20739977.0/4294967296.0,1,-nbitq), 
to_sfixed(-236579751.0/4294967296.0,1,-nbitq), 
to_sfixed(-153237909.0/4294967296.0,1,-nbitq), 
to_sfixed(445964863.0/4294967296.0,1,-nbitq), 
to_sfixed(-285533859.0/4294967296.0,1,-nbitq), 
to_sfixed(244078588.0/4294967296.0,1,-nbitq), 
to_sfixed(68656113.0/4294967296.0,1,-nbitq), 
to_sfixed(477539827.0/4294967296.0,1,-nbitq), 
to_sfixed(164710472.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(160342154.0/4294967296.0,1,-nbitq), 
to_sfixed(-1507495392.0/4294967296.0,1,-nbitq), 
to_sfixed(332265059.0/4294967296.0,1,-nbitq), 
to_sfixed(1053504323.0/4294967296.0,1,-nbitq), 
to_sfixed(-1078749888.0/4294967296.0,1,-nbitq), 
to_sfixed(-1053929384.0/4294967296.0,1,-nbitq), 
to_sfixed(-61553269.0/4294967296.0,1,-nbitq), 
to_sfixed(855654125.0/4294967296.0,1,-nbitq), 
to_sfixed(-620690707.0/4294967296.0,1,-nbitq), 
to_sfixed(425080458.0/4294967296.0,1,-nbitq), 
to_sfixed(-351862042.0/4294967296.0,1,-nbitq), 
to_sfixed(-60156262.0/4294967296.0,1,-nbitq), 
to_sfixed(-454355236.0/4294967296.0,1,-nbitq), 
to_sfixed(-76141234.0/4294967296.0,1,-nbitq), 
to_sfixed(-259788786.0/4294967296.0,1,-nbitq), 
to_sfixed(798016577.0/4294967296.0,1,-nbitq), 
to_sfixed(140586151.0/4294967296.0,1,-nbitq), 
to_sfixed(-225633371.0/4294967296.0,1,-nbitq), 
to_sfixed(-1107309905.0/4294967296.0,1,-nbitq), 
to_sfixed(-58672888.0/4294967296.0,1,-nbitq), 
to_sfixed(-339522934.0/4294967296.0,1,-nbitq), 
to_sfixed(171221155.0/4294967296.0,1,-nbitq), 
to_sfixed(-734605919.0/4294967296.0,1,-nbitq), 
to_sfixed(-84599732.0/4294967296.0,1,-nbitq), 
to_sfixed(177437184.0/4294967296.0,1,-nbitq), 
to_sfixed(-482286392.0/4294967296.0,1,-nbitq), 
to_sfixed(-199091327.0/4294967296.0,1,-nbitq), 
to_sfixed(-260717006.0/4294967296.0,1,-nbitq), 
to_sfixed(265573116.0/4294967296.0,1,-nbitq), 
to_sfixed(1455738872.0/4294967296.0,1,-nbitq), 
to_sfixed(39321810.0/4294967296.0,1,-nbitq), 
to_sfixed(153426096.0/4294967296.0,1,-nbitq), 
to_sfixed(-297562399.0/4294967296.0,1,-nbitq), 
to_sfixed(804987766.0/4294967296.0,1,-nbitq), 
to_sfixed(-599238337.0/4294967296.0,1,-nbitq), 
to_sfixed(-22950757.0/4294967296.0,1,-nbitq), 
to_sfixed(-492546558.0/4294967296.0,1,-nbitq), 
to_sfixed(705746855.0/4294967296.0,1,-nbitq), 
to_sfixed(-269613640.0/4294967296.0,1,-nbitq), 
to_sfixed(58279964.0/4294967296.0,1,-nbitq), 
to_sfixed(-646171232.0/4294967296.0,1,-nbitq), 
to_sfixed(20453770.0/4294967296.0,1,-nbitq), 
to_sfixed(-1560695177.0/4294967296.0,1,-nbitq), 
to_sfixed(-1048942951.0/4294967296.0,1,-nbitq), 
to_sfixed(603019797.0/4294967296.0,1,-nbitq), 
to_sfixed(-672475242.0/4294967296.0,1,-nbitq), 
to_sfixed(-394246823.0/4294967296.0,1,-nbitq), 
to_sfixed(684622057.0/4294967296.0,1,-nbitq), 
to_sfixed(147427635.0/4294967296.0,1,-nbitq), 
to_sfixed(-780136883.0/4294967296.0,1,-nbitq), 
to_sfixed(379848654.0/4294967296.0,1,-nbitq), 
to_sfixed(651666550.0/4294967296.0,1,-nbitq), 
to_sfixed(894295924.0/4294967296.0,1,-nbitq), 
to_sfixed(104402939.0/4294967296.0,1,-nbitq), 
to_sfixed(-1516117542.0/4294967296.0,1,-nbitq), 
to_sfixed(909766381.0/4294967296.0,1,-nbitq), 
to_sfixed(-189905284.0/4294967296.0,1,-nbitq), 
to_sfixed(532666193.0/4294967296.0,1,-nbitq), 
to_sfixed(363375886.0/4294967296.0,1,-nbitq), 
to_sfixed(361499181.0/4294967296.0,1,-nbitq), 
to_sfixed(376826678.0/4294967296.0,1,-nbitq), 
to_sfixed(-506518767.0/4294967296.0,1,-nbitq), 
to_sfixed(573756874.0/4294967296.0,1,-nbitq), 
to_sfixed(365582348.0/4294967296.0,1,-nbitq), 
to_sfixed(406194472.0/4294967296.0,1,-nbitq), 
to_sfixed(334578412.0/4294967296.0,1,-nbitq), 
to_sfixed(891506517.0/4294967296.0,1,-nbitq), 
to_sfixed(-741266482.0/4294967296.0,1,-nbitq), 
to_sfixed(98681472.0/4294967296.0,1,-nbitq), 
to_sfixed(524097099.0/4294967296.0,1,-nbitq), 
to_sfixed(-64899218.0/4294967296.0,1,-nbitq), 
to_sfixed(-200808543.0/4294967296.0,1,-nbitq), 
to_sfixed(-520096323.0/4294967296.0,1,-nbitq), 
to_sfixed(111447825.0/4294967296.0,1,-nbitq), 
to_sfixed(-132849297.0/4294967296.0,1,-nbitq), 
to_sfixed(94646020.0/4294967296.0,1,-nbitq), 
to_sfixed(892577371.0/4294967296.0,1,-nbitq), 
to_sfixed(166346175.0/4294967296.0,1,-nbitq), 
to_sfixed(-219233444.0/4294967296.0,1,-nbitq), 
to_sfixed(-51380896.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(7816857.0/4294967296.0,1,-nbitq), 
to_sfixed(-1404937133.0/4294967296.0,1,-nbitq), 
to_sfixed(-191101051.0/4294967296.0,1,-nbitq), 
to_sfixed(693097421.0/4294967296.0,1,-nbitq), 
to_sfixed(-77514619.0/4294967296.0,1,-nbitq), 
to_sfixed(-738328541.0/4294967296.0,1,-nbitq), 
to_sfixed(-304074965.0/4294967296.0,1,-nbitq), 
to_sfixed(861994610.0/4294967296.0,1,-nbitq), 
to_sfixed(-727677354.0/4294967296.0,1,-nbitq), 
to_sfixed(-44809926.0/4294967296.0,1,-nbitq), 
to_sfixed(117813766.0/4294967296.0,1,-nbitq), 
to_sfixed(317767717.0/4294967296.0,1,-nbitq), 
to_sfixed(-116404619.0/4294967296.0,1,-nbitq), 
to_sfixed(361780426.0/4294967296.0,1,-nbitq), 
to_sfixed(-205072803.0/4294967296.0,1,-nbitq), 
to_sfixed(-4275690.0/4294967296.0,1,-nbitq), 
to_sfixed(-119853239.0/4294967296.0,1,-nbitq), 
to_sfixed(199679260.0/4294967296.0,1,-nbitq), 
to_sfixed(-383953422.0/4294967296.0,1,-nbitq), 
to_sfixed(-407153983.0/4294967296.0,1,-nbitq), 
to_sfixed(148963100.0/4294967296.0,1,-nbitq), 
to_sfixed(-591430669.0/4294967296.0,1,-nbitq), 
to_sfixed(-621307814.0/4294967296.0,1,-nbitq), 
to_sfixed(-330264154.0/4294967296.0,1,-nbitq), 
to_sfixed(418475009.0/4294967296.0,1,-nbitq), 
to_sfixed(-1247949805.0/4294967296.0,1,-nbitq), 
to_sfixed(-407707607.0/4294967296.0,1,-nbitq), 
to_sfixed(126662159.0/4294967296.0,1,-nbitq), 
to_sfixed(-449047441.0/4294967296.0,1,-nbitq), 
to_sfixed(1464306562.0/4294967296.0,1,-nbitq), 
to_sfixed(-180420778.0/4294967296.0,1,-nbitq), 
to_sfixed(24145821.0/4294967296.0,1,-nbitq), 
to_sfixed(-710878669.0/4294967296.0,1,-nbitq), 
to_sfixed(195827236.0/4294967296.0,1,-nbitq), 
to_sfixed(-96081524.0/4294967296.0,1,-nbitq), 
to_sfixed(-201293225.0/4294967296.0,1,-nbitq), 
to_sfixed(-328828108.0/4294967296.0,1,-nbitq), 
to_sfixed(1045435103.0/4294967296.0,1,-nbitq), 
to_sfixed(168865818.0/4294967296.0,1,-nbitq), 
to_sfixed(121347776.0/4294967296.0,1,-nbitq), 
to_sfixed(2909756.0/4294967296.0,1,-nbitq), 
to_sfixed(-478943496.0/4294967296.0,1,-nbitq), 
to_sfixed(-1108641812.0/4294967296.0,1,-nbitq), 
to_sfixed(-1221663168.0/4294967296.0,1,-nbitq), 
to_sfixed(11831266.0/4294967296.0,1,-nbitq), 
to_sfixed(-190995035.0/4294967296.0,1,-nbitq), 
to_sfixed(245397140.0/4294967296.0,1,-nbitq), 
to_sfixed(436080794.0/4294967296.0,1,-nbitq), 
to_sfixed(-142542018.0/4294967296.0,1,-nbitq), 
to_sfixed(-69082456.0/4294967296.0,1,-nbitq), 
to_sfixed(95471811.0/4294967296.0,1,-nbitq), 
to_sfixed(782734442.0/4294967296.0,1,-nbitq), 
to_sfixed(414430442.0/4294967296.0,1,-nbitq), 
to_sfixed(-596199179.0/4294967296.0,1,-nbitq), 
to_sfixed(-1714340822.0/4294967296.0,1,-nbitq), 
to_sfixed(191959537.0/4294967296.0,1,-nbitq), 
to_sfixed(-2150768.0/4294967296.0,1,-nbitq), 
to_sfixed(879754907.0/4294967296.0,1,-nbitq), 
to_sfixed(-127194378.0/4294967296.0,1,-nbitq), 
to_sfixed(303451278.0/4294967296.0,1,-nbitq), 
to_sfixed(216929598.0/4294967296.0,1,-nbitq), 
to_sfixed(-6140346.0/4294967296.0,1,-nbitq), 
to_sfixed(14162719.0/4294967296.0,1,-nbitq), 
to_sfixed(420999536.0/4294967296.0,1,-nbitq), 
to_sfixed(-56889276.0/4294967296.0,1,-nbitq), 
to_sfixed(167020450.0/4294967296.0,1,-nbitq), 
to_sfixed(710629278.0/4294967296.0,1,-nbitq), 
to_sfixed(-116592325.0/4294967296.0,1,-nbitq), 
to_sfixed(382160192.0/4294967296.0,1,-nbitq), 
to_sfixed(741522090.0/4294967296.0,1,-nbitq), 
to_sfixed(-428966872.0/4294967296.0,1,-nbitq), 
to_sfixed(-123371822.0/4294967296.0,1,-nbitq), 
to_sfixed(87559686.0/4294967296.0,1,-nbitq), 
to_sfixed(179138209.0/4294967296.0,1,-nbitq), 
to_sfixed(119730481.0/4294967296.0,1,-nbitq), 
to_sfixed(-179882240.0/4294967296.0,1,-nbitq), 
to_sfixed(-234869458.0/4294967296.0,1,-nbitq), 
to_sfixed(-57965125.0/4294967296.0,1,-nbitq), 
to_sfixed(-378378834.0/4294967296.0,1,-nbitq), 
to_sfixed(-144226356.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-166115172.0/4294967296.0,1,-nbitq), 
to_sfixed(-17861441.0/4294967296.0,1,-nbitq), 
to_sfixed(52581850.0/4294967296.0,1,-nbitq), 
to_sfixed(-655101160.0/4294967296.0,1,-nbitq), 
to_sfixed(-755727908.0/4294967296.0,1,-nbitq), 
to_sfixed(-531899452.0/4294967296.0,1,-nbitq), 
to_sfixed(-24865946.0/4294967296.0,1,-nbitq), 
to_sfixed(291174382.0/4294967296.0,1,-nbitq), 
to_sfixed(73124978.0/4294967296.0,1,-nbitq), 
to_sfixed(423132969.0/4294967296.0,1,-nbitq), 
to_sfixed(-17080390.0/4294967296.0,1,-nbitq), 
to_sfixed(87831894.0/4294967296.0,1,-nbitq), 
to_sfixed(-16665779.0/4294967296.0,1,-nbitq), 
to_sfixed(564257561.0/4294967296.0,1,-nbitq), 
to_sfixed(60010553.0/4294967296.0,1,-nbitq), 
to_sfixed(475596495.0/4294967296.0,1,-nbitq), 
to_sfixed(-241588429.0/4294967296.0,1,-nbitq), 
to_sfixed(147494520.0/4294967296.0,1,-nbitq), 
to_sfixed(-301219961.0/4294967296.0,1,-nbitq), 
to_sfixed(94976308.0/4294967296.0,1,-nbitq), 
to_sfixed(-138163306.0/4294967296.0,1,-nbitq), 
to_sfixed(-595493867.0/4294967296.0,1,-nbitq), 
to_sfixed(-680775674.0/4294967296.0,1,-nbitq), 
to_sfixed(48010872.0/4294967296.0,1,-nbitq), 
to_sfixed(-216716933.0/4294967296.0,1,-nbitq), 
to_sfixed(-1151106317.0/4294967296.0,1,-nbitq), 
to_sfixed(-230792422.0/4294967296.0,1,-nbitq), 
to_sfixed(-166892958.0/4294967296.0,1,-nbitq), 
to_sfixed(-123397475.0/4294967296.0,1,-nbitq), 
to_sfixed(564182291.0/4294967296.0,1,-nbitq), 
to_sfixed(-100330072.0/4294967296.0,1,-nbitq), 
to_sfixed(-173733109.0/4294967296.0,1,-nbitq), 
to_sfixed(-181205652.0/4294967296.0,1,-nbitq), 
to_sfixed(-135828723.0/4294967296.0,1,-nbitq), 
to_sfixed(-623389333.0/4294967296.0,1,-nbitq), 
to_sfixed(-459571072.0/4294967296.0,1,-nbitq), 
to_sfixed(104492394.0/4294967296.0,1,-nbitq), 
to_sfixed(425189173.0/4294967296.0,1,-nbitq), 
to_sfixed(-208714169.0/4294967296.0,1,-nbitq), 
to_sfixed(160912030.0/4294967296.0,1,-nbitq), 
to_sfixed(297045705.0/4294967296.0,1,-nbitq), 
to_sfixed(-432942446.0/4294967296.0,1,-nbitq), 
to_sfixed(-546239837.0/4294967296.0,1,-nbitq), 
to_sfixed(-1278730235.0/4294967296.0,1,-nbitq), 
to_sfixed(-47350342.0/4294967296.0,1,-nbitq), 
to_sfixed(-809056270.0/4294967296.0,1,-nbitq), 
to_sfixed(-102607946.0/4294967296.0,1,-nbitq), 
to_sfixed(200088142.0/4294967296.0,1,-nbitq), 
to_sfixed(328504724.0/4294967296.0,1,-nbitq), 
to_sfixed(213228467.0/4294967296.0,1,-nbitq), 
to_sfixed(-90951225.0/4294967296.0,1,-nbitq), 
to_sfixed(196958931.0/4294967296.0,1,-nbitq), 
to_sfixed(260830675.0/4294967296.0,1,-nbitq), 
to_sfixed(-83057762.0/4294967296.0,1,-nbitq), 
to_sfixed(-810226707.0/4294967296.0,1,-nbitq), 
to_sfixed(-89549683.0/4294967296.0,1,-nbitq), 
to_sfixed(341673018.0/4294967296.0,1,-nbitq), 
to_sfixed(188741272.0/4294967296.0,1,-nbitq), 
to_sfixed(-224780203.0/4294967296.0,1,-nbitq), 
to_sfixed(-64741339.0/4294967296.0,1,-nbitq), 
to_sfixed(192508133.0/4294967296.0,1,-nbitq), 
to_sfixed(-90662999.0/4294967296.0,1,-nbitq), 
to_sfixed(215504309.0/4294967296.0,1,-nbitq), 
to_sfixed(258332013.0/4294967296.0,1,-nbitq), 
to_sfixed(-90628046.0/4294967296.0,1,-nbitq), 
to_sfixed(148857049.0/4294967296.0,1,-nbitq), 
to_sfixed(310582811.0/4294967296.0,1,-nbitq), 
to_sfixed(315716205.0/4294967296.0,1,-nbitq), 
to_sfixed(366719291.0/4294967296.0,1,-nbitq), 
to_sfixed(584656405.0/4294967296.0,1,-nbitq), 
to_sfixed(1784294.0/4294967296.0,1,-nbitq), 
to_sfixed(-390500174.0/4294967296.0,1,-nbitq), 
to_sfixed(637314115.0/4294967296.0,1,-nbitq), 
to_sfixed(104201574.0/4294967296.0,1,-nbitq), 
to_sfixed(146606111.0/4294967296.0,1,-nbitq), 
to_sfixed(408768040.0/4294967296.0,1,-nbitq), 
to_sfixed(-607525881.0/4294967296.0,1,-nbitq), 
to_sfixed(-117578638.0/4294967296.0,1,-nbitq), 
to_sfixed(-36075390.0/4294967296.0,1,-nbitq), 
to_sfixed(-106256982.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(154931421.0/4294967296.0,1,-nbitq), 
to_sfixed(-239757003.0/4294967296.0,1,-nbitq), 
to_sfixed(420814356.0/4294967296.0,1,-nbitq), 
to_sfixed(-411508845.0/4294967296.0,1,-nbitq), 
to_sfixed(-353690089.0/4294967296.0,1,-nbitq), 
to_sfixed(-956293224.0/4294967296.0,1,-nbitq), 
to_sfixed(-335762786.0/4294967296.0,1,-nbitq), 
to_sfixed(732607557.0/4294967296.0,1,-nbitq), 
to_sfixed(-548065807.0/4294967296.0,1,-nbitq), 
to_sfixed(160833353.0/4294967296.0,1,-nbitq), 
to_sfixed(281296916.0/4294967296.0,1,-nbitq), 
to_sfixed(-269074496.0/4294967296.0,1,-nbitq), 
to_sfixed(-250144060.0/4294967296.0,1,-nbitq), 
to_sfixed(65452114.0/4294967296.0,1,-nbitq), 
to_sfixed(-168867078.0/4294967296.0,1,-nbitq), 
to_sfixed(-39325158.0/4294967296.0,1,-nbitq), 
to_sfixed(-423436747.0/4294967296.0,1,-nbitq), 
to_sfixed(211268283.0/4294967296.0,1,-nbitq), 
to_sfixed(298749433.0/4294967296.0,1,-nbitq), 
to_sfixed(366227887.0/4294967296.0,1,-nbitq), 
to_sfixed(-107878408.0/4294967296.0,1,-nbitq), 
to_sfixed(-75653553.0/4294967296.0,1,-nbitq), 
to_sfixed(-491554257.0/4294967296.0,1,-nbitq), 
to_sfixed(439081563.0/4294967296.0,1,-nbitq), 
to_sfixed(110651038.0/4294967296.0,1,-nbitq), 
to_sfixed(-293099915.0/4294967296.0,1,-nbitq), 
to_sfixed(156370933.0/4294967296.0,1,-nbitq), 
to_sfixed(-121835479.0/4294967296.0,1,-nbitq), 
to_sfixed(280626444.0/4294967296.0,1,-nbitq), 
to_sfixed(200675642.0/4294967296.0,1,-nbitq), 
to_sfixed(-323688083.0/4294967296.0,1,-nbitq), 
to_sfixed(-100654622.0/4294967296.0,1,-nbitq), 
to_sfixed(-82528710.0/4294967296.0,1,-nbitq), 
to_sfixed(-202677358.0/4294967296.0,1,-nbitq), 
to_sfixed(-695038556.0/4294967296.0,1,-nbitq), 
to_sfixed(-577904239.0/4294967296.0,1,-nbitq), 
to_sfixed(-473194827.0/4294967296.0,1,-nbitq), 
to_sfixed(-346941111.0/4294967296.0,1,-nbitq), 
to_sfixed(-18548460.0/4294967296.0,1,-nbitq), 
to_sfixed(-182432813.0/4294967296.0,1,-nbitq), 
to_sfixed(-393412627.0/4294967296.0,1,-nbitq), 
to_sfixed(-168870230.0/4294967296.0,1,-nbitq), 
to_sfixed(78271138.0/4294967296.0,1,-nbitq), 
to_sfixed(-597746265.0/4294967296.0,1,-nbitq), 
to_sfixed(-133207113.0/4294967296.0,1,-nbitq), 
to_sfixed(-75199335.0/4294967296.0,1,-nbitq), 
to_sfixed(-328400397.0/4294967296.0,1,-nbitq), 
to_sfixed(-274169634.0/4294967296.0,1,-nbitq), 
to_sfixed(268691494.0/4294967296.0,1,-nbitq), 
to_sfixed(-179887003.0/4294967296.0,1,-nbitq), 
to_sfixed(270797167.0/4294967296.0,1,-nbitq), 
to_sfixed(370655763.0/4294967296.0,1,-nbitq), 
to_sfixed(267795608.0/4294967296.0,1,-nbitq), 
to_sfixed(108255184.0/4294967296.0,1,-nbitq), 
to_sfixed(20396661.0/4294967296.0,1,-nbitq), 
to_sfixed(-247564012.0/4294967296.0,1,-nbitq), 
to_sfixed(300229475.0/4294967296.0,1,-nbitq), 
to_sfixed(288661725.0/4294967296.0,1,-nbitq), 
to_sfixed(-107197972.0/4294967296.0,1,-nbitq), 
to_sfixed(-163374410.0/4294967296.0,1,-nbitq), 
to_sfixed(411930759.0/4294967296.0,1,-nbitq), 
to_sfixed(90731831.0/4294967296.0,1,-nbitq), 
to_sfixed(40264149.0/4294967296.0,1,-nbitq), 
to_sfixed(382159479.0/4294967296.0,1,-nbitq), 
to_sfixed(134357438.0/4294967296.0,1,-nbitq), 
to_sfixed(-198199314.0/4294967296.0,1,-nbitq), 
to_sfixed(508315261.0/4294967296.0,1,-nbitq), 
to_sfixed(-46717278.0/4294967296.0,1,-nbitq), 
to_sfixed(-328724935.0/4294967296.0,1,-nbitq), 
to_sfixed(81007086.0/4294967296.0,1,-nbitq), 
to_sfixed(179465832.0/4294967296.0,1,-nbitq), 
to_sfixed(108071216.0/4294967296.0,1,-nbitq), 
to_sfixed(149548780.0/4294967296.0,1,-nbitq), 
to_sfixed(265917836.0/4294967296.0,1,-nbitq), 
to_sfixed(-70949795.0/4294967296.0,1,-nbitq), 
to_sfixed(14318197.0/4294967296.0,1,-nbitq), 
to_sfixed(-596886573.0/4294967296.0,1,-nbitq), 
to_sfixed(-337545559.0/4294967296.0,1,-nbitq), 
to_sfixed(97390567.0/4294967296.0,1,-nbitq), 
to_sfixed(309452623.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(323866873.0/4294967296.0,1,-nbitq), 
to_sfixed(-305544472.0/4294967296.0,1,-nbitq), 
to_sfixed(670629870.0/4294967296.0,1,-nbitq), 
to_sfixed(80426146.0/4294967296.0,1,-nbitq), 
to_sfixed(80508180.0/4294967296.0,1,-nbitq), 
to_sfixed(-91984055.0/4294967296.0,1,-nbitq), 
to_sfixed(162477967.0/4294967296.0,1,-nbitq), 
to_sfixed(541033623.0/4294967296.0,1,-nbitq), 
to_sfixed(270551003.0/4294967296.0,1,-nbitq), 
to_sfixed(-176107151.0/4294967296.0,1,-nbitq), 
to_sfixed(301924074.0/4294967296.0,1,-nbitq), 
to_sfixed(41259901.0/4294967296.0,1,-nbitq), 
to_sfixed(132074148.0/4294967296.0,1,-nbitq), 
to_sfixed(145426750.0/4294967296.0,1,-nbitq), 
to_sfixed(-103202126.0/4294967296.0,1,-nbitq), 
to_sfixed(230101103.0/4294967296.0,1,-nbitq), 
to_sfixed(72795827.0/4294967296.0,1,-nbitq), 
to_sfixed(-69824969.0/4294967296.0,1,-nbitq), 
to_sfixed(-198361835.0/4294967296.0,1,-nbitq), 
to_sfixed(-369460896.0/4294967296.0,1,-nbitq), 
to_sfixed(-163660183.0/4294967296.0,1,-nbitq), 
to_sfixed(272739743.0/4294967296.0,1,-nbitq), 
to_sfixed(133288725.0/4294967296.0,1,-nbitq), 
to_sfixed(527003038.0/4294967296.0,1,-nbitq), 
to_sfixed(-93523162.0/4294967296.0,1,-nbitq), 
to_sfixed(-237830097.0/4294967296.0,1,-nbitq), 
to_sfixed(74121713.0/4294967296.0,1,-nbitq), 
to_sfixed(-9568933.0/4294967296.0,1,-nbitq), 
to_sfixed(64133416.0/4294967296.0,1,-nbitq), 
to_sfixed(84496545.0/4294967296.0,1,-nbitq), 
to_sfixed(-513062096.0/4294967296.0,1,-nbitq), 
to_sfixed(-202950891.0/4294967296.0,1,-nbitq), 
to_sfixed(141465674.0/4294967296.0,1,-nbitq), 
to_sfixed(-144684261.0/4294967296.0,1,-nbitq), 
to_sfixed(-280917344.0/4294967296.0,1,-nbitq), 
to_sfixed(185108653.0/4294967296.0,1,-nbitq), 
to_sfixed(-300473826.0/4294967296.0,1,-nbitq), 
to_sfixed(-382159153.0/4294967296.0,1,-nbitq), 
to_sfixed(189919366.0/4294967296.0,1,-nbitq), 
to_sfixed(-260757656.0/4294967296.0,1,-nbitq), 
to_sfixed(-473836301.0/4294967296.0,1,-nbitq), 
to_sfixed(55435366.0/4294967296.0,1,-nbitq), 
to_sfixed(-131154105.0/4294967296.0,1,-nbitq), 
to_sfixed(185197805.0/4294967296.0,1,-nbitq), 
to_sfixed(-247306530.0/4294967296.0,1,-nbitq), 
to_sfixed(-215516703.0/4294967296.0,1,-nbitq), 
to_sfixed(30202014.0/4294967296.0,1,-nbitq), 
to_sfixed(-400770168.0/4294967296.0,1,-nbitq), 
to_sfixed(42975500.0/4294967296.0,1,-nbitq), 
to_sfixed(225839303.0/4294967296.0,1,-nbitq), 
to_sfixed(-59726814.0/4294967296.0,1,-nbitq), 
to_sfixed(450004823.0/4294967296.0,1,-nbitq), 
to_sfixed(-437994372.0/4294967296.0,1,-nbitq), 
to_sfixed(282614985.0/4294967296.0,1,-nbitq), 
to_sfixed(4203536.0/4294967296.0,1,-nbitq), 
to_sfixed(336311730.0/4294967296.0,1,-nbitq), 
to_sfixed(-193174452.0/4294967296.0,1,-nbitq), 
to_sfixed(208597734.0/4294967296.0,1,-nbitq), 
to_sfixed(-50172878.0/4294967296.0,1,-nbitq), 
to_sfixed(-144416080.0/4294967296.0,1,-nbitq), 
to_sfixed(349022449.0/4294967296.0,1,-nbitq), 
to_sfixed(-127451581.0/4294967296.0,1,-nbitq), 
to_sfixed(-58693351.0/4294967296.0,1,-nbitq), 
to_sfixed(-344874497.0/4294967296.0,1,-nbitq), 
to_sfixed(-327209845.0/4294967296.0,1,-nbitq), 
to_sfixed(328051358.0/4294967296.0,1,-nbitq), 
to_sfixed(648134282.0/4294967296.0,1,-nbitq), 
to_sfixed(60954388.0/4294967296.0,1,-nbitq), 
to_sfixed(242316196.0/4294967296.0,1,-nbitq), 
to_sfixed(95259382.0/4294967296.0,1,-nbitq), 
to_sfixed(-145818834.0/4294967296.0,1,-nbitq), 
to_sfixed(-132822631.0/4294967296.0,1,-nbitq), 
to_sfixed(-220809117.0/4294967296.0,1,-nbitq), 
to_sfixed(267891194.0/4294967296.0,1,-nbitq), 
to_sfixed(-193382209.0/4294967296.0,1,-nbitq), 
to_sfixed(-534627751.0/4294967296.0,1,-nbitq), 
to_sfixed(-411598917.0/4294967296.0,1,-nbitq), 
to_sfixed(-346312119.0/4294967296.0,1,-nbitq), 
to_sfixed(320511247.0/4294967296.0,1,-nbitq), 
to_sfixed(293744016.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(244067872.0/4294967296.0,1,-nbitq), 
to_sfixed(-226228175.0/4294967296.0,1,-nbitq), 
to_sfixed(-201860577.0/4294967296.0,1,-nbitq), 
to_sfixed(-419368917.0/4294967296.0,1,-nbitq), 
to_sfixed(111556686.0/4294967296.0,1,-nbitq), 
to_sfixed(110211397.0/4294967296.0,1,-nbitq), 
to_sfixed(-317887079.0/4294967296.0,1,-nbitq), 
to_sfixed(-46219533.0/4294967296.0,1,-nbitq), 
to_sfixed(323048325.0/4294967296.0,1,-nbitq), 
to_sfixed(-5560833.0/4294967296.0,1,-nbitq), 
to_sfixed(-316191922.0/4294967296.0,1,-nbitq), 
to_sfixed(238726210.0/4294967296.0,1,-nbitq), 
to_sfixed(-60620151.0/4294967296.0,1,-nbitq), 
to_sfixed(-218582275.0/4294967296.0,1,-nbitq), 
to_sfixed(-250016081.0/4294967296.0,1,-nbitq), 
to_sfixed(-290415214.0/4294967296.0,1,-nbitq), 
to_sfixed(260915511.0/4294967296.0,1,-nbitq), 
to_sfixed(387770108.0/4294967296.0,1,-nbitq), 
to_sfixed(402629433.0/4294967296.0,1,-nbitq), 
to_sfixed(-439903673.0/4294967296.0,1,-nbitq), 
to_sfixed(135681750.0/4294967296.0,1,-nbitq), 
to_sfixed(290094253.0/4294967296.0,1,-nbitq), 
to_sfixed(-147523006.0/4294967296.0,1,-nbitq), 
to_sfixed(147150506.0/4294967296.0,1,-nbitq), 
to_sfixed(-286688980.0/4294967296.0,1,-nbitq), 
to_sfixed(462893845.0/4294967296.0,1,-nbitq), 
to_sfixed(451166844.0/4294967296.0,1,-nbitq), 
to_sfixed(-36362962.0/4294967296.0,1,-nbitq), 
to_sfixed(88830300.0/4294967296.0,1,-nbitq), 
to_sfixed(-137034121.0/4294967296.0,1,-nbitq), 
to_sfixed(112766007.0/4294967296.0,1,-nbitq), 
to_sfixed(-353824140.0/4294967296.0,1,-nbitq), 
to_sfixed(51017691.0/4294967296.0,1,-nbitq), 
to_sfixed(-226086043.0/4294967296.0,1,-nbitq), 
to_sfixed(282324416.0/4294967296.0,1,-nbitq), 
to_sfixed(-183556781.0/4294967296.0,1,-nbitq), 
to_sfixed(-217895907.0/4294967296.0,1,-nbitq), 
to_sfixed(355539421.0/4294967296.0,1,-nbitq), 
to_sfixed(-357959153.0/4294967296.0,1,-nbitq), 
to_sfixed(-9401296.0/4294967296.0,1,-nbitq), 
to_sfixed(114555567.0/4294967296.0,1,-nbitq), 
to_sfixed(343153898.0/4294967296.0,1,-nbitq), 
to_sfixed(-180275746.0/4294967296.0,1,-nbitq), 
to_sfixed(187973991.0/4294967296.0,1,-nbitq), 
to_sfixed(307632762.0/4294967296.0,1,-nbitq), 
to_sfixed(-130448861.0/4294967296.0,1,-nbitq), 
to_sfixed(-294515113.0/4294967296.0,1,-nbitq), 
to_sfixed(-325124227.0/4294967296.0,1,-nbitq), 
to_sfixed(-90695212.0/4294967296.0,1,-nbitq), 
to_sfixed(35903489.0/4294967296.0,1,-nbitq), 
to_sfixed(409852358.0/4294967296.0,1,-nbitq), 
to_sfixed(-610768.0/4294967296.0,1,-nbitq), 
to_sfixed(-403463069.0/4294967296.0,1,-nbitq), 
to_sfixed(-347129308.0/4294967296.0,1,-nbitq), 
to_sfixed(-51493860.0/4294967296.0,1,-nbitq), 
to_sfixed(75607781.0/4294967296.0,1,-nbitq), 
to_sfixed(180365668.0/4294967296.0,1,-nbitq), 
to_sfixed(-405603207.0/4294967296.0,1,-nbitq), 
to_sfixed(-360587226.0/4294967296.0,1,-nbitq), 
to_sfixed(138718385.0/4294967296.0,1,-nbitq), 
to_sfixed(279524455.0/4294967296.0,1,-nbitq), 
to_sfixed(283781965.0/4294967296.0,1,-nbitq), 
to_sfixed(153039164.0/4294967296.0,1,-nbitq), 
to_sfixed(20528026.0/4294967296.0,1,-nbitq), 
to_sfixed(-205064894.0/4294967296.0,1,-nbitq), 
to_sfixed(258830445.0/4294967296.0,1,-nbitq), 
to_sfixed(201973983.0/4294967296.0,1,-nbitq), 
to_sfixed(-189550418.0/4294967296.0,1,-nbitq), 
to_sfixed(-139151843.0/4294967296.0,1,-nbitq), 
to_sfixed(534070860.0/4294967296.0,1,-nbitq), 
to_sfixed(153304041.0/4294967296.0,1,-nbitq), 
to_sfixed(250426156.0/4294967296.0,1,-nbitq), 
to_sfixed(-104518649.0/4294967296.0,1,-nbitq), 
to_sfixed(-165182889.0/4294967296.0,1,-nbitq), 
to_sfixed(396123498.0/4294967296.0,1,-nbitq), 
to_sfixed(-231688059.0/4294967296.0,1,-nbitq), 
to_sfixed(-314326129.0/4294967296.0,1,-nbitq), 
to_sfixed(123615670.0/4294967296.0,1,-nbitq), 
to_sfixed(-263776892.0/4294967296.0,1,-nbitq), 
to_sfixed(-191176029.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(277872880.0/4294967296.0,1,-nbitq), 
to_sfixed(-47475953.0/4294967296.0,1,-nbitq), 
to_sfixed(393312507.0/4294967296.0,1,-nbitq), 
to_sfixed(-222726850.0/4294967296.0,1,-nbitq), 
to_sfixed(-11871568.0/4294967296.0,1,-nbitq), 
to_sfixed(-67199601.0/4294967296.0,1,-nbitq), 
to_sfixed(-191289539.0/4294967296.0,1,-nbitq), 
to_sfixed(-127048309.0/4294967296.0,1,-nbitq), 
to_sfixed(5761813.0/4294967296.0,1,-nbitq), 
to_sfixed(265305281.0/4294967296.0,1,-nbitq), 
to_sfixed(61580764.0/4294967296.0,1,-nbitq), 
to_sfixed(-302548420.0/4294967296.0,1,-nbitq), 
to_sfixed(-22018728.0/4294967296.0,1,-nbitq), 
to_sfixed(195295227.0/4294967296.0,1,-nbitq), 
to_sfixed(274764207.0/4294967296.0,1,-nbitq), 
to_sfixed(107863209.0/4294967296.0,1,-nbitq), 
to_sfixed(-329289021.0/4294967296.0,1,-nbitq), 
to_sfixed(-338782720.0/4294967296.0,1,-nbitq), 
to_sfixed(-294217783.0/4294967296.0,1,-nbitq), 
to_sfixed(30665355.0/4294967296.0,1,-nbitq), 
to_sfixed(-79024521.0/4294967296.0,1,-nbitq), 
to_sfixed(347375407.0/4294967296.0,1,-nbitq), 
to_sfixed(-162265242.0/4294967296.0,1,-nbitq), 
to_sfixed(13056957.0/4294967296.0,1,-nbitq), 
to_sfixed(307927724.0/4294967296.0,1,-nbitq), 
to_sfixed(-199520392.0/4294967296.0,1,-nbitq), 
to_sfixed(-43120384.0/4294967296.0,1,-nbitq), 
to_sfixed(47777030.0/4294967296.0,1,-nbitq), 
to_sfixed(220733506.0/4294967296.0,1,-nbitq), 
to_sfixed(-123247766.0/4294967296.0,1,-nbitq), 
to_sfixed(-407718087.0/4294967296.0,1,-nbitq), 
to_sfixed(88753445.0/4294967296.0,1,-nbitq), 
to_sfixed(517584667.0/4294967296.0,1,-nbitq), 
to_sfixed(-263526465.0/4294967296.0,1,-nbitq), 
to_sfixed(-224215169.0/4294967296.0,1,-nbitq), 
to_sfixed(62477944.0/4294967296.0,1,-nbitq), 
to_sfixed(99505287.0/4294967296.0,1,-nbitq), 
to_sfixed(-11227967.0/4294967296.0,1,-nbitq), 
to_sfixed(256161542.0/4294967296.0,1,-nbitq), 
to_sfixed(117128527.0/4294967296.0,1,-nbitq), 
to_sfixed(50631063.0/4294967296.0,1,-nbitq), 
to_sfixed(-285908236.0/4294967296.0,1,-nbitq), 
to_sfixed(-442612230.0/4294967296.0,1,-nbitq), 
to_sfixed(-285518544.0/4294967296.0,1,-nbitq), 
to_sfixed(-177423526.0/4294967296.0,1,-nbitq), 
to_sfixed(324658496.0/4294967296.0,1,-nbitq), 
to_sfixed(8972910.0/4294967296.0,1,-nbitq), 
to_sfixed(-588727077.0/4294967296.0,1,-nbitq), 
to_sfixed(50084535.0/4294967296.0,1,-nbitq), 
to_sfixed(-31075265.0/4294967296.0,1,-nbitq), 
to_sfixed(313060146.0/4294967296.0,1,-nbitq), 
to_sfixed(-308964443.0/4294967296.0,1,-nbitq), 
to_sfixed(-439456441.0/4294967296.0,1,-nbitq), 
to_sfixed(163325319.0/4294967296.0,1,-nbitq), 
to_sfixed(110456960.0/4294967296.0,1,-nbitq), 
to_sfixed(-327036347.0/4294967296.0,1,-nbitq), 
to_sfixed(132543660.0/4294967296.0,1,-nbitq), 
to_sfixed(-131775809.0/4294967296.0,1,-nbitq), 
to_sfixed(-251800700.0/4294967296.0,1,-nbitq), 
to_sfixed(-273641331.0/4294967296.0,1,-nbitq), 
to_sfixed(280550200.0/4294967296.0,1,-nbitq), 
to_sfixed(261228388.0/4294967296.0,1,-nbitq), 
to_sfixed(-511839963.0/4294967296.0,1,-nbitq), 
to_sfixed(48540463.0/4294967296.0,1,-nbitq), 
to_sfixed(-4357006.0/4294967296.0,1,-nbitq), 
to_sfixed(-420797251.0/4294967296.0,1,-nbitq), 
to_sfixed(760504396.0/4294967296.0,1,-nbitq), 
to_sfixed(253256964.0/4294967296.0,1,-nbitq), 
to_sfixed(253315986.0/4294967296.0,1,-nbitq), 
to_sfixed(670373942.0/4294967296.0,1,-nbitq), 
to_sfixed(326105614.0/4294967296.0,1,-nbitq), 
to_sfixed(349994357.0/4294967296.0,1,-nbitq), 
to_sfixed(130815732.0/4294967296.0,1,-nbitq), 
to_sfixed(-99065412.0/4294967296.0,1,-nbitq), 
to_sfixed(-265824924.0/4294967296.0,1,-nbitq), 
to_sfixed(53925143.0/4294967296.0,1,-nbitq), 
to_sfixed(293392368.0/4294967296.0,1,-nbitq), 
to_sfixed(212202966.0/4294967296.0,1,-nbitq), 
to_sfixed(143390914.0/4294967296.0,1,-nbitq), 
to_sfixed(-45846176.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-58908199.0/4294967296.0,1,-nbitq), 
to_sfixed(-502067681.0/4294967296.0,1,-nbitq), 
to_sfixed(-37636144.0/4294967296.0,1,-nbitq), 
to_sfixed(-714692439.0/4294967296.0,1,-nbitq), 
to_sfixed(-41755479.0/4294967296.0,1,-nbitq), 
to_sfixed(-328763563.0/4294967296.0,1,-nbitq), 
to_sfixed(312992508.0/4294967296.0,1,-nbitq), 
to_sfixed(534327073.0/4294967296.0,1,-nbitq), 
to_sfixed(-46159041.0/4294967296.0,1,-nbitq), 
to_sfixed(-215881760.0/4294967296.0,1,-nbitq), 
to_sfixed(-68201972.0/4294967296.0,1,-nbitq), 
to_sfixed(-351952525.0/4294967296.0,1,-nbitq), 
to_sfixed(-257439267.0/4294967296.0,1,-nbitq), 
to_sfixed(-8863636.0/4294967296.0,1,-nbitq), 
to_sfixed(54631669.0/4294967296.0,1,-nbitq), 
to_sfixed(-61164742.0/4294967296.0,1,-nbitq), 
to_sfixed(-163978057.0/4294967296.0,1,-nbitq), 
to_sfixed(58790965.0/4294967296.0,1,-nbitq), 
to_sfixed(-385271775.0/4294967296.0,1,-nbitq), 
to_sfixed(342800850.0/4294967296.0,1,-nbitq), 
to_sfixed(-339203684.0/4294967296.0,1,-nbitq), 
to_sfixed(-15147542.0/4294967296.0,1,-nbitq), 
to_sfixed(-45320113.0/4294967296.0,1,-nbitq), 
to_sfixed(516505361.0/4294967296.0,1,-nbitq), 
to_sfixed(132521037.0/4294967296.0,1,-nbitq), 
to_sfixed(-484401042.0/4294967296.0,1,-nbitq), 
to_sfixed(-99562841.0/4294967296.0,1,-nbitq), 
to_sfixed(-184540278.0/4294967296.0,1,-nbitq), 
to_sfixed(-199788639.0/4294967296.0,1,-nbitq), 
to_sfixed(426454126.0/4294967296.0,1,-nbitq), 
to_sfixed(-149824318.0/4294967296.0,1,-nbitq), 
to_sfixed(182527906.0/4294967296.0,1,-nbitq), 
to_sfixed(80697281.0/4294967296.0,1,-nbitq), 
to_sfixed(-198791056.0/4294967296.0,1,-nbitq), 
to_sfixed(258446768.0/4294967296.0,1,-nbitq), 
to_sfixed(-330811895.0/4294967296.0,1,-nbitq), 
to_sfixed(-179384456.0/4294967296.0,1,-nbitq), 
to_sfixed(-355203908.0/4294967296.0,1,-nbitq), 
to_sfixed(-1391932.0/4294967296.0,1,-nbitq), 
to_sfixed(412430117.0/4294967296.0,1,-nbitq), 
to_sfixed(-114446604.0/4294967296.0,1,-nbitq), 
to_sfixed(258196776.0/4294967296.0,1,-nbitq), 
to_sfixed(68468901.0/4294967296.0,1,-nbitq), 
to_sfixed(-264910789.0/4294967296.0,1,-nbitq), 
to_sfixed(162572494.0/4294967296.0,1,-nbitq), 
to_sfixed(-20478917.0/4294967296.0,1,-nbitq), 
to_sfixed(247607261.0/4294967296.0,1,-nbitq), 
to_sfixed(137288884.0/4294967296.0,1,-nbitq), 
to_sfixed(47520406.0/4294967296.0,1,-nbitq), 
to_sfixed(-459565434.0/4294967296.0,1,-nbitq), 
to_sfixed(-189617492.0/4294967296.0,1,-nbitq), 
to_sfixed(-47545034.0/4294967296.0,1,-nbitq), 
to_sfixed(-228355449.0/4294967296.0,1,-nbitq), 
to_sfixed(393694475.0/4294967296.0,1,-nbitq), 
to_sfixed(337429642.0/4294967296.0,1,-nbitq), 
to_sfixed(-206025847.0/4294967296.0,1,-nbitq), 
to_sfixed(385013597.0/4294967296.0,1,-nbitq), 
to_sfixed(242170743.0/4294967296.0,1,-nbitq), 
to_sfixed(-257201629.0/4294967296.0,1,-nbitq), 
to_sfixed(-139628449.0/4294967296.0,1,-nbitq), 
to_sfixed(-378589428.0/4294967296.0,1,-nbitq), 
to_sfixed(341238444.0/4294967296.0,1,-nbitq), 
to_sfixed(-152012561.0/4294967296.0,1,-nbitq), 
to_sfixed(-277446794.0/4294967296.0,1,-nbitq), 
to_sfixed(306411686.0/4294967296.0,1,-nbitq), 
to_sfixed(-265672375.0/4294967296.0,1,-nbitq), 
to_sfixed(-8408167.0/4294967296.0,1,-nbitq), 
to_sfixed(-6060870.0/4294967296.0,1,-nbitq), 
to_sfixed(282881386.0/4294967296.0,1,-nbitq), 
to_sfixed(704348080.0/4294967296.0,1,-nbitq), 
to_sfixed(209747605.0/4294967296.0,1,-nbitq), 
to_sfixed(142846068.0/4294967296.0,1,-nbitq), 
to_sfixed(-47328799.0/4294967296.0,1,-nbitq), 
to_sfixed(362426479.0/4294967296.0,1,-nbitq), 
to_sfixed(-248142353.0/4294967296.0,1,-nbitq), 
to_sfixed(-81778286.0/4294967296.0,1,-nbitq), 
to_sfixed(60154960.0/4294967296.0,1,-nbitq), 
to_sfixed(19966723.0/4294967296.0,1,-nbitq), 
to_sfixed(19345181.0/4294967296.0,1,-nbitq), 
to_sfixed(379713539.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(353744353.0/4294967296.0,1,-nbitq), 
to_sfixed(-347902536.0/4294967296.0,1,-nbitq), 
to_sfixed(374428223.0/4294967296.0,1,-nbitq), 
to_sfixed(-439518596.0/4294967296.0,1,-nbitq), 
to_sfixed(-197908123.0/4294967296.0,1,-nbitq), 
to_sfixed(-536761398.0/4294967296.0,1,-nbitq), 
to_sfixed(-125395520.0/4294967296.0,1,-nbitq), 
to_sfixed(658418075.0/4294967296.0,1,-nbitq), 
to_sfixed(222389254.0/4294967296.0,1,-nbitq), 
to_sfixed(-69788577.0/4294967296.0,1,-nbitq), 
to_sfixed(-106261306.0/4294967296.0,1,-nbitq), 
to_sfixed(-69183341.0/4294967296.0,1,-nbitq), 
to_sfixed(140824711.0/4294967296.0,1,-nbitq), 
to_sfixed(672051209.0/4294967296.0,1,-nbitq), 
to_sfixed(-57835949.0/4294967296.0,1,-nbitq), 
to_sfixed(884803818.0/4294967296.0,1,-nbitq), 
to_sfixed(-198000304.0/4294967296.0,1,-nbitq), 
to_sfixed(-45956502.0/4294967296.0,1,-nbitq), 
to_sfixed(549671478.0/4294967296.0,1,-nbitq), 
to_sfixed(346194261.0/4294967296.0,1,-nbitq), 
to_sfixed(348880983.0/4294967296.0,1,-nbitq), 
to_sfixed(-431905761.0/4294967296.0,1,-nbitq), 
to_sfixed(-1052343658.0/4294967296.0,1,-nbitq), 
to_sfixed(420471452.0/4294967296.0,1,-nbitq), 
to_sfixed(-285753604.0/4294967296.0,1,-nbitq), 
to_sfixed(-960653731.0/4294967296.0,1,-nbitq), 
to_sfixed(561388370.0/4294967296.0,1,-nbitq), 
to_sfixed(-415873016.0/4294967296.0,1,-nbitq), 
to_sfixed(39695193.0/4294967296.0,1,-nbitq), 
to_sfixed(180297839.0/4294967296.0,1,-nbitq), 
to_sfixed(212980403.0/4294967296.0,1,-nbitq), 
to_sfixed(609022032.0/4294967296.0,1,-nbitq), 
to_sfixed(-254147935.0/4294967296.0,1,-nbitq), 
to_sfixed(674581510.0/4294967296.0,1,-nbitq), 
to_sfixed(-166894494.0/4294967296.0,1,-nbitq), 
to_sfixed(-493016654.0/4294967296.0,1,-nbitq), 
to_sfixed(-40056802.0/4294967296.0,1,-nbitq), 
to_sfixed(119236743.0/4294967296.0,1,-nbitq), 
to_sfixed(54374455.0/4294967296.0,1,-nbitq), 
to_sfixed(-301595360.0/4294967296.0,1,-nbitq), 
to_sfixed(-478045644.0/4294967296.0,1,-nbitq), 
to_sfixed(-610396001.0/4294967296.0,1,-nbitq), 
to_sfixed(-730795139.0/4294967296.0,1,-nbitq), 
to_sfixed(-147511903.0/4294967296.0,1,-nbitq), 
to_sfixed(-661056990.0/4294967296.0,1,-nbitq), 
to_sfixed(608715923.0/4294967296.0,1,-nbitq), 
to_sfixed(268244070.0/4294967296.0,1,-nbitq), 
to_sfixed(-238906230.0/4294967296.0,1,-nbitq), 
to_sfixed(-24419907.0/4294967296.0,1,-nbitq), 
to_sfixed(-215172443.0/4294967296.0,1,-nbitq), 
to_sfixed(-373459508.0/4294967296.0,1,-nbitq), 
to_sfixed(-315205214.0/4294967296.0,1,-nbitq), 
to_sfixed(-228665447.0/4294967296.0,1,-nbitq), 
to_sfixed(-53193364.0/4294967296.0,1,-nbitq), 
to_sfixed(539698428.0/4294967296.0,1,-nbitq), 
to_sfixed(-28614603.0/4294967296.0,1,-nbitq), 
to_sfixed(98850203.0/4294967296.0,1,-nbitq), 
to_sfixed(-87180929.0/4294967296.0,1,-nbitq), 
to_sfixed(314400165.0/4294967296.0,1,-nbitq), 
to_sfixed(277405861.0/4294967296.0,1,-nbitq), 
to_sfixed(-410278298.0/4294967296.0,1,-nbitq), 
to_sfixed(-124413165.0/4294967296.0,1,-nbitq), 
to_sfixed(374834301.0/4294967296.0,1,-nbitq), 
to_sfixed(-561629646.0/4294967296.0,1,-nbitq), 
to_sfixed(-377009108.0/4294967296.0,1,-nbitq), 
to_sfixed(350357156.0/4294967296.0,1,-nbitq), 
to_sfixed(205992986.0/4294967296.0,1,-nbitq), 
to_sfixed(-96829187.0/4294967296.0,1,-nbitq), 
to_sfixed(405787443.0/4294967296.0,1,-nbitq), 
to_sfixed(560716660.0/4294967296.0,1,-nbitq), 
to_sfixed(248780693.0/4294967296.0,1,-nbitq), 
to_sfixed(64240465.0/4294967296.0,1,-nbitq), 
to_sfixed(108419550.0/4294967296.0,1,-nbitq), 
to_sfixed(121003773.0/4294967296.0,1,-nbitq), 
to_sfixed(-216697182.0/4294967296.0,1,-nbitq), 
to_sfixed(-118499126.0/4294967296.0,1,-nbitq), 
to_sfixed(-612228259.0/4294967296.0,1,-nbitq), 
to_sfixed(-139902073.0/4294967296.0,1,-nbitq), 
to_sfixed(58359621.0/4294967296.0,1,-nbitq), 
to_sfixed(-376427916.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(286214109.0/4294967296.0,1,-nbitq), 
to_sfixed(201634004.0/4294967296.0,1,-nbitq), 
to_sfixed(696485150.0/4294967296.0,1,-nbitq), 
to_sfixed(-1053786622.0/4294967296.0,1,-nbitq), 
to_sfixed(-372805982.0/4294967296.0,1,-nbitq), 
to_sfixed(-102326547.0/4294967296.0,1,-nbitq), 
to_sfixed(122470563.0/4294967296.0,1,-nbitq), 
to_sfixed(549806157.0/4294967296.0,1,-nbitq), 
to_sfixed(-430155809.0/4294967296.0,1,-nbitq), 
to_sfixed(215334868.0/4294967296.0,1,-nbitq), 
to_sfixed(324260642.0/4294967296.0,1,-nbitq), 
to_sfixed(-939450938.0/4294967296.0,1,-nbitq), 
to_sfixed(-13636411.0/4294967296.0,1,-nbitq), 
to_sfixed(1232370688.0/4294967296.0,1,-nbitq), 
to_sfixed(265242818.0/4294967296.0,1,-nbitq), 
to_sfixed(965121427.0/4294967296.0,1,-nbitq), 
to_sfixed(-71350762.0/4294967296.0,1,-nbitq), 
to_sfixed(-53115477.0/4294967296.0,1,-nbitq), 
to_sfixed(-89832757.0/4294967296.0,1,-nbitq), 
to_sfixed(1064837796.0/4294967296.0,1,-nbitq), 
to_sfixed(-303944520.0/4294967296.0,1,-nbitq), 
to_sfixed(-919585851.0/4294967296.0,1,-nbitq), 
to_sfixed(-1572584510.0/4294967296.0,1,-nbitq), 
to_sfixed(811824610.0/4294967296.0,1,-nbitq), 
to_sfixed(-74202071.0/4294967296.0,1,-nbitq), 
to_sfixed(-1235710824.0/4294967296.0,1,-nbitq), 
to_sfixed(188709184.0/4294967296.0,1,-nbitq), 
to_sfixed(-188370403.0/4294967296.0,1,-nbitq), 
to_sfixed(195183090.0/4294967296.0,1,-nbitq), 
to_sfixed(899113795.0/4294967296.0,1,-nbitq), 
to_sfixed(-329468814.0/4294967296.0,1,-nbitq), 
to_sfixed(135932061.0/4294967296.0,1,-nbitq), 
to_sfixed(576364355.0/4294967296.0,1,-nbitq), 
to_sfixed(219553893.0/4294967296.0,1,-nbitq), 
to_sfixed(-320201426.0/4294967296.0,1,-nbitq), 
to_sfixed(-20736884.0/4294967296.0,1,-nbitq), 
to_sfixed(-589915760.0/4294967296.0,1,-nbitq), 
to_sfixed(-159184932.0/4294967296.0,1,-nbitq), 
to_sfixed(-353941725.0/4294967296.0,1,-nbitq), 
to_sfixed(189158572.0/4294967296.0,1,-nbitq), 
to_sfixed(-244056998.0/4294967296.0,1,-nbitq), 
to_sfixed(-517497624.0/4294967296.0,1,-nbitq), 
to_sfixed(-310885471.0/4294967296.0,1,-nbitq), 
to_sfixed(-693449125.0/4294967296.0,1,-nbitq), 
to_sfixed(-648827907.0/4294967296.0,1,-nbitq), 
to_sfixed(-396202243.0/4294967296.0,1,-nbitq), 
to_sfixed(224424522.0/4294967296.0,1,-nbitq), 
to_sfixed(363419029.0/4294967296.0,1,-nbitq), 
to_sfixed(363631571.0/4294967296.0,1,-nbitq), 
to_sfixed(24399271.0/4294967296.0,1,-nbitq), 
to_sfixed(76313228.0/4294967296.0,1,-nbitq), 
to_sfixed(-924126513.0/4294967296.0,1,-nbitq), 
to_sfixed(-44969804.0/4294967296.0,1,-nbitq), 
to_sfixed(481662702.0/4294967296.0,1,-nbitq), 
to_sfixed(-236440303.0/4294967296.0,1,-nbitq), 
to_sfixed(-310863131.0/4294967296.0,1,-nbitq), 
to_sfixed(-197699692.0/4294967296.0,1,-nbitq), 
to_sfixed(-22121697.0/4294967296.0,1,-nbitq), 
to_sfixed(39494944.0/4294967296.0,1,-nbitq), 
to_sfixed(-322184714.0/4294967296.0,1,-nbitq), 
to_sfixed(147139385.0/4294967296.0,1,-nbitq), 
to_sfixed(482337548.0/4294967296.0,1,-nbitq), 
to_sfixed(1022015201.0/4294967296.0,1,-nbitq), 
to_sfixed(-482947381.0/4294967296.0,1,-nbitq), 
to_sfixed(103334812.0/4294967296.0,1,-nbitq), 
to_sfixed(-50926136.0/4294967296.0,1,-nbitq), 
to_sfixed(186285243.0/4294967296.0,1,-nbitq), 
to_sfixed(381837423.0/4294967296.0,1,-nbitq), 
to_sfixed(-27719904.0/4294967296.0,1,-nbitq), 
to_sfixed(330286467.0/4294967296.0,1,-nbitq), 
to_sfixed(799157162.0/4294967296.0,1,-nbitq), 
to_sfixed(-293799705.0/4294967296.0,1,-nbitq), 
to_sfixed(303653879.0/4294967296.0,1,-nbitq), 
to_sfixed(246434600.0/4294967296.0,1,-nbitq), 
to_sfixed(-68398111.0/4294967296.0,1,-nbitq), 
to_sfixed(365334019.0/4294967296.0,1,-nbitq), 
to_sfixed(-1334846354.0/4294967296.0,1,-nbitq), 
to_sfixed(-75409393.0/4294967296.0,1,-nbitq), 
to_sfixed(842538311.0/4294967296.0,1,-nbitq), 
to_sfixed(34687534.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-39508588.0/4294967296.0,1,-nbitq), 
to_sfixed(571857745.0/4294967296.0,1,-nbitq), 
to_sfixed(-57930255.0/4294967296.0,1,-nbitq), 
to_sfixed(-1483402830.0/4294967296.0,1,-nbitq), 
to_sfixed(-518151282.0/4294967296.0,1,-nbitq), 
to_sfixed(484705102.0/4294967296.0,1,-nbitq), 
to_sfixed(-427193135.0/4294967296.0,1,-nbitq), 
to_sfixed(88969150.0/4294967296.0,1,-nbitq), 
to_sfixed(-455244960.0/4294967296.0,1,-nbitq), 
to_sfixed(147467848.0/4294967296.0,1,-nbitq), 
to_sfixed(614402853.0/4294967296.0,1,-nbitq), 
to_sfixed(-1134299197.0/4294967296.0,1,-nbitq), 
to_sfixed(-213258027.0/4294967296.0,1,-nbitq), 
to_sfixed(1171806056.0/4294967296.0,1,-nbitq), 
to_sfixed(-371605509.0/4294967296.0,1,-nbitq), 
to_sfixed(1368622017.0/4294967296.0,1,-nbitq), 
to_sfixed(-389250389.0/4294967296.0,1,-nbitq), 
to_sfixed(-32630191.0/4294967296.0,1,-nbitq), 
to_sfixed(-169123138.0/4294967296.0,1,-nbitq), 
to_sfixed(1204410293.0/4294967296.0,1,-nbitq), 
to_sfixed(121797633.0/4294967296.0,1,-nbitq), 
to_sfixed(-241015574.0/4294967296.0,1,-nbitq), 
to_sfixed(-1232787911.0/4294967296.0,1,-nbitq), 
to_sfixed(974870840.0/4294967296.0,1,-nbitq), 
to_sfixed(-123358551.0/4294967296.0,1,-nbitq), 
to_sfixed(-1284304675.0/4294967296.0,1,-nbitq), 
to_sfixed(494463909.0/4294967296.0,1,-nbitq), 
to_sfixed(151420115.0/4294967296.0,1,-nbitq), 
to_sfixed(1102852736.0/4294967296.0,1,-nbitq), 
to_sfixed(820358876.0/4294967296.0,1,-nbitq), 
to_sfixed(-181606988.0/4294967296.0,1,-nbitq), 
to_sfixed(581488012.0/4294967296.0,1,-nbitq), 
to_sfixed(120687100.0/4294967296.0,1,-nbitq), 
to_sfixed(-379412161.0/4294967296.0,1,-nbitq), 
to_sfixed(277813023.0/4294967296.0,1,-nbitq), 
to_sfixed(-209766559.0/4294967296.0,1,-nbitq), 
to_sfixed(-653574642.0/4294967296.0,1,-nbitq), 
to_sfixed(-810438146.0/4294967296.0,1,-nbitq), 
to_sfixed(153351325.0/4294967296.0,1,-nbitq), 
to_sfixed(-69068910.0/4294967296.0,1,-nbitq), 
to_sfixed(-224883706.0/4294967296.0,1,-nbitq), 
to_sfixed(-511946766.0/4294967296.0,1,-nbitq), 
to_sfixed(111140286.0/4294967296.0,1,-nbitq), 
to_sfixed(-484689511.0/4294967296.0,1,-nbitq), 
to_sfixed(-634267640.0/4294967296.0,1,-nbitq), 
to_sfixed(-500711662.0/4294967296.0,1,-nbitq), 
to_sfixed(-264884643.0/4294967296.0,1,-nbitq), 
to_sfixed(151581726.0/4294967296.0,1,-nbitq), 
to_sfixed(400470162.0/4294967296.0,1,-nbitq), 
to_sfixed(-335672797.0/4294967296.0,1,-nbitq), 
to_sfixed(-194408093.0/4294967296.0,1,-nbitq), 
to_sfixed(-1138417039.0/4294967296.0,1,-nbitq), 
to_sfixed(409216343.0/4294967296.0,1,-nbitq), 
to_sfixed(564209377.0/4294967296.0,1,-nbitq), 
to_sfixed(-932187396.0/4294967296.0,1,-nbitq), 
to_sfixed(-409894690.0/4294967296.0,1,-nbitq), 
to_sfixed(295184276.0/4294967296.0,1,-nbitq), 
to_sfixed(-281986495.0/4294967296.0,1,-nbitq), 
to_sfixed(183564178.0/4294967296.0,1,-nbitq), 
to_sfixed(431098912.0/4294967296.0,1,-nbitq), 
to_sfixed(-80165088.0/4294967296.0,1,-nbitq), 
to_sfixed(-70770489.0/4294967296.0,1,-nbitq), 
to_sfixed(1060885350.0/4294967296.0,1,-nbitq), 
to_sfixed(-114379312.0/4294967296.0,1,-nbitq), 
to_sfixed(-10365387.0/4294967296.0,1,-nbitq), 
to_sfixed(337021536.0/4294967296.0,1,-nbitq), 
to_sfixed(242204070.0/4294967296.0,1,-nbitq), 
to_sfixed(62464185.0/4294967296.0,1,-nbitq), 
to_sfixed(387740789.0/4294967296.0,1,-nbitq), 
to_sfixed(93489144.0/4294967296.0,1,-nbitq), 
to_sfixed(511512763.0/4294967296.0,1,-nbitq), 
to_sfixed(-218521755.0/4294967296.0,1,-nbitq), 
to_sfixed(370253480.0/4294967296.0,1,-nbitq), 
to_sfixed(256274378.0/4294967296.0,1,-nbitq), 
to_sfixed(-175712272.0/4294967296.0,1,-nbitq), 
to_sfixed(217554139.0/4294967296.0,1,-nbitq), 
to_sfixed(-1973942011.0/4294967296.0,1,-nbitq), 
to_sfixed(109369733.0/4294967296.0,1,-nbitq), 
to_sfixed(-127471875.0/4294967296.0,1,-nbitq), 
to_sfixed(3541901.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-535590161.0/4294967296.0,1,-nbitq), 
to_sfixed(336400202.0/4294967296.0,1,-nbitq), 
to_sfixed(-606984940.0/4294967296.0,1,-nbitq), 
to_sfixed(-1088764368.0/4294967296.0,1,-nbitq), 
to_sfixed(212532210.0/4294967296.0,1,-nbitq), 
to_sfixed(1775559724.0/4294967296.0,1,-nbitq), 
to_sfixed(450975620.0/4294967296.0,1,-nbitq), 
to_sfixed(1031502764.0/4294967296.0,1,-nbitq), 
to_sfixed(-562789526.0/4294967296.0,1,-nbitq), 
to_sfixed(-142265302.0/4294967296.0,1,-nbitq), 
to_sfixed(-188999061.0/4294967296.0,1,-nbitq), 
to_sfixed(-767851612.0/4294967296.0,1,-nbitq), 
to_sfixed(-414005144.0/4294967296.0,1,-nbitq), 
to_sfixed(236243946.0/4294967296.0,1,-nbitq), 
to_sfixed(-205842486.0/4294967296.0,1,-nbitq), 
to_sfixed(849849273.0/4294967296.0,1,-nbitq), 
to_sfixed(-269501569.0/4294967296.0,1,-nbitq), 
to_sfixed(283913380.0/4294967296.0,1,-nbitq), 
to_sfixed(-448801293.0/4294967296.0,1,-nbitq), 
to_sfixed(1218905787.0/4294967296.0,1,-nbitq), 
to_sfixed(-52113918.0/4294967296.0,1,-nbitq), 
to_sfixed(-307008987.0/4294967296.0,1,-nbitq), 
to_sfixed(-543723018.0/4294967296.0,1,-nbitq), 
to_sfixed(-145968712.0/4294967296.0,1,-nbitq), 
to_sfixed(460162002.0/4294967296.0,1,-nbitq), 
to_sfixed(-735839962.0/4294967296.0,1,-nbitq), 
to_sfixed(634751185.0/4294967296.0,1,-nbitq), 
to_sfixed(386847134.0/4294967296.0,1,-nbitq), 
to_sfixed(965022655.0/4294967296.0,1,-nbitq), 
to_sfixed(493643188.0/4294967296.0,1,-nbitq), 
to_sfixed(180174613.0/4294967296.0,1,-nbitq), 
to_sfixed(612684072.0/4294967296.0,1,-nbitq), 
to_sfixed(219543485.0/4294967296.0,1,-nbitq), 
to_sfixed(87628536.0/4294967296.0,1,-nbitq), 
to_sfixed(73216833.0/4294967296.0,1,-nbitq), 
to_sfixed(-1360906415.0/4294967296.0,1,-nbitq), 
to_sfixed(-780878404.0/4294967296.0,1,-nbitq), 
to_sfixed(116222064.0/4294967296.0,1,-nbitq), 
to_sfixed(-159850712.0/4294967296.0,1,-nbitq), 
to_sfixed(147081985.0/4294967296.0,1,-nbitq), 
to_sfixed(-92883292.0/4294967296.0,1,-nbitq), 
to_sfixed(-444563779.0/4294967296.0,1,-nbitq), 
to_sfixed(205740849.0/4294967296.0,1,-nbitq), 
to_sfixed(8031525.0/4294967296.0,1,-nbitq), 
to_sfixed(-280383363.0/4294967296.0,1,-nbitq), 
to_sfixed(91751658.0/4294967296.0,1,-nbitq), 
to_sfixed(-22054201.0/4294967296.0,1,-nbitq), 
to_sfixed(900478983.0/4294967296.0,1,-nbitq), 
to_sfixed(90597109.0/4294967296.0,1,-nbitq), 
to_sfixed(-30710731.0/4294967296.0,1,-nbitq), 
to_sfixed(-784251425.0/4294967296.0,1,-nbitq), 
to_sfixed(-1626981541.0/4294967296.0,1,-nbitq), 
to_sfixed(576971977.0/4294967296.0,1,-nbitq), 
to_sfixed(1148605817.0/4294967296.0,1,-nbitq), 
to_sfixed(-728524357.0/4294967296.0,1,-nbitq), 
to_sfixed(-1289121599.0/4294967296.0,1,-nbitq), 
to_sfixed(-76942815.0/4294967296.0,1,-nbitq), 
to_sfixed(-1002969580.0/4294967296.0,1,-nbitq), 
to_sfixed(-117273320.0/4294967296.0,1,-nbitq), 
to_sfixed(299545224.0/4294967296.0,1,-nbitq), 
to_sfixed(33952518.0/4294967296.0,1,-nbitq), 
to_sfixed(124678344.0/4294967296.0,1,-nbitq), 
to_sfixed(996121777.0/4294967296.0,1,-nbitq), 
to_sfixed(219410300.0/4294967296.0,1,-nbitq), 
to_sfixed(98457776.0/4294967296.0,1,-nbitq), 
to_sfixed(401259837.0/4294967296.0,1,-nbitq), 
to_sfixed(-313141136.0/4294967296.0,1,-nbitq), 
to_sfixed(696650062.0/4294967296.0,1,-nbitq), 
to_sfixed(-118761317.0/4294967296.0,1,-nbitq), 
to_sfixed(3350610.0/4294967296.0,1,-nbitq), 
to_sfixed(775841194.0/4294967296.0,1,-nbitq), 
to_sfixed(353211239.0/4294967296.0,1,-nbitq), 
to_sfixed(-9062813.0/4294967296.0,1,-nbitq), 
to_sfixed(87464931.0/4294967296.0,1,-nbitq), 
to_sfixed(-134338948.0/4294967296.0,1,-nbitq), 
to_sfixed(151580638.0/4294967296.0,1,-nbitq), 
to_sfixed(-1545650637.0/4294967296.0,1,-nbitq), 
to_sfixed(167470138.0/4294967296.0,1,-nbitq), 
to_sfixed(63120536.0/4294967296.0,1,-nbitq), 
to_sfixed(-7736095.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-690802911.0/4294967296.0,1,-nbitq), 
to_sfixed(259065810.0/4294967296.0,1,-nbitq), 
to_sfixed(-355960382.0/4294967296.0,1,-nbitq), 
to_sfixed(129915932.0/4294967296.0,1,-nbitq), 
to_sfixed(79574780.0/4294967296.0,1,-nbitq), 
to_sfixed(2035908467.0/4294967296.0,1,-nbitq), 
to_sfixed(72330845.0/4294967296.0,1,-nbitq), 
to_sfixed(1591378337.0/4294967296.0,1,-nbitq), 
to_sfixed(-538677298.0/4294967296.0,1,-nbitq), 
to_sfixed(310373971.0/4294967296.0,1,-nbitq), 
to_sfixed(-411125596.0/4294967296.0,1,-nbitq), 
to_sfixed(-2302769434.0/4294967296.0,1,-nbitq), 
to_sfixed(-604715244.0/4294967296.0,1,-nbitq), 
to_sfixed(927202696.0/4294967296.0,1,-nbitq), 
to_sfixed(405774290.0/4294967296.0,1,-nbitq), 
to_sfixed(695992786.0/4294967296.0,1,-nbitq), 
to_sfixed(313969399.0/4294967296.0,1,-nbitq), 
to_sfixed(-268334585.0/4294967296.0,1,-nbitq), 
to_sfixed(-187792603.0/4294967296.0,1,-nbitq), 
to_sfixed(1256551295.0/4294967296.0,1,-nbitq), 
to_sfixed(69298058.0/4294967296.0,1,-nbitq), 
to_sfixed(-436382436.0/4294967296.0,1,-nbitq), 
to_sfixed(-396795107.0/4294967296.0,1,-nbitq), 
to_sfixed(831954597.0/4294967296.0,1,-nbitq), 
to_sfixed(435629835.0/4294967296.0,1,-nbitq), 
to_sfixed(-1175752901.0/4294967296.0,1,-nbitq), 
to_sfixed(461159904.0/4294967296.0,1,-nbitq), 
to_sfixed(183704587.0/4294967296.0,1,-nbitq), 
to_sfixed(437844811.0/4294967296.0,1,-nbitq), 
to_sfixed(1108758613.0/4294967296.0,1,-nbitq), 
to_sfixed(529066939.0/4294967296.0,1,-nbitq), 
to_sfixed(510128811.0/4294967296.0,1,-nbitq), 
to_sfixed(618343570.0/4294967296.0,1,-nbitq), 
to_sfixed(370793774.0/4294967296.0,1,-nbitq), 
to_sfixed(-306046733.0/4294967296.0,1,-nbitq), 
to_sfixed(-2002091975.0/4294967296.0,1,-nbitq), 
to_sfixed(-1134809429.0/4294967296.0,1,-nbitq), 
to_sfixed(182249686.0/4294967296.0,1,-nbitq), 
to_sfixed(175942596.0/4294967296.0,1,-nbitq), 
to_sfixed(204120571.0/4294967296.0,1,-nbitq), 
to_sfixed(-254103356.0/4294967296.0,1,-nbitq), 
to_sfixed(-547354961.0/4294967296.0,1,-nbitq), 
to_sfixed(-223527845.0/4294967296.0,1,-nbitq), 
to_sfixed(-1125771598.0/4294967296.0,1,-nbitq), 
to_sfixed(-155994541.0/4294967296.0,1,-nbitq), 
to_sfixed(140128781.0/4294967296.0,1,-nbitq), 
to_sfixed(-143778231.0/4294967296.0,1,-nbitq), 
to_sfixed(964133135.0/4294967296.0,1,-nbitq), 
to_sfixed(389594346.0/4294967296.0,1,-nbitq), 
to_sfixed(-584673684.0/4294967296.0,1,-nbitq), 
to_sfixed(50112945.0/4294967296.0,1,-nbitq), 
to_sfixed(-1330607898.0/4294967296.0,1,-nbitq), 
to_sfixed(1113582219.0/4294967296.0,1,-nbitq), 
to_sfixed(531059426.0/4294967296.0,1,-nbitq), 
to_sfixed(519951448.0/4294967296.0,1,-nbitq), 
to_sfixed(-1483005753.0/4294967296.0,1,-nbitq), 
to_sfixed(-303590276.0/4294967296.0,1,-nbitq), 
to_sfixed(-941903725.0/4294967296.0,1,-nbitq), 
to_sfixed(172087161.0/4294967296.0,1,-nbitq), 
to_sfixed(39049618.0/4294967296.0,1,-nbitq), 
to_sfixed(-374659861.0/4294967296.0,1,-nbitq), 
to_sfixed(422833832.0/4294967296.0,1,-nbitq), 
to_sfixed(1543086952.0/4294967296.0,1,-nbitq), 
to_sfixed(-14377485.0/4294967296.0,1,-nbitq), 
to_sfixed(-26254734.0/4294967296.0,1,-nbitq), 
to_sfixed(268657950.0/4294967296.0,1,-nbitq), 
to_sfixed(-1008380315.0/4294967296.0,1,-nbitq), 
to_sfixed(92119776.0/4294967296.0,1,-nbitq), 
to_sfixed(6477069.0/4294967296.0,1,-nbitq), 
to_sfixed(-410018251.0/4294967296.0,1,-nbitq), 
to_sfixed(782595020.0/4294967296.0,1,-nbitq), 
to_sfixed(211457120.0/4294967296.0,1,-nbitq), 
to_sfixed(320813123.0/4294967296.0,1,-nbitq), 
to_sfixed(385946853.0/4294967296.0,1,-nbitq), 
to_sfixed(15134238.0/4294967296.0,1,-nbitq), 
to_sfixed(1020036978.0/4294967296.0,1,-nbitq), 
to_sfixed(-481877425.0/4294967296.0,1,-nbitq), 
to_sfixed(739244485.0/4294967296.0,1,-nbitq), 
to_sfixed(-698087565.0/4294967296.0,1,-nbitq), 
to_sfixed(408584799.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-573754881.0/4294967296.0,1,-nbitq), 
to_sfixed(-101785055.0/4294967296.0,1,-nbitq), 
to_sfixed(95244649.0/4294967296.0,1,-nbitq), 
to_sfixed(476568278.0/4294967296.0,1,-nbitq), 
to_sfixed(-126602372.0/4294967296.0,1,-nbitq), 
to_sfixed(1935116380.0/4294967296.0,1,-nbitq), 
to_sfixed(228370319.0/4294967296.0,1,-nbitq), 
to_sfixed(1537604875.0/4294967296.0,1,-nbitq), 
to_sfixed(-1090230104.0/4294967296.0,1,-nbitq), 
to_sfixed(-233467775.0/4294967296.0,1,-nbitq), 
to_sfixed(-1036071481.0/4294967296.0,1,-nbitq), 
to_sfixed(-2766997678.0/4294967296.0,1,-nbitq), 
to_sfixed(30520272.0/4294967296.0,1,-nbitq), 
to_sfixed(1687366585.0/4294967296.0,1,-nbitq), 
to_sfixed(-211766157.0/4294967296.0,1,-nbitq), 
to_sfixed(702724579.0/4294967296.0,1,-nbitq), 
to_sfixed(-136178672.0/4294967296.0,1,-nbitq), 
to_sfixed(128609018.0/4294967296.0,1,-nbitq), 
to_sfixed(1667581445.0/4294967296.0,1,-nbitq), 
to_sfixed(1035570756.0/4294967296.0,1,-nbitq), 
to_sfixed(-170949344.0/4294967296.0,1,-nbitq), 
to_sfixed(-391143557.0/4294967296.0,1,-nbitq), 
to_sfixed(-166062032.0/4294967296.0,1,-nbitq), 
to_sfixed(1495696424.0/4294967296.0,1,-nbitq), 
to_sfixed(54932791.0/4294967296.0,1,-nbitq), 
to_sfixed(-1705416039.0/4294967296.0,1,-nbitq), 
to_sfixed(180931581.0/4294967296.0,1,-nbitq), 
to_sfixed(297043292.0/4294967296.0,1,-nbitq), 
to_sfixed(187655583.0/4294967296.0,1,-nbitq), 
to_sfixed(1110411551.0/4294967296.0,1,-nbitq), 
to_sfixed(387252032.0/4294967296.0,1,-nbitq), 
to_sfixed(-266162979.0/4294967296.0,1,-nbitq), 
to_sfixed(-518243978.0/4294967296.0,1,-nbitq), 
to_sfixed(462474320.0/4294967296.0,1,-nbitq), 
to_sfixed(-476921387.0/4294967296.0,1,-nbitq), 
to_sfixed(-147899819.0/4294967296.0,1,-nbitq), 
to_sfixed(-785129202.0/4294967296.0,1,-nbitq), 
to_sfixed(120218298.0/4294967296.0,1,-nbitq), 
to_sfixed(-163495232.0/4294967296.0,1,-nbitq), 
to_sfixed(87342915.0/4294967296.0,1,-nbitq), 
to_sfixed(45488562.0/4294967296.0,1,-nbitq), 
to_sfixed(95957463.0/4294967296.0,1,-nbitq), 
to_sfixed(-320996379.0/4294967296.0,1,-nbitq), 
to_sfixed(-718423756.0/4294967296.0,1,-nbitq), 
to_sfixed(-119916940.0/4294967296.0,1,-nbitq), 
to_sfixed(140155015.0/4294967296.0,1,-nbitq), 
to_sfixed(297559931.0/4294967296.0,1,-nbitq), 
to_sfixed(958757427.0/4294967296.0,1,-nbitq), 
to_sfixed(267406729.0/4294967296.0,1,-nbitq), 
to_sfixed(-980385148.0/4294967296.0,1,-nbitq), 
to_sfixed(-820563096.0/4294967296.0,1,-nbitq), 
to_sfixed(-777803895.0/4294967296.0,1,-nbitq), 
to_sfixed(866513517.0/4294967296.0,1,-nbitq), 
to_sfixed(-462333088.0/4294967296.0,1,-nbitq), 
to_sfixed(306487005.0/4294967296.0,1,-nbitq), 
to_sfixed(-1018608821.0/4294967296.0,1,-nbitq), 
to_sfixed(368706406.0/4294967296.0,1,-nbitq), 
to_sfixed(-612167170.0/4294967296.0,1,-nbitq), 
to_sfixed(174326919.0/4294967296.0,1,-nbitq), 
to_sfixed(-339014012.0/4294967296.0,1,-nbitq), 
to_sfixed(-148127821.0/4294967296.0,1,-nbitq), 
to_sfixed(436622469.0/4294967296.0,1,-nbitq), 
to_sfixed(1175080106.0/4294967296.0,1,-nbitq), 
to_sfixed(106532503.0/4294967296.0,1,-nbitq), 
to_sfixed(46659524.0/4294967296.0,1,-nbitq), 
to_sfixed(322367710.0/4294967296.0,1,-nbitq), 
to_sfixed(-1406692968.0/4294967296.0,1,-nbitq), 
to_sfixed(-157780783.0/4294967296.0,1,-nbitq), 
to_sfixed(6944219.0/4294967296.0,1,-nbitq), 
to_sfixed(-1253147222.0/4294967296.0,1,-nbitq), 
to_sfixed(397493405.0/4294967296.0,1,-nbitq), 
to_sfixed(-68515088.0/4294967296.0,1,-nbitq), 
to_sfixed(404830706.0/4294967296.0,1,-nbitq), 
to_sfixed(-100735113.0/4294967296.0,1,-nbitq), 
to_sfixed(364108572.0/4294967296.0,1,-nbitq), 
to_sfixed(-487759068.0/4294967296.0,1,-nbitq), 
to_sfixed(-610421047.0/4294967296.0,1,-nbitq), 
to_sfixed(609284128.0/4294967296.0,1,-nbitq), 
to_sfixed(-1062837021.0/4294967296.0,1,-nbitq), 
to_sfixed(-187680368.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(15432732.0/4294967296.0,1,-nbitq), 
to_sfixed(-2849909.0/4294967296.0,1,-nbitq), 
to_sfixed(301780877.0/4294967296.0,1,-nbitq), 
to_sfixed(579709394.0/4294967296.0,1,-nbitq), 
to_sfixed(-6443896.0/4294967296.0,1,-nbitq), 
to_sfixed(-125991414.0/4294967296.0,1,-nbitq), 
to_sfixed(546083244.0/4294967296.0,1,-nbitq), 
to_sfixed(1488840541.0/4294967296.0,1,-nbitq), 
to_sfixed(-1327557433.0/4294967296.0,1,-nbitq), 
to_sfixed(201917897.0/4294967296.0,1,-nbitq), 
to_sfixed(-1259694050.0/4294967296.0,1,-nbitq), 
to_sfixed(-1920585387.0/4294967296.0,1,-nbitq), 
to_sfixed(-774951489.0/4294967296.0,1,-nbitq), 
to_sfixed(741865767.0/4294967296.0,1,-nbitq), 
to_sfixed(392375157.0/4294967296.0,1,-nbitq), 
to_sfixed(950714301.0/4294967296.0,1,-nbitq), 
to_sfixed(-63865460.0/4294967296.0,1,-nbitq), 
to_sfixed(-136862871.0/4294967296.0,1,-nbitq), 
to_sfixed(1852427294.0/4294967296.0,1,-nbitq), 
to_sfixed(787033717.0/4294967296.0,1,-nbitq), 
to_sfixed(-341292821.0/4294967296.0,1,-nbitq), 
to_sfixed(123523617.0/4294967296.0,1,-nbitq), 
to_sfixed(-258620970.0/4294967296.0,1,-nbitq), 
to_sfixed(832140719.0/4294967296.0,1,-nbitq), 
to_sfixed(-138180722.0/4294967296.0,1,-nbitq), 
to_sfixed(-1561400199.0/4294967296.0,1,-nbitq), 
to_sfixed(-485877643.0/4294967296.0,1,-nbitq), 
to_sfixed(1025165316.0/4294967296.0,1,-nbitq), 
to_sfixed(872009899.0/4294967296.0,1,-nbitq), 
to_sfixed(1218503906.0/4294967296.0,1,-nbitq), 
to_sfixed(-207024981.0/4294967296.0,1,-nbitq), 
to_sfixed(-211849996.0/4294967296.0,1,-nbitq), 
to_sfixed(-300306355.0/4294967296.0,1,-nbitq), 
to_sfixed(586051104.0/4294967296.0,1,-nbitq), 
to_sfixed(-132731696.0/4294967296.0,1,-nbitq), 
to_sfixed(98776018.0/4294967296.0,1,-nbitq), 
to_sfixed(33529601.0/4294967296.0,1,-nbitq), 
to_sfixed(437872703.0/4294967296.0,1,-nbitq), 
to_sfixed(-369699628.0/4294967296.0,1,-nbitq), 
to_sfixed(-301142031.0/4294967296.0,1,-nbitq), 
to_sfixed(-455190091.0/4294967296.0,1,-nbitq), 
to_sfixed(359304686.0/4294967296.0,1,-nbitq), 
to_sfixed(-216388243.0/4294967296.0,1,-nbitq), 
to_sfixed(230479352.0/4294967296.0,1,-nbitq), 
to_sfixed(-226880004.0/4294967296.0,1,-nbitq), 
to_sfixed(-59324606.0/4294967296.0,1,-nbitq), 
to_sfixed(-408834352.0/4294967296.0,1,-nbitq), 
to_sfixed(1523590602.0/4294967296.0,1,-nbitq), 
to_sfixed(281537828.0/4294967296.0,1,-nbitq), 
to_sfixed(-325498703.0/4294967296.0,1,-nbitq), 
to_sfixed(-889440856.0/4294967296.0,1,-nbitq), 
to_sfixed(359837889.0/4294967296.0,1,-nbitq), 
to_sfixed(1370916356.0/4294967296.0,1,-nbitq), 
to_sfixed(46942669.0/4294967296.0,1,-nbitq), 
to_sfixed(553988179.0/4294967296.0,1,-nbitq), 
to_sfixed(-400012738.0/4294967296.0,1,-nbitq), 
to_sfixed(-141144057.0/4294967296.0,1,-nbitq), 
to_sfixed(-726653515.0/4294967296.0,1,-nbitq), 
to_sfixed(-210465233.0/4294967296.0,1,-nbitq), 
to_sfixed(137852869.0/4294967296.0,1,-nbitq), 
to_sfixed(204348409.0/4294967296.0,1,-nbitq), 
to_sfixed(-1447373206.0/4294967296.0,1,-nbitq), 
to_sfixed(974500201.0/4294967296.0,1,-nbitq), 
to_sfixed(-533514191.0/4294967296.0,1,-nbitq), 
to_sfixed(207769704.0/4294967296.0,1,-nbitq), 
to_sfixed(-158275151.0/4294967296.0,1,-nbitq), 
to_sfixed(-2026050718.0/4294967296.0,1,-nbitq), 
to_sfixed(-1333171294.0/4294967296.0,1,-nbitq), 
to_sfixed(-140883228.0/4294967296.0,1,-nbitq), 
to_sfixed(-1300505863.0/4294967296.0,1,-nbitq), 
to_sfixed(943893046.0/4294967296.0,1,-nbitq), 
to_sfixed(289541934.0/4294967296.0,1,-nbitq), 
to_sfixed(352237367.0/4294967296.0,1,-nbitq), 
to_sfixed(129534038.0/4294967296.0,1,-nbitq), 
to_sfixed(364188931.0/4294967296.0,1,-nbitq), 
to_sfixed(-62086899.0/4294967296.0,1,-nbitq), 
to_sfixed(-1060966391.0/4294967296.0,1,-nbitq), 
to_sfixed(329404736.0/4294967296.0,1,-nbitq), 
to_sfixed(-1130334743.0/4294967296.0,1,-nbitq), 
to_sfixed(266128773.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-54320058.0/4294967296.0,1,-nbitq), 
to_sfixed(229053352.0/4294967296.0,1,-nbitq), 
to_sfixed(-581629969.0/4294967296.0,1,-nbitq), 
to_sfixed(-131185440.0/4294967296.0,1,-nbitq), 
to_sfixed(1002662684.0/4294967296.0,1,-nbitq), 
to_sfixed(-837533319.0/4294967296.0,1,-nbitq), 
to_sfixed(272413470.0/4294967296.0,1,-nbitq), 
to_sfixed(-410227379.0/4294967296.0,1,-nbitq), 
to_sfixed(-2248325749.0/4294967296.0,1,-nbitq), 
to_sfixed(-116021716.0/4294967296.0,1,-nbitq), 
to_sfixed(-1433030454.0/4294967296.0,1,-nbitq), 
to_sfixed(-858876016.0/4294967296.0,1,-nbitq), 
to_sfixed(-343570382.0/4294967296.0,1,-nbitq), 
to_sfixed(1418768935.0/4294967296.0,1,-nbitq), 
to_sfixed(-94431253.0/4294967296.0,1,-nbitq), 
to_sfixed(1353745534.0/4294967296.0,1,-nbitq), 
to_sfixed(-407417725.0/4294967296.0,1,-nbitq), 
to_sfixed(-323386776.0/4294967296.0,1,-nbitq), 
to_sfixed(1624196178.0/4294967296.0,1,-nbitq), 
to_sfixed(188103151.0/4294967296.0,1,-nbitq), 
to_sfixed(-347942854.0/4294967296.0,1,-nbitq), 
to_sfixed(-211924530.0/4294967296.0,1,-nbitq), 
to_sfixed(-71795986.0/4294967296.0,1,-nbitq), 
to_sfixed(343292925.0/4294967296.0,1,-nbitq), 
to_sfixed(-36136799.0/4294967296.0,1,-nbitq), 
to_sfixed(-1036772994.0/4294967296.0,1,-nbitq), 
to_sfixed(-347445222.0/4294967296.0,1,-nbitq), 
to_sfixed(982024030.0/4294967296.0,1,-nbitq), 
to_sfixed(1210324802.0/4294967296.0,1,-nbitq), 
to_sfixed(1483201889.0/4294967296.0,1,-nbitq), 
to_sfixed(75462224.0/4294967296.0,1,-nbitq), 
to_sfixed(485751568.0/4294967296.0,1,-nbitq), 
to_sfixed(-250794435.0/4294967296.0,1,-nbitq), 
to_sfixed(1460704446.0/4294967296.0,1,-nbitq), 
to_sfixed(32002201.0/4294967296.0,1,-nbitq), 
to_sfixed(-158163601.0/4294967296.0,1,-nbitq), 
to_sfixed(409222101.0/4294967296.0,1,-nbitq), 
to_sfixed(819704256.0/4294967296.0,1,-nbitq), 
to_sfixed(-742981221.0/4294967296.0,1,-nbitq), 
to_sfixed(-186125292.0/4294967296.0,1,-nbitq), 
to_sfixed(-234334998.0/4294967296.0,1,-nbitq), 
to_sfixed(-162674558.0/4294967296.0,1,-nbitq), 
to_sfixed(-684079121.0/4294967296.0,1,-nbitq), 
to_sfixed(396579168.0/4294967296.0,1,-nbitq), 
to_sfixed(-40364646.0/4294967296.0,1,-nbitq), 
to_sfixed(92303807.0/4294967296.0,1,-nbitq), 
to_sfixed(-140300328.0/4294967296.0,1,-nbitq), 
to_sfixed(612133994.0/4294967296.0,1,-nbitq), 
to_sfixed(334723991.0/4294967296.0,1,-nbitq), 
to_sfixed(-910364226.0/4294967296.0,1,-nbitq), 
to_sfixed(-739724114.0/4294967296.0,1,-nbitq), 
to_sfixed(-7370697.0/4294967296.0,1,-nbitq), 
to_sfixed(1817160718.0/4294967296.0,1,-nbitq), 
to_sfixed(432574027.0/4294967296.0,1,-nbitq), 
to_sfixed(1626013165.0/4294967296.0,1,-nbitq), 
to_sfixed(-737725349.0/4294967296.0,1,-nbitq), 
to_sfixed(435980872.0/4294967296.0,1,-nbitq), 
to_sfixed(-1357537256.0/4294967296.0,1,-nbitq), 
to_sfixed(-14082796.0/4294967296.0,1,-nbitq), 
to_sfixed(-167589899.0/4294967296.0,1,-nbitq), 
to_sfixed(276548630.0/4294967296.0,1,-nbitq), 
to_sfixed(-1733207899.0/4294967296.0,1,-nbitq), 
to_sfixed(164050677.0/4294967296.0,1,-nbitq), 
to_sfixed(-212048535.0/4294967296.0,1,-nbitq), 
to_sfixed(-300806539.0/4294967296.0,1,-nbitq), 
to_sfixed(-36979732.0/4294967296.0,1,-nbitq), 
to_sfixed(764145376.0/4294967296.0,1,-nbitq), 
to_sfixed(-1439482214.0/4294967296.0,1,-nbitq), 
to_sfixed(-113921567.0/4294967296.0,1,-nbitq), 
to_sfixed(-1365129443.0/4294967296.0,1,-nbitq), 
to_sfixed(1232098150.0/4294967296.0,1,-nbitq), 
to_sfixed(-142335331.0/4294967296.0,1,-nbitq), 
to_sfixed(236900569.0/4294967296.0,1,-nbitq), 
to_sfixed(-137242957.0/4294967296.0,1,-nbitq), 
to_sfixed(-203258997.0/4294967296.0,1,-nbitq), 
to_sfixed(158043214.0/4294967296.0,1,-nbitq), 
to_sfixed(-374960825.0/4294967296.0,1,-nbitq), 
to_sfixed(512989914.0/4294967296.0,1,-nbitq), 
to_sfixed(-142206154.0/4294967296.0,1,-nbitq), 
to_sfixed(-49078818.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(56121541.0/4294967296.0,1,-nbitq), 
to_sfixed(-412195554.0/4294967296.0,1,-nbitq), 
to_sfixed(-955828705.0/4294967296.0,1,-nbitq), 
to_sfixed(260558166.0/4294967296.0,1,-nbitq), 
to_sfixed(2005822279.0/4294967296.0,1,-nbitq), 
to_sfixed(-705524368.0/4294967296.0,1,-nbitq), 
to_sfixed(2756042.0/4294967296.0,1,-nbitq), 
to_sfixed(-1495706444.0/4294967296.0,1,-nbitq), 
to_sfixed(-2000342174.0/4294967296.0,1,-nbitq), 
to_sfixed(302455027.0/4294967296.0,1,-nbitq), 
to_sfixed(-1367122555.0/4294967296.0,1,-nbitq), 
to_sfixed(113203050.0/4294967296.0,1,-nbitq), 
to_sfixed(-1457672976.0/4294967296.0,1,-nbitq), 
to_sfixed(53905925.0/4294967296.0,1,-nbitq), 
to_sfixed(260432624.0/4294967296.0,1,-nbitq), 
to_sfixed(1973092953.0/4294967296.0,1,-nbitq), 
to_sfixed(96380847.0/4294967296.0,1,-nbitq), 
to_sfixed(-113107179.0/4294967296.0,1,-nbitq), 
to_sfixed(941718416.0/4294967296.0,1,-nbitq), 
to_sfixed(653294755.0/4294967296.0,1,-nbitq), 
to_sfixed(377922816.0/4294967296.0,1,-nbitq), 
to_sfixed(-1297412968.0/4294967296.0,1,-nbitq), 
to_sfixed(-100575436.0/4294967296.0,1,-nbitq), 
to_sfixed(1213835605.0/4294967296.0,1,-nbitq), 
to_sfixed(249628551.0/4294967296.0,1,-nbitq), 
to_sfixed(-1727298325.0/4294967296.0,1,-nbitq), 
to_sfixed(-345824702.0/4294967296.0,1,-nbitq), 
to_sfixed(873485195.0/4294967296.0,1,-nbitq), 
to_sfixed(-1376255149.0/4294967296.0,1,-nbitq), 
to_sfixed(1431112811.0/4294967296.0,1,-nbitq), 
to_sfixed(1471830597.0/4294967296.0,1,-nbitq), 
to_sfixed(217752362.0/4294967296.0,1,-nbitq), 
to_sfixed(-734709808.0/4294967296.0,1,-nbitq), 
to_sfixed(1182293323.0/4294967296.0,1,-nbitq), 
to_sfixed(469588472.0/4294967296.0,1,-nbitq), 
to_sfixed(874935233.0/4294967296.0,1,-nbitq), 
to_sfixed(282576607.0/4294967296.0,1,-nbitq), 
to_sfixed(613929830.0/4294967296.0,1,-nbitq), 
to_sfixed(-216212484.0/4294967296.0,1,-nbitq), 
to_sfixed(-266753572.0/4294967296.0,1,-nbitq), 
to_sfixed(-992667819.0/4294967296.0,1,-nbitq), 
to_sfixed(-476259799.0/4294967296.0,1,-nbitq), 
to_sfixed(-1186827399.0/4294967296.0,1,-nbitq), 
to_sfixed(296952475.0/4294967296.0,1,-nbitq), 
to_sfixed(38012726.0/4294967296.0,1,-nbitq), 
to_sfixed(-327589188.0/4294967296.0,1,-nbitq), 
to_sfixed(222990761.0/4294967296.0,1,-nbitq), 
to_sfixed(-55151339.0/4294967296.0,1,-nbitq), 
to_sfixed(-407528626.0/4294967296.0,1,-nbitq), 
to_sfixed(-1092881693.0/4294967296.0,1,-nbitq), 
to_sfixed(-581882138.0/4294967296.0,1,-nbitq), 
to_sfixed(307741691.0/4294967296.0,1,-nbitq), 
to_sfixed(1356294616.0/4294967296.0,1,-nbitq), 
to_sfixed(-527764420.0/4294967296.0,1,-nbitq), 
to_sfixed(2199794836.0/4294967296.0,1,-nbitq), 
to_sfixed(-671919892.0/4294967296.0,1,-nbitq), 
to_sfixed(117356363.0/4294967296.0,1,-nbitq), 
to_sfixed(-329724344.0/4294967296.0,1,-nbitq), 
to_sfixed(-167252413.0/4294967296.0,1,-nbitq), 
to_sfixed(152301542.0/4294967296.0,1,-nbitq), 
to_sfixed(77767917.0/4294967296.0,1,-nbitq), 
to_sfixed(-1332134964.0/4294967296.0,1,-nbitq), 
to_sfixed(-1157388987.0/4294967296.0,1,-nbitq), 
to_sfixed(-265125268.0/4294967296.0,1,-nbitq), 
to_sfixed(-71013309.0/4294967296.0,1,-nbitq), 
to_sfixed(-3491787.0/4294967296.0,1,-nbitq), 
to_sfixed(1827495460.0/4294967296.0,1,-nbitq), 
to_sfixed(-1018232550.0/4294967296.0,1,-nbitq), 
to_sfixed(7446697.0/4294967296.0,1,-nbitq), 
to_sfixed(-890036647.0/4294967296.0,1,-nbitq), 
to_sfixed(1100061994.0/4294967296.0,1,-nbitq), 
to_sfixed(-7821965.0/4294967296.0,1,-nbitq), 
to_sfixed(-375476973.0/4294967296.0,1,-nbitq), 
to_sfixed(59436386.0/4294967296.0,1,-nbitq), 
to_sfixed(-306812919.0/4294967296.0,1,-nbitq), 
to_sfixed(987918464.0/4294967296.0,1,-nbitq), 
to_sfixed(-543223507.0/4294967296.0,1,-nbitq), 
to_sfixed(616116936.0/4294967296.0,1,-nbitq), 
to_sfixed(862567200.0/4294967296.0,1,-nbitq), 
to_sfixed(-224214470.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-188994358.0/4294967296.0,1,-nbitq), 
to_sfixed(-707567230.0/4294967296.0,1,-nbitq), 
to_sfixed(-496825129.0/4294967296.0,1,-nbitq), 
to_sfixed(-66764281.0/4294967296.0,1,-nbitq), 
to_sfixed(2517142863.0/4294967296.0,1,-nbitq), 
to_sfixed(-410251609.0/4294967296.0,1,-nbitq), 
to_sfixed(116222238.0/4294967296.0,1,-nbitq), 
to_sfixed(-983917609.0/4294967296.0,1,-nbitq), 
to_sfixed(-2318991618.0/4294967296.0,1,-nbitq), 
to_sfixed(-385711379.0/4294967296.0,1,-nbitq), 
to_sfixed(-1079406653.0/4294967296.0,1,-nbitq), 
to_sfixed(674352865.0/4294967296.0,1,-nbitq), 
to_sfixed(-172103721.0/4294967296.0,1,-nbitq), 
to_sfixed(-708699717.0/4294967296.0,1,-nbitq), 
to_sfixed(386024172.0/4294967296.0,1,-nbitq), 
to_sfixed(896219480.0/4294967296.0,1,-nbitq), 
to_sfixed(3211034.0/4294967296.0,1,-nbitq), 
to_sfixed(233495525.0/4294967296.0,1,-nbitq), 
to_sfixed(-109168586.0/4294967296.0,1,-nbitq), 
to_sfixed(80598840.0/4294967296.0,1,-nbitq), 
to_sfixed(-96612381.0/4294967296.0,1,-nbitq), 
to_sfixed(-1514771026.0/4294967296.0,1,-nbitq), 
to_sfixed(1039221937.0/4294967296.0,1,-nbitq), 
to_sfixed(1722000713.0/4294967296.0,1,-nbitq), 
to_sfixed(-127569075.0/4294967296.0,1,-nbitq), 
to_sfixed(-936686702.0/4294967296.0,1,-nbitq), 
to_sfixed(-276498683.0/4294967296.0,1,-nbitq), 
to_sfixed(204314432.0/4294967296.0,1,-nbitq), 
to_sfixed(-2347003620.0/4294967296.0,1,-nbitq), 
to_sfixed(1048082307.0/4294967296.0,1,-nbitq), 
to_sfixed(1831031808.0/4294967296.0,1,-nbitq), 
to_sfixed(-16574187.0/4294967296.0,1,-nbitq), 
to_sfixed(-314891627.0/4294967296.0,1,-nbitq), 
to_sfixed(576206090.0/4294967296.0,1,-nbitq), 
to_sfixed(269376818.0/4294967296.0,1,-nbitq), 
to_sfixed(2164068744.0/4294967296.0,1,-nbitq), 
to_sfixed(81114345.0/4294967296.0,1,-nbitq), 
to_sfixed(520681169.0/4294967296.0,1,-nbitq), 
to_sfixed(350205694.0/4294967296.0,1,-nbitq), 
to_sfixed(-52741689.0/4294967296.0,1,-nbitq), 
to_sfixed(181282568.0/4294967296.0,1,-nbitq), 
to_sfixed(-799540796.0/4294967296.0,1,-nbitq), 
to_sfixed(-1188810828.0/4294967296.0,1,-nbitq), 
to_sfixed(1365992819.0/4294967296.0,1,-nbitq), 
to_sfixed(-366841429.0/4294967296.0,1,-nbitq), 
to_sfixed(-1070448249.0/4294967296.0,1,-nbitq), 
to_sfixed(117524644.0/4294967296.0,1,-nbitq), 
to_sfixed(338181828.0/4294967296.0,1,-nbitq), 
to_sfixed(217365678.0/4294967296.0,1,-nbitq), 
to_sfixed(-623730871.0/4294967296.0,1,-nbitq), 
to_sfixed(-1062942483.0/4294967296.0,1,-nbitq), 
to_sfixed(-62997681.0/4294967296.0,1,-nbitq), 
to_sfixed(1077798380.0/4294967296.0,1,-nbitq), 
to_sfixed(-259499758.0/4294967296.0,1,-nbitq), 
to_sfixed(2280108768.0/4294967296.0,1,-nbitq), 
to_sfixed(-567099326.0/4294967296.0,1,-nbitq), 
to_sfixed(32066058.0/4294967296.0,1,-nbitq), 
to_sfixed(-1364574238.0/4294967296.0,1,-nbitq), 
to_sfixed(-150118452.0/4294967296.0,1,-nbitq), 
to_sfixed(73523789.0/4294967296.0,1,-nbitq), 
to_sfixed(324739567.0/4294967296.0,1,-nbitq), 
to_sfixed(-68664043.0/4294967296.0,1,-nbitq), 
to_sfixed(-1506901551.0/4294967296.0,1,-nbitq), 
to_sfixed(-608043443.0/4294967296.0,1,-nbitq), 
to_sfixed(187063424.0/4294967296.0,1,-nbitq), 
to_sfixed(-195317695.0/4294967296.0,1,-nbitq), 
to_sfixed(301597771.0/4294967296.0,1,-nbitq), 
to_sfixed(177089506.0/4294967296.0,1,-nbitq), 
to_sfixed(104299287.0/4294967296.0,1,-nbitq), 
to_sfixed(-44334477.0/4294967296.0,1,-nbitq), 
to_sfixed(1230049842.0/4294967296.0,1,-nbitq), 
to_sfixed(-140135772.0/4294967296.0,1,-nbitq), 
to_sfixed(-711676264.0/4294967296.0,1,-nbitq), 
to_sfixed(-297923913.0/4294967296.0,1,-nbitq), 
to_sfixed(170440169.0/4294967296.0,1,-nbitq), 
to_sfixed(667547178.0/4294967296.0,1,-nbitq), 
to_sfixed(103774309.0/4294967296.0,1,-nbitq), 
to_sfixed(713449674.0/4294967296.0,1,-nbitq), 
to_sfixed(1323345442.0/4294967296.0,1,-nbitq), 
to_sfixed(16194008.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(370290091.0/4294967296.0,1,-nbitq), 
to_sfixed(59717123.0/4294967296.0,1,-nbitq), 
to_sfixed(195297172.0/4294967296.0,1,-nbitq), 
to_sfixed(-911903719.0/4294967296.0,1,-nbitq), 
to_sfixed(1595287046.0/4294967296.0,1,-nbitq), 
to_sfixed(418889469.0/4294967296.0,1,-nbitq), 
to_sfixed(527353399.0/4294967296.0,1,-nbitq), 
to_sfixed(-208364209.0/4294967296.0,1,-nbitq), 
to_sfixed(-2277442942.0/4294967296.0,1,-nbitq), 
to_sfixed(35014749.0/4294967296.0,1,-nbitq), 
to_sfixed(-54075023.0/4294967296.0,1,-nbitq), 
to_sfixed(1011350960.0/4294967296.0,1,-nbitq), 
to_sfixed(-798636087.0/4294967296.0,1,-nbitq), 
to_sfixed(-1290884539.0/4294967296.0,1,-nbitq), 
to_sfixed(-85696371.0/4294967296.0,1,-nbitq), 
to_sfixed(315685594.0/4294967296.0,1,-nbitq), 
to_sfixed(220469039.0/4294967296.0,1,-nbitq), 
to_sfixed(-381446359.0/4294967296.0,1,-nbitq), 
to_sfixed(-1600714718.0/4294967296.0,1,-nbitq), 
to_sfixed(-535699203.0/4294967296.0,1,-nbitq), 
to_sfixed(-215832470.0/4294967296.0,1,-nbitq), 
to_sfixed(-756480793.0/4294967296.0,1,-nbitq), 
to_sfixed(1592785235.0/4294967296.0,1,-nbitq), 
to_sfixed(-558989352.0/4294967296.0,1,-nbitq), 
to_sfixed(-186564668.0/4294967296.0,1,-nbitq), 
to_sfixed(191053825.0/4294967296.0,1,-nbitq), 
to_sfixed(-452126555.0/4294967296.0,1,-nbitq), 
to_sfixed(-728085818.0/4294967296.0,1,-nbitq), 
to_sfixed(-563372634.0/4294967296.0,1,-nbitq), 
to_sfixed(931468953.0/4294967296.0,1,-nbitq), 
to_sfixed(310004854.0/4294967296.0,1,-nbitq), 
to_sfixed(297912646.0/4294967296.0,1,-nbitq), 
to_sfixed(-679416143.0/4294967296.0,1,-nbitq), 
to_sfixed(243162269.0/4294967296.0,1,-nbitq), 
to_sfixed(643451960.0/4294967296.0,1,-nbitq), 
to_sfixed(554920674.0/4294967296.0,1,-nbitq), 
to_sfixed(612322204.0/4294967296.0,1,-nbitq), 
to_sfixed(-903613315.0/4294967296.0,1,-nbitq), 
to_sfixed(696611153.0/4294967296.0,1,-nbitq), 
to_sfixed(187499190.0/4294967296.0,1,-nbitq), 
to_sfixed(730740338.0/4294967296.0,1,-nbitq), 
to_sfixed(-113965367.0/4294967296.0,1,-nbitq), 
to_sfixed(-620425802.0/4294967296.0,1,-nbitq), 
to_sfixed(2025690622.0/4294967296.0,1,-nbitq), 
to_sfixed(-991093928.0/4294967296.0,1,-nbitq), 
to_sfixed(-775152693.0/4294967296.0,1,-nbitq), 
to_sfixed(152363463.0/4294967296.0,1,-nbitq), 
to_sfixed(562661382.0/4294967296.0,1,-nbitq), 
to_sfixed(54019495.0/4294967296.0,1,-nbitq), 
to_sfixed(-1010974938.0/4294967296.0,1,-nbitq), 
to_sfixed(-1106141253.0/4294967296.0,1,-nbitq), 
to_sfixed(-241745631.0/4294967296.0,1,-nbitq), 
to_sfixed(93209796.0/4294967296.0,1,-nbitq), 
to_sfixed(-1265258633.0/4294967296.0,1,-nbitq), 
to_sfixed(-769025113.0/4294967296.0,1,-nbitq), 
to_sfixed(747821737.0/4294967296.0,1,-nbitq), 
to_sfixed(-1144442204.0/4294967296.0,1,-nbitq), 
to_sfixed(-1015737773.0/4294967296.0,1,-nbitq), 
to_sfixed(-378386634.0/4294967296.0,1,-nbitq), 
to_sfixed(12770541.0/4294967296.0,1,-nbitq), 
to_sfixed(-193162219.0/4294967296.0,1,-nbitq), 
to_sfixed(79777033.0/4294967296.0,1,-nbitq), 
to_sfixed(-434435446.0/4294967296.0,1,-nbitq), 
to_sfixed(-58598257.0/4294967296.0,1,-nbitq), 
to_sfixed(288019810.0/4294967296.0,1,-nbitq), 
to_sfixed(35325756.0/4294967296.0,1,-nbitq), 
to_sfixed(694381679.0/4294967296.0,1,-nbitq), 
to_sfixed(1151320894.0/4294967296.0,1,-nbitq), 
to_sfixed(-133167642.0/4294967296.0,1,-nbitq), 
to_sfixed(554089724.0/4294967296.0,1,-nbitq), 
to_sfixed(1823442662.0/4294967296.0,1,-nbitq), 
to_sfixed(-6293082.0/4294967296.0,1,-nbitq), 
to_sfixed(-899569881.0/4294967296.0,1,-nbitq), 
to_sfixed(-108907930.0/4294967296.0,1,-nbitq), 
to_sfixed(336673555.0/4294967296.0,1,-nbitq), 
to_sfixed(-42558151.0/4294967296.0,1,-nbitq), 
to_sfixed(277548807.0/4294967296.0,1,-nbitq), 
to_sfixed(88540959.0/4294967296.0,1,-nbitq), 
to_sfixed(815860724.0/4294967296.0,1,-nbitq), 
to_sfixed(-87169726.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(94654624.0/4294967296.0,1,-nbitq), 
to_sfixed(442843863.0/4294967296.0,1,-nbitq), 
to_sfixed(287612294.0/4294967296.0,1,-nbitq), 
to_sfixed(-449786567.0/4294967296.0,1,-nbitq), 
to_sfixed(366019151.0/4294967296.0,1,-nbitq), 
to_sfixed(1096623439.0/4294967296.0,1,-nbitq), 
to_sfixed(-59894893.0/4294967296.0,1,-nbitq), 
to_sfixed(364747943.0/4294967296.0,1,-nbitq), 
to_sfixed(-1757850146.0/4294967296.0,1,-nbitq), 
to_sfixed(228460476.0/4294967296.0,1,-nbitq), 
to_sfixed(-484735327.0/4294967296.0,1,-nbitq), 
to_sfixed(1501657563.0/4294967296.0,1,-nbitq), 
to_sfixed(-627917157.0/4294967296.0,1,-nbitq), 
to_sfixed(-2138402906.0/4294967296.0,1,-nbitq), 
to_sfixed(-136397521.0/4294967296.0,1,-nbitq), 
to_sfixed(477051000.0/4294967296.0,1,-nbitq), 
to_sfixed(-221674305.0/4294967296.0,1,-nbitq), 
to_sfixed(187325562.0/4294967296.0,1,-nbitq), 
to_sfixed(-1955271434.0/4294967296.0,1,-nbitq), 
to_sfixed(-700238404.0/4294967296.0,1,-nbitq), 
to_sfixed(292082334.0/4294967296.0,1,-nbitq), 
to_sfixed(-401594176.0/4294967296.0,1,-nbitq), 
to_sfixed(1296356564.0/4294967296.0,1,-nbitq), 
to_sfixed(-1186763738.0/4294967296.0,1,-nbitq), 
to_sfixed(100481632.0/4294967296.0,1,-nbitq), 
to_sfixed(242419310.0/4294967296.0,1,-nbitq), 
to_sfixed(-80219414.0/4294967296.0,1,-nbitq), 
to_sfixed(-1055515766.0/4294967296.0,1,-nbitq), 
to_sfixed(965053490.0/4294967296.0,1,-nbitq), 
to_sfixed(464904600.0/4294967296.0,1,-nbitq), 
to_sfixed(-2111823513.0/4294967296.0,1,-nbitq), 
to_sfixed(-401363286.0/4294967296.0,1,-nbitq), 
to_sfixed(-140079544.0/4294967296.0,1,-nbitq), 
to_sfixed(8081392.0/4294967296.0,1,-nbitq), 
to_sfixed(1038270854.0/4294967296.0,1,-nbitq), 
to_sfixed(137025635.0/4294967296.0,1,-nbitq), 
to_sfixed(581724321.0/4294967296.0,1,-nbitq), 
to_sfixed(-699070280.0/4294967296.0,1,-nbitq), 
to_sfixed(216497836.0/4294967296.0,1,-nbitq), 
to_sfixed(-158616123.0/4294967296.0,1,-nbitq), 
to_sfixed(992667588.0/4294967296.0,1,-nbitq), 
to_sfixed(541824790.0/4294967296.0,1,-nbitq), 
to_sfixed(-566532482.0/4294967296.0,1,-nbitq), 
to_sfixed(2591173628.0/4294967296.0,1,-nbitq), 
to_sfixed(127318333.0/4294967296.0,1,-nbitq), 
to_sfixed(-190853770.0/4294967296.0,1,-nbitq), 
to_sfixed(-360227382.0/4294967296.0,1,-nbitq), 
to_sfixed(707279670.0/4294967296.0,1,-nbitq), 
to_sfixed(-491201259.0/4294967296.0,1,-nbitq), 
to_sfixed(-307174823.0/4294967296.0,1,-nbitq), 
to_sfixed(-653408847.0/4294967296.0,1,-nbitq), 
to_sfixed(339136678.0/4294967296.0,1,-nbitq), 
to_sfixed(134461224.0/4294967296.0,1,-nbitq), 
to_sfixed(-1144570140.0/4294967296.0,1,-nbitq), 
to_sfixed(-1604753762.0/4294967296.0,1,-nbitq), 
to_sfixed(341936766.0/4294967296.0,1,-nbitq), 
to_sfixed(-1467163403.0/4294967296.0,1,-nbitq), 
to_sfixed(127837000.0/4294967296.0,1,-nbitq), 
to_sfixed(370064122.0/4294967296.0,1,-nbitq), 
to_sfixed(-327292583.0/4294967296.0,1,-nbitq), 
to_sfixed(-199891248.0/4294967296.0,1,-nbitq), 
to_sfixed(1075084920.0/4294967296.0,1,-nbitq), 
to_sfixed(-353988387.0/4294967296.0,1,-nbitq), 
to_sfixed(-465216801.0/4294967296.0,1,-nbitq), 
to_sfixed(-484813371.0/4294967296.0,1,-nbitq), 
to_sfixed(159841144.0/4294967296.0,1,-nbitq), 
to_sfixed(1420178135.0/4294967296.0,1,-nbitq), 
to_sfixed(1437307492.0/4294967296.0,1,-nbitq), 
to_sfixed(333365218.0/4294967296.0,1,-nbitq), 
to_sfixed(1008914264.0/4294967296.0,1,-nbitq), 
to_sfixed(2592961060.0/4294967296.0,1,-nbitq), 
to_sfixed(-217217482.0/4294967296.0,1,-nbitq), 
to_sfixed(-1659257907.0/4294967296.0,1,-nbitq), 
to_sfixed(125031216.0/4294967296.0,1,-nbitq), 
to_sfixed(-16638193.0/4294967296.0,1,-nbitq), 
to_sfixed(-801948115.0/4294967296.0,1,-nbitq), 
to_sfixed(391409319.0/4294967296.0,1,-nbitq), 
to_sfixed(-53980204.0/4294967296.0,1,-nbitq), 
to_sfixed(920571232.0/4294967296.0,1,-nbitq), 
to_sfixed(-314018125.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-68304999.0/4294967296.0,1,-nbitq), 
to_sfixed(1111102047.0/4294967296.0,1,-nbitq), 
to_sfixed(-1550550639.0/4294967296.0,1,-nbitq), 
to_sfixed(983471500.0/4294967296.0,1,-nbitq), 
to_sfixed(-1881278628.0/4294967296.0,1,-nbitq), 
to_sfixed(1381295185.0/4294967296.0,1,-nbitq), 
to_sfixed(-470394823.0/4294967296.0,1,-nbitq), 
to_sfixed(645744821.0/4294967296.0,1,-nbitq), 
to_sfixed(-1694396262.0/4294967296.0,1,-nbitq), 
to_sfixed(-94062942.0/4294967296.0,1,-nbitq), 
to_sfixed(-253238410.0/4294967296.0,1,-nbitq), 
to_sfixed(1193939375.0/4294967296.0,1,-nbitq), 
to_sfixed(-423265518.0/4294967296.0,1,-nbitq), 
to_sfixed(-2983161471.0/4294967296.0,1,-nbitq), 
to_sfixed(-283231321.0/4294967296.0,1,-nbitq), 
to_sfixed(482357153.0/4294967296.0,1,-nbitq), 
to_sfixed(-253533882.0/4294967296.0,1,-nbitq), 
to_sfixed(-342035851.0/4294967296.0,1,-nbitq), 
to_sfixed(-1767802752.0/4294967296.0,1,-nbitq), 
to_sfixed(-640128987.0/4294967296.0,1,-nbitq), 
to_sfixed(-35342113.0/4294967296.0,1,-nbitq), 
to_sfixed(-584866514.0/4294967296.0,1,-nbitq), 
to_sfixed(-440000231.0/4294967296.0,1,-nbitq), 
to_sfixed(-517047882.0/4294967296.0,1,-nbitq), 
to_sfixed(96186466.0/4294967296.0,1,-nbitq), 
to_sfixed(320683529.0/4294967296.0,1,-nbitq), 
to_sfixed(-171682230.0/4294967296.0,1,-nbitq), 
to_sfixed(-301327120.0/4294967296.0,1,-nbitq), 
to_sfixed(117652329.0/4294967296.0,1,-nbitq), 
to_sfixed(1104302286.0/4294967296.0,1,-nbitq), 
to_sfixed(-2497102629.0/4294967296.0,1,-nbitq), 
to_sfixed(-878592860.0/4294967296.0,1,-nbitq), 
to_sfixed(-228068319.0/4294967296.0,1,-nbitq), 
to_sfixed(-295298513.0/4294967296.0,1,-nbitq), 
to_sfixed(156716720.0/4294967296.0,1,-nbitq), 
to_sfixed(-186675627.0/4294967296.0,1,-nbitq), 
to_sfixed(271119236.0/4294967296.0,1,-nbitq), 
to_sfixed(-356199190.0/4294967296.0,1,-nbitq), 
to_sfixed(581003262.0/4294967296.0,1,-nbitq), 
to_sfixed(296636412.0/4294967296.0,1,-nbitq), 
to_sfixed(1127573447.0/4294967296.0,1,-nbitq), 
to_sfixed(1237276459.0/4294967296.0,1,-nbitq), 
to_sfixed(-611496188.0/4294967296.0,1,-nbitq), 
to_sfixed(425764495.0/4294967296.0,1,-nbitq), 
to_sfixed(215494028.0/4294967296.0,1,-nbitq), 
to_sfixed(-226056416.0/4294967296.0,1,-nbitq), 
to_sfixed(-224333653.0/4294967296.0,1,-nbitq), 
to_sfixed(542695335.0/4294967296.0,1,-nbitq), 
to_sfixed(85657805.0/4294967296.0,1,-nbitq), 
to_sfixed(1502514523.0/4294967296.0,1,-nbitq), 
to_sfixed(-482138753.0/4294967296.0,1,-nbitq), 
to_sfixed(609006347.0/4294967296.0,1,-nbitq), 
to_sfixed(174892809.0/4294967296.0,1,-nbitq), 
to_sfixed(81924068.0/4294967296.0,1,-nbitq), 
to_sfixed(-702241754.0/4294967296.0,1,-nbitq), 
to_sfixed(325105476.0/4294967296.0,1,-nbitq), 
to_sfixed(-1151363844.0/4294967296.0,1,-nbitq), 
to_sfixed(10800435.0/4294967296.0,1,-nbitq), 
to_sfixed(-306388129.0/4294967296.0,1,-nbitq), 
to_sfixed(-192906306.0/4294967296.0,1,-nbitq), 
to_sfixed(254204544.0/4294967296.0,1,-nbitq), 
to_sfixed(1036385766.0/4294967296.0,1,-nbitq), 
to_sfixed(672193522.0/4294967296.0,1,-nbitq), 
to_sfixed(-207141785.0/4294967296.0,1,-nbitq), 
to_sfixed(-358539760.0/4294967296.0,1,-nbitq), 
to_sfixed(456768596.0/4294967296.0,1,-nbitq), 
to_sfixed(-915339234.0/4294967296.0,1,-nbitq), 
to_sfixed(329824920.0/4294967296.0,1,-nbitq), 
to_sfixed(221646890.0/4294967296.0,1,-nbitq), 
to_sfixed(1914451998.0/4294967296.0,1,-nbitq), 
to_sfixed(1742080203.0/4294967296.0,1,-nbitq), 
to_sfixed(84637625.0/4294967296.0,1,-nbitq), 
to_sfixed(-1461090962.0/4294967296.0,1,-nbitq), 
to_sfixed(201305081.0/4294967296.0,1,-nbitq), 
to_sfixed(-94036576.0/4294967296.0,1,-nbitq), 
to_sfixed(-1165156037.0/4294967296.0,1,-nbitq), 
to_sfixed(332360065.0/4294967296.0,1,-nbitq), 
to_sfixed(660325603.0/4294967296.0,1,-nbitq), 
to_sfixed(273875803.0/4294967296.0,1,-nbitq), 
to_sfixed(346817204.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-273056988.0/4294967296.0,1,-nbitq), 
to_sfixed(760718689.0/4294967296.0,1,-nbitq), 
to_sfixed(-1237769198.0/4294967296.0,1,-nbitq), 
to_sfixed(2635532944.0/4294967296.0,1,-nbitq), 
to_sfixed(-2463896042.0/4294967296.0,1,-nbitq), 
to_sfixed(1561133886.0/4294967296.0,1,-nbitq), 
to_sfixed(-358896611.0/4294967296.0,1,-nbitq), 
to_sfixed(697869073.0/4294967296.0,1,-nbitq), 
to_sfixed(-980245454.0/4294967296.0,1,-nbitq), 
to_sfixed(26689863.0/4294967296.0,1,-nbitq), 
to_sfixed(461261078.0/4294967296.0,1,-nbitq), 
to_sfixed(632022052.0/4294967296.0,1,-nbitq), 
to_sfixed(900947721.0/4294967296.0,1,-nbitq), 
to_sfixed(-2609812941.0/4294967296.0,1,-nbitq), 
to_sfixed(131690956.0/4294967296.0,1,-nbitq), 
to_sfixed(117047831.0/4294967296.0,1,-nbitq), 
to_sfixed(-339135987.0/4294967296.0,1,-nbitq), 
to_sfixed(-129875577.0/4294967296.0,1,-nbitq), 
to_sfixed(-2123972742.0/4294967296.0,1,-nbitq), 
to_sfixed(-241984824.0/4294967296.0,1,-nbitq), 
to_sfixed(-351167343.0/4294967296.0,1,-nbitq), 
to_sfixed(287212466.0/4294967296.0,1,-nbitq), 
to_sfixed(-182077337.0/4294967296.0,1,-nbitq), 
to_sfixed(-520972589.0/4294967296.0,1,-nbitq), 
to_sfixed(-179022199.0/4294967296.0,1,-nbitq), 
to_sfixed(1219956802.0/4294967296.0,1,-nbitq), 
to_sfixed(-266992293.0/4294967296.0,1,-nbitq), 
to_sfixed(48745019.0/4294967296.0,1,-nbitq), 
to_sfixed(-685551645.0/4294967296.0,1,-nbitq), 
to_sfixed(2200570220.0/4294967296.0,1,-nbitq), 
to_sfixed(-832482105.0/4294967296.0,1,-nbitq), 
to_sfixed(1019338234.0/4294967296.0,1,-nbitq), 
to_sfixed(999393658.0/4294967296.0,1,-nbitq), 
to_sfixed(116673636.0/4294967296.0,1,-nbitq), 
to_sfixed(-1046993435.0/4294967296.0,1,-nbitq), 
to_sfixed(-1138373659.0/4294967296.0,1,-nbitq), 
to_sfixed(-515980928.0/4294967296.0,1,-nbitq), 
to_sfixed(-609021210.0/4294967296.0,1,-nbitq), 
to_sfixed(672292650.0/4294967296.0,1,-nbitq), 
to_sfixed(58307483.0/4294967296.0,1,-nbitq), 
to_sfixed(-791653172.0/4294967296.0,1,-nbitq), 
to_sfixed(1498927530.0/4294967296.0,1,-nbitq), 
to_sfixed(-1101472759.0/4294967296.0,1,-nbitq), 
to_sfixed(-441934734.0/4294967296.0,1,-nbitq), 
to_sfixed(-541090615.0/4294967296.0,1,-nbitq), 
to_sfixed(-1225938375.0/4294967296.0,1,-nbitq), 
to_sfixed(164016147.0/4294967296.0,1,-nbitq), 
to_sfixed(785073096.0/4294967296.0,1,-nbitq), 
to_sfixed(-525673726.0/4294967296.0,1,-nbitq), 
to_sfixed(12366685.0/4294967296.0,1,-nbitq), 
to_sfixed(339135273.0/4294967296.0,1,-nbitq), 
to_sfixed(710149263.0/4294967296.0,1,-nbitq), 
to_sfixed(-217433468.0/4294967296.0,1,-nbitq), 
to_sfixed(553026521.0/4294967296.0,1,-nbitq), 
to_sfixed(-1099184575.0/4294967296.0,1,-nbitq), 
to_sfixed(246128256.0/4294967296.0,1,-nbitq), 
to_sfixed(-1007773480.0/4294967296.0,1,-nbitq), 
to_sfixed(12530850.0/4294967296.0,1,-nbitq), 
to_sfixed(-26928953.0/4294967296.0,1,-nbitq), 
to_sfixed(-272148471.0/4294967296.0,1,-nbitq), 
to_sfixed(-306972608.0/4294967296.0,1,-nbitq), 
to_sfixed(804667742.0/4294967296.0,1,-nbitq), 
to_sfixed(134753900.0/4294967296.0,1,-nbitq), 
to_sfixed(72097744.0/4294967296.0,1,-nbitq), 
to_sfixed(-290272596.0/4294967296.0,1,-nbitq), 
to_sfixed(-241326908.0/4294967296.0,1,-nbitq), 
to_sfixed(-2855279402.0/4294967296.0,1,-nbitq), 
to_sfixed(-1170516833.0/4294967296.0,1,-nbitq), 
to_sfixed(2090344.0/4294967296.0,1,-nbitq), 
to_sfixed(1028653570.0/4294967296.0,1,-nbitq), 
to_sfixed(526025407.0/4294967296.0,1,-nbitq), 
to_sfixed(-179100819.0/4294967296.0,1,-nbitq), 
to_sfixed(-852531796.0/4294967296.0,1,-nbitq), 
to_sfixed(285687716.0/4294967296.0,1,-nbitq), 
to_sfixed(446214345.0/4294967296.0,1,-nbitq), 
to_sfixed(797167731.0/4294967296.0,1,-nbitq), 
to_sfixed(214046530.0/4294967296.0,1,-nbitq), 
to_sfixed(386111436.0/4294967296.0,1,-nbitq), 
to_sfixed(313961741.0/4294967296.0,1,-nbitq), 
to_sfixed(-343205064.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-419983383.0/4294967296.0,1,-nbitq), 
to_sfixed(444889570.0/4294967296.0,1,-nbitq), 
to_sfixed(-524039221.0/4294967296.0,1,-nbitq), 
to_sfixed(1988875686.0/4294967296.0,1,-nbitq), 
to_sfixed(-2267373176.0/4294967296.0,1,-nbitq), 
to_sfixed(1359485466.0/4294967296.0,1,-nbitq), 
to_sfixed(101250077.0/4294967296.0,1,-nbitq), 
to_sfixed(-147167085.0/4294967296.0,1,-nbitq), 
to_sfixed(-732769114.0/4294967296.0,1,-nbitq), 
to_sfixed(-23692985.0/4294967296.0,1,-nbitq), 
to_sfixed(-57457550.0/4294967296.0,1,-nbitq), 
to_sfixed(807261880.0/4294967296.0,1,-nbitq), 
to_sfixed(473492477.0/4294967296.0,1,-nbitq), 
to_sfixed(-1479006511.0/4294967296.0,1,-nbitq), 
to_sfixed(261521657.0/4294967296.0,1,-nbitq), 
to_sfixed(48674868.0/4294967296.0,1,-nbitq), 
to_sfixed(154801105.0/4294967296.0,1,-nbitq), 
to_sfixed(245043922.0/4294967296.0,1,-nbitq), 
to_sfixed(-1601329617.0/4294967296.0,1,-nbitq), 
to_sfixed(-147277882.0/4294967296.0,1,-nbitq), 
to_sfixed(146946967.0/4294967296.0,1,-nbitq), 
to_sfixed(253715656.0/4294967296.0,1,-nbitq), 
to_sfixed(-527445707.0/4294967296.0,1,-nbitq), 
to_sfixed(-362372809.0/4294967296.0,1,-nbitq), 
to_sfixed(-189797941.0/4294967296.0,1,-nbitq), 
to_sfixed(614322047.0/4294967296.0,1,-nbitq), 
to_sfixed(92441580.0/4294967296.0,1,-nbitq), 
to_sfixed(115474350.0/4294967296.0,1,-nbitq), 
to_sfixed(-700333370.0/4294967296.0,1,-nbitq), 
to_sfixed(2064775607.0/4294967296.0,1,-nbitq), 
to_sfixed(-543805962.0/4294967296.0,1,-nbitq), 
to_sfixed(1001060942.0/4294967296.0,1,-nbitq), 
to_sfixed(542872643.0/4294967296.0,1,-nbitq), 
to_sfixed(264311841.0/4294967296.0,1,-nbitq), 
to_sfixed(-37493821.0/4294967296.0,1,-nbitq), 
to_sfixed(-858255372.0/4294967296.0,1,-nbitq), 
to_sfixed(-1198956474.0/4294967296.0,1,-nbitq), 
to_sfixed(-358907542.0/4294967296.0,1,-nbitq), 
to_sfixed(265640804.0/4294967296.0,1,-nbitq), 
to_sfixed(559203352.0/4294967296.0,1,-nbitq), 
to_sfixed(-920794035.0/4294967296.0,1,-nbitq), 
to_sfixed(1130788108.0/4294967296.0,1,-nbitq), 
to_sfixed(-1618260064.0/4294967296.0,1,-nbitq), 
to_sfixed(-418205721.0/4294967296.0,1,-nbitq), 
to_sfixed(-704744401.0/4294967296.0,1,-nbitq), 
to_sfixed(-2096896291.0/4294967296.0,1,-nbitq), 
to_sfixed(-151022421.0/4294967296.0,1,-nbitq), 
to_sfixed(1273602853.0/4294967296.0,1,-nbitq), 
to_sfixed(-682716149.0/4294967296.0,1,-nbitq), 
to_sfixed(145576747.0/4294967296.0,1,-nbitq), 
to_sfixed(480531577.0/4294967296.0,1,-nbitq), 
to_sfixed(-70443850.0/4294967296.0,1,-nbitq), 
to_sfixed(76181727.0/4294967296.0,1,-nbitq), 
to_sfixed(644135206.0/4294967296.0,1,-nbitq), 
to_sfixed(-1888845020.0/4294967296.0,1,-nbitq), 
to_sfixed(230873194.0/4294967296.0,1,-nbitq), 
to_sfixed(-739584234.0/4294967296.0,1,-nbitq), 
to_sfixed(593137694.0/4294967296.0,1,-nbitq), 
to_sfixed(282221063.0/4294967296.0,1,-nbitq), 
to_sfixed(-64808708.0/4294967296.0,1,-nbitq), 
to_sfixed(38845383.0/4294967296.0,1,-nbitq), 
to_sfixed(826547723.0/4294967296.0,1,-nbitq), 
to_sfixed(604055637.0/4294967296.0,1,-nbitq), 
to_sfixed(469730560.0/4294967296.0,1,-nbitq), 
to_sfixed(138450425.0/4294967296.0,1,-nbitq), 
to_sfixed(272809656.0/4294967296.0,1,-nbitq), 
to_sfixed(-1469009119.0/4294967296.0,1,-nbitq), 
to_sfixed(-532219817.0/4294967296.0,1,-nbitq), 
to_sfixed(49179459.0/4294967296.0,1,-nbitq), 
to_sfixed(735641565.0/4294967296.0,1,-nbitq), 
to_sfixed(993065643.0/4294967296.0,1,-nbitq), 
to_sfixed(-419076907.0/4294967296.0,1,-nbitq), 
to_sfixed(-1589699704.0/4294967296.0,1,-nbitq), 
to_sfixed(-246412585.0/4294967296.0,1,-nbitq), 
to_sfixed(267532908.0/4294967296.0,1,-nbitq), 
to_sfixed(973566836.0/4294967296.0,1,-nbitq), 
to_sfixed(388483294.0/4294967296.0,1,-nbitq), 
to_sfixed(457031075.0/4294967296.0,1,-nbitq), 
to_sfixed(71759549.0/4294967296.0,1,-nbitq), 
to_sfixed(-265911909.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-551080222.0/4294967296.0,1,-nbitq), 
to_sfixed(92534589.0/4294967296.0,1,-nbitq), 
to_sfixed(-894594002.0/4294967296.0,1,-nbitq), 
to_sfixed(1947250053.0/4294967296.0,1,-nbitq), 
to_sfixed(-1001642416.0/4294967296.0,1,-nbitq), 
to_sfixed(954609524.0/4294967296.0,1,-nbitq), 
to_sfixed(-91971675.0/4294967296.0,1,-nbitq), 
to_sfixed(-412438197.0/4294967296.0,1,-nbitq), 
to_sfixed(-939979985.0/4294967296.0,1,-nbitq), 
to_sfixed(287316128.0/4294967296.0,1,-nbitq), 
to_sfixed(285799667.0/4294967296.0,1,-nbitq), 
to_sfixed(707835779.0/4294967296.0,1,-nbitq), 
to_sfixed(317592650.0/4294967296.0,1,-nbitq), 
to_sfixed(-1193491725.0/4294967296.0,1,-nbitq), 
to_sfixed(-146536491.0/4294967296.0,1,-nbitq), 
to_sfixed(468964526.0/4294967296.0,1,-nbitq), 
to_sfixed(-45589860.0/4294967296.0,1,-nbitq), 
to_sfixed(232513099.0/4294967296.0,1,-nbitq), 
to_sfixed(-1286870266.0/4294967296.0,1,-nbitq), 
to_sfixed(-287985358.0/4294967296.0,1,-nbitq), 
to_sfixed(128150219.0/4294967296.0,1,-nbitq), 
to_sfixed(-431894876.0/4294967296.0,1,-nbitq), 
to_sfixed(-1377221161.0/4294967296.0,1,-nbitq), 
to_sfixed(-924917083.0/4294967296.0,1,-nbitq), 
to_sfixed(244411128.0/4294967296.0,1,-nbitq), 
to_sfixed(-508993997.0/4294967296.0,1,-nbitq), 
to_sfixed(-13946348.0/4294967296.0,1,-nbitq), 
to_sfixed(876476138.0/4294967296.0,1,-nbitq), 
to_sfixed(-118897022.0/4294967296.0,1,-nbitq), 
to_sfixed(1706099884.0/4294967296.0,1,-nbitq), 
to_sfixed(330398540.0/4294967296.0,1,-nbitq), 
to_sfixed(684796966.0/4294967296.0,1,-nbitq), 
to_sfixed(267496296.0/4294967296.0,1,-nbitq), 
to_sfixed(-60835004.0/4294967296.0,1,-nbitq), 
to_sfixed(-298424473.0/4294967296.0,1,-nbitq), 
to_sfixed(-133493728.0/4294967296.0,1,-nbitq), 
to_sfixed(-1273709659.0/4294967296.0,1,-nbitq), 
to_sfixed(-169685102.0/4294967296.0,1,-nbitq), 
to_sfixed(-3896808.0/4294967296.0,1,-nbitq), 
to_sfixed(597578587.0/4294967296.0,1,-nbitq), 
to_sfixed(-1355251969.0/4294967296.0,1,-nbitq), 
to_sfixed(1062372382.0/4294967296.0,1,-nbitq), 
to_sfixed(-1469919296.0/4294967296.0,1,-nbitq), 
to_sfixed(-782709102.0/4294967296.0,1,-nbitq), 
to_sfixed(-598754017.0/4294967296.0,1,-nbitq), 
to_sfixed(-2085192461.0/4294967296.0,1,-nbitq), 
to_sfixed(-355108005.0/4294967296.0,1,-nbitq), 
to_sfixed(899579129.0/4294967296.0,1,-nbitq), 
to_sfixed(-206199106.0/4294967296.0,1,-nbitq), 
to_sfixed(234698461.0/4294967296.0,1,-nbitq), 
to_sfixed(740536803.0/4294967296.0,1,-nbitq), 
to_sfixed(370109500.0/4294967296.0,1,-nbitq), 
to_sfixed(1543886788.0/4294967296.0,1,-nbitq), 
to_sfixed(758687418.0/4294967296.0,1,-nbitq), 
to_sfixed(-901356618.0/4294967296.0,1,-nbitq), 
to_sfixed(574843964.0/4294967296.0,1,-nbitq), 
to_sfixed(-186129081.0/4294967296.0,1,-nbitq), 
to_sfixed(557101880.0/4294967296.0,1,-nbitq), 
to_sfixed(-313311174.0/4294967296.0,1,-nbitq), 
to_sfixed(14872142.0/4294967296.0,1,-nbitq), 
to_sfixed(293706002.0/4294967296.0,1,-nbitq), 
to_sfixed(226930880.0/4294967296.0,1,-nbitq), 
to_sfixed(742076082.0/4294967296.0,1,-nbitq), 
to_sfixed(75064214.0/4294967296.0,1,-nbitq), 
to_sfixed(79269384.0/4294967296.0,1,-nbitq), 
to_sfixed(-30698619.0/4294967296.0,1,-nbitq), 
to_sfixed(-889405357.0/4294967296.0,1,-nbitq), 
to_sfixed(-460041467.0/4294967296.0,1,-nbitq), 
to_sfixed(-235620748.0/4294967296.0,1,-nbitq), 
to_sfixed(701738351.0/4294967296.0,1,-nbitq), 
to_sfixed(558998386.0/4294967296.0,1,-nbitq), 
to_sfixed(73595062.0/4294967296.0,1,-nbitq), 
to_sfixed(-1124961505.0/4294967296.0,1,-nbitq), 
to_sfixed(-289073519.0/4294967296.0,1,-nbitq), 
to_sfixed(82016661.0/4294967296.0,1,-nbitq), 
to_sfixed(426229143.0/4294967296.0,1,-nbitq), 
to_sfixed(516354567.0/4294967296.0,1,-nbitq), 
to_sfixed(-225527555.0/4294967296.0,1,-nbitq), 
to_sfixed(-234927095.0/4294967296.0,1,-nbitq), 
to_sfixed(105653600.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(66071299.0/4294967296.0,1,-nbitq), 
to_sfixed(-758295772.0/4294967296.0,1,-nbitq), 
to_sfixed(-433449827.0/4294967296.0,1,-nbitq), 
to_sfixed(1817409248.0/4294967296.0,1,-nbitq), 
to_sfixed(-1060549214.0/4294967296.0,1,-nbitq), 
to_sfixed(566918969.0/4294967296.0,1,-nbitq), 
to_sfixed(-59857026.0/4294967296.0,1,-nbitq), 
to_sfixed(266678869.0/4294967296.0,1,-nbitq), 
to_sfixed(-568440762.0/4294967296.0,1,-nbitq), 
to_sfixed(-165813123.0/4294967296.0,1,-nbitq), 
to_sfixed(-267111188.0/4294967296.0,1,-nbitq), 
to_sfixed(466934698.0/4294967296.0,1,-nbitq), 
to_sfixed(695504741.0/4294967296.0,1,-nbitq), 
to_sfixed(-603676368.0/4294967296.0,1,-nbitq), 
to_sfixed(153049497.0/4294967296.0,1,-nbitq), 
to_sfixed(260519329.0/4294967296.0,1,-nbitq), 
to_sfixed(160672111.0/4294967296.0,1,-nbitq), 
to_sfixed(42781605.0/4294967296.0,1,-nbitq), 
to_sfixed(-800883278.0/4294967296.0,1,-nbitq), 
to_sfixed(-642105898.0/4294967296.0,1,-nbitq), 
to_sfixed(372654127.0/4294967296.0,1,-nbitq), 
to_sfixed(-258951527.0/4294967296.0,1,-nbitq), 
to_sfixed(-1824427471.0/4294967296.0,1,-nbitq), 
to_sfixed(-572067762.0/4294967296.0,1,-nbitq), 
to_sfixed(-124166813.0/4294967296.0,1,-nbitq), 
to_sfixed(-378207378.0/4294967296.0,1,-nbitq), 
to_sfixed(-241920340.0/4294967296.0,1,-nbitq), 
to_sfixed(1221354215.0/4294967296.0,1,-nbitq), 
to_sfixed(-465033375.0/4294967296.0,1,-nbitq), 
to_sfixed(1597835645.0/4294967296.0,1,-nbitq), 
to_sfixed(1433123717.0/4294967296.0,1,-nbitq), 
to_sfixed(1244447778.0/4294967296.0,1,-nbitq), 
to_sfixed(-33351054.0/4294967296.0,1,-nbitq), 
to_sfixed(387708360.0/4294967296.0,1,-nbitq), 
to_sfixed(561445083.0/4294967296.0,1,-nbitq), 
to_sfixed(259444042.0/4294967296.0,1,-nbitq), 
to_sfixed(-999380301.0/4294967296.0,1,-nbitq), 
to_sfixed(-199936084.0/4294967296.0,1,-nbitq), 
to_sfixed(-220826654.0/4294967296.0,1,-nbitq), 
to_sfixed(620671246.0/4294967296.0,1,-nbitq), 
to_sfixed(-497824672.0/4294967296.0,1,-nbitq), 
to_sfixed(1091103448.0/4294967296.0,1,-nbitq), 
to_sfixed(-1220989098.0/4294967296.0,1,-nbitq), 
to_sfixed(-150810946.0/4294967296.0,1,-nbitq), 
to_sfixed(-845880447.0/4294967296.0,1,-nbitq), 
to_sfixed(-1848076623.0/4294967296.0,1,-nbitq), 
to_sfixed(146990456.0/4294967296.0,1,-nbitq), 
to_sfixed(398796431.0/4294967296.0,1,-nbitq), 
to_sfixed(46865652.0/4294967296.0,1,-nbitq), 
to_sfixed(-293467423.0/4294967296.0,1,-nbitq), 
to_sfixed(589471162.0/4294967296.0,1,-nbitq), 
to_sfixed(-726162989.0/4294967296.0,1,-nbitq), 
to_sfixed(1825200129.0/4294967296.0,1,-nbitq), 
to_sfixed(171326429.0/4294967296.0,1,-nbitq), 
to_sfixed(-1915241845.0/4294967296.0,1,-nbitq), 
to_sfixed(323034519.0/4294967296.0,1,-nbitq), 
to_sfixed(276394755.0/4294967296.0,1,-nbitq), 
to_sfixed(455323008.0/4294967296.0,1,-nbitq), 
to_sfixed(-209354711.0/4294967296.0,1,-nbitq), 
to_sfixed(359987452.0/4294967296.0,1,-nbitq), 
to_sfixed(16144589.0/4294967296.0,1,-nbitq), 
to_sfixed(-293256598.0/4294967296.0,1,-nbitq), 
to_sfixed(-3138533.0/4294967296.0,1,-nbitq), 
to_sfixed(206212804.0/4294967296.0,1,-nbitq), 
to_sfixed(585756263.0/4294967296.0,1,-nbitq), 
to_sfixed(97260236.0/4294967296.0,1,-nbitq), 
to_sfixed(316516483.0/4294967296.0,1,-nbitq), 
to_sfixed(-246169693.0/4294967296.0,1,-nbitq), 
to_sfixed(126450965.0/4294967296.0,1,-nbitq), 
to_sfixed(563062345.0/4294967296.0,1,-nbitq), 
to_sfixed(642378153.0/4294967296.0,1,-nbitq), 
to_sfixed(484995450.0/4294967296.0,1,-nbitq), 
to_sfixed(-709618746.0/4294967296.0,1,-nbitq), 
to_sfixed(305187208.0/4294967296.0,1,-nbitq), 
to_sfixed(-117737383.0/4294967296.0,1,-nbitq), 
to_sfixed(152012220.0/4294967296.0,1,-nbitq), 
to_sfixed(206737362.0/4294967296.0,1,-nbitq), 
to_sfixed(108291360.0/4294967296.0,1,-nbitq), 
to_sfixed(209780450.0/4294967296.0,1,-nbitq), 
to_sfixed(-192362971.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(73844690.0/4294967296.0,1,-nbitq), 
to_sfixed(-471037459.0/4294967296.0,1,-nbitq), 
to_sfixed(-182260745.0/4294967296.0,1,-nbitq), 
to_sfixed(1963506424.0/4294967296.0,1,-nbitq), 
to_sfixed(-831461582.0/4294967296.0,1,-nbitq), 
to_sfixed(-1391517694.0/4294967296.0,1,-nbitq), 
to_sfixed(-236545148.0/4294967296.0,1,-nbitq), 
to_sfixed(514368035.0/4294967296.0,1,-nbitq), 
to_sfixed(-569756121.0/4294967296.0,1,-nbitq), 
to_sfixed(-235361090.0/4294967296.0,1,-nbitq), 
to_sfixed(-333020408.0/4294967296.0,1,-nbitq), 
to_sfixed(651550158.0/4294967296.0,1,-nbitq), 
to_sfixed(49757177.0/4294967296.0,1,-nbitq), 
to_sfixed(-1731999165.0/4294967296.0,1,-nbitq), 
to_sfixed(170727340.0/4294967296.0,1,-nbitq), 
to_sfixed(785784865.0/4294967296.0,1,-nbitq), 
to_sfixed(-68260461.0/4294967296.0,1,-nbitq), 
to_sfixed(14012620.0/4294967296.0,1,-nbitq), 
to_sfixed(-1105182143.0/4294967296.0,1,-nbitq), 
to_sfixed(77924863.0/4294967296.0,1,-nbitq), 
to_sfixed(-185271671.0/4294967296.0,1,-nbitq), 
to_sfixed(-360479368.0/4294967296.0,1,-nbitq), 
to_sfixed(-1099443717.0/4294967296.0,1,-nbitq), 
to_sfixed(-1619636381.0/4294967296.0,1,-nbitq), 
to_sfixed(-213827987.0/4294967296.0,1,-nbitq), 
to_sfixed(-784349194.0/4294967296.0,1,-nbitq), 
to_sfixed(-250313867.0/4294967296.0,1,-nbitq), 
to_sfixed(572302538.0/4294967296.0,1,-nbitq), 
to_sfixed(-698296759.0/4294967296.0,1,-nbitq), 
to_sfixed(1543987846.0/4294967296.0,1,-nbitq), 
to_sfixed(1822148069.0/4294967296.0,1,-nbitq), 
to_sfixed(1147995015.0/4294967296.0,1,-nbitq), 
to_sfixed(24404897.0/4294967296.0,1,-nbitq), 
to_sfixed(755549751.0/4294967296.0,1,-nbitq), 
to_sfixed(-659531963.0/4294967296.0,1,-nbitq), 
to_sfixed(-276535338.0/4294967296.0,1,-nbitq), 
to_sfixed(-564957650.0/4294967296.0,1,-nbitq), 
to_sfixed(-388847614.0/4294967296.0,1,-nbitq), 
to_sfixed(435697911.0/4294967296.0,1,-nbitq), 
to_sfixed(-79785211.0/4294967296.0,1,-nbitq), 
to_sfixed(2188251.0/4294967296.0,1,-nbitq), 
to_sfixed(-408123918.0/4294967296.0,1,-nbitq), 
to_sfixed(-840121512.0/4294967296.0,1,-nbitq), 
to_sfixed(-87653713.0/4294967296.0,1,-nbitq), 
to_sfixed(-958651368.0/4294967296.0,1,-nbitq), 
to_sfixed(-698178343.0/4294967296.0,1,-nbitq), 
to_sfixed(-120604028.0/4294967296.0,1,-nbitq), 
to_sfixed(776462729.0/4294967296.0,1,-nbitq), 
to_sfixed(3469669.0/4294967296.0,1,-nbitq), 
to_sfixed(-776875998.0/4294967296.0,1,-nbitq), 
to_sfixed(817965726.0/4294967296.0,1,-nbitq), 
to_sfixed(-781086237.0/4294967296.0,1,-nbitq), 
to_sfixed(1456898390.0/4294967296.0,1,-nbitq), 
to_sfixed(-232813818.0/4294967296.0,1,-nbitq), 
to_sfixed(-511106472.0/4294967296.0,1,-nbitq), 
to_sfixed(433646515.0/4294967296.0,1,-nbitq), 
to_sfixed(432927730.0/4294967296.0,1,-nbitq), 
to_sfixed(853939438.0/4294967296.0,1,-nbitq), 
to_sfixed(-89032872.0/4294967296.0,1,-nbitq), 
to_sfixed(-92501334.0/4294967296.0,1,-nbitq), 
to_sfixed(257131687.0/4294967296.0,1,-nbitq), 
to_sfixed(-500788756.0/4294967296.0,1,-nbitq), 
to_sfixed(338346194.0/4294967296.0,1,-nbitq), 
to_sfixed(703605180.0/4294967296.0,1,-nbitq), 
to_sfixed(-24139465.0/4294967296.0,1,-nbitq), 
to_sfixed(-68902639.0/4294967296.0,1,-nbitq), 
to_sfixed(1069849386.0/4294967296.0,1,-nbitq), 
to_sfixed(9994150.0/4294967296.0,1,-nbitq), 
to_sfixed(222849833.0/4294967296.0,1,-nbitq), 
to_sfixed(739277477.0/4294967296.0,1,-nbitq), 
to_sfixed(522003168.0/4294967296.0,1,-nbitq), 
to_sfixed(322840488.0/4294967296.0,1,-nbitq), 
to_sfixed(-55254315.0/4294967296.0,1,-nbitq), 
to_sfixed(331593337.0/4294967296.0,1,-nbitq), 
to_sfixed(3479917.0/4294967296.0,1,-nbitq), 
to_sfixed(497619203.0/4294967296.0,1,-nbitq), 
to_sfixed(131013295.0/4294967296.0,1,-nbitq), 
to_sfixed(-115509876.0/4294967296.0,1,-nbitq), 
to_sfixed(-49029752.0/4294967296.0,1,-nbitq), 
to_sfixed(-207537191.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-371965395.0/4294967296.0,1,-nbitq), 
to_sfixed(-698680414.0/4294967296.0,1,-nbitq), 
to_sfixed(188536419.0/4294967296.0,1,-nbitq), 
to_sfixed(299512329.0/4294967296.0,1,-nbitq), 
to_sfixed(-657150587.0/4294967296.0,1,-nbitq), 
to_sfixed(-1519991655.0/4294967296.0,1,-nbitq), 
to_sfixed(366950082.0/4294967296.0,1,-nbitq), 
to_sfixed(659617142.0/4294967296.0,1,-nbitq), 
to_sfixed(-661905990.0/4294967296.0,1,-nbitq), 
to_sfixed(-331552328.0/4294967296.0,1,-nbitq), 
to_sfixed(175013119.0/4294967296.0,1,-nbitq), 
to_sfixed(-80469705.0/4294967296.0,1,-nbitq), 
to_sfixed(-279041675.0/4294967296.0,1,-nbitq), 
to_sfixed(-345945067.0/4294967296.0,1,-nbitq), 
to_sfixed(-79260882.0/4294967296.0,1,-nbitq), 
to_sfixed(214808303.0/4294967296.0,1,-nbitq), 
to_sfixed(-83547597.0/4294967296.0,1,-nbitq), 
to_sfixed(294265186.0/4294967296.0,1,-nbitq), 
to_sfixed(-150091497.0/4294967296.0,1,-nbitq), 
to_sfixed(131970420.0/4294967296.0,1,-nbitq), 
to_sfixed(18523529.0/4294967296.0,1,-nbitq), 
to_sfixed(-309196842.0/4294967296.0,1,-nbitq), 
to_sfixed(-743157368.0/4294967296.0,1,-nbitq), 
to_sfixed(-546032411.0/4294967296.0,1,-nbitq), 
to_sfixed(-82272322.0/4294967296.0,1,-nbitq), 
to_sfixed(-1179055495.0/4294967296.0,1,-nbitq), 
to_sfixed(53362728.0/4294967296.0,1,-nbitq), 
to_sfixed(239609773.0/4294967296.0,1,-nbitq), 
to_sfixed(-13149920.0/4294967296.0,1,-nbitq), 
to_sfixed(705946672.0/4294967296.0,1,-nbitq), 
to_sfixed(-208998108.0/4294967296.0,1,-nbitq), 
to_sfixed(670114536.0/4294967296.0,1,-nbitq), 
to_sfixed(279420344.0/4294967296.0,1,-nbitq), 
to_sfixed(965325466.0/4294967296.0,1,-nbitq), 
to_sfixed(-356201157.0/4294967296.0,1,-nbitq), 
to_sfixed(151928414.0/4294967296.0,1,-nbitq), 
to_sfixed(-11205692.0/4294967296.0,1,-nbitq), 
to_sfixed(125045003.0/4294967296.0,1,-nbitq), 
to_sfixed(-263758576.0/4294967296.0,1,-nbitq), 
to_sfixed(32062758.0/4294967296.0,1,-nbitq), 
to_sfixed(-621018435.0/4294967296.0,1,-nbitq), 
to_sfixed(-126726855.0/4294967296.0,1,-nbitq), 
to_sfixed(-843573911.0/4294967296.0,1,-nbitq), 
to_sfixed(-445026974.0/4294967296.0,1,-nbitq), 
to_sfixed(-437273488.0/4294967296.0,1,-nbitq), 
to_sfixed(-415315419.0/4294967296.0,1,-nbitq), 
to_sfixed(305667668.0/4294967296.0,1,-nbitq), 
to_sfixed(816569795.0/4294967296.0,1,-nbitq), 
to_sfixed(-312106320.0/4294967296.0,1,-nbitq), 
to_sfixed(-781391480.0/4294967296.0,1,-nbitq), 
to_sfixed(735941668.0/4294967296.0,1,-nbitq), 
to_sfixed(-157821393.0/4294967296.0,1,-nbitq), 
to_sfixed(1006262387.0/4294967296.0,1,-nbitq), 
to_sfixed(135146320.0/4294967296.0,1,-nbitq), 
to_sfixed(-1266201824.0/4294967296.0,1,-nbitq), 
to_sfixed(24901608.0/4294967296.0,1,-nbitq), 
to_sfixed(531202993.0/4294967296.0,1,-nbitq), 
to_sfixed(667802514.0/4294967296.0,1,-nbitq), 
to_sfixed(16472487.0/4294967296.0,1,-nbitq), 
to_sfixed(301795457.0/4294967296.0,1,-nbitq), 
to_sfixed(221466371.0/4294967296.0,1,-nbitq), 
to_sfixed(-408205139.0/4294967296.0,1,-nbitq), 
to_sfixed(161956980.0/4294967296.0,1,-nbitq), 
to_sfixed(453807804.0/4294967296.0,1,-nbitq), 
to_sfixed(116229513.0/4294967296.0,1,-nbitq), 
to_sfixed(-23308511.0/4294967296.0,1,-nbitq), 
to_sfixed(655674516.0/4294967296.0,1,-nbitq), 
to_sfixed(-856795396.0/4294967296.0,1,-nbitq), 
to_sfixed(66469048.0/4294967296.0,1,-nbitq), 
to_sfixed(621958393.0/4294967296.0,1,-nbitq), 
to_sfixed(-47863836.0/4294967296.0,1,-nbitq), 
to_sfixed(412565572.0/4294967296.0,1,-nbitq), 
to_sfixed(297868426.0/4294967296.0,1,-nbitq), 
to_sfixed(161048623.0/4294967296.0,1,-nbitq), 
to_sfixed(432784307.0/4294967296.0,1,-nbitq), 
to_sfixed(-77939218.0/4294967296.0,1,-nbitq), 
to_sfixed(508422578.0/4294967296.0,1,-nbitq), 
to_sfixed(43210771.0/4294967296.0,1,-nbitq), 
to_sfixed(866612051.0/4294967296.0,1,-nbitq), 
to_sfixed(136040651.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-369334348.0/4294967296.0,1,-nbitq), 
to_sfixed(-58713691.0/4294967296.0,1,-nbitq), 
to_sfixed(-224922137.0/4294967296.0,1,-nbitq), 
to_sfixed(-323725968.0/4294967296.0,1,-nbitq), 
to_sfixed(-836484232.0/4294967296.0,1,-nbitq), 
to_sfixed(-832083360.0/4294967296.0,1,-nbitq), 
to_sfixed(167800509.0/4294967296.0,1,-nbitq), 
to_sfixed(1061226363.0/4294967296.0,1,-nbitq), 
to_sfixed(-1021778508.0/4294967296.0,1,-nbitq), 
to_sfixed(4672203.0/4294967296.0,1,-nbitq), 
to_sfixed(214691575.0/4294967296.0,1,-nbitq), 
to_sfixed(103744310.0/4294967296.0,1,-nbitq), 
to_sfixed(-592746006.0/4294967296.0,1,-nbitq), 
to_sfixed(-939410347.0/4294967296.0,1,-nbitq), 
to_sfixed(-336663662.0/4294967296.0,1,-nbitq), 
to_sfixed(103665807.0/4294967296.0,1,-nbitq), 
to_sfixed(-122870303.0/4294967296.0,1,-nbitq), 
to_sfixed(332726664.0/4294967296.0,1,-nbitq), 
to_sfixed(-603436859.0/4294967296.0,1,-nbitq), 
to_sfixed(-443954523.0/4294967296.0,1,-nbitq), 
to_sfixed(-195136481.0/4294967296.0,1,-nbitq), 
to_sfixed(-424957719.0/4294967296.0,1,-nbitq), 
to_sfixed(-707605830.0/4294967296.0,1,-nbitq), 
to_sfixed(-537946283.0/4294967296.0,1,-nbitq), 
to_sfixed(-90021150.0/4294967296.0,1,-nbitq), 
to_sfixed(-1151814829.0/4294967296.0,1,-nbitq), 
to_sfixed(530272045.0/4294967296.0,1,-nbitq), 
to_sfixed(-312849513.0/4294967296.0,1,-nbitq), 
to_sfixed(-425362995.0/4294967296.0,1,-nbitq), 
to_sfixed(1071771537.0/4294967296.0,1,-nbitq), 
to_sfixed(-138825494.0/4294967296.0,1,-nbitq), 
to_sfixed(77179905.0/4294967296.0,1,-nbitq), 
to_sfixed(-516636982.0/4294967296.0,1,-nbitq), 
to_sfixed(290582645.0/4294967296.0,1,-nbitq), 
to_sfixed(-500541301.0/4294967296.0,1,-nbitq), 
to_sfixed(-27468103.0/4294967296.0,1,-nbitq), 
to_sfixed(-123141855.0/4294967296.0,1,-nbitq), 
to_sfixed(1069064129.0/4294967296.0,1,-nbitq), 
to_sfixed(-230691562.0/4294967296.0,1,-nbitq), 
to_sfixed(175782470.0/4294967296.0,1,-nbitq), 
to_sfixed(-128282904.0/4294967296.0,1,-nbitq), 
to_sfixed(-118403893.0/4294967296.0,1,-nbitq), 
to_sfixed(-890168188.0/4294967296.0,1,-nbitq), 
to_sfixed(-1040987071.0/4294967296.0,1,-nbitq), 
to_sfixed(-456976649.0/4294967296.0,1,-nbitq), 
to_sfixed(-795248472.0/4294967296.0,1,-nbitq), 
to_sfixed(-200031715.0/4294967296.0,1,-nbitq), 
to_sfixed(401111333.0/4294967296.0,1,-nbitq), 
to_sfixed(314044925.0/4294967296.0,1,-nbitq), 
to_sfixed(-86930642.0/4294967296.0,1,-nbitq), 
to_sfixed(516182553.0/4294967296.0,1,-nbitq), 
to_sfixed(98479354.0/4294967296.0,1,-nbitq), 
to_sfixed(892614130.0/4294967296.0,1,-nbitq), 
to_sfixed(-1042962819.0/4294967296.0,1,-nbitq), 
to_sfixed(-1247215911.0/4294967296.0,1,-nbitq), 
to_sfixed(-67872182.0/4294967296.0,1,-nbitq), 
to_sfixed(667079119.0/4294967296.0,1,-nbitq), 
to_sfixed(397918784.0/4294967296.0,1,-nbitq), 
to_sfixed(-376929124.0/4294967296.0,1,-nbitq), 
to_sfixed(-344873045.0/4294967296.0,1,-nbitq), 
to_sfixed(157563368.0/4294967296.0,1,-nbitq), 
to_sfixed(-272075217.0/4294967296.0,1,-nbitq), 
to_sfixed(649357427.0/4294967296.0,1,-nbitq), 
to_sfixed(446846633.0/4294967296.0,1,-nbitq), 
to_sfixed(-163531817.0/4294967296.0,1,-nbitq), 
to_sfixed(42426478.0/4294967296.0,1,-nbitq), 
to_sfixed(510022211.0/4294967296.0,1,-nbitq), 
to_sfixed(-278839855.0/4294967296.0,1,-nbitq), 
to_sfixed(38162948.0/4294967296.0,1,-nbitq), 
to_sfixed(649100026.0/4294967296.0,1,-nbitq), 
to_sfixed(-292155586.0/4294967296.0,1,-nbitq), 
to_sfixed(-217194215.0/4294967296.0,1,-nbitq), 
to_sfixed(323364791.0/4294967296.0,1,-nbitq), 
to_sfixed(382192516.0/4294967296.0,1,-nbitq), 
to_sfixed(419279502.0/4294967296.0,1,-nbitq), 
to_sfixed(63816092.0/4294967296.0,1,-nbitq), 
to_sfixed(-106616111.0/4294967296.0,1,-nbitq), 
to_sfixed(-225179438.0/4294967296.0,1,-nbitq), 
to_sfixed(489776609.0/4294967296.0,1,-nbitq), 
to_sfixed(133031619.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(76365602.0/4294967296.0,1,-nbitq), 
to_sfixed(99812452.0/4294967296.0,1,-nbitq), 
to_sfixed(77168510.0/4294967296.0,1,-nbitq), 
to_sfixed(-619051282.0/4294967296.0,1,-nbitq), 
to_sfixed(-332491810.0/4294967296.0,1,-nbitq), 
to_sfixed(-718102912.0/4294967296.0,1,-nbitq), 
to_sfixed(-71458962.0/4294967296.0,1,-nbitq), 
to_sfixed(636914714.0/4294967296.0,1,-nbitq), 
to_sfixed(-50346196.0/4294967296.0,1,-nbitq), 
to_sfixed(40630278.0/4294967296.0,1,-nbitq), 
to_sfixed(-176835487.0/4294967296.0,1,-nbitq), 
to_sfixed(-287834741.0/4294967296.0,1,-nbitq), 
to_sfixed(-452217620.0/4294967296.0,1,-nbitq), 
to_sfixed(-86296445.0/4294967296.0,1,-nbitq), 
to_sfixed(164559785.0/4294967296.0,1,-nbitq), 
to_sfixed(400983436.0/4294967296.0,1,-nbitq), 
to_sfixed(-374761282.0/4294967296.0,1,-nbitq), 
to_sfixed(-94935166.0/4294967296.0,1,-nbitq), 
to_sfixed(-390813970.0/4294967296.0,1,-nbitq), 
to_sfixed(-331769440.0/4294967296.0,1,-nbitq), 
to_sfixed(171411216.0/4294967296.0,1,-nbitq), 
to_sfixed(-367222372.0/4294967296.0,1,-nbitq), 
to_sfixed(-215903579.0/4294967296.0,1,-nbitq), 
to_sfixed(16215591.0/4294967296.0,1,-nbitq), 
to_sfixed(-161845183.0/4294967296.0,1,-nbitq), 
to_sfixed(-1006289008.0/4294967296.0,1,-nbitq), 
to_sfixed(631978951.0/4294967296.0,1,-nbitq), 
to_sfixed(-187173640.0/4294967296.0,1,-nbitq), 
to_sfixed(-175057487.0/4294967296.0,1,-nbitq), 
to_sfixed(743636401.0/4294967296.0,1,-nbitq), 
to_sfixed(-241630819.0/4294967296.0,1,-nbitq), 
to_sfixed(43189169.0/4294967296.0,1,-nbitq), 
to_sfixed(-319412949.0/4294967296.0,1,-nbitq), 
to_sfixed(255690424.0/4294967296.0,1,-nbitq), 
to_sfixed(-797130847.0/4294967296.0,1,-nbitq), 
to_sfixed(-121686993.0/4294967296.0,1,-nbitq), 
to_sfixed(-261541234.0/4294967296.0,1,-nbitq), 
to_sfixed(140617056.0/4294967296.0,1,-nbitq), 
to_sfixed(-235258101.0/4294967296.0,1,-nbitq), 
to_sfixed(-118359084.0/4294967296.0,1,-nbitq), 
to_sfixed(292793124.0/4294967296.0,1,-nbitq), 
to_sfixed(-302953192.0/4294967296.0,1,-nbitq), 
to_sfixed(-432983235.0/4294967296.0,1,-nbitq), 
to_sfixed(-1040395478.0/4294967296.0,1,-nbitq), 
to_sfixed(-276617609.0/4294967296.0,1,-nbitq), 
to_sfixed(-673931636.0/4294967296.0,1,-nbitq), 
to_sfixed(-44569287.0/4294967296.0,1,-nbitq), 
to_sfixed(248198258.0/4294967296.0,1,-nbitq), 
to_sfixed(148453562.0/4294967296.0,1,-nbitq), 
to_sfixed(101098393.0/4294967296.0,1,-nbitq), 
to_sfixed(198428443.0/4294967296.0,1,-nbitq), 
to_sfixed(-49869301.0/4294967296.0,1,-nbitq), 
to_sfixed(890981881.0/4294967296.0,1,-nbitq), 
to_sfixed(-209877611.0/4294967296.0,1,-nbitq), 
to_sfixed(-305507954.0/4294967296.0,1,-nbitq), 
to_sfixed(-240223889.0/4294967296.0,1,-nbitq), 
to_sfixed(409898630.0/4294967296.0,1,-nbitq), 
to_sfixed(94489647.0/4294967296.0,1,-nbitq), 
to_sfixed(207961900.0/4294967296.0,1,-nbitq), 
to_sfixed(-271172273.0/4294967296.0,1,-nbitq), 
to_sfixed(7850155.0/4294967296.0,1,-nbitq), 
to_sfixed(23069547.0/4294967296.0,1,-nbitq), 
to_sfixed(396258487.0/4294967296.0,1,-nbitq), 
to_sfixed(483585126.0/4294967296.0,1,-nbitq), 
to_sfixed(78925472.0/4294967296.0,1,-nbitq), 
to_sfixed(-244421707.0/4294967296.0,1,-nbitq), 
to_sfixed(848590213.0/4294967296.0,1,-nbitq), 
to_sfixed(-346366837.0/4294967296.0,1,-nbitq), 
to_sfixed(-31771755.0/4294967296.0,1,-nbitq), 
to_sfixed(605419828.0/4294967296.0,1,-nbitq), 
to_sfixed(-194915743.0/4294967296.0,1,-nbitq), 
to_sfixed(254559163.0/4294967296.0,1,-nbitq), 
to_sfixed(728002979.0/4294967296.0,1,-nbitq), 
to_sfixed(-111593786.0/4294967296.0,1,-nbitq), 
to_sfixed(-146413796.0/4294967296.0,1,-nbitq), 
to_sfixed(152763567.0/4294967296.0,1,-nbitq), 
to_sfixed(-792683671.0/4294967296.0,1,-nbitq), 
to_sfixed(-139726182.0/4294967296.0,1,-nbitq), 
to_sfixed(-52080143.0/4294967296.0,1,-nbitq), 
to_sfixed(-53450857.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(300403075.0/4294967296.0,1,-nbitq), 
to_sfixed(-223472445.0/4294967296.0,1,-nbitq), 
to_sfixed(797163826.0/4294967296.0,1,-nbitq), 
to_sfixed(-688338622.0/4294967296.0,1,-nbitq), 
to_sfixed(-184495160.0/4294967296.0,1,-nbitq), 
to_sfixed(-836551768.0/4294967296.0,1,-nbitq), 
to_sfixed(-121112814.0/4294967296.0,1,-nbitq), 
to_sfixed(29370800.0/4294967296.0,1,-nbitq), 
to_sfixed(-515482714.0/4294967296.0,1,-nbitq), 
to_sfixed(434578721.0/4294967296.0,1,-nbitq), 
to_sfixed(465276625.0/4294967296.0,1,-nbitq), 
to_sfixed(-128084236.0/4294967296.0,1,-nbitq), 
to_sfixed(169296677.0/4294967296.0,1,-nbitq), 
to_sfixed(161075107.0/4294967296.0,1,-nbitq), 
to_sfixed(248720759.0/4294967296.0,1,-nbitq), 
to_sfixed(440779166.0/4294967296.0,1,-nbitq), 
to_sfixed(-260078368.0/4294967296.0,1,-nbitq), 
to_sfixed(-17699234.0/4294967296.0,1,-nbitq), 
to_sfixed(559371285.0/4294967296.0,1,-nbitq), 
to_sfixed(-72889287.0/4294967296.0,1,-nbitq), 
to_sfixed(-178280035.0/4294967296.0,1,-nbitq), 
to_sfixed(-58501023.0/4294967296.0,1,-nbitq), 
to_sfixed(-111933170.0/4294967296.0,1,-nbitq), 
to_sfixed(341826489.0/4294967296.0,1,-nbitq), 
to_sfixed(136406793.0/4294967296.0,1,-nbitq), 
to_sfixed(-868952275.0/4294967296.0,1,-nbitq), 
to_sfixed(66944442.0/4294967296.0,1,-nbitq), 
to_sfixed(-260829695.0/4294967296.0,1,-nbitq), 
to_sfixed(399741888.0/4294967296.0,1,-nbitq), 
to_sfixed(409242494.0/4294967296.0,1,-nbitq), 
to_sfixed(13242821.0/4294967296.0,1,-nbitq), 
to_sfixed(95481071.0/4294967296.0,1,-nbitq), 
to_sfixed(102715362.0/4294967296.0,1,-nbitq), 
to_sfixed(-329390018.0/4294967296.0,1,-nbitq), 
to_sfixed(-270754306.0/4294967296.0,1,-nbitq), 
to_sfixed(68402525.0/4294967296.0,1,-nbitq), 
to_sfixed(36781573.0/4294967296.0,1,-nbitq), 
to_sfixed(-24767129.0/4294967296.0,1,-nbitq), 
to_sfixed(-93383325.0/4294967296.0,1,-nbitq), 
to_sfixed(218481761.0/4294967296.0,1,-nbitq), 
to_sfixed(315058086.0/4294967296.0,1,-nbitq), 
to_sfixed(-55110808.0/4294967296.0,1,-nbitq), 
to_sfixed(-439589673.0/4294967296.0,1,-nbitq), 
to_sfixed(-804932066.0/4294967296.0,1,-nbitq), 
to_sfixed(348431386.0/4294967296.0,1,-nbitq), 
to_sfixed(-812311798.0/4294967296.0,1,-nbitq), 
to_sfixed(144546632.0/4294967296.0,1,-nbitq), 
to_sfixed(-399440002.0/4294967296.0,1,-nbitq), 
to_sfixed(-264455178.0/4294967296.0,1,-nbitq), 
to_sfixed(171030083.0/4294967296.0,1,-nbitq), 
to_sfixed(231434606.0/4294967296.0,1,-nbitq), 
to_sfixed(-70378143.0/4294967296.0,1,-nbitq), 
to_sfixed(50363516.0/4294967296.0,1,-nbitq), 
to_sfixed(-355139365.0/4294967296.0,1,-nbitq), 
to_sfixed(-367655207.0/4294967296.0,1,-nbitq), 
to_sfixed(128500800.0/4294967296.0,1,-nbitq), 
to_sfixed(464491136.0/4294967296.0,1,-nbitq), 
to_sfixed(146986578.0/4294967296.0,1,-nbitq), 
to_sfixed(-319809044.0/4294967296.0,1,-nbitq), 
to_sfixed(177258418.0/4294967296.0,1,-nbitq), 
to_sfixed(175370924.0/4294967296.0,1,-nbitq), 
to_sfixed(-242409797.0/4294967296.0,1,-nbitq), 
to_sfixed(70498934.0/4294967296.0,1,-nbitq), 
to_sfixed(48987245.0/4294967296.0,1,-nbitq), 
to_sfixed(352592348.0/4294967296.0,1,-nbitq), 
to_sfixed(-182511471.0/4294967296.0,1,-nbitq), 
to_sfixed(274025476.0/4294967296.0,1,-nbitq), 
to_sfixed(-76191693.0/4294967296.0,1,-nbitq), 
to_sfixed(165257896.0/4294967296.0,1,-nbitq), 
to_sfixed(561985978.0/4294967296.0,1,-nbitq), 
to_sfixed(-53963561.0/4294967296.0,1,-nbitq), 
to_sfixed(221687847.0/4294967296.0,1,-nbitq), 
to_sfixed(365565825.0/4294967296.0,1,-nbitq), 
to_sfixed(112365961.0/4294967296.0,1,-nbitq), 
to_sfixed(384911717.0/4294967296.0,1,-nbitq), 
to_sfixed(99052577.0/4294967296.0,1,-nbitq), 
to_sfixed(55593104.0/4294967296.0,1,-nbitq), 
to_sfixed(229995261.0/4294967296.0,1,-nbitq), 
to_sfixed(142696545.0/4294967296.0,1,-nbitq), 
to_sfixed(-114953644.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(169693450.0/4294967296.0,1,-nbitq), 
to_sfixed(165587057.0/4294967296.0,1,-nbitq), 
to_sfixed(-77171112.0/4294967296.0,1,-nbitq), 
to_sfixed(-648162857.0/4294967296.0,1,-nbitq), 
to_sfixed(-164173135.0/4294967296.0,1,-nbitq), 
to_sfixed(-749903183.0/4294967296.0,1,-nbitq), 
to_sfixed(-166594778.0/4294967296.0,1,-nbitq), 
to_sfixed(-107595745.0/4294967296.0,1,-nbitq), 
to_sfixed(33655738.0/4294967296.0,1,-nbitq), 
to_sfixed(285234671.0/4294967296.0,1,-nbitq), 
to_sfixed(351878197.0/4294967296.0,1,-nbitq), 
to_sfixed(-216641004.0/4294967296.0,1,-nbitq), 
to_sfixed(-238992595.0/4294967296.0,1,-nbitq), 
to_sfixed(266974534.0/4294967296.0,1,-nbitq), 
to_sfixed(-49687483.0/4294967296.0,1,-nbitq), 
to_sfixed(179467676.0/4294967296.0,1,-nbitq), 
to_sfixed(256303575.0/4294967296.0,1,-nbitq), 
to_sfixed(-134129282.0/4294967296.0,1,-nbitq), 
to_sfixed(202377626.0/4294967296.0,1,-nbitq), 
to_sfixed(-411645406.0/4294967296.0,1,-nbitq), 
to_sfixed(-363278193.0/4294967296.0,1,-nbitq), 
to_sfixed(-76301639.0/4294967296.0,1,-nbitq), 
to_sfixed(-68313802.0/4294967296.0,1,-nbitq), 
to_sfixed(133943742.0/4294967296.0,1,-nbitq), 
to_sfixed(33145204.0/4294967296.0,1,-nbitq), 
to_sfixed(-349849332.0/4294967296.0,1,-nbitq), 
to_sfixed(522217545.0/4294967296.0,1,-nbitq), 
to_sfixed(-252920361.0/4294967296.0,1,-nbitq), 
to_sfixed(29937233.0/4294967296.0,1,-nbitq), 
to_sfixed(46294217.0/4294967296.0,1,-nbitq), 
to_sfixed(91607473.0/4294967296.0,1,-nbitq), 
to_sfixed(-336151882.0/4294967296.0,1,-nbitq), 
to_sfixed(435608140.0/4294967296.0,1,-nbitq), 
to_sfixed(-221929374.0/4294967296.0,1,-nbitq), 
to_sfixed(223971771.0/4294967296.0,1,-nbitq), 
to_sfixed(-566636164.0/4294967296.0,1,-nbitq), 
to_sfixed(-254326307.0/4294967296.0,1,-nbitq), 
to_sfixed(183331966.0/4294967296.0,1,-nbitq), 
to_sfixed(158139079.0/4294967296.0,1,-nbitq), 
to_sfixed(-85441516.0/4294967296.0,1,-nbitq), 
to_sfixed(65756125.0/4294967296.0,1,-nbitq), 
to_sfixed(90149603.0/4294967296.0,1,-nbitq), 
to_sfixed(245597846.0/4294967296.0,1,-nbitq), 
to_sfixed(-12477860.0/4294967296.0,1,-nbitq), 
to_sfixed(327653446.0/4294967296.0,1,-nbitq), 
to_sfixed(-62201590.0/4294967296.0,1,-nbitq), 
to_sfixed(-271884473.0/4294967296.0,1,-nbitq), 
to_sfixed(125831611.0/4294967296.0,1,-nbitq), 
to_sfixed(208559440.0/4294967296.0,1,-nbitq), 
to_sfixed(-326912277.0/4294967296.0,1,-nbitq), 
to_sfixed(-177024544.0/4294967296.0,1,-nbitq), 
to_sfixed(-19979649.0/4294967296.0,1,-nbitq), 
to_sfixed(-39923790.0/4294967296.0,1,-nbitq), 
to_sfixed(218909029.0/4294967296.0,1,-nbitq), 
to_sfixed(70701438.0/4294967296.0,1,-nbitq), 
to_sfixed(22369813.0/4294967296.0,1,-nbitq), 
to_sfixed(71498587.0/4294967296.0,1,-nbitq), 
to_sfixed(-109416844.0/4294967296.0,1,-nbitq), 
to_sfixed(309098641.0/4294967296.0,1,-nbitq), 
to_sfixed(143507241.0/4294967296.0,1,-nbitq), 
to_sfixed(391749274.0/4294967296.0,1,-nbitq), 
to_sfixed(-335094126.0/4294967296.0,1,-nbitq), 
to_sfixed(21113056.0/4294967296.0,1,-nbitq), 
to_sfixed(-158705250.0/4294967296.0,1,-nbitq), 
to_sfixed(270655198.0/4294967296.0,1,-nbitq), 
to_sfixed(-167217765.0/4294967296.0,1,-nbitq), 
to_sfixed(403032861.0/4294967296.0,1,-nbitq), 
to_sfixed(-338382981.0/4294967296.0,1,-nbitq), 
to_sfixed(-44747708.0/4294967296.0,1,-nbitq), 
to_sfixed(112417007.0/4294967296.0,1,-nbitq), 
to_sfixed(-42772497.0/4294967296.0,1,-nbitq), 
to_sfixed(-337981170.0/4294967296.0,1,-nbitq), 
to_sfixed(-204661693.0/4294967296.0,1,-nbitq), 
to_sfixed(286408101.0/4294967296.0,1,-nbitq), 
to_sfixed(-62330818.0/4294967296.0,1,-nbitq), 
to_sfixed(-383164675.0/4294967296.0,1,-nbitq), 
to_sfixed(210980684.0/4294967296.0,1,-nbitq), 
to_sfixed(-395022774.0/4294967296.0,1,-nbitq), 
to_sfixed(7262633.0/4294967296.0,1,-nbitq), 
to_sfixed(-338715252.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(54860893.0/4294967296.0,1,-nbitq), 
to_sfixed(-498974043.0/4294967296.0,1,-nbitq), 
to_sfixed(229192609.0/4294967296.0,1,-nbitq), 
to_sfixed(68352785.0/4294967296.0,1,-nbitq), 
to_sfixed(425734187.0/4294967296.0,1,-nbitq), 
to_sfixed(-144052590.0/4294967296.0,1,-nbitq), 
to_sfixed(290609275.0/4294967296.0,1,-nbitq), 
to_sfixed(-194904836.0/4294967296.0,1,-nbitq), 
to_sfixed(-8074800.0/4294967296.0,1,-nbitq), 
to_sfixed(449714453.0/4294967296.0,1,-nbitq), 
to_sfixed(323479367.0/4294967296.0,1,-nbitq), 
to_sfixed(392505344.0/4294967296.0,1,-nbitq), 
to_sfixed(-240273164.0/4294967296.0,1,-nbitq), 
to_sfixed(269059250.0/4294967296.0,1,-nbitq), 
to_sfixed(-310411599.0/4294967296.0,1,-nbitq), 
to_sfixed(45805059.0/4294967296.0,1,-nbitq), 
to_sfixed(-278049158.0/4294967296.0,1,-nbitq), 
to_sfixed(-111246068.0/4294967296.0,1,-nbitq), 
to_sfixed(502656275.0/4294967296.0,1,-nbitq), 
to_sfixed(-217754572.0/4294967296.0,1,-nbitq), 
to_sfixed(-193218757.0/4294967296.0,1,-nbitq), 
to_sfixed(-28580447.0/4294967296.0,1,-nbitq), 
to_sfixed(-82461104.0/4294967296.0,1,-nbitq), 
to_sfixed(-277157291.0/4294967296.0,1,-nbitq), 
to_sfixed(-255543857.0/4294967296.0,1,-nbitq), 
to_sfixed(113076662.0/4294967296.0,1,-nbitq), 
to_sfixed(-313733563.0/4294967296.0,1,-nbitq), 
to_sfixed(-287643118.0/4294967296.0,1,-nbitq), 
to_sfixed(-7895349.0/4294967296.0,1,-nbitq), 
to_sfixed(267784731.0/4294967296.0,1,-nbitq), 
to_sfixed(-415219218.0/4294967296.0,1,-nbitq), 
to_sfixed(-273482319.0/4294967296.0,1,-nbitq), 
to_sfixed(-236000277.0/4294967296.0,1,-nbitq), 
to_sfixed(90529279.0/4294967296.0,1,-nbitq), 
to_sfixed(154844529.0/4294967296.0,1,-nbitq), 
to_sfixed(-397915539.0/4294967296.0,1,-nbitq), 
to_sfixed(311333790.0/4294967296.0,1,-nbitq), 
to_sfixed(2157120.0/4294967296.0,1,-nbitq), 
to_sfixed(-2531121.0/4294967296.0,1,-nbitq), 
to_sfixed(120260317.0/4294967296.0,1,-nbitq), 
to_sfixed(-61633268.0/4294967296.0,1,-nbitq), 
to_sfixed(301373230.0/4294967296.0,1,-nbitq), 
to_sfixed(169312751.0/4294967296.0,1,-nbitq), 
to_sfixed(-264261853.0/4294967296.0,1,-nbitq), 
to_sfixed(306521726.0/4294967296.0,1,-nbitq), 
to_sfixed(249927216.0/4294967296.0,1,-nbitq), 
to_sfixed(171559612.0/4294967296.0,1,-nbitq), 
to_sfixed(-291628064.0/4294967296.0,1,-nbitq), 
to_sfixed(-88781589.0/4294967296.0,1,-nbitq), 
to_sfixed(-181344060.0/4294967296.0,1,-nbitq), 
to_sfixed(290746299.0/4294967296.0,1,-nbitq), 
to_sfixed(-10284190.0/4294967296.0,1,-nbitq), 
to_sfixed(27854538.0/4294967296.0,1,-nbitq), 
to_sfixed(440207954.0/4294967296.0,1,-nbitq), 
to_sfixed(427295471.0/4294967296.0,1,-nbitq), 
to_sfixed(-49562917.0/4294967296.0,1,-nbitq), 
to_sfixed(277684811.0/4294967296.0,1,-nbitq), 
to_sfixed(-378295212.0/4294967296.0,1,-nbitq), 
to_sfixed(298188342.0/4294967296.0,1,-nbitq), 
to_sfixed(426671919.0/4294967296.0,1,-nbitq), 
to_sfixed(222032515.0/4294967296.0,1,-nbitq), 
to_sfixed(-110368917.0/4294967296.0,1,-nbitq), 
to_sfixed(277141420.0/4294967296.0,1,-nbitq), 
to_sfixed(32944963.0/4294967296.0,1,-nbitq), 
to_sfixed(104771177.0/4294967296.0,1,-nbitq), 
to_sfixed(243122520.0/4294967296.0,1,-nbitq), 
to_sfixed(243137143.0/4294967296.0,1,-nbitq), 
to_sfixed(-190347379.0/4294967296.0,1,-nbitq), 
to_sfixed(300304285.0/4294967296.0,1,-nbitq), 
to_sfixed(-230985089.0/4294967296.0,1,-nbitq), 
to_sfixed(-38912164.0/4294967296.0,1,-nbitq), 
to_sfixed(-200401855.0/4294967296.0,1,-nbitq), 
to_sfixed(-220993465.0/4294967296.0,1,-nbitq), 
to_sfixed(-328223848.0/4294967296.0,1,-nbitq), 
to_sfixed(147254841.0/4294967296.0,1,-nbitq), 
to_sfixed(-409227756.0/4294967296.0,1,-nbitq), 
to_sfixed(-221914577.0/4294967296.0,1,-nbitq), 
to_sfixed(-230836506.0/4294967296.0,1,-nbitq), 
to_sfixed(-503723373.0/4294967296.0,1,-nbitq), 
to_sfixed(-359402215.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-330686541.0/4294967296.0,1,-nbitq), 
to_sfixed(-139401319.0/4294967296.0,1,-nbitq), 
to_sfixed(-188338471.0/4294967296.0,1,-nbitq), 
to_sfixed(-502984732.0/4294967296.0,1,-nbitq), 
to_sfixed(-39105813.0/4294967296.0,1,-nbitq), 
to_sfixed(-33650468.0/4294967296.0,1,-nbitq), 
to_sfixed(-374902998.0/4294967296.0,1,-nbitq), 
to_sfixed(177473505.0/4294967296.0,1,-nbitq), 
to_sfixed(-445915703.0/4294967296.0,1,-nbitq), 
to_sfixed(341075096.0/4294967296.0,1,-nbitq), 
to_sfixed(61096556.0/4294967296.0,1,-nbitq), 
to_sfixed(-144400272.0/4294967296.0,1,-nbitq), 
to_sfixed(-27119166.0/4294967296.0,1,-nbitq), 
to_sfixed(-190776018.0/4294967296.0,1,-nbitq), 
to_sfixed(-48028110.0/4294967296.0,1,-nbitq), 
to_sfixed(-333227120.0/4294967296.0,1,-nbitq), 
to_sfixed(-168941369.0/4294967296.0,1,-nbitq), 
to_sfixed(308772963.0/4294967296.0,1,-nbitq), 
to_sfixed(-304052332.0/4294967296.0,1,-nbitq), 
to_sfixed(-283708540.0/4294967296.0,1,-nbitq), 
to_sfixed(248850690.0/4294967296.0,1,-nbitq), 
to_sfixed(-253838528.0/4294967296.0,1,-nbitq), 
to_sfixed(-94324068.0/4294967296.0,1,-nbitq), 
to_sfixed(-60873225.0/4294967296.0,1,-nbitq), 
to_sfixed(-66315573.0/4294967296.0,1,-nbitq), 
to_sfixed(512673981.0/4294967296.0,1,-nbitq), 
to_sfixed(-236621516.0/4294967296.0,1,-nbitq), 
to_sfixed(118738703.0/4294967296.0,1,-nbitq), 
to_sfixed(-13422510.0/4294967296.0,1,-nbitq), 
to_sfixed(392722037.0/4294967296.0,1,-nbitq), 
to_sfixed(-103985349.0/4294967296.0,1,-nbitq), 
to_sfixed(-160569447.0/4294967296.0,1,-nbitq), 
to_sfixed(235105312.0/4294967296.0,1,-nbitq), 
to_sfixed(15894900.0/4294967296.0,1,-nbitq), 
to_sfixed(57412771.0/4294967296.0,1,-nbitq), 
to_sfixed(-259851513.0/4294967296.0,1,-nbitq), 
to_sfixed(-267979915.0/4294967296.0,1,-nbitq), 
to_sfixed(177487329.0/4294967296.0,1,-nbitq), 
to_sfixed(-225551207.0/4294967296.0,1,-nbitq), 
to_sfixed(261947545.0/4294967296.0,1,-nbitq), 
to_sfixed(7317995.0/4294967296.0,1,-nbitq), 
to_sfixed(367086939.0/4294967296.0,1,-nbitq), 
to_sfixed(-142988315.0/4294967296.0,1,-nbitq), 
to_sfixed(-217977763.0/4294967296.0,1,-nbitq), 
to_sfixed(-347097866.0/4294967296.0,1,-nbitq), 
to_sfixed(-257868444.0/4294967296.0,1,-nbitq), 
to_sfixed(-235002174.0/4294967296.0,1,-nbitq), 
to_sfixed(82694316.0/4294967296.0,1,-nbitq), 
to_sfixed(-256070235.0/4294967296.0,1,-nbitq), 
to_sfixed(345316956.0/4294967296.0,1,-nbitq), 
to_sfixed(-13863583.0/4294967296.0,1,-nbitq), 
to_sfixed(-77404277.0/4294967296.0,1,-nbitq), 
to_sfixed(-469044300.0/4294967296.0,1,-nbitq), 
to_sfixed(-26858037.0/4294967296.0,1,-nbitq), 
to_sfixed(-67394462.0/4294967296.0,1,-nbitq), 
to_sfixed(109955517.0/4294967296.0,1,-nbitq), 
to_sfixed(334356635.0/4294967296.0,1,-nbitq), 
to_sfixed(134799408.0/4294967296.0,1,-nbitq), 
to_sfixed(-342387918.0/4294967296.0,1,-nbitq), 
to_sfixed(92589794.0/4294967296.0,1,-nbitq), 
to_sfixed(292192711.0/4294967296.0,1,-nbitq), 
to_sfixed(419747462.0/4294967296.0,1,-nbitq), 
to_sfixed(327276584.0/4294967296.0,1,-nbitq), 
to_sfixed(59887470.0/4294967296.0,1,-nbitq), 
to_sfixed(-176296799.0/4294967296.0,1,-nbitq), 
to_sfixed(123918685.0/4294967296.0,1,-nbitq), 
to_sfixed(129054050.0/4294967296.0,1,-nbitq), 
to_sfixed(-77433596.0/4294967296.0,1,-nbitq), 
to_sfixed(-113451881.0/4294967296.0,1,-nbitq), 
to_sfixed(600912062.0/4294967296.0,1,-nbitq), 
to_sfixed(-97799038.0/4294967296.0,1,-nbitq), 
to_sfixed(-373802745.0/4294967296.0,1,-nbitq), 
to_sfixed(-303845586.0/4294967296.0,1,-nbitq), 
to_sfixed(-24581102.0/4294967296.0,1,-nbitq), 
to_sfixed(-137473414.0/4294967296.0,1,-nbitq), 
to_sfixed(243983187.0/4294967296.0,1,-nbitq), 
to_sfixed(-261560355.0/4294967296.0,1,-nbitq), 
to_sfixed(167921770.0/4294967296.0,1,-nbitq), 
to_sfixed(98745809.0/4294967296.0,1,-nbitq), 
to_sfixed(-378746598.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(304718104.0/4294967296.0,1,-nbitq), 
to_sfixed(-38489767.0/4294967296.0,1,-nbitq), 
to_sfixed(490352889.0/4294967296.0,1,-nbitq), 
to_sfixed(-527498946.0/4294967296.0,1,-nbitq), 
to_sfixed(117512712.0/4294967296.0,1,-nbitq), 
to_sfixed(66547238.0/4294967296.0,1,-nbitq), 
to_sfixed(-271791555.0/4294967296.0,1,-nbitq), 
to_sfixed(339760158.0/4294967296.0,1,-nbitq), 
to_sfixed(-474087192.0/4294967296.0,1,-nbitq), 
to_sfixed(-184776136.0/4294967296.0,1,-nbitq), 
to_sfixed(-8502126.0/4294967296.0,1,-nbitq), 
to_sfixed(241504260.0/4294967296.0,1,-nbitq), 
to_sfixed(475975956.0/4294967296.0,1,-nbitq), 
to_sfixed(593404428.0/4294967296.0,1,-nbitq), 
to_sfixed(135495716.0/4294967296.0,1,-nbitq), 
to_sfixed(227059545.0/4294967296.0,1,-nbitq), 
to_sfixed(-376091785.0/4294967296.0,1,-nbitq), 
to_sfixed(-247430228.0/4294967296.0,1,-nbitq), 
to_sfixed(-92542275.0/4294967296.0,1,-nbitq), 
to_sfixed(258508932.0/4294967296.0,1,-nbitq), 
to_sfixed(-243799283.0/4294967296.0,1,-nbitq), 
to_sfixed(-90514121.0/4294967296.0,1,-nbitq), 
to_sfixed(-222674865.0/4294967296.0,1,-nbitq), 
to_sfixed(19004736.0/4294967296.0,1,-nbitq), 
to_sfixed(228025468.0/4294967296.0,1,-nbitq), 
to_sfixed(-161843818.0/4294967296.0,1,-nbitq), 
to_sfixed(25743408.0/4294967296.0,1,-nbitq), 
to_sfixed(-176660717.0/4294967296.0,1,-nbitq), 
to_sfixed(57624968.0/4294967296.0,1,-nbitq), 
to_sfixed(14262556.0/4294967296.0,1,-nbitq), 
to_sfixed(60080899.0/4294967296.0,1,-nbitq), 
to_sfixed(-260012321.0/4294967296.0,1,-nbitq), 
to_sfixed(-60987778.0/4294967296.0,1,-nbitq), 
to_sfixed(-310910896.0/4294967296.0,1,-nbitq), 
to_sfixed(-274190380.0/4294967296.0,1,-nbitq), 
to_sfixed(41430233.0/4294967296.0,1,-nbitq), 
to_sfixed(97776046.0/4294967296.0,1,-nbitq), 
to_sfixed(416076205.0/4294967296.0,1,-nbitq), 
to_sfixed(-328473836.0/4294967296.0,1,-nbitq), 
to_sfixed(460497073.0/4294967296.0,1,-nbitq), 
to_sfixed(-594707250.0/4294967296.0,1,-nbitq), 
to_sfixed(-44147086.0/4294967296.0,1,-nbitq), 
to_sfixed(-567068589.0/4294967296.0,1,-nbitq), 
to_sfixed(-14403617.0/4294967296.0,1,-nbitq), 
to_sfixed(-309851057.0/4294967296.0,1,-nbitq), 
to_sfixed(-121480752.0/4294967296.0,1,-nbitq), 
to_sfixed(-95586278.0/4294967296.0,1,-nbitq), 
to_sfixed(-359150552.0/4294967296.0,1,-nbitq), 
to_sfixed(-183099088.0/4294967296.0,1,-nbitq), 
to_sfixed(210411843.0/4294967296.0,1,-nbitq), 
to_sfixed(4153431.0/4294967296.0,1,-nbitq), 
to_sfixed(153569605.0/4294967296.0,1,-nbitq), 
to_sfixed(29394161.0/4294967296.0,1,-nbitq), 
to_sfixed(88499470.0/4294967296.0,1,-nbitq), 
to_sfixed(-118339331.0/4294967296.0,1,-nbitq), 
to_sfixed(57422071.0/4294967296.0,1,-nbitq), 
to_sfixed(62661045.0/4294967296.0,1,-nbitq), 
to_sfixed(42287588.0/4294967296.0,1,-nbitq), 
to_sfixed(268027420.0/4294967296.0,1,-nbitq), 
to_sfixed(-219062668.0/4294967296.0,1,-nbitq), 
to_sfixed(50368686.0/4294967296.0,1,-nbitq), 
to_sfixed(430972589.0/4294967296.0,1,-nbitq), 
to_sfixed(-137341449.0/4294967296.0,1,-nbitq), 
to_sfixed(208973054.0/4294967296.0,1,-nbitq), 
to_sfixed(-417472721.0/4294967296.0,1,-nbitq), 
to_sfixed(291822912.0/4294967296.0,1,-nbitq), 
to_sfixed(321720282.0/4294967296.0,1,-nbitq), 
to_sfixed(363407189.0/4294967296.0,1,-nbitq), 
to_sfixed(-66738935.0/4294967296.0,1,-nbitq), 
to_sfixed(751587890.0/4294967296.0,1,-nbitq), 
to_sfixed(453675154.0/4294967296.0,1,-nbitq), 
to_sfixed(285625296.0/4294967296.0,1,-nbitq), 
to_sfixed(-51880801.0/4294967296.0,1,-nbitq), 
to_sfixed(9494562.0/4294967296.0,1,-nbitq), 
to_sfixed(510209005.0/4294967296.0,1,-nbitq), 
to_sfixed(-159133998.0/4294967296.0,1,-nbitq), 
to_sfixed(117826022.0/4294967296.0,1,-nbitq), 
to_sfixed(-481267975.0/4294967296.0,1,-nbitq), 
to_sfixed(-99933844.0/4294967296.0,1,-nbitq), 
to_sfixed(104208125.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-54231126.0/4294967296.0,1,-nbitq), 
to_sfixed(-89940553.0/4294967296.0,1,-nbitq), 
to_sfixed(829134064.0/4294967296.0,1,-nbitq), 
to_sfixed(-553201526.0/4294967296.0,1,-nbitq), 
to_sfixed(-405126801.0/4294967296.0,1,-nbitq), 
to_sfixed(-226449262.0/4294967296.0,1,-nbitq), 
to_sfixed(57821412.0/4294967296.0,1,-nbitq), 
to_sfixed(337756637.0/4294967296.0,1,-nbitq), 
to_sfixed(-632495318.0/4294967296.0,1,-nbitq), 
to_sfixed(420902420.0/4294967296.0,1,-nbitq), 
to_sfixed(-181840248.0/4294967296.0,1,-nbitq), 
to_sfixed(-66522076.0/4294967296.0,1,-nbitq), 
to_sfixed(679920666.0/4294967296.0,1,-nbitq), 
to_sfixed(1072719597.0/4294967296.0,1,-nbitq), 
to_sfixed(-11632102.0/4294967296.0,1,-nbitq), 
to_sfixed(641869807.0/4294967296.0,1,-nbitq), 
to_sfixed(-71720949.0/4294967296.0,1,-nbitq), 
to_sfixed(330056871.0/4294967296.0,1,-nbitq), 
to_sfixed(-226033546.0/4294967296.0,1,-nbitq), 
to_sfixed(51878528.0/4294967296.0,1,-nbitq), 
to_sfixed(341007605.0/4294967296.0,1,-nbitq), 
to_sfixed(-571573413.0/4294967296.0,1,-nbitq), 
to_sfixed(-424609385.0/4294967296.0,1,-nbitq), 
to_sfixed(-73860019.0/4294967296.0,1,-nbitq), 
to_sfixed(383147625.0/4294967296.0,1,-nbitq), 
to_sfixed(-1124321285.0/4294967296.0,1,-nbitq), 
to_sfixed(74384537.0/4294967296.0,1,-nbitq), 
to_sfixed(103835819.0/4294967296.0,1,-nbitq), 
to_sfixed(206888702.0/4294967296.0,1,-nbitq), 
to_sfixed(53794480.0/4294967296.0,1,-nbitq), 
to_sfixed(-33869713.0/4294967296.0,1,-nbitq), 
to_sfixed(-99919513.0/4294967296.0,1,-nbitq), 
to_sfixed(-53112971.0/4294967296.0,1,-nbitq), 
to_sfixed(552451493.0/4294967296.0,1,-nbitq), 
to_sfixed(-131226699.0/4294967296.0,1,-nbitq), 
to_sfixed(-391233517.0/4294967296.0,1,-nbitq), 
to_sfixed(13634282.0/4294967296.0,1,-nbitq), 
to_sfixed(383845894.0/4294967296.0,1,-nbitq), 
to_sfixed(-363476897.0/4294967296.0,1,-nbitq), 
to_sfixed(123339830.0/4294967296.0,1,-nbitq), 
to_sfixed(-173871805.0/4294967296.0,1,-nbitq), 
to_sfixed(-187545679.0/4294967296.0,1,-nbitq), 
to_sfixed(-792679390.0/4294967296.0,1,-nbitq), 
to_sfixed(-220732231.0/4294967296.0,1,-nbitq), 
to_sfixed(-238922634.0/4294967296.0,1,-nbitq), 
to_sfixed(-183550235.0/4294967296.0,1,-nbitq), 
to_sfixed(-241155317.0/4294967296.0,1,-nbitq), 
to_sfixed(383880883.0/4294967296.0,1,-nbitq), 
to_sfixed(-179427821.0/4294967296.0,1,-nbitq), 
to_sfixed(-445350071.0/4294967296.0,1,-nbitq), 
to_sfixed(-202856011.0/4294967296.0,1,-nbitq), 
to_sfixed(-777927237.0/4294967296.0,1,-nbitq), 
to_sfixed(-281143414.0/4294967296.0,1,-nbitq), 
to_sfixed(51714369.0/4294967296.0,1,-nbitq), 
to_sfixed(468854553.0/4294967296.0,1,-nbitq), 
to_sfixed(24497876.0/4294967296.0,1,-nbitq), 
to_sfixed(38463588.0/4294967296.0,1,-nbitq), 
to_sfixed(187418925.0/4294967296.0,1,-nbitq), 
to_sfixed(-328531049.0/4294967296.0,1,-nbitq), 
to_sfixed(64534064.0/4294967296.0,1,-nbitq), 
to_sfixed(-44018390.0/4294967296.0,1,-nbitq), 
to_sfixed(51819428.0/4294967296.0,1,-nbitq), 
to_sfixed(767363249.0/4294967296.0,1,-nbitq), 
to_sfixed(-3050091.0/4294967296.0,1,-nbitq), 
to_sfixed(-344248371.0/4294967296.0,1,-nbitq), 
to_sfixed(-240872815.0/4294967296.0,1,-nbitq), 
to_sfixed(55144823.0/4294967296.0,1,-nbitq), 
to_sfixed(112452143.0/4294967296.0,1,-nbitq), 
to_sfixed(-337092805.0/4294967296.0,1,-nbitq), 
to_sfixed(249469147.0/4294967296.0,1,-nbitq), 
to_sfixed(579534536.0/4294967296.0,1,-nbitq), 
to_sfixed(182506839.0/4294967296.0,1,-nbitq), 
to_sfixed(258765369.0/4294967296.0,1,-nbitq), 
to_sfixed(-197016689.0/4294967296.0,1,-nbitq), 
to_sfixed(228683740.0/4294967296.0,1,-nbitq), 
to_sfixed(55269769.0/4294967296.0,1,-nbitq), 
to_sfixed(-970713508.0/4294967296.0,1,-nbitq), 
to_sfixed(-287087011.0/4294967296.0,1,-nbitq), 
to_sfixed(729923865.0/4294967296.0,1,-nbitq), 
to_sfixed(-326636634.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-126684811.0/4294967296.0,1,-nbitq), 
to_sfixed(194363334.0/4294967296.0,1,-nbitq), 
to_sfixed(1263735776.0/4294967296.0,1,-nbitq), 
to_sfixed(-1912863389.0/4294967296.0,1,-nbitq), 
to_sfixed(-1260866226.0/4294967296.0,1,-nbitq), 
to_sfixed(-497046411.0/4294967296.0,1,-nbitq), 
to_sfixed(-325266518.0/4294967296.0,1,-nbitq), 
to_sfixed(-111774740.0/4294967296.0,1,-nbitq), 
to_sfixed(-887585801.0/4294967296.0,1,-nbitq), 
to_sfixed(167262041.0/4294967296.0,1,-nbitq), 
to_sfixed(207724462.0/4294967296.0,1,-nbitq), 
to_sfixed(-406436934.0/4294967296.0,1,-nbitq), 
to_sfixed(1009169561.0/4294967296.0,1,-nbitq), 
to_sfixed(956471987.0/4294967296.0,1,-nbitq), 
to_sfixed(386725147.0/4294967296.0,1,-nbitq), 
to_sfixed(1299841405.0/4294967296.0,1,-nbitq), 
to_sfixed(-26606045.0/4294967296.0,1,-nbitq), 
to_sfixed(-338111501.0/4294967296.0,1,-nbitq), 
to_sfixed(75429273.0/4294967296.0,1,-nbitq), 
to_sfixed(1124213589.0/4294967296.0,1,-nbitq), 
to_sfixed(-417980062.0/4294967296.0,1,-nbitq), 
to_sfixed(-339282479.0/4294967296.0,1,-nbitq), 
to_sfixed(-1547046828.0/4294967296.0,1,-nbitq), 
to_sfixed(938866115.0/4294967296.0,1,-nbitq), 
to_sfixed(374658086.0/4294967296.0,1,-nbitq), 
to_sfixed(-1038350558.0/4294967296.0,1,-nbitq), 
to_sfixed(402373406.0/4294967296.0,1,-nbitq), 
to_sfixed(-11333903.0/4294967296.0,1,-nbitq), 
to_sfixed(126532457.0/4294967296.0,1,-nbitq), 
to_sfixed(1174218022.0/4294967296.0,1,-nbitq), 
to_sfixed(134439821.0/4294967296.0,1,-nbitq), 
to_sfixed(195133909.0/4294967296.0,1,-nbitq), 
to_sfixed(-230460702.0/4294967296.0,1,-nbitq), 
to_sfixed(487077756.0/4294967296.0,1,-nbitq), 
to_sfixed(-368435205.0/4294967296.0,1,-nbitq), 
to_sfixed(-84553058.0/4294967296.0,1,-nbitq), 
to_sfixed(-455284555.0/4294967296.0,1,-nbitq), 
to_sfixed(-456981232.0/4294967296.0,1,-nbitq), 
to_sfixed(20232687.0/4294967296.0,1,-nbitq), 
to_sfixed(-314136681.0/4294967296.0,1,-nbitq), 
to_sfixed(-567199149.0/4294967296.0,1,-nbitq), 
to_sfixed(-336917114.0/4294967296.0,1,-nbitq), 
to_sfixed(-58424867.0/4294967296.0,1,-nbitq), 
to_sfixed(169798086.0/4294967296.0,1,-nbitq), 
to_sfixed(-721428722.0/4294967296.0,1,-nbitq), 
to_sfixed(-216660638.0/4294967296.0,1,-nbitq), 
to_sfixed(-253851057.0/4294967296.0,1,-nbitq), 
to_sfixed(-39414557.0/4294967296.0,1,-nbitq), 
to_sfixed(36499696.0/4294967296.0,1,-nbitq), 
to_sfixed(84003803.0/4294967296.0,1,-nbitq), 
to_sfixed(19950965.0/4294967296.0,1,-nbitq), 
to_sfixed(-1382344451.0/4294967296.0,1,-nbitq), 
to_sfixed(-27401265.0/4294967296.0,1,-nbitq), 
to_sfixed(-94934682.0/4294967296.0,1,-nbitq), 
to_sfixed(56119420.0/4294967296.0,1,-nbitq), 
to_sfixed(-350194874.0/4294967296.0,1,-nbitq), 
to_sfixed(-162507129.0/4294967296.0,1,-nbitq), 
to_sfixed(79906475.0/4294967296.0,1,-nbitq), 
to_sfixed(-378079.0/4294967296.0,1,-nbitq), 
to_sfixed(137170360.0/4294967296.0,1,-nbitq), 
to_sfixed(-397972575.0/4294967296.0,1,-nbitq), 
to_sfixed(305027771.0/4294967296.0,1,-nbitq), 
to_sfixed(618836802.0/4294967296.0,1,-nbitq), 
to_sfixed(35989764.0/4294967296.0,1,-nbitq), 
to_sfixed(51092919.0/4294967296.0,1,-nbitq), 
to_sfixed(-86072409.0/4294967296.0,1,-nbitq), 
to_sfixed(47674533.0/4294967296.0,1,-nbitq), 
to_sfixed(144752110.0/4294967296.0,1,-nbitq), 
to_sfixed(-60338854.0/4294967296.0,1,-nbitq), 
to_sfixed(571025103.0/4294967296.0,1,-nbitq), 
to_sfixed(512488264.0/4294967296.0,1,-nbitq), 
to_sfixed(-240183972.0/4294967296.0,1,-nbitq), 
to_sfixed(-55889662.0/4294967296.0,1,-nbitq), 
to_sfixed(-31924277.0/4294967296.0,1,-nbitq), 
to_sfixed(536608347.0/4294967296.0,1,-nbitq), 
to_sfixed(-132737419.0/4294967296.0,1,-nbitq), 
to_sfixed(-545190852.0/4294967296.0,1,-nbitq), 
to_sfixed(259348816.0/4294967296.0,1,-nbitq), 
to_sfixed(1081678908.0/4294967296.0,1,-nbitq), 
to_sfixed(-336859481.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-98520066.0/4294967296.0,1,-nbitq), 
to_sfixed(308583181.0/4294967296.0,1,-nbitq), 
to_sfixed(428600539.0/4294967296.0,1,-nbitq), 
to_sfixed(-1837208307.0/4294967296.0,1,-nbitq), 
to_sfixed(-929881680.0/4294967296.0,1,-nbitq), 
to_sfixed(688754501.0/4294967296.0,1,-nbitq), 
to_sfixed(-433185619.0/4294967296.0,1,-nbitq), 
to_sfixed(323722123.0/4294967296.0,1,-nbitq), 
to_sfixed(-546226900.0/4294967296.0,1,-nbitq), 
to_sfixed(-156197823.0/4294967296.0,1,-nbitq), 
to_sfixed(-149486027.0/4294967296.0,1,-nbitq), 
to_sfixed(-268284983.0/4294967296.0,1,-nbitq), 
to_sfixed(983751991.0/4294967296.0,1,-nbitq), 
to_sfixed(1257732877.0/4294967296.0,1,-nbitq), 
to_sfixed(-189970634.0/4294967296.0,1,-nbitq), 
to_sfixed(1467990694.0/4294967296.0,1,-nbitq), 
to_sfixed(-338853711.0/4294967296.0,1,-nbitq), 
to_sfixed(-401749484.0/4294967296.0,1,-nbitq), 
to_sfixed(-718160267.0/4294967296.0,1,-nbitq), 
to_sfixed(1272809987.0/4294967296.0,1,-nbitq), 
to_sfixed(220205546.0/4294967296.0,1,-nbitq), 
to_sfixed(-306266882.0/4294967296.0,1,-nbitq), 
to_sfixed(-1162105671.0/4294967296.0,1,-nbitq), 
to_sfixed(646785591.0/4294967296.0,1,-nbitq), 
to_sfixed(-300740902.0/4294967296.0,1,-nbitq), 
to_sfixed(-1769100069.0/4294967296.0,1,-nbitq), 
to_sfixed(25974979.0/4294967296.0,1,-nbitq), 
to_sfixed(567595252.0/4294967296.0,1,-nbitq), 
to_sfixed(542477767.0/4294967296.0,1,-nbitq), 
to_sfixed(1303711325.0/4294967296.0,1,-nbitq), 
to_sfixed(-370964505.0/4294967296.0,1,-nbitq), 
to_sfixed(86444394.0/4294967296.0,1,-nbitq), 
to_sfixed(-87640978.0/4294967296.0,1,-nbitq), 
to_sfixed(328386512.0/4294967296.0,1,-nbitq), 
to_sfixed(-427795398.0/4294967296.0,1,-nbitq), 
to_sfixed(85391106.0/4294967296.0,1,-nbitq), 
to_sfixed(-289236294.0/4294967296.0,1,-nbitq), 
to_sfixed(-847311592.0/4294967296.0,1,-nbitq), 
to_sfixed(-253225330.0/4294967296.0,1,-nbitq), 
to_sfixed(-215324458.0/4294967296.0,1,-nbitq), 
to_sfixed(-452016918.0/4294967296.0,1,-nbitq), 
to_sfixed(-398480751.0/4294967296.0,1,-nbitq), 
to_sfixed(129789307.0/4294967296.0,1,-nbitq), 
to_sfixed(416316030.0/4294967296.0,1,-nbitq), 
to_sfixed(-1039288496.0/4294967296.0,1,-nbitq), 
to_sfixed(-685554857.0/4294967296.0,1,-nbitq), 
to_sfixed(178295364.0/4294967296.0,1,-nbitq), 
to_sfixed(336071086.0/4294967296.0,1,-nbitq), 
to_sfixed(248364173.0/4294967296.0,1,-nbitq), 
to_sfixed(49663724.0/4294967296.0,1,-nbitq), 
to_sfixed(-583123975.0/4294967296.0,1,-nbitq), 
to_sfixed(-1478047094.0/4294967296.0,1,-nbitq), 
to_sfixed(297358402.0/4294967296.0,1,-nbitq), 
to_sfixed(83590353.0/4294967296.0,1,-nbitq), 
to_sfixed(-120819319.0/4294967296.0,1,-nbitq), 
to_sfixed(-775235096.0/4294967296.0,1,-nbitq), 
to_sfixed(-384252382.0/4294967296.0,1,-nbitq), 
to_sfixed(-998732495.0/4294967296.0,1,-nbitq), 
to_sfixed(337230880.0/4294967296.0,1,-nbitq), 
to_sfixed(379009157.0/4294967296.0,1,-nbitq), 
to_sfixed(-69863738.0/4294967296.0,1,-nbitq), 
to_sfixed(312820380.0/4294967296.0,1,-nbitq), 
to_sfixed(816586259.0/4294967296.0,1,-nbitq), 
to_sfixed(-395134062.0/4294967296.0,1,-nbitq), 
to_sfixed(-397430030.0/4294967296.0,1,-nbitq), 
to_sfixed(360865094.0/4294967296.0,1,-nbitq), 
to_sfixed(-21171230.0/4294967296.0,1,-nbitq), 
to_sfixed(288228365.0/4294967296.0,1,-nbitq), 
to_sfixed(49201858.0/4294967296.0,1,-nbitq), 
to_sfixed(116206255.0/4294967296.0,1,-nbitq), 
to_sfixed(1187490945.0/4294967296.0,1,-nbitq), 
to_sfixed(130014682.0/4294967296.0,1,-nbitq), 
to_sfixed(470488435.0/4294967296.0,1,-nbitq), 
to_sfixed(-222979465.0/4294967296.0,1,-nbitq), 
to_sfixed(416187296.0/4294967296.0,1,-nbitq), 
to_sfixed(649428723.0/4294967296.0,1,-nbitq), 
to_sfixed(-1443328891.0/4294967296.0,1,-nbitq), 
to_sfixed(456216507.0/4294967296.0,1,-nbitq), 
to_sfixed(915080197.0/4294967296.0,1,-nbitq), 
to_sfixed(285217481.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-42454111.0/4294967296.0,1,-nbitq), 
to_sfixed(653356713.0/4294967296.0,1,-nbitq), 
to_sfixed(-657646573.0/4294967296.0,1,-nbitq), 
to_sfixed(-1494341977.0/4294967296.0,1,-nbitq), 
to_sfixed(314038328.0/4294967296.0,1,-nbitq), 
to_sfixed(1718362042.0/4294967296.0,1,-nbitq), 
to_sfixed(82304104.0/4294967296.0,1,-nbitq), 
to_sfixed(649364911.0/4294967296.0,1,-nbitq), 
to_sfixed(-1113031770.0/4294967296.0,1,-nbitq), 
to_sfixed(-61707673.0/4294967296.0,1,-nbitq), 
to_sfixed(-277660548.0/4294967296.0,1,-nbitq), 
to_sfixed(-843189677.0/4294967296.0,1,-nbitq), 
to_sfixed(-76491891.0/4294967296.0,1,-nbitq), 
to_sfixed(1516852549.0/4294967296.0,1,-nbitq), 
to_sfixed(370933823.0/4294967296.0,1,-nbitq), 
to_sfixed(1368091632.0/4294967296.0,1,-nbitq), 
to_sfixed(286337283.0/4294967296.0,1,-nbitq), 
to_sfixed(276010372.0/4294967296.0,1,-nbitq), 
to_sfixed(-521478244.0/4294967296.0,1,-nbitq), 
to_sfixed(694637738.0/4294967296.0,1,-nbitq), 
to_sfixed(312967088.0/4294967296.0,1,-nbitq), 
to_sfixed(-441243537.0/4294967296.0,1,-nbitq), 
to_sfixed(-794600406.0/4294967296.0,1,-nbitq), 
to_sfixed(762991592.0/4294967296.0,1,-nbitq), 
to_sfixed(459621870.0/4294967296.0,1,-nbitq), 
to_sfixed(-655146304.0/4294967296.0,1,-nbitq), 
to_sfixed(-292136588.0/4294967296.0,1,-nbitq), 
to_sfixed(2465864.0/4294967296.0,1,-nbitq), 
to_sfixed(700371660.0/4294967296.0,1,-nbitq), 
to_sfixed(556343990.0/4294967296.0,1,-nbitq), 
to_sfixed(-262407906.0/4294967296.0,1,-nbitq), 
to_sfixed(720925802.0/4294967296.0,1,-nbitq), 
to_sfixed(132959083.0/4294967296.0,1,-nbitq), 
to_sfixed(551797347.0/4294967296.0,1,-nbitq), 
to_sfixed(198524955.0/4294967296.0,1,-nbitq), 
to_sfixed(-1006259471.0/4294967296.0,1,-nbitq), 
to_sfixed(-77667008.0/4294967296.0,1,-nbitq), 
to_sfixed(520850281.0/4294967296.0,1,-nbitq), 
to_sfixed(-371653518.0/4294967296.0,1,-nbitq), 
to_sfixed(395020905.0/4294967296.0,1,-nbitq), 
to_sfixed(-587610394.0/4294967296.0,1,-nbitq), 
to_sfixed(-609636269.0/4294967296.0,1,-nbitq), 
to_sfixed(269144880.0/4294967296.0,1,-nbitq), 
to_sfixed(360226468.0/4294967296.0,1,-nbitq), 
to_sfixed(-480667268.0/4294967296.0,1,-nbitq), 
to_sfixed(-472539082.0/4294967296.0,1,-nbitq), 
to_sfixed(-111396425.0/4294967296.0,1,-nbitq), 
to_sfixed(705391676.0/4294967296.0,1,-nbitq), 
to_sfixed(245798847.0/4294967296.0,1,-nbitq), 
to_sfixed(-591849495.0/4294967296.0,1,-nbitq), 
to_sfixed(-244225181.0/4294967296.0,1,-nbitq), 
to_sfixed(-1390646235.0/4294967296.0,1,-nbitq), 
to_sfixed(471160000.0/4294967296.0,1,-nbitq), 
to_sfixed(286841335.0/4294967296.0,1,-nbitq), 
to_sfixed(290231486.0/4294967296.0,1,-nbitq), 
to_sfixed(-1043191718.0/4294967296.0,1,-nbitq), 
to_sfixed(-387040792.0/4294967296.0,1,-nbitq), 
to_sfixed(-879182979.0/4294967296.0,1,-nbitq), 
to_sfixed(-388536462.0/4294967296.0,1,-nbitq), 
to_sfixed(-72923775.0/4294967296.0,1,-nbitq), 
to_sfixed(-312917064.0/4294967296.0,1,-nbitq), 
to_sfixed(552551710.0/4294967296.0,1,-nbitq), 
to_sfixed(1119325016.0/4294967296.0,1,-nbitq), 
to_sfixed(-88884608.0/4294967296.0,1,-nbitq), 
to_sfixed(-177086211.0/4294967296.0,1,-nbitq), 
to_sfixed(-254542258.0/4294967296.0,1,-nbitq), 
to_sfixed(172612613.0/4294967296.0,1,-nbitq), 
to_sfixed(644261563.0/4294967296.0,1,-nbitq), 
to_sfixed(-9171534.0/4294967296.0,1,-nbitq), 
to_sfixed(-406393251.0/4294967296.0,1,-nbitq), 
to_sfixed(818932836.0/4294967296.0,1,-nbitq), 
to_sfixed(-283216251.0/4294967296.0,1,-nbitq), 
to_sfixed(-327388344.0/4294967296.0,1,-nbitq), 
to_sfixed(-348221045.0/4294967296.0,1,-nbitq), 
to_sfixed(-17800617.0/4294967296.0,1,-nbitq), 
to_sfixed(93944964.0/4294967296.0,1,-nbitq), 
to_sfixed(-1512768455.0/4294967296.0,1,-nbitq), 
to_sfixed(40924149.0/4294967296.0,1,-nbitq), 
to_sfixed(211415967.0/4294967296.0,1,-nbitq), 
to_sfixed(220809363.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-308057938.0/4294967296.0,1,-nbitq), 
to_sfixed(-365193996.0/4294967296.0,1,-nbitq), 
to_sfixed(-1630100386.0/4294967296.0,1,-nbitq), 
to_sfixed(-1684927496.0/4294967296.0,1,-nbitq), 
to_sfixed(-274466827.0/4294967296.0,1,-nbitq), 
to_sfixed(2313721225.0/4294967296.0,1,-nbitq), 
to_sfixed(279178469.0/4294967296.0,1,-nbitq), 
to_sfixed(1116383564.0/4294967296.0,1,-nbitq), 
to_sfixed(-1662738558.0/4294967296.0,1,-nbitq), 
to_sfixed(-209793088.0/4294967296.0,1,-nbitq), 
to_sfixed(-588623767.0/4294967296.0,1,-nbitq), 
to_sfixed(-1759913967.0/4294967296.0,1,-nbitq), 
to_sfixed(28185277.0/4294967296.0,1,-nbitq), 
to_sfixed(1438336628.0/4294967296.0,1,-nbitq), 
to_sfixed(-242030594.0/4294967296.0,1,-nbitq), 
to_sfixed(1279907565.0/4294967296.0,1,-nbitq), 
to_sfixed(-3060819.0/4294967296.0,1,-nbitq), 
to_sfixed(281328064.0/4294967296.0,1,-nbitq), 
to_sfixed(340578593.0/4294967296.0,1,-nbitq), 
to_sfixed(671104180.0/4294967296.0,1,-nbitq), 
to_sfixed(-117948668.0/4294967296.0,1,-nbitq), 
to_sfixed(-968148553.0/4294967296.0,1,-nbitq), 
to_sfixed(-876729556.0/4294967296.0,1,-nbitq), 
to_sfixed(1031296548.0/4294967296.0,1,-nbitq), 
to_sfixed(200239446.0/4294967296.0,1,-nbitq), 
to_sfixed(-923481136.0/4294967296.0,1,-nbitq), 
to_sfixed(613295877.0/4294967296.0,1,-nbitq), 
to_sfixed(236445642.0/4294967296.0,1,-nbitq), 
to_sfixed(234720204.0/4294967296.0,1,-nbitq), 
to_sfixed(1018536199.0/4294967296.0,1,-nbitq), 
to_sfixed(574658397.0/4294967296.0,1,-nbitq), 
to_sfixed(-80792047.0/4294967296.0,1,-nbitq), 
to_sfixed(-415781013.0/4294967296.0,1,-nbitq), 
to_sfixed(12595233.0/4294967296.0,1,-nbitq), 
to_sfixed(390620171.0/4294967296.0,1,-nbitq), 
to_sfixed(-665254355.0/4294967296.0,1,-nbitq), 
to_sfixed(147017876.0/4294967296.0,1,-nbitq), 
to_sfixed(995076368.0/4294967296.0,1,-nbitq), 
to_sfixed(101647072.0/4294967296.0,1,-nbitq), 
to_sfixed(-276537493.0/4294967296.0,1,-nbitq), 
to_sfixed(-248508755.0/4294967296.0,1,-nbitq), 
to_sfixed(-671875692.0/4294967296.0,1,-nbitq), 
to_sfixed(-115897160.0/4294967296.0,1,-nbitq), 
to_sfixed(-191569191.0/4294967296.0,1,-nbitq), 
to_sfixed(-870663684.0/4294967296.0,1,-nbitq), 
to_sfixed(-127921731.0/4294967296.0,1,-nbitq), 
to_sfixed(337692965.0/4294967296.0,1,-nbitq), 
to_sfixed(1284380885.0/4294967296.0,1,-nbitq), 
to_sfixed(67020739.0/4294967296.0,1,-nbitq), 
to_sfixed(-1273295264.0/4294967296.0,1,-nbitq), 
to_sfixed(-221883876.0/4294967296.0,1,-nbitq), 
to_sfixed(-2132237192.0/4294967296.0,1,-nbitq), 
to_sfixed(1005156626.0/4294967296.0,1,-nbitq), 
to_sfixed(-116088492.0/4294967296.0,1,-nbitq), 
to_sfixed(1067234949.0/4294967296.0,1,-nbitq), 
to_sfixed(-1054259231.0/4294967296.0,1,-nbitq), 
to_sfixed(-35734740.0/4294967296.0,1,-nbitq), 
to_sfixed(-1085325494.0/4294967296.0,1,-nbitq), 
to_sfixed(-180224457.0/4294967296.0,1,-nbitq), 
to_sfixed(-349135678.0/4294967296.0,1,-nbitq), 
to_sfixed(216412180.0/4294967296.0,1,-nbitq), 
to_sfixed(-10811109.0/4294967296.0,1,-nbitq), 
to_sfixed(1022061878.0/4294967296.0,1,-nbitq), 
to_sfixed(-718415540.0/4294967296.0,1,-nbitq), 
to_sfixed(-149621335.0/4294967296.0,1,-nbitq), 
to_sfixed(294045762.0/4294967296.0,1,-nbitq), 
to_sfixed(-646945245.0/4294967296.0,1,-nbitq), 
to_sfixed(662030663.0/4294967296.0,1,-nbitq), 
to_sfixed(60061854.0/4294967296.0,1,-nbitq), 
to_sfixed(-896650948.0/4294967296.0,1,-nbitq), 
to_sfixed(924051551.0/4294967296.0,1,-nbitq), 
to_sfixed(-232433383.0/4294967296.0,1,-nbitq), 
to_sfixed(63800089.0/4294967296.0,1,-nbitq), 
to_sfixed(138702704.0/4294967296.0,1,-nbitq), 
to_sfixed(101938963.0/4294967296.0,1,-nbitq), 
to_sfixed(455293511.0/4294967296.0,1,-nbitq), 
to_sfixed(-672105935.0/4294967296.0,1,-nbitq), 
to_sfixed(489134708.0/4294967296.0,1,-nbitq), 
to_sfixed(-514203323.0/4294967296.0,1,-nbitq), 
to_sfixed(-349938969.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-389813858.0/4294967296.0,1,-nbitq), 
to_sfixed(474854269.0/4294967296.0,1,-nbitq), 
to_sfixed(-1392517361.0/4294967296.0,1,-nbitq), 
to_sfixed(-286228428.0/4294967296.0,1,-nbitq), 
to_sfixed(-118245790.0/4294967296.0,1,-nbitq), 
to_sfixed(2141691251.0/4294967296.0,1,-nbitq), 
to_sfixed(156122696.0/4294967296.0,1,-nbitq), 
to_sfixed(1631529139.0/4294967296.0,1,-nbitq), 
to_sfixed(-1961172056.0/4294967296.0,1,-nbitq), 
to_sfixed(-62637105.0/4294967296.0,1,-nbitq), 
to_sfixed(475249770.0/4294967296.0,1,-nbitq), 
to_sfixed(-1391455418.0/4294967296.0,1,-nbitq), 
to_sfixed(617840430.0/4294967296.0,1,-nbitq), 
to_sfixed(1563415673.0/4294967296.0,1,-nbitq), 
to_sfixed(11754735.0/4294967296.0,1,-nbitq), 
to_sfixed(1051677905.0/4294967296.0,1,-nbitq), 
to_sfixed(-335594625.0/4294967296.0,1,-nbitq), 
to_sfixed(31659643.0/4294967296.0,1,-nbitq), 
to_sfixed(559671062.0/4294967296.0,1,-nbitq), 
to_sfixed(900405064.0/4294967296.0,1,-nbitq), 
to_sfixed(-111752394.0/4294967296.0,1,-nbitq), 
to_sfixed(-139881383.0/4294967296.0,1,-nbitq), 
to_sfixed(-386620735.0/4294967296.0,1,-nbitq), 
to_sfixed(1715636714.0/4294967296.0,1,-nbitq), 
to_sfixed(-85693293.0/4294967296.0,1,-nbitq), 
to_sfixed(-1235632180.0/4294967296.0,1,-nbitq), 
to_sfixed(748446756.0/4294967296.0,1,-nbitq), 
to_sfixed(-326031701.0/4294967296.0,1,-nbitq), 
to_sfixed(121784883.0/4294967296.0,1,-nbitq), 
to_sfixed(1504798693.0/4294967296.0,1,-nbitq), 
to_sfixed(7561315.0/4294967296.0,1,-nbitq), 
to_sfixed(92413464.0/4294967296.0,1,-nbitq), 
to_sfixed(-444097800.0/4294967296.0,1,-nbitq), 
to_sfixed(-65265141.0/4294967296.0,1,-nbitq), 
to_sfixed(45502497.0/4294967296.0,1,-nbitq), 
to_sfixed(26760734.0/4294967296.0,1,-nbitq), 
to_sfixed(371533986.0/4294967296.0,1,-nbitq), 
to_sfixed(212591391.0/4294967296.0,1,-nbitq), 
to_sfixed(18542955.0/4294967296.0,1,-nbitq), 
to_sfixed(155887748.0/4294967296.0,1,-nbitq), 
to_sfixed(-397218653.0/4294967296.0,1,-nbitq), 
to_sfixed(62214894.0/4294967296.0,1,-nbitq), 
to_sfixed(-758855056.0/4294967296.0,1,-nbitq), 
to_sfixed(-465928435.0/4294967296.0,1,-nbitq), 
to_sfixed(-1082295323.0/4294967296.0,1,-nbitq), 
to_sfixed(-210972582.0/4294967296.0,1,-nbitq), 
to_sfixed(191801359.0/4294967296.0,1,-nbitq), 
to_sfixed(1478430761.0/4294967296.0,1,-nbitq), 
to_sfixed(750862801.0/4294967296.0,1,-nbitq), 
to_sfixed(-1610961278.0/4294967296.0,1,-nbitq), 
to_sfixed(-50895731.0/4294967296.0,1,-nbitq), 
to_sfixed(-1009236010.0/4294967296.0,1,-nbitq), 
to_sfixed(1177322084.0/4294967296.0,1,-nbitq), 
to_sfixed(-34910471.0/4294967296.0,1,-nbitq), 
to_sfixed(1564311259.0/4294967296.0,1,-nbitq), 
to_sfixed(-684830859.0/4294967296.0,1,-nbitq), 
to_sfixed(-256220721.0/4294967296.0,1,-nbitq), 
to_sfixed(-535220642.0/4294967296.0,1,-nbitq), 
to_sfixed(-338095924.0/4294967296.0,1,-nbitq), 
to_sfixed(-218782553.0/4294967296.0,1,-nbitq), 
to_sfixed(263113031.0/4294967296.0,1,-nbitq), 
to_sfixed(-286202527.0/4294967296.0,1,-nbitq), 
to_sfixed(631616271.0/4294967296.0,1,-nbitq), 
to_sfixed(-522713245.0/4294967296.0,1,-nbitq), 
to_sfixed(-70424359.0/4294967296.0,1,-nbitq), 
to_sfixed(-474639891.0/4294967296.0,1,-nbitq), 
to_sfixed(-1703737458.0/4294967296.0,1,-nbitq), 
to_sfixed(44441407.0/4294967296.0,1,-nbitq), 
to_sfixed(93633406.0/4294967296.0,1,-nbitq), 
to_sfixed(-414572435.0/4294967296.0,1,-nbitq), 
to_sfixed(1961923809.0/4294967296.0,1,-nbitq), 
to_sfixed(120624736.0/4294967296.0,1,-nbitq), 
to_sfixed(34291741.0/4294967296.0,1,-nbitq), 
to_sfixed(-162578170.0/4294967296.0,1,-nbitq), 
to_sfixed(-98754962.0/4294967296.0,1,-nbitq), 
to_sfixed(328435517.0/4294967296.0,1,-nbitq), 
to_sfixed(-1202263669.0/4294967296.0,1,-nbitq), 
to_sfixed(732675783.0/4294967296.0,1,-nbitq), 
to_sfixed(-1612921213.0/4294967296.0,1,-nbitq), 
to_sfixed(321009433.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(268515238.0/4294967296.0,1,-nbitq), 
to_sfixed(1110882952.0/4294967296.0,1,-nbitq), 
to_sfixed(-404133403.0/4294967296.0,1,-nbitq), 
to_sfixed(-213829853.0/4294967296.0,1,-nbitq), 
to_sfixed(90189668.0/4294967296.0,1,-nbitq), 
to_sfixed(-81175753.0/4294967296.0,1,-nbitq), 
to_sfixed(584010863.0/4294967296.0,1,-nbitq), 
to_sfixed(1897171717.0/4294967296.0,1,-nbitq), 
to_sfixed(-1301695552.0/4294967296.0,1,-nbitq), 
to_sfixed(-257917458.0/4294967296.0,1,-nbitq), 
to_sfixed(87203672.0/4294967296.0,1,-nbitq), 
to_sfixed(-1970976974.0/4294967296.0,1,-nbitq), 
to_sfixed(327962015.0/4294967296.0,1,-nbitq), 
to_sfixed(1748202973.0/4294967296.0,1,-nbitq), 
to_sfixed(-64707172.0/4294967296.0,1,-nbitq), 
to_sfixed(1022499428.0/4294967296.0,1,-nbitq), 
to_sfixed(-280103705.0/4294967296.0,1,-nbitq), 
to_sfixed(112790893.0/4294967296.0,1,-nbitq), 
to_sfixed(675478151.0/4294967296.0,1,-nbitq), 
to_sfixed(439541591.0/4294967296.0,1,-nbitq), 
to_sfixed(328672823.0/4294967296.0,1,-nbitq), 
to_sfixed(-224963431.0/4294967296.0,1,-nbitq), 
to_sfixed(181849028.0/4294967296.0,1,-nbitq), 
to_sfixed(926128807.0/4294967296.0,1,-nbitq), 
to_sfixed(121147285.0/4294967296.0,1,-nbitq), 
to_sfixed(-1332054499.0/4294967296.0,1,-nbitq), 
to_sfixed(-225317614.0/4294967296.0,1,-nbitq), 
to_sfixed(586471283.0/4294967296.0,1,-nbitq), 
to_sfixed(983184025.0/4294967296.0,1,-nbitq), 
to_sfixed(1584730557.0/4294967296.0,1,-nbitq), 
to_sfixed(-206795977.0/4294967296.0,1,-nbitq), 
to_sfixed(-552663368.0/4294967296.0,1,-nbitq), 
to_sfixed(-700097162.0/4294967296.0,1,-nbitq), 
to_sfixed(-38971065.0/4294967296.0,1,-nbitq), 
to_sfixed(364598358.0/4294967296.0,1,-nbitq), 
to_sfixed(671113379.0/4294967296.0,1,-nbitq), 
to_sfixed(925737978.0/4294967296.0,1,-nbitq), 
to_sfixed(823090442.0/4294967296.0,1,-nbitq), 
to_sfixed(-333649762.0/4294967296.0,1,-nbitq), 
to_sfixed(569806006.0/4294967296.0,1,-nbitq), 
to_sfixed(-1132680399.0/4294967296.0,1,-nbitq), 
to_sfixed(-224583322.0/4294967296.0,1,-nbitq), 
to_sfixed(-349607531.0/4294967296.0,1,-nbitq), 
to_sfixed(-320976495.0/4294967296.0,1,-nbitq), 
to_sfixed(-519629765.0/4294967296.0,1,-nbitq), 
to_sfixed(53000564.0/4294967296.0,1,-nbitq), 
to_sfixed(-69901781.0/4294967296.0,1,-nbitq), 
to_sfixed(1410586399.0/4294967296.0,1,-nbitq), 
to_sfixed(435975542.0/4294967296.0,1,-nbitq), 
to_sfixed(-1445640508.0/4294967296.0,1,-nbitq), 
to_sfixed(-249381022.0/4294967296.0,1,-nbitq), 
to_sfixed(-1231376463.0/4294967296.0,1,-nbitq), 
to_sfixed(1117484861.0/4294967296.0,1,-nbitq), 
to_sfixed(-661184803.0/4294967296.0,1,-nbitq), 
to_sfixed(1371288802.0/4294967296.0,1,-nbitq), 
to_sfixed(-437952506.0/4294967296.0,1,-nbitq), 
to_sfixed(7596144.0/4294967296.0,1,-nbitq), 
to_sfixed(-1323634580.0/4294967296.0,1,-nbitq), 
to_sfixed(178255297.0/4294967296.0,1,-nbitq), 
to_sfixed(-113912101.0/4294967296.0,1,-nbitq), 
to_sfixed(60590400.0/4294967296.0,1,-nbitq), 
to_sfixed(-98346573.0/4294967296.0,1,-nbitq), 
to_sfixed(600228281.0/4294967296.0,1,-nbitq), 
to_sfixed(119157830.0/4294967296.0,1,-nbitq), 
to_sfixed(323128774.0/4294967296.0,1,-nbitq), 
to_sfixed(-407915727.0/4294967296.0,1,-nbitq), 
to_sfixed(-2657215009.0/4294967296.0,1,-nbitq), 
to_sfixed(-297818798.0/4294967296.0,1,-nbitq), 
to_sfixed(71831497.0/4294967296.0,1,-nbitq), 
to_sfixed(-873506645.0/4294967296.0,1,-nbitq), 
to_sfixed(1727070173.0/4294967296.0,1,-nbitq), 
to_sfixed(393389046.0/4294967296.0,1,-nbitq), 
to_sfixed(426239021.0/4294967296.0,1,-nbitq), 
to_sfixed(373607718.0/4294967296.0,1,-nbitq), 
to_sfixed(396899525.0/4294967296.0,1,-nbitq), 
to_sfixed(-509088958.0/4294967296.0,1,-nbitq), 
to_sfixed(-917189637.0/4294967296.0,1,-nbitq), 
to_sfixed(189088413.0/4294967296.0,1,-nbitq), 
to_sfixed(-1664866618.0/4294967296.0,1,-nbitq), 
to_sfixed(346275049.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(457360561.0/4294967296.0,1,-nbitq), 
to_sfixed(1162864705.0/4294967296.0,1,-nbitq), 
to_sfixed(-1244564981.0/4294967296.0,1,-nbitq), 
to_sfixed(-614633668.0/4294967296.0,1,-nbitq), 
to_sfixed(487407260.0/4294967296.0,1,-nbitq), 
to_sfixed(-1696253856.0/4294967296.0,1,-nbitq), 
to_sfixed(7072954.0/4294967296.0,1,-nbitq), 
to_sfixed(-845019527.0/4294967296.0,1,-nbitq), 
to_sfixed(-874724575.0/4294967296.0,1,-nbitq), 
to_sfixed(-280384011.0/4294967296.0,1,-nbitq), 
to_sfixed(-324183077.0/4294967296.0,1,-nbitq), 
to_sfixed(-1810035297.0/4294967296.0,1,-nbitq), 
to_sfixed(210786800.0/4294967296.0,1,-nbitq), 
to_sfixed(1087412480.0/4294967296.0,1,-nbitq), 
to_sfixed(189275119.0/4294967296.0,1,-nbitq), 
to_sfixed(1005285131.0/4294967296.0,1,-nbitq), 
to_sfixed(-192750920.0/4294967296.0,1,-nbitq), 
to_sfixed(72458238.0/4294967296.0,1,-nbitq), 
to_sfixed(255162113.0/4294967296.0,1,-nbitq), 
to_sfixed(255172975.0/4294967296.0,1,-nbitq), 
to_sfixed(70591719.0/4294967296.0,1,-nbitq), 
to_sfixed(-1027393160.0/4294967296.0,1,-nbitq), 
to_sfixed(-436346308.0/4294967296.0,1,-nbitq), 
to_sfixed(468140670.0/4294967296.0,1,-nbitq), 
to_sfixed(36374608.0/4294967296.0,1,-nbitq), 
to_sfixed(-569494904.0/4294967296.0,1,-nbitq), 
to_sfixed(-662017909.0/4294967296.0,1,-nbitq), 
to_sfixed(1508398501.0/4294967296.0,1,-nbitq), 
to_sfixed(1344768161.0/4294967296.0,1,-nbitq), 
to_sfixed(1259170848.0/4294967296.0,1,-nbitq), 
to_sfixed(96687060.0/4294967296.0,1,-nbitq), 
to_sfixed(244678797.0/4294967296.0,1,-nbitq), 
to_sfixed(-537890105.0/4294967296.0,1,-nbitq), 
to_sfixed(1061690771.0/4294967296.0,1,-nbitq), 
to_sfixed(657162749.0/4294967296.0,1,-nbitq), 
to_sfixed(-230249886.0/4294967296.0,1,-nbitq), 
to_sfixed(518811643.0/4294967296.0,1,-nbitq), 
to_sfixed(1546372880.0/4294967296.0,1,-nbitq), 
to_sfixed(-466365228.0/4294967296.0,1,-nbitq), 
to_sfixed(63167643.0/4294967296.0,1,-nbitq), 
to_sfixed(-378060223.0/4294967296.0,1,-nbitq), 
to_sfixed(-13904822.0/4294967296.0,1,-nbitq), 
to_sfixed(-796466504.0/4294967296.0,1,-nbitq), 
to_sfixed(-365422340.0/4294967296.0,1,-nbitq), 
to_sfixed(-879865563.0/4294967296.0,1,-nbitq), 
to_sfixed(-1097569999.0/4294967296.0,1,-nbitq), 
to_sfixed(127863379.0/4294967296.0,1,-nbitq), 
to_sfixed(1218020299.0/4294967296.0,1,-nbitq), 
to_sfixed(230733260.0/4294967296.0,1,-nbitq), 
to_sfixed(-1631638765.0/4294967296.0,1,-nbitq), 
to_sfixed(-827240268.0/4294967296.0,1,-nbitq), 
to_sfixed(-724988645.0/4294967296.0,1,-nbitq), 
to_sfixed(1848058674.0/4294967296.0,1,-nbitq), 
to_sfixed(244515998.0/4294967296.0,1,-nbitq), 
to_sfixed(1721261203.0/4294967296.0,1,-nbitq), 
to_sfixed(-54635726.0/4294967296.0,1,-nbitq), 
to_sfixed(424661613.0/4294967296.0,1,-nbitq), 
to_sfixed(-928074175.0/4294967296.0,1,-nbitq), 
to_sfixed(174748522.0/4294967296.0,1,-nbitq), 
to_sfixed(-291338090.0/4294967296.0,1,-nbitq), 
to_sfixed(-210474051.0/4294967296.0,1,-nbitq), 
to_sfixed(186972014.0/4294967296.0,1,-nbitq), 
to_sfixed(-1475779001.0/4294967296.0,1,-nbitq), 
to_sfixed(-595725011.0/4294967296.0,1,-nbitq), 
to_sfixed(-213073929.0/4294967296.0,1,-nbitq), 
to_sfixed(90663497.0/4294967296.0,1,-nbitq), 
to_sfixed(-469111449.0/4294967296.0,1,-nbitq), 
to_sfixed(-818732301.0/4294967296.0,1,-nbitq), 
to_sfixed(389899273.0/4294967296.0,1,-nbitq), 
to_sfixed(-571486688.0/4294967296.0,1,-nbitq), 
to_sfixed(1416018571.0/4294967296.0,1,-nbitq), 
to_sfixed(125602130.0/4294967296.0,1,-nbitq), 
to_sfixed(82750518.0/4294967296.0,1,-nbitq), 
to_sfixed(-18699358.0/4294967296.0,1,-nbitq), 
to_sfixed(113390500.0/4294967296.0,1,-nbitq), 
to_sfixed(-1678888868.0/4294967296.0,1,-nbitq), 
to_sfixed(-749946845.0/4294967296.0,1,-nbitq), 
to_sfixed(545303994.0/4294967296.0,1,-nbitq), 
to_sfixed(-967121924.0/4294967296.0,1,-nbitq), 
to_sfixed(221525855.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(342248595.0/4294967296.0,1,-nbitq), 
to_sfixed(321149610.0/4294967296.0,1,-nbitq), 
to_sfixed(-1559389947.0/4294967296.0,1,-nbitq), 
to_sfixed(-883231242.0/4294967296.0,1,-nbitq), 
to_sfixed(1691626636.0/4294967296.0,1,-nbitq), 
to_sfixed(-467247019.0/4294967296.0,1,-nbitq), 
to_sfixed(653161226.0/4294967296.0,1,-nbitq), 
to_sfixed(-1772770962.0/4294967296.0,1,-nbitq), 
to_sfixed(-851971161.0/4294967296.0,1,-nbitq), 
to_sfixed(44225733.0/4294967296.0,1,-nbitq), 
to_sfixed(-677540317.0/4294967296.0,1,-nbitq), 
to_sfixed(-1454266359.0/4294967296.0,1,-nbitq), 
to_sfixed(-352221363.0/4294967296.0,1,-nbitq), 
to_sfixed(-230079290.0/4294967296.0,1,-nbitq), 
to_sfixed(240442388.0/4294967296.0,1,-nbitq), 
to_sfixed(643481307.0/4294967296.0,1,-nbitq), 
to_sfixed(259845634.0/4294967296.0,1,-nbitq), 
to_sfixed(88301934.0/4294967296.0,1,-nbitq), 
to_sfixed(263693836.0/4294967296.0,1,-nbitq), 
to_sfixed(152260524.0/4294967296.0,1,-nbitq), 
to_sfixed(-181775262.0/4294967296.0,1,-nbitq), 
to_sfixed(-1538260328.0/4294967296.0,1,-nbitq), 
to_sfixed(-498254771.0/4294967296.0,1,-nbitq), 
to_sfixed(725511438.0/4294967296.0,1,-nbitq), 
to_sfixed(-183257891.0/4294967296.0,1,-nbitq), 
to_sfixed(-767527748.0/4294967296.0,1,-nbitq), 
to_sfixed(-230735477.0/4294967296.0,1,-nbitq), 
to_sfixed(1703999951.0/4294967296.0,1,-nbitq), 
to_sfixed(-1866352546.0/4294967296.0,1,-nbitq), 
to_sfixed(322141305.0/4294967296.0,1,-nbitq), 
to_sfixed(1551873766.0/4294967296.0,1,-nbitq), 
to_sfixed(478161005.0/4294967296.0,1,-nbitq), 
to_sfixed(-806800887.0/4294967296.0,1,-nbitq), 
to_sfixed(1794514638.0/4294967296.0,1,-nbitq), 
to_sfixed(510686962.0/4294967296.0,1,-nbitq), 
to_sfixed(1296177171.0/4294967296.0,1,-nbitq), 
to_sfixed(478677537.0/4294967296.0,1,-nbitq), 
to_sfixed(1353862878.0/4294967296.0,1,-nbitq), 
to_sfixed(86540657.0/4294967296.0,1,-nbitq), 
to_sfixed(-144974844.0/4294967296.0,1,-nbitq), 
to_sfixed(-506799086.0/4294967296.0,1,-nbitq), 
to_sfixed(-913414205.0/4294967296.0,1,-nbitq), 
to_sfixed(-915788721.0/4294967296.0,1,-nbitq), 
to_sfixed(-548366184.0/4294967296.0,1,-nbitq), 
to_sfixed(-321672656.0/4294967296.0,1,-nbitq), 
to_sfixed(-43447665.0/4294967296.0,1,-nbitq), 
to_sfixed(-5060640.0/4294967296.0,1,-nbitq), 
to_sfixed(298578101.0/4294967296.0,1,-nbitq), 
to_sfixed(-33150958.0/4294967296.0,1,-nbitq), 
to_sfixed(-1100017415.0/4294967296.0,1,-nbitq), 
to_sfixed(-521327769.0/4294967296.0,1,-nbitq), 
to_sfixed(348167796.0/4294967296.0,1,-nbitq), 
to_sfixed(1956465674.0/4294967296.0,1,-nbitq), 
to_sfixed(-648462171.0/4294967296.0,1,-nbitq), 
to_sfixed(2458796689.0/4294967296.0,1,-nbitq), 
to_sfixed(-349645948.0/4294967296.0,1,-nbitq), 
to_sfixed(492441269.0/4294967296.0,1,-nbitq), 
to_sfixed(-352932702.0/4294967296.0,1,-nbitq), 
to_sfixed(-243875113.0/4294967296.0,1,-nbitq), 
to_sfixed(395817364.0/4294967296.0,1,-nbitq), 
to_sfixed(236944969.0/4294967296.0,1,-nbitq), 
to_sfixed(-252105121.0/4294967296.0,1,-nbitq), 
to_sfixed(-2235395411.0/4294967296.0,1,-nbitq), 
to_sfixed(-1132366680.0/4294967296.0,1,-nbitq), 
to_sfixed(-171318456.0/4294967296.0,1,-nbitq), 
to_sfixed(49933341.0/4294967296.0,1,-nbitq), 
to_sfixed(1696809711.0/4294967296.0,1,-nbitq), 
to_sfixed(-984114859.0/4294967296.0,1,-nbitq), 
to_sfixed(348991731.0/4294967296.0,1,-nbitq), 
to_sfixed(1340137777.0/4294967296.0,1,-nbitq), 
to_sfixed(404203262.0/4294967296.0,1,-nbitq), 
to_sfixed(175497689.0/4294967296.0,1,-nbitq), 
to_sfixed(6754571.0/4294967296.0,1,-nbitq), 
to_sfixed(359560881.0/4294967296.0,1,-nbitq), 
to_sfixed(255120771.0/4294967296.0,1,-nbitq), 
to_sfixed(-745580723.0/4294967296.0,1,-nbitq), 
to_sfixed(-69494614.0/4294967296.0,1,-nbitq), 
to_sfixed(678757987.0/4294967296.0,1,-nbitq), 
to_sfixed(-1005618019.0/4294967296.0,1,-nbitq), 
to_sfixed(-357699952.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(7284479.0/4294967296.0,1,-nbitq), 
to_sfixed(-458522544.0/4294967296.0,1,-nbitq), 
to_sfixed(-298315747.0/4294967296.0,1,-nbitq), 
to_sfixed(-1891723329.0/4294967296.0,1,-nbitq), 
to_sfixed(1653935142.0/4294967296.0,1,-nbitq), 
to_sfixed(-247935728.0/4294967296.0,1,-nbitq), 
to_sfixed(524167515.0/4294967296.0,1,-nbitq), 
to_sfixed(-1494526046.0/4294967296.0,1,-nbitq), 
to_sfixed(-2020719815.0/4294967296.0,1,-nbitq), 
to_sfixed(-71730841.0/4294967296.0,1,-nbitq), 
to_sfixed(-838334789.0/4294967296.0,1,-nbitq), 
to_sfixed(32762687.0/4294967296.0,1,-nbitq), 
to_sfixed(35622097.0/4294967296.0,1,-nbitq), 
to_sfixed(381263305.0/4294967296.0,1,-nbitq), 
to_sfixed(-49595746.0/4294967296.0,1,-nbitq), 
to_sfixed(-71474758.0/4294967296.0,1,-nbitq), 
to_sfixed(292219533.0/4294967296.0,1,-nbitq), 
to_sfixed(385935285.0/4294967296.0,1,-nbitq), 
to_sfixed(383452262.0/4294967296.0,1,-nbitq), 
to_sfixed(-300356873.0/4294967296.0,1,-nbitq), 
to_sfixed(197843743.0/4294967296.0,1,-nbitq), 
to_sfixed(-1917970934.0/4294967296.0,1,-nbitq), 
to_sfixed(910110478.0/4294967296.0,1,-nbitq), 
to_sfixed(2242214153.0/4294967296.0,1,-nbitq), 
to_sfixed(73281832.0/4294967296.0,1,-nbitq), 
to_sfixed(-864230006.0/4294967296.0,1,-nbitq), 
to_sfixed(-371310709.0/4294967296.0,1,-nbitq), 
to_sfixed(-48236584.0/4294967296.0,1,-nbitq), 
to_sfixed(-2300902598.0/4294967296.0,1,-nbitq), 
to_sfixed(581925438.0/4294967296.0,1,-nbitq), 
to_sfixed(2045104002.0/4294967296.0,1,-nbitq), 
to_sfixed(-206890017.0/4294967296.0,1,-nbitq), 
to_sfixed(-1041893962.0/4294967296.0,1,-nbitq), 
to_sfixed(984636727.0/4294967296.0,1,-nbitq), 
to_sfixed(-586414594.0/4294967296.0,1,-nbitq), 
to_sfixed(1827254138.0/4294967296.0,1,-nbitq), 
to_sfixed(422206212.0/4294967296.0,1,-nbitq), 
to_sfixed(915293248.0/4294967296.0,1,-nbitq), 
to_sfixed(-161839680.0/4294967296.0,1,-nbitq), 
to_sfixed(-102113295.0/4294967296.0,1,-nbitq), 
to_sfixed(418271297.0/4294967296.0,1,-nbitq), 
to_sfixed(-682242472.0/4294967296.0,1,-nbitq), 
to_sfixed(-203069455.0/4294967296.0,1,-nbitq), 
to_sfixed(-181608532.0/4294967296.0,1,-nbitq), 
to_sfixed(-1057128530.0/4294967296.0,1,-nbitq), 
to_sfixed(-244517600.0/4294967296.0,1,-nbitq), 
to_sfixed(195758032.0/4294967296.0,1,-nbitq), 
to_sfixed(688823337.0/4294967296.0,1,-nbitq), 
to_sfixed(-117819742.0/4294967296.0,1,-nbitq), 
to_sfixed(-1002683652.0/4294967296.0,1,-nbitq), 
to_sfixed(-595540385.0/4294967296.0,1,-nbitq), 
to_sfixed(-259443571.0/4294967296.0,1,-nbitq), 
to_sfixed(1097786798.0/4294967296.0,1,-nbitq), 
to_sfixed(-891179617.0/4294967296.0,1,-nbitq), 
to_sfixed(1297200330.0/4294967296.0,1,-nbitq), 
to_sfixed(-1132001558.0/4294967296.0,1,-nbitq), 
to_sfixed(415440793.0/4294967296.0,1,-nbitq), 
to_sfixed(-369178057.0/4294967296.0,1,-nbitq), 
to_sfixed(-167953867.0/4294967296.0,1,-nbitq), 
to_sfixed(-293174653.0/4294967296.0,1,-nbitq), 
to_sfixed(-256388999.0/4294967296.0,1,-nbitq), 
to_sfixed(-331620532.0/4294967296.0,1,-nbitq), 
to_sfixed(-1535476233.0/4294967296.0,1,-nbitq), 
to_sfixed(-626953710.0/4294967296.0,1,-nbitq), 
to_sfixed(-388884038.0/4294967296.0,1,-nbitq), 
to_sfixed(308115278.0/4294967296.0,1,-nbitq), 
to_sfixed(24976974.0/4294967296.0,1,-nbitq), 
to_sfixed(600272287.0/4294967296.0,1,-nbitq), 
to_sfixed(88841020.0/4294967296.0,1,-nbitq), 
to_sfixed(681804101.0/4294967296.0,1,-nbitq), 
to_sfixed(739445222.0/4294967296.0,1,-nbitq), 
to_sfixed(-162240818.0/4294967296.0,1,-nbitq), 
to_sfixed(-453295752.0/4294967296.0,1,-nbitq), 
to_sfixed(-198299718.0/4294967296.0,1,-nbitq), 
to_sfixed(-16681623.0/4294967296.0,1,-nbitq), 
to_sfixed(224338434.0/4294967296.0,1,-nbitq), 
to_sfixed(-1317070033.0/4294967296.0,1,-nbitq), 
to_sfixed(163980818.0/4294967296.0,1,-nbitq), 
to_sfixed(-375115924.0/4294967296.0,1,-nbitq), 
to_sfixed(1676106.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(334122462.0/4294967296.0,1,-nbitq), 
to_sfixed(-108182392.0/4294967296.0,1,-nbitq), 
to_sfixed(-123813590.0/4294967296.0,1,-nbitq), 
to_sfixed(-1054817375.0/4294967296.0,1,-nbitq), 
to_sfixed(2222357698.0/4294967296.0,1,-nbitq), 
to_sfixed(413730116.0/4294967296.0,1,-nbitq), 
to_sfixed(311866568.0/4294967296.0,1,-nbitq), 
to_sfixed(-280239357.0/4294967296.0,1,-nbitq), 
to_sfixed(-2100883877.0/4294967296.0,1,-nbitq), 
to_sfixed(365996978.0/4294967296.0,1,-nbitq), 
to_sfixed(-483660730.0/4294967296.0,1,-nbitq), 
to_sfixed(1460555827.0/4294967296.0,1,-nbitq), 
to_sfixed(1098655028.0/4294967296.0,1,-nbitq), 
to_sfixed(241508946.0/4294967296.0,1,-nbitq), 
to_sfixed(-405277972.0/4294967296.0,1,-nbitq), 
to_sfixed(-285643318.0/4294967296.0,1,-nbitq), 
to_sfixed(143651082.0/4294967296.0,1,-nbitq), 
to_sfixed(348365761.0/4294967296.0,1,-nbitq), 
to_sfixed(-1438979072.0/4294967296.0,1,-nbitq), 
to_sfixed(-866693726.0/4294967296.0,1,-nbitq), 
to_sfixed(-76007996.0/4294967296.0,1,-nbitq), 
to_sfixed(-660799326.0/4294967296.0,1,-nbitq), 
to_sfixed(1664175200.0/4294967296.0,1,-nbitq), 
to_sfixed(-97118839.0/4294967296.0,1,-nbitq), 
to_sfixed(-354295476.0/4294967296.0,1,-nbitq), 
to_sfixed(-504533989.0/4294967296.0,1,-nbitq), 
to_sfixed(-140522097.0/4294967296.0,1,-nbitq), 
to_sfixed(-1048927832.0/4294967296.0,1,-nbitq), 
to_sfixed(-1172000387.0/4294967296.0,1,-nbitq), 
to_sfixed(530017438.0/4294967296.0,1,-nbitq), 
to_sfixed(251823627.0/4294967296.0,1,-nbitq), 
to_sfixed(-534150343.0/4294967296.0,1,-nbitq), 
to_sfixed(-1279928958.0/4294967296.0,1,-nbitq), 
to_sfixed(1091568953.0/4294967296.0,1,-nbitq), 
to_sfixed(-119811430.0/4294967296.0,1,-nbitq), 
to_sfixed(588804759.0/4294967296.0,1,-nbitq), 
to_sfixed(20258245.0/4294967296.0,1,-nbitq), 
to_sfixed(-42940437.0/4294967296.0,1,-nbitq), 
to_sfixed(115515882.0/4294967296.0,1,-nbitq), 
to_sfixed(-216824692.0/4294967296.0,1,-nbitq), 
to_sfixed(1432500593.0/4294967296.0,1,-nbitq), 
to_sfixed(480717178.0/4294967296.0,1,-nbitq), 
to_sfixed(-63445012.0/4294967296.0,1,-nbitq), 
to_sfixed(564854198.0/4294967296.0,1,-nbitq), 
to_sfixed(-1039004296.0/4294967296.0,1,-nbitq), 
to_sfixed(268402791.0/4294967296.0,1,-nbitq), 
to_sfixed(88549424.0/4294967296.0,1,-nbitq), 
to_sfixed(787193620.0/4294967296.0,1,-nbitq), 
to_sfixed(-690526822.0/4294967296.0,1,-nbitq), 
to_sfixed(-1381354926.0/4294967296.0,1,-nbitq), 
to_sfixed(-24426181.0/4294967296.0,1,-nbitq), 
to_sfixed(224661224.0/4294967296.0,1,-nbitq), 
to_sfixed(823260093.0/4294967296.0,1,-nbitq), 
to_sfixed(-761853699.0/4294967296.0,1,-nbitq), 
to_sfixed(-1680075770.0/4294967296.0,1,-nbitq), 
to_sfixed(-119908842.0/4294967296.0,1,-nbitq), 
to_sfixed(-576366813.0/4294967296.0,1,-nbitq), 
to_sfixed(-466936583.0/4294967296.0,1,-nbitq), 
to_sfixed(22534547.0/4294967296.0,1,-nbitq), 
to_sfixed(16935396.0/4294967296.0,1,-nbitq), 
to_sfixed(-144756884.0/4294967296.0,1,-nbitq), 
to_sfixed(-654342064.0/4294967296.0,1,-nbitq), 
to_sfixed(-608249030.0/4294967296.0,1,-nbitq), 
to_sfixed(-531238231.0/4294967296.0,1,-nbitq), 
to_sfixed(64354585.0/4294967296.0,1,-nbitq), 
to_sfixed(-138093867.0/4294967296.0,1,-nbitq), 
to_sfixed(474830017.0/4294967296.0,1,-nbitq), 
to_sfixed(928942719.0/4294967296.0,1,-nbitq), 
to_sfixed(-367908506.0/4294967296.0,1,-nbitq), 
to_sfixed(1264678426.0/4294967296.0,1,-nbitq), 
to_sfixed(1076479881.0/4294967296.0,1,-nbitq), 
to_sfixed(-690784659.0/4294967296.0,1,-nbitq), 
to_sfixed(-277695207.0/4294967296.0,1,-nbitq), 
to_sfixed(-93699931.0/4294967296.0,1,-nbitq), 
to_sfixed(-326112044.0/4294967296.0,1,-nbitq), 
to_sfixed(-285699166.0/4294967296.0,1,-nbitq), 
to_sfixed(-683225772.0/4294967296.0,1,-nbitq), 
to_sfixed(137743255.0/4294967296.0,1,-nbitq), 
to_sfixed(386729057.0/4294967296.0,1,-nbitq), 
to_sfixed(27346381.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(300091343.0/4294967296.0,1,-nbitq), 
to_sfixed(552237958.0/4294967296.0,1,-nbitq), 
to_sfixed(-186556391.0/4294967296.0,1,-nbitq), 
to_sfixed(38276756.0/4294967296.0,1,-nbitq), 
to_sfixed(1425735512.0/4294967296.0,1,-nbitq), 
to_sfixed(1694698084.0/4294967296.0,1,-nbitq), 
to_sfixed(-180114243.0/4294967296.0,1,-nbitq), 
to_sfixed(600737431.0/4294967296.0,1,-nbitq), 
to_sfixed(-2110948533.0/4294967296.0,1,-nbitq), 
to_sfixed(-358170584.0/4294967296.0,1,-nbitq), 
to_sfixed(-318889270.0/4294967296.0,1,-nbitq), 
to_sfixed(1403902766.0/4294967296.0,1,-nbitq), 
to_sfixed(1016600143.0/4294967296.0,1,-nbitq), 
to_sfixed(-901047946.0/4294967296.0,1,-nbitq), 
to_sfixed(156325632.0/4294967296.0,1,-nbitq), 
to_sfixed(126715596.0/4294967296.0,1,-nbitq), 
to_sfixed(-146730301.0/4294967296.0,1,-nbitq), 
to_sfixed(-230187063.0/4294967296.0,1,-nbitq), 
to_sfixed(-2281074597.0/4294967296.0,1,-nbitq), 
to_sfixed(-1107841258.0/4294967296.0,1,-nbitq), 
to_sfixed(311040825.0/4294967296.0,1,-nbitq), 
to_sfixed(-69305127.0/4294967296.0,1,-nbitq), 
to_sfixed(709618675.0/4294967296.0,1,-nbitq), 
to_sfixed(-2347523131.0/4294967296.0,1,-nbitq), 
to_sfixed(-266607032.0/4294967296.0,1,-nbitq), 
to_sfixed(-89129468.0/4294967296.0,1,-nbitq), 
to_sfixed(-821261597.0/4294967296.0,1,-nbitq), 
to_sfixed(-749115125.0/4294967296.0,1,-nbitq), 
to_sfixed(1140019756.0/4294967296.0,1,-nbitq), 
to_sfixed(1553255050.0/4294967296.0,1,-nbitq), 
to_sfixed(-2281868656.0/4294967296.0,1,-nbitq), 
to_sfixed(-1171469658.0/4294967296.0,1,-nbitq), 
to_sfixed(-1035581222.0/4294967296.0,1,-nbitq), 
to_sfixed(754432413.0/4294967296.0,1,-nbitq), 
to_sfixed(945148390.0/4294967296.0,1,-nbitq), 
to_sfixed(-810544130.0/4294967296.0,1,-nbitq), 
to_sfixed(-298226279.0/4294967296.0,1,-nbitq), 
to_sfixed(-686907456.0/4294967296.0,1,-nbitq), 
to_sfixed(112805999.0/4294967296.0,1,-nbitq), 
to_sfixed(-216928065.0/4294967296.0,1,-nbitq), 
to_sfixed(857499661.0/4294967296.0,1,-nbitq), 
to_sfixed(1128641275.0/4294967296.0,1,-nbitq), 
to_sfixed(-653473975.0/4294967296.0,1,-nbitq), 
to_sfixed(334008791.0/4294967296.0,1,-nbitq), 
to_sfixed(-1026534336.0/4294967296.0,1,-nbitq), 
to_sfixed(-1231408097.0/4294967296.0,1,-nbitq), 
to_sfixed(332789362.0/4294967296.0,1,-nbitq), 
to_sfixed(630739356.0/4294967296.0,1,-nbitq), 
to_sfixed(-210071717.0/4294967296.0,1,-nbitq), 
to_sfixed(-108096589.0/4294967296.0,1,-nbitq), 
to_sfixed(-539206474.0/4294967296.0,1,-nbitq), 
to_sfixed(334476666.0/4294967296.0,1,-nbitq), 
to_sfixed(1336620410.0/4294967296.0,1,-nbitq), 
to_sfixed(-869989977.0/4294967296.0,1,-nbitq), 
to_sfixed(-1580082083.0/4294967296.0,1,-nbitq), 
to_sfixed(-390380884.0/4294967296.0,1,-nbitq), 
to_sfixed(-652946703.0/4294967296.0,1,-nbitq), 
to_sfixed(959018538.0/4294967296.0,1,-nbitq), 
to_sfixed(-122063206.0/4294967296.0,1,-nbitq), 
to_sfixed(-338283247.0/4294967296.0,1,-nbitq), 
to_sfixed(-228327665.0/4294967296.0,1,-nbitq), 
to_sfixed(-884249426.0/4294967296.0,1,-nbitq), 
to_sfixed(1379816916.0/4294967296.0,1,-nbitq), 
to_sfixed(439424858.0/4294967296.0,1,-nbitq), 
to_sfixed(-694887124.0/4294967296.0,1,-nbitq), 
to_sfixed(-62692672.0/4294967296.0,1,-nbitq), 
to_sfixed(1079483190.0/4294967296.0,1,-nbitq), 
to_sfixed(1418554918.0/4294967296.0,1,-nbitq), 
to_sfixed(289661517.0/4294967296.0,1,-nbitq), 
to_sfixed(1399565102.0/4294967296.0,1,-nbitq), 
to_sfixed(1709297498.0/4294967296.0,1,-nbitq), 
to_sfixed(-166605249.0/4294967296.0,1,-nbitq), 
to_sfixed(-2038448483.0/4294967296.0,1,-nbitq), 
to_sfixed(402688311.0/4294967296.0,1,-nbitq), 
to_sfixed(-117265773.0/4294967296.0,1,-nbitq), 
to_sfixed(383638325.0/4294967296.0,1,-nbitq), 
to_sfixed(-1570147380.0/4294967296.0,1,-nbitq), 
to_sfixed(152574629.0/4294967296.0,1,-nbitq), 
to_sfixed(513567231.0/4294967296.0,1,-nbitq), 
to_sfixed(-169732949.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-136423698.0/4294967296.0,1,-nbitq), 
to_sfixed(804787603.0/4294967296.0,1,-nbitq), 
to_sfixed(-1452518646.0/4294967296.0,1,-nbitq), 
to_sfixed(123692180.0/4294967296.0,1,-nbitq), 
to_sfixed(-452639465.0/4294967296.0,1,-nbitq), 
to_sfixed(1433205642.0/4294967296.0,1,-nbitq), 
to_sfixed(-536958101.0/4294967296.0,1,-nbitq), 
to_sfixed(363284589.0/4294967296.0,1,-nbitq), 
to_sfixed(-942745281.0/4294967296.0,1,-nbitq), 
to_sfixed(-9494683.0/4294967296.0,1,-nbitq), 
to_sfixed(-480431117.0/4294967296.0,1,-nbitq), 
to_sfixed(1377364679.0/4294967296.0,1,-nbitq), 
to_sfixed(887347598.0/4294967296.0,1,-nbitq), 
to_sfixed(-1326772434.0/4294967296.0,1,-nbitq), 
to_sfixed(-78066653.0/4294967296.0,1,-nbitq), 
to_sfixed(243137081.0/4294967296.0,1,-nbitq), 
to_sfixed(32596399.0/4294967296.0,1,-nbitq), 
to_sfixed(287633932.0/4294967296.0,1,-nbitq), 
to_sfixed(-2059507100.0/4294967296.0,1,-nbitq), 
to_sfixed(-994387398.0/4294967296.0,1,-nbitq), 
to_sfixed(297253153.0/4294967296.0,1,-nbitq), 
to_sfixed(338271164.0/4294967296.0,1,-nbitq), 
to_sfixed(283414794.0/4294967296.0,1,-nbitq), 
to_sfixed(-1621723134.0/4294967296.0,1,-nbitq), 
to_sfixed(61252161.0/4294967296.0,1,-nbitq), 
to_sfixed(157711929.0/4294967296.0,1,-nbitq), 
to_sfixed(-814430927.0/4294967296.0,1,-nbitq), 
to_sfixed(-392325571.0/4294967296.0,1,-nbitq), 
to_sfixed(-190414857.0/4294967296.0,1,-nbitq), 
to_sfixed(1552184185.0/4294967296.0,1,-nbitq), 
to_sfixed(-3224363757.0/4294967296.0,1,-nbitq), 
to_sfixed(-181383107.0/4294967296.0,1,-nbitq), 
to_sfixed(-296830275.0/4294967296.0,1,-nbitq), 
to_sfixed(82750492.0/4294967296.0,1,-nbitq), 
to_sfixed(-62677178.0/4294967296.0,1,-nbitq), 
to_sfixed(-1167905852.0/4294967296.0,1,-nbitq), 
to_sfixed(389621901.0/4294967296.0,1,-nbitq), 
to_sfixed(-688703171.0/4294967296.0,1,-nbitq), 
to_sfixed(227918485.0/4294967296.0,1,-nbitq), 
to_sfixed(405137726.0/4294967296.0,1,-nbitq), 
to_sfixed(566331023.0/4294967296.0,1,-nbitq), 
to_sfixed(847778424.0/4294967296.0,1,-nbitq), 
to_sfixed(-155772107.0/4294967296.0,1,-nbitq), 
to_sfixed(-755403773.0/4294967296.0,1,-nbitq), 
to_sfixed(-759429283.0/4294967296.0,1,-nbitq), 
to_sfixed(-1661365452.0/4294967296.0,1,-nbitq), 
to_sfixed(267607478.0/4294967296.0,1,-nbitq), 
to_sfixed(219360157.0/4294967296.0,1,-nbitq), 
to_sfixed(-811979362.0/4294967296.0,1,-nbitq), 
to_sfixed(1068751121.0/4294967296.0,1,-nbitq), 
to_sfixed(-817675602.0/4294967296.0,1,-nbitq), 
to_sfixed(148652729.0/4294967296.0,1,-nbitq), 
to_sfixed(894297426.0/4294967296.0,1,-nbitq), 
to_sfixed(283595482.0/4294967296.0,1,-nbitq), 
to_sfixed(-1049590729.0/4294967296.0,1,-nbitq), 
to_sfixed(-1340355505.0/4294967296.0,1,-nbitq), 
to_sfixed(-544422059.0/4294967296.0,1,-nbitq), 
to_sfixed(181877472.0/4294967296.0,1,-nbitq), 
to_sfixed(337929640.0/4294967296.0,1,-nbitq), 
to_sfixed(426303858.0/4294967296.0,1,-nbitq), 
to_sfixed(177613131.0/4294967296.0,1,-nbitq), 
to_sfixed(-705079706.0/4294967296.0,1,-nbitq), 
to_sfixed(956241887.0/4294967296.0,1,-nbitq), 
to_sfixed(276735604.0/4294967296.0,1,-nbitq), 
to_sfixed(-325446686.0/4294967296.0,1,-nbitq), 
to_sfixed(385645829.0/4294967296.0,1,-nbitq), 
to_sfixed(-793793727.0/4294967296.0,1,-nbitq), 
to_sfixed(384628834.0/4294967296.0,1,-nbitq), 
to_sfixed(-136756128.0/4294967296.0,1,-nbitq), 
to_sfixed(830364224.0/4294967296.0,1,-nbitq), 
to_sfixed(514690800.0/4294967296.0,1,-nbitq), 
to_sfixed(-251915877.0/4294967296.0,1,-nbitq), 
to_sfixed(-1161348859.0/4294967296.0,1,-nbitq), 
to_sfixed(152918421.0/4294967296.0,1,-nbitq), 
to_sfixed(223848141.0/4294967296.0,1,-nbitq), 
to_sfixed(-234099225.0/4294967296.0,1,-nbitq), 
to_sfixed(-2475634518.0/4294967296.0,1,-nbitq), 
to_sfixed(453472041.0/4294967296.0,1,-nbitq), 
to_sfixed(301843369.0/4294967296.0,1,-nbitq), 
to_sfixed(262637222.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-401299768.0/4294967296.0,1,-nbitq), 
to_sfixed(1681142505.0/4294967296.0,1,-nbitq), 
to_sfixed(-1728617986.0/4294967296.0,1,-nbitq), 
to_sfixed(765362245.0/4294967296.0,1,-nbitq), 
to_sfixed(-1039983592.0/4294967296.0,1,-nbitq), 
to_sfixed(1056545538.0/4294967296.0,1,-nbitq), 
to_sfixed(224883350.0/4294967296.0,1,-nbitq), 
to_sfixed(727419851.0/4294967296.0,1,-nbitq), 
to_sfixed(-795497932.0/4294967296.0,1,-nbitq), 
to_sfixed(76704065.0/4294967296.0,1,-nbitq), 
to_sfixed(-416256516.0/4294967296.0,1,-nbitq), 
to_sfixed(668244923.0/4294967296.0,1,-nbitq), 
to_sfixed(851283173.0/4294967296.0,1,-nbitq), 
to_sfixed(-2062666490.0/4294967296.0,1,-nbitq), 
to_sfixed(-194966185.0/4294967296.0,1,-nbitq), 
to_sfixed(-257118700.0/4294967296.0,1,-nbitq), 
to_sfixed(98968240.0/4294967296.0,1,-nbitq), 
to_sfixed(236307190.0/4294967296.0,1,-nbitq), 
to_sfixed(-1454536043.0/4294967296.0,1,-nbitq), 
to_sfixed(16572959.0/4294967296.0,1,-nbitq), 
to_sfixed(22948975.0/4294967296.0,1,-nbitq), 
to_sfixed(692808861.0/4294967296.0,1,-nbitq), 
to_sfixed(649078902.0/4294967296.0,1,-nbitq), 
to_sfixed(-716908731.0/4294967296.0,1,-nbitq), 
to_sfixed(345424960.0/4294967296.0,1,-nbitq), 
to_sfixed(1425353425.0/4294967296.0,1,-nbitq), 
to_sfixed(-284172741.0/4294967296.0,1,-nbitq), 
to_sfixed(-646815386.0/4294967296.0,1,-nbitq), 
to_sfixed(-444889737.0/4294967296.0,1,-nbitq), 
to_sfixed(1434097781.0/4294967296.0,1,-nbitq), 
to_sfixed(-958729599.0/4294967296.0,1,-nbitq), 
to_sfixed(1806143291.0/4294967296.0,1,-nbitq), 
to_sfixed(-8257568.0/4294967296.0,1,-nbitq), 
to_sfixed(-497451365.0/4294967296.0,1,-nbitq), 
to_sfixed(-799824485.0/4294967296.0,1,-nbitq), 
to_sfixed(-885134743.0/4294967296.0,1,-nbitq), 
to_sfixed(-389075341.0/4294967296.0,1,-nbitq), 
to_sfixed(-915195468.0/4294967296.0,1,-nbitq), 
to_sfixed(299051283.0/4294967296.0,1,-nbitq), 
to_sfixed(123493198.0/4294967296.0,1,-nbitq), 
to_sfixed(-119015280.0/4294967296.0,1,-nbitq), 
to_sfixed(69901998.0/4294967296.0,1,-nbitq), 
to_sfixed(-961801226.0/4294967296.0,1,-nbitq), 
to_sfixed(-934656340.0/4294967296.0,1,-nbitq), 
to_sfixed(-669301600.0/4294967296.0,1,-nbitq), 
to_sfixed(-1329274996.0/4294967296.0,1,-nbitq), 
to_sfixed(226904336.0/4294967296.0,1,-nbitq), 
to_sfixed(764221150.0/4294967296.0,1,-nbitq), 
to_sfixed(-336802574.0/4294967296.0,1,-nbitq), 
to_sfixed(907197920.0/4294967296.0,1,-nbitq), 
to_sfixed(-100014797.0/4294967296.0,1,-nbitq), 
to_sfixed(-447284674.0/4294967296.0,1,-nbitq), 
to_sfixed(330573429.0/4294967296.0,1,-nbitq), 
to_sfixed(705373435.0/4294967296.0,1,-nbitq), 
to_sfixed(-1266119377.0/4294967296.0,1,-nbitq), 
to_sfixed(-1191914105.0/4294967296.0,1,-nbitq), 
to_sfixed(311363937.0/4294967296.0,1,-nbitq), 
to_sfixed(-233840777.0/4294967296.0,1,-nbitq), 
to_sfixed(-236863538.0/4294967296.0,1,-nbitq), 
to_sfixed(-306557321.0/4294967296.0,1,-nbitq), 
to_sfixed(-317410754.0/4294967296.0,1,-nbitq), 
to_sfixed(-650264302.0/4294967296.0,1,-nbitq), 
to_sfixed(528611028.0/4294967296.0,1,-nbitq), 
to_sfixed(324121015.0/4294967296.0,1,-nbitq), 
to_sfixed(-129671511.0/4294967296.0,1,-nbitq), 
to_sfixed(258488866.0/4294967296.0,1,-nbitq), 
to_sfixed(-2297131464.0/4294967296.0,1,-nbitq), 
to_sfixed(-452282310.0/4294967296.0,1,-nbitq), 
to_sfixed(385061993.0/4294967296.0,1,-nbitq), 
to_sfixed(649147659.0/4294967296.0,1,-nbitq), 
to_sfixed(433537135.0/4294967296.0,1,-nbitq), 
to_sfixed(-3082719.0/4294967296.0,1,-nbitq), 
to_sfixed(-752585001.0/4294967296.0,1,-nbitq), 
to_sfixed(-45589414.0/4294967296.0,1,-nbitq), 
to_sfixed(261466473.0/4294967296.0,1,-nbitq), 
to_sfixed(426203940.0/4294967296.0,1,-nbitq), 
to_sfixed(-1425774849.0/4294967296.0,1,-nbitq), 
to_sfixed(594639528.0/4294967296.0,1,-nbitq), 
to_sfixed(-41909779.0/4294967296.0,1,-nbitq), 
to_sfixed(-73207890.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-288784036.0/4294967296.0,1,-nbitq), 
to_sfixed(1567315244.0/4294967296.0,1,-nbitq), 
to_sfixed(-1187320602.0/4294967296.0,1,-nbitq), 
to_sfixed(1380321240.0/4294967296.0,1,-nbitq), 
to_sfixed(-1929390113.0/4294967296.0,1,-nbitq), 
to_sfixed(1187332702.0/4294967296.0,1,-nbitq), 
to_sfixed(196403565.0/4294967296.0,1,-nbitq), 
to_sfixed(-463921564.0/4294967296.0,1,-nbitq), 
to_sfixed(-774519505.0/4294967296.0,1,-nbitq), 
to_sfixed(-337823370.0/4294967296.0,1,-nbitq), 
to_sfixed(-16026653.0/4294967296.0,1,-nbitq), 
to_sfixed(-187119802.0/4294967296.0,1,-nbitq), 
to_sfixed(1018058763.0/4294967296.0,1,-nbitq), 
to_sfixed(-2683566949.0/4294967296.0,1,-nbitq), 
to_sfixed(62277716.0/4294967296.0,1,-nbitq), 
to_sfixed(-653934700.0/4294967296.0,1,-nbitq), 
to_sfixed(-47183355.0/4294967296.0,1,-nbitq), 
to_sfixed(-99358662.0/4294967296.0,1,-nbitq), 
to_sfixed(-1406665747.0/4294967296.0,1,-nbitq), 
to_sfixed(-245749491.0/4294967296.0,1,-nbitq), 
to_sfixed(161309736.0/4294967296.0,1,-nbitq), 
to_sfixed(327739434.0/4294967296.0,1,-nbitq), 
to_sfixed(-245514011.0/4294967296.0,1,-nbitq), 
to_sfixed(-1651335293.0/4294967296.0,1,-nbitq), 
to_sfixed(-333293149.0/4294967296.0,1,-nbitq), 
to_sfixed(1304186554.0/4294967296.0,1,-nbitq), 
to_sfixed(-470273808.0/4294967296.0,1,-nbitq), 
to_sfixed(-574026212.0/4294967296.0,1,-nbitq), 
to_sfixed(-389083853.0/4294967296.0,1,-nbitq), 
to_sfixed(1509894875.0/4294967296.0,1,-nbitq), 
to_sfixed(-835004260.0/4294967296.0,1,-nbitq), 
to_sfixed(1945470165.0/4294967296.0,1,-nbitq), 
to_sfixed(207559499.0/4294967296.0,1,-nbitq), 
to_sfixed(-119887948.0/4294967296.0,1,-nbitq), 
to_sfixed(-93938252.0/4294967296.0,1,-nbitq), 
to_sfixed(-1180869296.0/4294967296.0,1,-nbitq), 
to_sfixed(-867575127.0/4294967296.0,1,-nbitq), 
to_sfixed(-615096139.0/4294967296.0,1,-nbitq), 
to_sfixed(-34040712.0/4294967296.0,1,-nbitq), 
to_sfixed(-145919875.0/4294967296.0,1,-nbitq), 
to_sfixed(-645682650.0/4294967296.0,1,-nbitq), 
to_sfixed(359983067.0/4294967296.0,1,-nbitq), 
to_sfixed(-1328742260.0/4294967296.0,1,-nbitq), 
to_sfixed(-1399312511.0/4294967296.0,1,-nbitq), 
to_sfixed(-785094419.0/4294967296.0,1,-nbitq), 
to_sfixed(-1793875136.0/4294967296.0,1,-nbitq), 
to_sfixed(8982686.0/4294967296.0,1,-nbitq), 
to_sfixed(1152667393.0/4294967296.0,1,-nbitq), 
to_sfixed(-513983826.0/4294967296.0,1,-nbitq), 
to_sfixed(1706101896.0/4294967296.0,1,-nbitq), 
to_sfixed(-144077536.0/4294967296.0,1,-nbitq), 
to_sfixed(-300935062.0/4294967296.0,1,-nbitq), 
to_sfixed(1244553128.0/4294967296.0,1,-nbitq), 
to_sfixed(-148214041.0/4294967296.0,1,-nbitq), 
to_sfixed(-958969739.0/4294967296.0,1,-nbitq), 
to_sfixed(-800954588.0/4294967296.0,1,-nbitq), 
to_sfixed(2734980.0/4294967296.0,1,-nbitq), 
to_sfixed(470687365.0/4294967296.0,1,-nbitq), 
to_sfixed(-267070131.0/4294967296.0,1,-nbitq), 
to_sfixed(294154025.0/4294967296.0,1,-nbitq), 
to_sfixed(-445866978.0/4294967296.0,1,-nbitq), 
to_sfixed(825541166.0/4294967296.0,1,-nbitq), 
to_sfixed(282928415.0/4294967296.0,1,-nbitq), 
to_sfixed(847802305.0/4294967296.0,1,-nbitq), 
to_sfixed(157604924.0/4294967296.0,1,-nbitq), 
to_sfixed(255902943.0/4294967296.0,1,-nbitq), 
to_sfixed(-2013619387.0/4294967296.0,1,-nbitq), 
to_sfixed(-383101271.0/4294967296.0,1,-nbitq), 
to_sfixed(204796694.0/4294967296.0,1,-nbitq), 
to_sfixed(1207752294.0/4294967296.0,1,-nbitq), 
to_sfixed(490594055.0/4294967296.0,1,-nbitq), 
to_sfixed(-689709193.0/4294967296.0,1,-nbitq), 
to_sfixed(-719780188.0/4294967296.0,1,-nbitq), 
to_sfixed(400204511.0/4294967296.0,1,-nbitq), 
to_sfixed(-33934187.0/4294967296.0,1,-nbitq), 
to_sfixed(163178335.0/4294967296.0,1,-nbitq), 
to_sfixed(-970852435.0/4294967296.0,1,-nbitq), 
to_sfixed(173994644.0/4294967296.0,1,-nbitq), 
to_sfixed(-569275109.0/4294967296.0,1,-nbitq), 
to_sfixed(290289172.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-403245634.0/4294967296.0,1,-nbitq), 
to_sfixed(585543135.0/4294967296.0,1,-nbitq), 
to_sfixed(-384452516.0/4294967296.0,1,-nbitq), 
to_sfixed(998180562.0/4294967296.0,1,-nbitq), 
to_sfixed(-2348658256.0/4294967296.0,1,-nbitq), 
to_sfixed(290812014.0/4294967296.0,1,-nbitq), 
to_sfixed(-188724300.0/4294967296.0,1,-nbitq), 
to_sfixed(-413988479.0/4294967296.0,1,-nbitq), 
to_sfixed(-703984650.0/4294967296.0,1,-nbitq), 
to_sfixed(168298371.0/4294967296.0,1,-nbitq), 
to_sfixed(182575827.0/4294967296.0,1,-nbitq), 
to_sfixed(267152509.0/4294967296.0,1,-nbitq), 
to_sfixed(151997429.0/4294967296.0,1,-nbitq), 
to_sfixed(-1585594261.0/4294967296.0,1,-nbitq), 
to_sfixed(-164801851.0/4294967296.0,1,-nbitq), 
to_sfixed(-72632186.0/4294967296.0,1,-nbitq), 
to_sfixed(-296882297.0/4294967296.0,1,-nbitq), 
to_sfixed(-96059786.0/4294967296.0,1,-nbitq), 
to_sfixed(-823599161.0/4294967296.0,1,-nbitq), 
to_sfixed(-423481723.0/4294967296.0,1,-nbitq), 
to_sfixed(-332854631.0/4294967296.0,1,-nbitq), 
to_sfixed(61944523.0/4294967296.0,1,-nbitq), 
to_sfixed(-1866793813.0/4294967296.0,1,-nbitq), 
to_sfixed(-1117026450.0/4294967296.0,1,-nbitq), 
to_sfixed(-145625857.0/4294967296.0,1,-nbitq), 
to_sfixed(653572876.0/4294967296.0,1,-nbitq), 
to_sfixed(-654614364.0/4294967296.0,1,-nbitq), 
to_sfixed(624720442.0/4294967296.0,1,-nbitq), 
to_sfixed(-657285411.0/4294967296.0,1,-nbitq), 
to_sfixed(1206484235.0/4294967296.0,1,-nbitq), 
to_sfixed(-417264376.0/4294967296.0,1,-nbitq), 
to_sfixed(1607385973.0/4294967296.0,1,-nbitq), 
to_sfixed(-40032986.0/4294967296.0,1,-nbitq), 
to_sfixed(8410078.0/4294967296.0,1,-nbitq), 
to_sfixed(77672453.0/4294967296.0,1,-nbitq), 
to_sfixed(-280563125.0/4294967296.0,1,-nbitq), 
to_sfixed(-1416700993.0/4294967296.0,1,-nbitq), 
to_sfixed(-274283843.0/4294967296.0,1,-nbitq), 
to_sfixed(312226559.0/4294967296.0,1,-nbitq), 
to_sfixed(329055125.0/4294967296.0,1,-nbitq), 
to_sfixed(-432660437.0/4294967296.0,1,-nbitq), 
to_sfixed(224093587.0/4294967296.0,1,-nbitq), 
to_sfixed(-796474663.0/4294967296.0,1,-nbitq), 
to_sfixed(-1197101724.0/4294967296.0,1,-nbitq), 
to_sfixed(-504604700.0/4294967296.0,1,-nbitq), 
to_sfixed(-912819745.0/4294967296.0,1,-nbitq), 
to_sfixed(247145610.0/4294967296.0,1,-nbitq), 
to_sfixed(1411888285.0/4294967296.0,1,-nbitq), 
to_sfixed(-219871454.0/4294967296.0,1,-nbitq), 
to_sfixed(869578623.0/4294967296.0,1,-nbitq), 
to_sfixed(-25967668.0/4294967296.0,1,-nbitq), 
to_sfixed(-425864151.0/4294967296.0,1,-nbitq), 
to_sfixed(1302077865.0/4294967296.0,1,-nbitq), 
to_sfixed(530729995.0/4294967296.0,1,-nbitq), 
to_sfixed(-965689908.0/4294967296.0,1,-nbitq), 
to_sfixed(128423748.0/4294967296.0,1,-nbitq), 
to_sfixed(515303854.0/4294967296.0,1,-nbitq), 
to_sfixed(208859194.0/4294967296.0,1,-nbitq), 
to_sfixed(387899723.0/4294967296.0,1,-nbitq), 
to_sfixed(-316882522.0/4294967296.0,1,-nbitq), 
to_sfixed(-89667971.0/4294967296.0,1,-nbitq), 
to_sfixed(1080300254.0/4294967296.0,1,-nbitq), 
to_sfixed(475586355.0/4294967296.0,1,-nbitq), 
to_sfixed(57192395.0/4294967296.0,1,-nbitq), 
to_sfixed(122051912.0/4294967296.0,1,-nbitq), 
to_sfixed(31042066.0/4294967296.0,1,-nbitq), 
to_sfixed(-876957281.0/4294967296.0,1,-nbitq), 
to_sfixed(-245289223.0/4294967296.0,1,-nbitq), 
to_sfixed(-261285783.0/4294967296.0,1,-nbitq), 
to_sfixed(463593455.0/4294967296.0,1,-nbitq), 
to_sfixed(692452935.0/4294967296.0,1,-nbitq), 
to_sfixed(153515354.0/4294967296.0,1,-nbitq), 
to_sfixed(-617279267.0/4294967296.0,1,-nbitq), 
to_sfixed(-262767343.0/4294967296.0,1,-nbitq), 
to_sfixed(-108702529.0/4294967296.0,1,-nbitq), 
to_sfixed(925975478.0/4294967296.0,1,-nbitq), 
to_sfixed(-578008250.0/4294967296.0,1,-nbitq), 
to_sfixed(266587795.0/4294967296.0,1,-nbitq), 
to_sfixed(-272097921.0/4294967296.0,1,-nbitq), 
to_sfixed(-42187278.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(129938964.0/4294967296.0,1,-nbitq), 
to_sfixed(660586343.0/4294967296.0,1,-nbitq), 
to_sfixed(-1884630530.0/4294967296.0,1,-nbitq), 
to_sfixed(591370556.0/4294967296.0,1,-nbitq), 
to_sfixed(-1735690216.0/4294967296.0,1,-nbitq), 
to_sfixed(-222534437.0/4294967296.0,1,-nbitq), 
to_sfixed(-203571502.0/4294967296.0,1,-nbitq), 
to_sfixed(3261633.0/4294967296.0,1,-nbitq), 
to_sfixed(-1761458010.0/4294967296.0,1,-nbitq), 
to_sfixed(-223123371.0/4294967296.0,1,-nbitq), 
to_sfixed(-363893316.0/4294967296.0,1,-nbitq), 
to_sfixed(-201844184.0/4294967296.0,1,-nbitq), 
to_sfixed(-15192500.0/4294967296.0,1,-nbitq), 
to_sfixed(-579262369.0/4294967296.0,1,-nbitq), 
to_sfixed(-21446545.0/4294967296.0,1,-nbitq), 
to_sfixed(-16732157.0/4294967296.0,1,-nbitq), 
to_sfixed(45709881.0/4294967296.0,1,-nbitq), 
to_sfixed(-211778200.0/4294967296.0,1,-nbitq), 
to_sfixed(-420017607.0/4294967296.0,1,-nbitq), 
to_sfixed(-347165676.0/4294967296.0,1,-nbitq), 
to_sfixed(-314206947.0/4294967296.0,1,-nbitq), 
to_sfixed(-860646794.0/4294967296.0,1,-nbitq), 
to_sfixed(-2059670653.0/4294967296.0,1,-nbitq), 
to_sfixed(-1536683715.0/4294967296.0,1,-nbitq), 
to_sfixed(268803060.0/4294967296.0,1,-nbitq), 
to_sfixed(212434043.0/4294967296.0,1,-nbitq), 
to_sfixed(-302989219.0/4294967296.0,1,-nbitq), 
to_sfixed(1134565713.0/4294967296.0,1,-nbitq), 
to_sfixed(-830185233.0/4294967296.0,1,-nbitq), 
to_sfixed(1346031943.0/4294967296.0,1,-nbitq), 
to_sfixed(389321355.0/4294967296.0,1,-nbitq), 
to_sfixed(1196073455.0/4294967296.0,1,-nbitq), 
to_sfixed(-466413713.0/4294967296.0,1,-nbitq), 
to_sfixed(304977466.0/4294967296.0,1,-nbitq), 
to_sfixed(922836451.0/4294967296.0,1,-nbitq), 
to_sfixed(34677444.0/4294967296.0,1,-nbitq), 
to_sfixed(-1340200903.0/4294967296.0,1,-nbitq), 
to_sfixed(355257900.0/4294967296.0,1,-nbitq), 
to_sfixed(211191535.0/4294967296.0,1,-nbitq), 
to_sfixed(-58632428.0/4294967296.0,1,-nbitq), 
to_sfixed(69978571.0/4294967296.0,1,-nbitq), 
to_sfixed(105153773.0/4294967296.0,1,-nbitq), 
to_sfixed(-1751825390.0/4294967296.0,1,-nbitq), 
to_sfixed(-1545181169.0/4294967296.0,1,-nbitq), 
to_sfixed(-944493223.0/4294967296.0,1,-nbitq), 
to_sfixed(-1943484216.0/4294967296.0,1,-nbitq), 
to_sfixed(287955427.0/4294967296.0,1,-nbitq), 
to_sfixed(887782092.0/4294967296.0,1,-nbitq), 
to_sfixed(160548279.0/4294967296.0,1,-nbitq), 
to_sfixed(1056491385.0/4294967296.0,1,-nbitq), 
to_sfixed(124579148.0/4294967296.0,1,-nbitq), 
to_sfixed(-566689319.0/4294967296.0,1,-nbitq), 
to_sfixed(1003492161.0/4294967296.0,1,-nbitq), 
to_sfixed(-76600061.0/4294967296.0,1,-nbitq), 
to_sfixed(-1111367649.0/4294967296.0,1,-nbitq), 
to_sfixed(202983995.0/4294967296.0,1,-nbitq), 
to_sfixed(494723456.0/4294967296.0,1,-nbitq), 
to_sfixed(517200174.0/4294967296.0,1,-nbitq), 
to_sfixed(318202027.0/4294967296.0,1,-nbitq), 
to_sfixed(-123782070.0/4294967296.0,1,-nbitq), 
to_sfixed(-71444635.0/4294967296.0,1,-nbitq), 
to_sfixed(12584678.0/4294967296.0,1,-nbitq), 
to_sfixed(1031265564.0/4294967296.0,1,-nbitq), 
to_sfixed(524365123.0/4294967296.0,1,-nbitq), 
to_sfixed(55126225.0/4294967296.0,1,-nbitq), 
to_sfixed(467932577.0/4294967296.0,1,-nbitq), 
to_sfixed(-33623318.0/4294967296.0,1,-nbitq), 
to_sfixed(-979143906.0/4294967296.0,1,-nbitq), 
to_sfixed(129603652.0/4294967296.0,1,-nbitq), 
to_sfixed(648501812.0/4294967296.0,1,-nbitq), 
to_sfixed(345413857.0/4294967296.0,1,-nbitq), 
to_sfixed(193220340.0/4294967296.0,1,-nbitq), 
to_sfixed(42565856.0/4294967296.0,1,-nbitq), 
to_sfixed(-362555389.0/4294967296.0,1,-nbitq), 
to_sfixed(-199650658.0/4294967296.0,1,-nbitq), 
to_sfixed(545881053.0/4294967296.0,1,-nbitq), 
to_sfixed(-1344901966.0/4294967296.0,1,-nbitq), 
to_sfixed(-100570015.0/4294967296.0,1,-nbitq), 
to_sfixed(-159082000.0/4294967296.0,1,-nbitq), 
to_sfixed(-293732499.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(3491557.0/4294967296.0,1,-nbitq), 
to_sfixed(367238888.0/4294967296.0,1,-nbitq), 
to_sfixed(-773854580.0/4294967296.0,1,-nbitq), 
to_sfixed(776684414.0/4294967296.0,1,-nbitq), 
to_sfixed(-1535418223.0/4294967296.0,1,-nbitq), 
to_sfixed(-743111232.0/4294967296.0,1,-nbitq), 
to_sfixed(-60420869.0/4294967296.0,1,-nbitq), 
to_sfixed(131719924.0/4294967296.0,1,-nbitq), 
to_sfixed(-1166864346.0/4294967296.0,1,-nbitq), 
to_sfixed(-306702019.0/4294967296.0,1,-nbitq), 
to_sfixed(210294250.0/4294967296.0,1,-nbitq), 
to_sfixed(767410992.0/4294967296.0,1,-nbitq), 
to_sfixed(651461987.0/4294967296.0,1,-nbitq), 
to_sfixed(-1407616766.0/4294967296.0,1,-nbitq), 
to_sfixed(173429592.0/4294967296.0,1,-nbitq), 
to_sfixed(211582922.0/4294967296.0,1,-nbitq), 
to_sfixed(333716241.0/4294967296.0,1,-nbitq), 
to_sfixed(333012257.0/4294967296.0,1,-nbitq), 
to_sfixed(-253910612.0/4294967296.0,1,-nbitq), 
to_sfixed(243505673.0/4294967296.0,1,-nbitq), 
to_sfixed(-267121981.0/4294967296.0,1,-nbitq), 
to_sfixed(-489561459.0/4294967296.0,1,-nbitq), 
to_sfixed(-1840596904.0/4294967296.0,1,-nbitq), 
to_sfixed(-1290762272.0/4294967296.0,1,-nbitq), 
to_sfixed(-58163645.0/4294967296.0,1,-nbitq), 
to_sfixed(-797244261.0/4294967296.0,1,-nbitq), 
to_sfixed(-90273501.0/4294967296.0,1,-nbitq), 
to_sfixed(358294221.0/4294967296.0,1,-nbitq), 
to_sfixed(-529901519.0/4294967296.0,1,-nbitq), 
to_sfixed(1028074808.0/4294967296.0,1,-nbitq), 
to_sfixed(1895770772.0/4294967296.0,1,-nbitq), 
to_sfixed(840388609.0/4294967296.0,1,-nbitq), 
to_sfixed(405941003.0/4294967296.0,1,-nbitq), 
to_sfixed(731742297.0/4294967296.0,1,-nbitq), 
to_sfixed(-9523938.0/4294967296.0,1,-nbitq), 
to_sfixed(285248192.0/4294967296.0,1,-nbitq), 
to_sfixed(-246465060.0/4294967296.0,1,-nbitq), 
to_sfixed(230431887.0/4294967296.0,1,-nbitq), 
to_sfixed(-35305148.0/4294967296.0,1,-nbitq), 
to_sfixed(-164126593.0/4294967296.0,1,-nbitq), 
to_sfixed(-130742182.0/4294967296.0,1,-nbitq), 
to_sfixed(95675946.0/4294967296.0,1,-nbitq), 
to_sfixed(-1054664973.0/4294967296.0,1,-nbitq), 
to_sfixed(-1362923.0/4294967296.0,1,-nbitq), 
to_sfixed(-1312248587.0/4294967296.0,1,-nbitq), 
to_sfixed(-68120895.0/4294967296.0,1,-nbitq), 
to_sfixed(-42542324.0/4294967296.0,1,-nbitq), 
to_sfixed(802803467.0/4294967296.0,1,-nbitq), 
to_sfixed(416714980.0/4294967296.0,1,-nbitq), 
to_sfixed(-284693563.0/4294967296.0,1,-nbitq), 
to_sfixed(-124993392.0/4294967296.0,1,-nbitq), 
to_sfixed(-1041013939.0/4294967296.0,1,-nbitq), 
to_sfixed(1796026186.0/4294967296.0,1,-nbitq), 
to_sfixed(244490201.0/4294967296.0,1,-nbitq), 
to_sfixed(-606096367.0/4294967296.0,1,-nbitq), 
to_sfixed(-93358615.0/4294967296.0,1,-nbitq), 
to_sfixed(457014143.0/4294967296.0,1,-nbitq), 
to_sfixed(257612023.0/4294967296.0,1,-nbitq), 
to_sfixed(-275368935.0/4294967296.0,1,-nbitq), 
to_sfixed(168739213.0/4294967296.0,1,-nbitq), 
to_sfixed(23551034.0/4294967296.0,1,-nbitq), 
to_sfixed(-676159792.0/4294967296.0,1,-nbitq), 
to_sfixed(487883511.0/4294967296.0,1,-nbitq), 
to_sfixed(275977135.0/4294967296.0,1,-nbitq), 
to_sfixed(551806632.0/4294967296.0,1,-nbitq), 
to_sfixed(374385149.0/4294967296.0,1,-nbitq), 
to_sfixed(397817167.0/4294967296.0,1,-nbitq), 
to_sfixed(268159541.0/4294967296.0,1,-nbitq), 
to_sfixed(-196629120.0/4294967296.0,1,-nbitq), 
to_sfixed(255662635.0/4294967296.0,1,-nbitq), 
to_sfixed(682687240.0/4294967296.0,1,-nbitq), 
to_sfixed(251282086.0/4294967296.0,1,-nbitq), 
to_sfixed(-490159804.0/4294967296.0,1,-nbitq), 
to_sfixed(-106286592.0/4294967296.0,1,-nbitq), 
to_sfixed(152324242.0/4294967296.0,1,-nbitq), 
to_sfixed(493374317.0/4294967296.0,1,-nbitq), 
to_sfixed(-485309055.0/4294967296.0,1,-nbitq), 
to_sfixed(-21839909.0/4294967296.0,1,-nbitq), 
to_sfixed(47270377.0/4294967296.0,1,-nbitq), 
to_sfixed(209239297.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-209296811.0/4294967296.0,1,-nbitq), 
to_sfixed(385263618.0/4294967296.0,1,-nbitq), 
to_sfixed(-784585445.0/4294967296.0,1,-nbitq), 
to_sfixed(231839720.0/4294967296.0,1,-nbitq), 
to_sfixed(-1097678878.0/4294967296.0,1,-nbitq), 
to_sfixed(-906823094.0/4294967296.0,1,-nbitq), 
to_sfixed(296445958.0/4294967296.0,1,-nbitq), 
to_sfixed(918124834.0/4294967296.0,1,-nbitq), 
to_sfixed(-1077726318.0/4294967296.0,1,-nbitq), 
to_sfixed(33480827.0/4294967296.0,1,-nbitq), 
to_sfixed(412848314.0/4294967296.0,1,-nbitq), 
to_sfixed(-466705319.0/4294967296.0,1,-nbitq), 
to_sfixed(-60112903.0/4294967296.0,1,-nbitq), 
to_sfixed(-487359731.0/4294967296.0,1,-nbitq), 
to_sfixed(8128087.0/4294967296.0,1,-nbitq), 
to_sfixed(650760931.0/4294967296.0,1,-nbitq), 
to_sfixed(-426896763.0/4294967296.0,1,-nbitq), 
to_sfixed(-429966282.0/4294967296.0,1,-nbitq), 
to_sfixed(-110655335.0/4294967296.0,1,-nbitq), 
to_sfixed(-259094728.0/4294967296.0,1,-nbitq), 
to_sfixed(216614689.0/4294967296.0,1,-nbitq), 
to_sfixed(-390236102.0/4294967296.0,1,-nbitq), 
to_sfixed(-995526361.0/4294967296.0,1,-nbitq), 
to_sfixed(-611668025.0/4294967296.0,1,-nbitq), 
to_sfixed(-302672442.0/4294967296.0,1,-nbitq), 
to_sfixed(-1469761183.0/4294967296.0,1,-nbitq), 
to_sfixed(-24760543.0/4294967296.0,1,-nbitq), 
to_sfixed(456924880.0/4294967296.0,1,-nbitq), 
to_sfixed(69404391.0/4294967296.0,1,-nbitq), 
to_sfixed(650255941.0/4294967296.0,1,-nbitq), 
to_sfixed(228210490.0/4294967296.0,1,-nbitq), 
to_sfixed(669802862.0/4294967296.0,1,-nbitq), 
to_sfixed(311244647.0/4294967296.0,1,-nbitq), 
to_sfixed(933547938.0/4294967296.0,1,-nbitq), 
to_sfixed(-356110724.0/4294967296.0,1,-nbitq), 
to_sfixed(-77952134.0/4294967296.0,1,-nbitq), 
to_sfixed(-291455925.0/4294967296.0,1,-nbitq), 
to_sfixed(459804722.0/4294967296.0,1,-nbitq), 
to_sfixed(361048582.0/4294967296.0,1,-nbitq), 
to_sfixed(119799044.0/4294967296.0,1,-nbitq), 
to_sfixed(-550194040.0/4294967296.0,1,-nbitq), 
to_sfixed(-425775871.0/4294967296.0,1,-nbitq), 
to_sfixed(-710252569.0/4294967296.0,1,-nbitq), 
to_sfixed(-534264477.0/4294967296.0,1,-nbitq), 
to_sfixed(-1037557926.0/4294967296.0,1,-nbitq), 
to_sfixed(-750654066.0/4294967296.0,1,-nbitq), 
to_sfixed(305565842.0/4294967296.0,1,-nbitq), 
to_sfixed(829145798.0/4294967296.0,1,-nbitq), 
to_sfixed(-240368075.0/4294967296.0,1,-nbitq), 
to_sfixed(-538420269.0/4294967296.0,1,-nbitq), 
to_sfixed(435207349.0/4294967296.0,1,-nbitq), 
to_sfixed(-245319000.0/4294967296.0,1,-nbitq), 
to_sfixed(1117854108.0/4294967296.0,1,-nbitq), 
to_sfixed(-313620545.0/4294967296.0,1,-nbitq), 
to_sfixed(-783591145.0/4294967296.0,1,-nbitq), 
to_sfixed(141746134.0/4294967296.0,1,-nbitq), 
to_sfixed(734595783.0/4294967296.0,1,-nbitq), 
to_sfixed(431802029.0/4294967296.0,1,-nbitq), 
to_sfixed(-384711720.0/4294967296.0,1,-nbitq), 
to_sfixed(405078273.0/4294967296.0,1,-nbitq), 
to_sfixed(189523087.0/4294967296.0,1,-nbitq), 
to_sfixed(-672316856.0/4294967296.0,1,-nbitq), 
to_sfixed(247105695.0/4294967296.0,1,-nbitq), 
to_sfixed(-196645567.0/4294967296.0,1,-nbitq), 
to_sfixed(-235953031.0/4294967296.0,1,-nbitq), 
to_sfixed(-162326547.0/4294967296.0,1,-nbitq), 
to_sfixed(897652173.0/4294967296.0,1,-nbitq), 
to_sfixed(-561252662.0/4294967296.0,1,-nbitq), 
to_sfixed(-70515694.0/4294967296.0,1,-nbitq), 
to_sfixed(319576088.0/4294967296.0,1,-nbitq), 
to_sfixed(-41350870.0/4294967296.0,1,-nbitq), 
to_sfixed(319969463.0/4294967296.0,1,-nbitq), 
to_sfixed(-59895129.0/4294967296.0,1,-nbitq), 
to_sfixed(-147122127.0/4294967296.0,1,-nbitq), 
to_sfixed(439221521.0/4294967296.0,1,-nbitq), 
to_sfixed(544396139.0/4294967296.0,1,-nbitq), 
to_sfixed(-32379364.0/4294967296.0,1,-nbitq), 
to_sfixed(-293165165.0/4294967296.0,1,-nbitq), 
to_sfixed(-47802321.0/4294967296.0,1,-nbitq), 
to_sfixed(-88724218.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-149901187.0/4294967296.0,1,-nbitq), 
to_sfixed(692889389.0/4294967296.0,1,-nbitq), 
to_sfixed(-826604084.0/4294967296.0,1,-nbitq), 
to_sfixed(-716325277.0/4294967296.0,1,-nbitq), 
to_sfixed(-692018902.0/4294967296.0,1,-nbitq), 
to_sfixed(-336273971.0/4294967296.0,1,-nbitq), 
to_sfixed(115974478.0/4294967296.0,1,-nbitq), 
to_sfixed(910663361.0/4294967296.0,1,-nbitq), 
to_sfixed(-1083481353.0/4294967296.0,1,-nbitq), 
to_sfixed(225709144.0/4294967296.0,1,-nbitq), 
to_sfixed(416517741.0/4294967296.0,1,-nbitq), 
to_sfixed(-838781982.0/4294967296.0,1,-nbitq), 
to_sfixed(118144962.0/4294967296.0,1,-nbitq), 
to_sfixed(-385642096.0/4294967296.0,1,-nbitq), 
to_sfixed(46119418.0/4294967296.0,1,-nbitq), 
to_sfixed(-85652604.0/4294967296.0,1,-nbitq), 
to_sfixed(-250243232.0/4294967296.0,1,-nbitq), 
to_sfixed(-381246866.0/4294967296.0,1,-nbitq), 
to_sfixed(-237355773.0/4294967296.0,1,-nbitq), 
to_sfixed(-220621472.0/4294967296.0,1,-nbitq), 
to_sfixed(-283627099.0/4294967296.0,1,-nbitq), 
to_sfixed(-555675567.0/4294967296.0,1,-nbitq), 
to_sfixed(-957977556.0/4294967296.0,1,-nbitq), 
to_sfixed(-1038561195.0/4294967296.0,1,-nbitq), 
to_sfixed(415449794.0/4294967296.0,1,-nbitq), 
to_sfixed(-1398067950.0/4294967296.0,1,-nbitq), 
to_sfixed(509397316.0/4294967296.0,1,-nbitq), 
to_sfixed(352629660.0/4294967296.0,1,-nbitq), 
to_sfixed(-119297997.0/4294967296.0,1,-nbitq), 
to_sfixed(635101262.0/4294967296.0,1,-nbitq), 
to_sfixed(60438538.0/4294967296.0,1,-nbitq), 
to_sfixed(247783165.0/4294967296.0,1,-nbitq), 
to_sfixed(-151340809.0/4294967296.0,1,-nbitq), 
to_sfixed(97116361.0/4294967296.0,1,-nbitq), 
to_sfixed(-706260802.0/4294967296.0,1,-nbitq), 
to_sfixed(155695180.0/4294967296.0,1,-nbitq), 
to_sfixed(80240906.0/4294967296.0,1,-nbitq), 
to_sfixed(-46786753.0/4294967296.0,1,-nbitq), 
to_sfixed(260585872.0/4294967296.0,1,-nbitq), 
to_sfixed(232923348.0/4294967296.0,1,-nbitq), 
to_sfixed(433194244.0/4294967296.0,1,-nbitq), 
to_sfixed(-1263237620.0/4294967296.0,1,-nbitq), 
to_sfixed(-333247343.0/4294967296.0,1,-nbitq), 
to_sfixed(-1143547448.0/4294967296.0,1,-nbitq), 
to_sfixed(-463509040.0/4294967296.0,1,-nbitq), 
to_sfixed(-694527081.0/4294967296.0,1,-nbitq), 
to_sfixed(123640283.0/4294967296.0,1,-nbitq), 
to_sfixed(-442039183.0/4294967296.0,1,-nbitq), 
to_sfixed(-188263240.0/4294967296.0,1,-nbitq), 
to_sfixed(267715179.0/4294967296.0,1,-nbitq), 
to_sfixed(724341258.0/4294967296.0,1,-nbitq), 
to_sfixed(-345992000.0/4294967296.0,1,-nbitq), 
to_sfixed(831053683.0/4294967296.0,1,-nbitq), 
to_sfixed(-405319630.0/4294967296.0,1,-nbitq), 
to_sfixed(-705224449.0/4294967296.0,1,-nbitq), 
to_sfixed(-75852205.0/4294967296.0,1,-nbitq), 
to_sfixed(874458362.0/4294967296.0,1,-nbitq), 
to_sfixed(212557140.0/4294967296.0,1,-nbitq), 
to_sfixed(395898422.0/4294967296.0,1,-nbitq), 
to_sfixed(-272281528.0/4294967296.0,1,-nbitq), 
to_sfixed(138838730.0/4294967296.0,1,-nbitq), 
to_sfixed(-223140443.0/4294967296.0,1,-nbitq), 
to_sfixed(255227209.0/4294967296.0,1,-nbitq), 
to_sfixed(-40430248.0/4294967296.0,1,-nbitq), 
to_sfixed(-116168168.0/4294967296.0,1,-nbitq), 
to_sfixed(-241390789.0/4294967296.0,1,-nbitq), 
to_sfixed(-234521956.0/4294967296.0,1,-nbitq), 
to_sfixed(-185590315.0/4294967296.0,1,-nbitq), 
to_sfixed(364038906.0/4294967296.0,1,-nbitq), 
to_sfixed(289665443.0/4294967296.0,1,-nbitq), 
to_sfixed(-328743327.0/4294967296.0,1,-nbitq), 
to_sfixed(198260592.0/4294967296.0,1,-nbitq), 
to_sfixed(1028911425.0/4294967296.0,1,-nbitq), 
to_sfixed(392805233.0/4294967296.0,1,-nbitq), 
to_sfixed(167436850.0/4294967296.0,1,-nbitq), 
to_sfixed(-127156247.0/4294967296.0,1,-nbitq), 
to_sfixed(-848165934.0/4294967296.0,1,-nbitq), 
to_sfixed(-18661570.0/4294967296.0,1,-nbitq), 
to_sfixed(682606423.0/4294967296.0,1,-nbitq), 
to_sfixed(169167001.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(169073695.0/4294967296.0,1,-nbitq), 
to_sfixed(342847478.0/4294967296.0,1,-nbitq), 
to_sfixed(-142331682.0/4294967296.0,1,-nbitq), 
to_sfixed(-670167464.0/4294967296.0,1,-nbitq), 
to_sfixed(-95240515.0/4294967296.0,1,-nbitq), 
to_sfixed(-837494477.0/4294967296.0,1,-nbitq), 
to_sfixed(3105437.0/4294967296.0,1,-nbitq), 
to_sfixed(501435413.0/4294967296.0,1,-nbitq), 
to_sfixed(-807766212.0/4294967296.0,1,-nbitq), 
to_sfixed(91981237.0/4294967296.0,1,-nbitq), 
to_sfixed(540985472.0/4294967296.0,1,-nbitq), 
to_sfixed(-59815627.0/4294967296.0,1,-nbitq), 
to_sfixed(-253309619.0/4294967296.0,1,-nbitq), 
to_sfixed(-158278785.0/4294967296.0,1,-nbitq), 
to_sfixed(-190692801.0/4294967296.0,1,-nbitq), 
to_sfixed(186945822.0/4294967296.0,1,-nbitq), 
to_sfixed(-139737972.0/4294967296.0,1,-nbitq), 
to_sfixed(79692360.0/4294967296.0,1,-nbitq), 
to_sfixed(219558648.0/4294967296.0,1,-nbitq), 
to_sfixed(2944279.0/4294967296.0,1,-nbitq), 
to_sfixed(-329609574.0/4294967296.0,1,-nbitq), 
to_sfixed(25979308.0/4294967296.0,1,-nbitq), 
to_sfixed(-351113559.0/4294967296.0,1,-nbitq), 
to_sfixed(-405447042.0/4294967296.0,1,-nbitq), 
to_sfixed(-101648359.0/4294967296.0,1,-nbitq), 
to_sfixed(-880923050.0/4294967296.0,1,-nbitq), 
to_sfixed(822392578.0/4294967296.0,1,-nbitq), 
to_sfixed(322538872.0/4294967296.0,1,-nbitq), 
to_sfixed(20991530.0/4294967296.0,1,-nbitq), 
to_sfixed(291850316.0/4294967296.0,1,-nbitq), 
to_sfixed(-451506662.0/4294967296.0,1,-nbitq), 
to_sfixed(-195864488.0/4294967296.0,1,-nbitq), 
to_sfixed(-11048440.0/4294967296.0,1,-nbitq), 
to_sfixed(-16315441.0/4294967296.0,1,-nbitq), 
to_sfixed(-189964024.0/4294967296.0,1,-nbitq), 
to_sfixed(-37345785.0/4294967296.0,1,-nbitq), 
to_sfixed(-448094307.0/4294967296.0,1,-nbitq), 
to_sfixed(-89560490.0/4294967296.0,1,-nbitq), 
to_sfixed(-270409557.0/4294967296.0,1,-nbitq), 
to_sfixed(76766222.0/4294967296.0,1,-nbitq), 
to_sfixed(-43748544.0/4294967296.0,1,-nbitq), 
to_sfixed(-107774141.0/4294967296.0,1,-nbitq), 
to_sfixed(-478525504.0/4294967296.0,1,-nbitq), 
to_sfixed(-1191547123.0/4294967296.0,1,-nbitq), 
to_sfixed(-834256392.0/4294967296.0,1,-nbitq), 
to_sfixed(-547954683.0/4294967296.0,1,-nbitq), 
to_sfixed(-400388668.0/4294967296.0,1,-nbitq), 
to_sfixed(46163683.0/4294967296.0,1,-nbitq), 
to_sfixed(-433589198.0/4294967296.0,1,-nbitq), 
to_sfixed(-113697512.0/4294967296.0,1,-nbitq), 
to_sfixed(-37731621.0/4294967296.0,1,-nbitq), 
to_sfixed(241025758.0/4294967296.0,1,-nbitq), 
to_sfixed(925854245.0/4294967296.0,1,-nbitq), 
to_sfixed(-655933681.0/4294967296.0,1,-nbitq), 
to_sfixed(-370795173.0/4294967296.0,1,-nbitq), 
to_sfixed(856043.0/4294967296.0,1,-nbitq), 
to_sfixed(482130201.0/4294967296.0,1,-nbitq), 
to_sfixed(613043135.0/4294967296.0,1,-nbitq), 
to_sfixed(100433208.0/4294967296.0,1,-nbitq), 
to_sfixed(-283063007.0/4294967296.0,1,-nbitq), 
to_sfixed(-104503758.0/4294967296.0,1,-nbitq), 
to_sfixed(-291412202.0/4294967296.0,1,-nbitq), 
to_sfixed(196071099.0/4294967296.0,1,-nbitq), 
to_sfixed(64711436.0/4294967296.0,1,-nbitq), 
to_sfixed(4345029.0/4294967296.0,1,-nbitq), 
to_sfixed(199179032.0/4294967296.0,1,-nbitq), 
to_sfixed(716274806.0/4294967296.0,1,-nbitq), 
to_sfixed(268184959.0/4294967296.0,1,-nbitq), 
to_sfixed(-206263631.0/4294967296.0,1,-nbitq), 
to_sfixed(333419799.0/4294967296.0,1,-nbitq), 
to_sfixed(-141656041.0/4294967296.0,1,-nbitq), 
to_sfixed(-423735072.0/4294967296.0,1,-nbitq), 
to_sfixed(898011036.0/4294967296.0,1,-nbitq), 
to_sfixed(124321052.0/4294967296.0,1,-nbitq), 
to_sfixed(225537581.0/4294967296.0,1,-nbitq), 
to_sfixed(-102276408.0/4294967296.0,1,-nbitq), 
to_sfixed(-696930181.0/4294967296.0,1,-nbitq), 
to_sfixed(-310361880.0/4294967296.0,1,-nbitq), 
to_sfixed(514577044.0/4294967296.0,1,-nbitq), 
to_sfixed(378036105.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-437697.0/4294967296.0,1,-nbitq), 
to_sfixed(37619110.0/4294967296.0,1,-nbitq), 
to_sfixed(-48865524.0/4294967296.0,1,-nbitq), 
to_sfixed(-713058796.0/4294967296.0,1,-nbitq), 
to_sfixed(109053923.0/4294967296.0,1,-nbitq), 
to_sfixed(-817469140.0/4294967296.0,1,-nbitq), 
to_sfixed(338809905.0/4294967296.0,1,-nbitq), 
to_sfixed(-25631086.0/4294967296.0,1,-nbitq), 
to_sfixed(115479492.0/4294967296.0,1,-nbitq), 
to_sfixed(-80174262.0/4294967296.0,1,-nbitq), 
to_sfixed(546875875.0/4294967296.0,1,-nbitq), 
to_sfixed(-377369690.0/4294967296.0,1,-nbitq), 
to_sfixed(74064157.0/4294967296.0,1,-nbitq), 
to_sfixed(-68563274.0/4294967296.0,1,-nbitq), 
to_sfixed(360952098.0/4294967296.0,1,-nbitq), 
to_sfixed(328001438.0/4294967296.0,1,-nbitq), 
to_sfixed(203809533.0/4294967296.0,1,-nbitq), 
to_sfixed(312088832.0/4294967296.0,1,-nbitq), 
to_sfixed(174947820.0/4294967296.0,1,-nbitq), 
to_sfixed(-237403445.0/4294967296.0,1,-nbitq), 
to_sfixed(16352205.0/4294967296.0,1,-nbitq), 
to_sfixed(-155206461.0/4294967296.0,1,-nbitq), 
to_sfixed(-209050495.0/4294967296.0,1,-nbitq), 
to_sfixed(-139878136.0/4294967296.0,1,-nbitq), 
to_sfixed(58603397.0/4294967296.0,1,-nbitq), 
to_sfixed(-470022361.0/4294967296.0,1,-nbitq), 
to_sfixed(499350080.0/4294967296.0,1,-nbitq), 
to_sfixed(-360082783.0/4294967296.0,1,-nbitq), 
to_sfixed(484014368.0/4294967296.0,1,-nbitq), 
to_sfixed(528288727.0/4294967296.0,1,-nbitq), 
to_sfixed(-598233218.0/4294967296.0,1,-nbitq), 
to_sfixed(44795964.0/4294967296.0,1,-nbitq), 
to_sfixed(-15592325.0/4294967296.0,1,-nbitq), 
to_sfixed(143008353.0/4294967296.0,1,-nbitq), 
to_sfixed(-645395766.0/4294967296.0,1,-nbitq), 
to_sfixed(-581791304.0/4294967296.0,1,-nbitq), 
to_sfixed(-71234721.0/4294967296.0,1,-nbitq), 
to_sfixed(212491549.0/4294967296.0,1,-nbitq), 
to_sfixed(-181335662.0/4294967296.0,1,-nbitq), 
to_sfixed(17933710.0/4294967296.0,1,-nbitq), 
to_sfixed(-44698299.0/4294967296.0,1,-nbitq), 
to_sfixed(-299419413.0/4294967296.0,1,-nbitq), 
to_sfixed(166870787.0/4294967296.0,1,-nbitq), 
to_sfixed(-895511621.0/4294967296.0,1,-nbitq), 
to_sfixed(-60478231.0/4294967296.0,1,-nbitq), 
to_sfixed(-186918856.0/4294967296.0,1,-nbitq), 
to_sfixed(39032801.0/4294967296.0,1,-nbitq), 
to_sfixed(-224390354.0/4294967296.0,1,-nbitq), 
to_sfixed(-44309840.0/4294967296.0,1,-nbitq), 
to_sfixed(378530359.0/4294967296.0,1,-nbitq), 
to_sfixed(467967813.0/4294967296.0,1,-nbitq), 
to_sfixed(-239743368.0/4294967296.0,1,-nbitq), 
to_sfixed(83699794.0/4294967296.0,1,-nbitq), 
to_sfixed(97513196.0/4294967296.0,1,-nbitq), 
to_sfixed(-23698692.0/4294967296.0,1,-nbitq), 
to_sfixed(-369162007.0/4294967296.0,1,-nbitq), 
to_sfixed(-197698961.0/4294967296.0,1,-nbitq), 
to_sfixed(-131787247.0/4294967296.0,1,-nbitq), 
to_sfixed(373442133.0/4294967296.0,1,-nbitq), 
to_sfixed(310246147.0/4294967296.0,1,-nbitq), 
to_sfixed(-11359497.0/4294967296.0,1,-nbitq), 
to_sfixed(270631081.0/4294967296.0,1,-nbitq), 
to_sfixed(-233914777.0/4294967296.0,1,-nbitq), 
to_sfixed(-186045519.0/4294967296.0,1,-nbitq), 
to_sfixed(205076749.0/4294967296.0,1,-nbitq), 
to_sfixed(241226424.0/4294967296.0,1,-nbitq), 
to_sfixed(204888442.0/4294967296.0,1,-nbitq), 
to_sfixed(-110575091.0/4294967296.0,1,-nbitq), 
to_sfixed(69150374.0/4294967296.0,1,-nbitq), 
to_sfixed(-41209821.0/4294967296.0,1,-nbitq), 
to_sfixed(-482816325.0/4294967296.0,1,-nbitq), 
to_sfixed(-457844885.0/4294967296.0,1,-nbitq), 
to_sfixed(182113939.0/4294967296.0,1,-nbitq), 
to_sfixed(272650264.0/4294967296.0,1,-nbitq), 
to_sfixed(462021740.0/4294967296.0,1,-nbitq), 
to_sfixed(-78739672.0/4294967296.0,1,-nbitq), 
to_sfixed(-409758248.0/4294967296.0,1,-nbitq), 
to_sfixed(-22587447.0/4294967296.0,1,-nbitq), 
to_sfixed(413688645.0/4294967296.0,1,-nbitq), 
to_sfixed(-256614209.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(242271983.0/4294967296.0,1,-nbitq), 
to_sfixed(-192454131.0/4294967296.0,1,-nbitq), 
to_sfixed(661673430.0/4294967296.0,1,-nbitq), 
to_sfixed(-342310625.0/4294967296.0,1,-nbitq), 
to_sfixed(60665341.0/4294967296.0,1,-nbitq), 
to_sfixed(-97495039.0/4294967296.0,1,-nbitq), 
to_sfixed(-257285434.0/4294967296.0,1,-nbitq), 
to_sfixed(-186815180.0/4294967296.0,1,-nbitq), 
to_sfixed(-338904088.0/4294967296.0,1,-nbitq), 
to_sfixed(368850805.0/4294967296.0,1,-nbitq), 
to_sfixed(15509583.0/4294967296.0,1,-nbitq), 
to_sfixed(-410588571.0/4294967296.0,1,-nbitq), 
to_sfixed(397994332.0/4294967296.0,1,-nbitq), 
to_sfixed(256619302.0/4294967296.0,1,-nbitq), 
to_sfixed(-189911522.0/4294967296.0,1,-nbitq), 
to_sfixed(287520484.0/4294967296.0,1,-nbitq), 
to_sfixed(-301187455.0/4294967296.0,1,-nbitq), 
to_sfixed(295129061.0/4294967296.0,1,-nbitq), 
to_sfixed(-258581357.0/4294967296.0,1,-nbitq), 
to_sfixed(296541245.0/4294967296.0,1,-nbitq), 
to_sfixed(-217462602.0/4294967296.0,1,-nbitq), 
to_sfixed(-193235902.0/4294967296.0,1,-nbitq), 
to_sfixed(-366378420.0/4294967296.0,1,-nbitq), 
to_sfixed(-242857385.0/4294967296.0,1,-nbitq), 
to_sfixed(191725756.0/4294967296.0,1,-nbitq), 
to_sfixed(218792869.0/4294967296.0,1,-nbitq), 
to_sfixed(-10205197.0/4294967296.0,1,-nbitq), 
to_sfixed(-303275902.0/4294967296.0,1,-nbitq), 
to_sfixed(634135911.0/4294967296.0,1,-nbitq), 
to_sfixed(363783247.0/4294967296.0,1,-nbitq), 
to_sfixed(-430248556.0/4294967296.0,1,-nbitq), 
to_sfixed(111293276.0/4294967296.0,1,-nbitq), 
to_sfixed(19018117.0/4294967296.0,1,-nbitq), 
to_sfixed(39442872.0/4294967296.0,1,-nbitq), 
to_sfixed(-391769262.0/4294967296.0,1,-nbitq), 
to_sfixed(168193650.0/4294967296.0,1,-nbitq), 
to_sfixed(-261365569.0/4294967296.0,1,-nbitq), 
to_sfixed(185977601.0/4294967296.0,1,-nbitq), 
to_sfixed(196178046.0/4294967296.0,1,-nbitq), 
to_sfixed(330114140.0/4294967296.0,1,-nbitq), 
to_sfixed(-275991399.0/4294967296.0,1,-nbitq), 
to_sfixed(-167556950.0/4294967296.0,1,-nbitq), 
to_sfixed(-7463070.0/4294967296.0,1,-nbitq), 
to_sfixed(-92166837.0/4294967296.0,1,-nbitq), 
to_sfixed(-93698945.0/4294967296.0,1,-nbitq), 
to_sfixed(-532132245.0/4294967296.0,1,-nbitq), 
to_sfixed(-358448469.0/4294967296.0,1,-nbitq), 
to_sfixed(-495169669.0/4294967296.0,1,-nbitq), 
to_sfixed(29073695.0/4294967296.0,1,-nbitq), 
to_sfixed(-134096069.0/4294967296.0,1,-nbitq), 
to_sfixed(-339160350.0/4294967296.0,1,-nbitq), 
to_sfixed(231832621.0/4294967296.0,1,-nbitq), 
to_sfixed(-138753692.0/4294967296.0,1,-nbitq), 
to_sfixed(-122644086.0/4294967296.0,1,-nbitq), 
to_sfixed(91793653.0/4294967296.0,1,-nbitq), 
to_sfixed(-275050949.0/4294967296.0,1,-nbitq), 
to_sfixed(137309839.0/4294967296.0,1,-nbitq), 
to_sfixed(298325124.0/4294967296.0,1,-nbitq), 
to_sfixed(-81193873.0/4294967296.0,1,-nbitq), 
to_sfixed(217427320.0/4294967296.0,1,-nbitq), 
to_sfixed(120642289.0/4294967296.0,1,-nbitq), 
to_sfixed(-406100156.0/4294967296.0,1,-nbitq), 
to_sfixed(-205555794.0/4294967296.0,1,-nbitq), 
to_sfixed(-352432054.0/4294967296.0,1,-nbitq), 
to_sfixed(-317059133.0/4294967296.0,1,-nbitq), 
to_sfixed(-29018303.0/4294967296.0,1,-nbitq), 
to_sfixed(145392708.0/4294967296.0,1,-nbitq), 
to_sfixed(331864363.0/4294967296.0,1,-nbitq), 
to_sfixed(-155497900.0/4294967296.0,1,-nbitq), 
to_sfixed(-128486300.0/4294967296.0,1,-nbitq), 
to_sfixed(45857083.0/4294967296.0,1,-nbitq), 
to_sfixed(128551775.0/4294967296.0,1,-nbitq), 
to_sfixed(-67364941.0/4294967296.0,1,-nbitq), 
to_sfixed(352083577.0/4294967296.0,1,-nbitq), 
to_sfixed(202417116.0/4294967296.0,1,-nbitq), 
to_sfixed(-474176708.0/4294967296.0,1,-nbitq), 
to_sfixed(-374698539.0/4294967296.0,1,-nbitq), 
to_sfixed(274879637.0/4294967296.0,1,-nbitq), 
to_sfixed(-305863145.0/4294967296.0,1,-nbitq), 
to_sfixed(-219003546.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(247860966.0/4294967296.0,1,-nbitq), 
to_sfixed(-169075555.0/4294967296.0,1,-nbitq), 
to_sfixed(193350628.0/4294967296.0,1,-nbitq), 
to_sfixed(32686791.0/4294967296.0,1,-nbitq), 
to_sfixed(166439563.0/4294967296.0,1,-nbitq), 
to_sfixed(-489113819.0/4294967296.0,1,-nbitq), 
to_sfixed(72059873.0/4294967296.0,1,-nbitq), 
to_sfixed(-54792679.0/4294967296.0,1,-nbitq), 
to_sfixed(169326661.0/4294967296.0,1,-nbitq), 
to_sfixed(-92623519.0/4294967296.0,1,-nbitq), 
to_sfixed(213234171.0/4294967296.0,1,-nbitq), 
to_sfixed(-251798702.0/4294967296.0,1,-nbitq), 
to_sfixed(145576652.0/4294967296.0,1,-nbitq), 
to_sfixed(387255725.0/4294967296.0,1,-nbitq), 
to_sfixed(-306706892.0/4294967296.0,1,-nbitq), 
to_sfixed(277671194.0/4294967296.0,1,-nbitq), 
to_sfixed(-391773760.0/4294967296.0,1,-nbitq), 
to_sfixed(-94073019.0/4294967296.0,1,-nbitq), 
to_sfixed(427638965.0/4294967296.0,1,-nbitq), 
to_sfixed(-99777382.0/4294967296.0,1,-nbitq), 
to_sfixed(-121436018.0/4294967296.0,1,-nbitq), 
to_sfixed(-105995363.0/4294967296.0,1,-nbitq), 
to_sfixed(-32207694.0/4294967296.0,1,-nbitq), 
to_sfixed(139396547.0/4294967296.0,1,-nbitq), 
to_sfixed(270355954.0/4294967296.0,1,-nbitq), 
to_sfixed(209498078.0/4294967296.0,1,-nbitq), 
to_sfixed(136290005.0/4294967296.0,1,-nbitq), 
to_sfixed(-96673754.0/4294967296.0,1,-nbitq), 
to_sfixed(374027954.0/4294967296.0,1,-nbitq), 
to_sfixed(23788680.0/4294967296.0,1,-nbitq), 
to_sfixed(-367781745.0/4294967296.0,1,-nbitq), 
to_sfixed(-83110306.0/4294967296.0,1,-nbitq), 
to_sfixed(40267108.0/4294967296.0,1,-nbitq), 
to_sfixed(-525761461.0/4294967296.0,1,-nbitq), 
to_sfixed(186506569.0/4294967296.0,1,-nbitq), 
to_sfixed(291888616.0/4294967296.0,1,-nbitq), 
to_sfixed(146142696.0/4294967296.0,1,-nbitq), 
to_sfixed(-5869623.0/4294967296.0,1,-nbitq), 
to_sfixed(1818999.0/4294967296.0,1,-nbitq), 
to_sfixed(62158095.0/4294967296.0,1,-nbitq), 
to_sfixed(-402461776.0/4294967296.0,1,-nbitq), 
to_sfixed(-150006459.0/4294967296.0,1,-nbitq), 
to_sfixed(-294202440.0/4294967296.0,1,-nbitq), 
to_sfixed(-143760154.0/4294967296.0,1,-nbitq), 
to_sfixed(149837579.0/4294967296.0,1,-nbitq), 
to_sfixed(-337620308.0/4294967296.0,1,-nbitq), 
to_sfixed(-252681353.0/4294967296.0,1,-nbitq), 
to_sfixed(-80105277.0/4294967296.0,1,-nbitq), 
to_sfixed(-127322367.0/4294967296.0,1,-nbitq), 
to_sfixed(56794614.0/4294967296.0,1,-nbitq), 
to_sfixed(-301520842.0/4294967296.0,1,-nbitq), 
to_sfixed(23217196.0/4294967296.0,1,-nbitq), 
to_sfixed(8670985.0/4294967296.0,1,-nbitq), 
to_sfixed(11839664.0/4294967296.0,1,-nbitq), 
to_sfixed(475913796.0/4294967296.0,1,-nbitq), 
to_sfixed(-202598553.0/4294967296.0,1,-nbitq), 
to_sfixed(188860213.0/4294967296.0,1,-nbitq), 
to_sfixed(-338976367.0/4294967296.0,1,-nbitq), 
to_sfixed(384590082.0/4294967296.0,1,-nbitq), 
to_sfixed(84070770.0/4294967296.0,1,-nbitq), 
to_sfixed(-183993849.0/4294967296.0,1,-nbitq), 
to_sfixed(139788612.0/4294967296.0,1,-nbitq), 
to_sfixed(-38330495.0/4294967296.0,1,-nbitq), 
to_sfixed(-172442672.0/4294967296.0,1,-nbitq), 
to_sfixed(323187566.0/4294967296.0,1,-nbitq), 
to_sfixed(327284005.0/4294967296.0,1,-nbitq), 
to_sfixed(550014382.0/4294967296.0,1,-nbitq), 
to_sfixed(-136750533.0/4294967296.0,1,-nbitq), 
to_sfixed(42195240.0/4294967296.0,1,-nbitq), 
to_sfixed(381837245.0/4294967296.0,1,-nbitq), 
to_sfixed(319431835.0/4294967296.0,1,-nbitq), 
to_sfixed(-187202118.0/4294967296.0,1,-nbitq), 
to_sfixed(66865397.0/4294967296.0,1,-nbitq), 
to_sfixed(337674187.0/4294967296.0,1,-nbitq), 
to_sfixed(453327082.0/4294967296.0,1,-nbitq), 
to_sfixed(-340448380.0/4294967296.0,1,-nbitq), 
to_sfixed(129030923.0/4294967296.0,1,-nbitq), 
to_sfixed(-309258160.0/4294967296.0,1,-nbitq), 
to_sfixed(-55295420.0/4294967296.0,1,-nbitq), 
to_sfixed(-144640447.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(333881853.0/4294967296.0,1,-nbitq), 
to_sfixed(210957711.0/4294967296.0,1,-nbitq), 
to_sfixed(379309183.0/4294967296.0,1,-nbitq), 
to_sfixed(-475172636.0/4294967296.0,1,-nbitq), 
to_sfixed(84014859.0/4294967296.0,1,-nbitq), 
to_sfixed(-301430696.0/4294967296.0,1,-nbitq), 
to_sfixed(152766303.0/4294967296.0,1,-nbitq), 
to_sfixed(251889548.0/4294967296.0,1,-nbitq), 
to_sfixed(229618873.0/4294967296.0,1,-nbitq), 
to_sfixed(131622162.0/4294967296.0,1,-nbitq), 
to_sfixed(112030951.0/4294967296.0,1,-nbitq), 
to_sfixed(-68315648.0/4294967296.0,1,-nbitq), 
to_sfixed(434793162.0/4294967296.0,1,-nbitq), 
to_sfixed(371970614.0/4294967296.0,1,-nbitq), 
to_sfixed(-24389228.0/4294967296.0,1,-nbitq), 
to_sfixed(404769987.0/4294967296.0,1,-nbitq), 
to_sfixed(316634718.0/4294967296.0,1,-nbitq), 
to_sfixed(276211974.0/4294967296.0,1,-nbitq), 
to_sfixed(14129858.0/4294967296.0,1,-nbitq), 
to_sfixed(267402416.0/4294967296.0,1,-nbitq), 
to_sfixed(174159316.0/4294967296.0,1,-nbitq), 
to_sfixed(102264401.0/4294967296.0,1,-nbitq), 
to_sfixed(-302215837.0/4294967296.0,1,-nbitq), 
to_sfixed(382020819.0/4294967296.0,1,-nbitq), 
to_sfixed(-124762428.0/4294967296.0,1,-nbitq), 
to_sfixed(-15841222.0/4294967296.0,1,-nbitq), 
to_sfixed(400227587.0/4294967296.0,1,-nbitq), 
to_sfixed(-118861528.0/4294967296.0,1,-nbitq), 
to_sfixed(284597905.0/4294967296.0,1,-nbitq), 
to_sfixed(-336776399.0/4294967296.0,1,-nbitq), 
to_sfixed(185855165.0/4294967296.0,1,-nbitq), 
to_sfixed(-476292691.0/4294967296.0,1,-nbitq), 
to_sfixed(-267480964.0/4294967296.0,1,-nbitq), 
to_sfixed(-139681684.0/4294967296.0,1,-nbitq), 
to_sfixed(355158596.0/4294967296.0,1,-nbitq), 
to_sfixed(129114152.0/4294967296.0,1,-nbitq), 
to_sfixed(378164856.0/4294967296.0,1,-nbitq), 
to_sfixed(-354883736.0/4294967296.0,1,-nbitq), 
to_sfixed(296252117.0/4294967296.0,1,-nbitq), 
to_sfixed(-100293266.0/4294967296.0,1,-nbitq), 
to_sfixed(-135364944.0/4294967296.0,1,-nbitq), 
to_sfixed(268064003.0/4294967296.0,1,-nbitq), 
to_sfixed(-278266410.0/4294967296.0,1,-nbitq), 
to_sfixed(124618377.0/4294967296.0,1,-nbitq), 
to_sfixed(223471010.0/4294967296.0,1,-nbitq), 
to_sfixed(-160947583.0/4294967296.0,1,-nbitq), 
to_sfixed(237993757.0/4294967296.0,1,-nbitq), 
to_sfixed(-307336239.0/4294967296.0,1,-nbitq), 
to_sfixed(-428034106.0/4294967296.0,1,-nbitq), 
to_sfixed(-210559486.0/4294967296.0,1,-nbitq), 
to_sfixed(-347516562.0/4294967296.0,1,-nbitq), 
to_sfixed(203406844.0/4294967296.0,1,-nbitq), 
to_sfixed(-4785948.0/4294967296.0,1,-nbitq), 
to_sfixed(411648542.0/4294967296.0,1,-nbitq), 
to_sfixed(180957893.0/4294967296.0,1,-nbitq), 
to_sfixed(-431187883.0/4294967296.0,1,-nbitq), 
to_sfixed(-337556044.0/4294967296.0,1,-nbitq), 
to_sfixed(-443191185.0/4294967296.0,1,-nbitq), 
to_sfixed(-326791392.0/4294967296.0,1,-nbitq), 
to_sfixed(-109989261.0/4294967296.0,1,-nbitq), 
to_sfixed(-114448350.0/4294967296.0,1,-nbitq), 
to_sfixed(-46605894.0/4294967296.0,1,-nbitq), 
to_sfixed(-327299261.0/4294967296.0,1,-nbitq), 
to_sfixed(289359869.0/4294967296.0,1,-nbitq), 
to_sfixed(372973934.0/4294967296.0,1,-nbitq), 
to_sfixed(-241201601.0/4294967296.0,1,-nbitq), 
to_sfixed(356374123.0/4294967296.0,1,-nbitq), 
to_sfixed(-127233862.0/4294967296.0,1,-nbitq), 
to_sfixed(-4657247.0/4294967296.0,1,-nbitq), 
to_sfixed(173509383.0/4294967296.0,1,-nbitq), 
to_sfixed(19487956.0/4294967296.0,1,-nbitq), 
to_sfixed(-87524345.0/4294967296.0,1,-nbitq), 
to_sfixed(260608592.0/4294967296.0,1,-nbitq), 
to_sfixed(-336885540.0/4294967296.0,1,-nbitq), 
to_sfixed(512186158.0/4294967296.0,1,-nbitq), 
to_sfixed(-109593040.0/4294967296.0,1,-nbitq), 
to_sfixed(-259244394.0/4294967296.0,1,-nbitq), 
to_sfixed(-329083475.0/4294967296.0,1,-nbitq), 
to_sfixed(219394478.0/4294967296.0,1,-nbitq), 
to_sfixed(354155579.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-54713305.0/4294967296.0,1,-nbitq), 
to_sfixed(199338943.0/4294967296.0,1,-nbitq), 
to_sfixed(523273112.0/4294967296.0,1,-nbitq), 
to_sfixed(-626563534.0/4294967296.0,1,-nbitq), 
to_sfixed(315699894.0/4294967296.0,1,-nbitq), 
to_sfixed(-547642109.0/4294967296.0,1,-nbitq), 
to_sfixed(373836396.0/4294967296.0,1,-nbitq), 
to_sfixed(8536422.0/4294967296.0,1,-nbitq), 
to_sfixed(103880132.0/4294967296.0,1,-nbitq), 
to_sfixed(-85606236.0/4294967296.0,1,-nbitq), 
to_sfixed(-477124368.0/4294967296.0,1,-nbitq), 
to_sfixed(-96891171.0/4294967296.0,1,-nbitq), 
to_sfixed(318615107.0/4294967296.0,1,-nbitq), 
to_sfixed(201905758.0/4294967296.0,1,-nbitq), 
to_sfixed(314955540.0/4294967296.0,1,-nbitq), 
to_sfixed(-107840460.0/4294967296.0,1,-nbitq), 
to_sfixed(-147737305.0/4294967296.0,1,-nbitq), 
to_sfixed(-151234493.0/4294967296.0,1,-nbitq), 
to_sfixed(190231011.0/4294967296.0,1,-nbitq), 
to_sfixed(-56989089.0/4294967296.0,1,-nbitq), 
to_sfixed(211523243.0/4294967296.0,1,-nbitq), 
to_sfixed(-244252556.0/4294967296.0,1,-nbitq), 
to_sfixed(223701160.0/4294967296.0,1,-nbitq), 
to_sfixed(120076702.0/4294967296.0,1,-nbitq), 
to_sfixed(-56181784.0/4294967296.0,1,-nbitq), 
to_sfixed(-356088841.0/4294967296.0,1,-nbitq), 
to_sfixed(-37962174.0/4294967296.0,1,-nbitq), 
to_sfixed(-520489696.0/4294967296.0,1,-nbitq), 
to_sfixed(154157311.0/4294967296.0,1,-nbitq), 
to_sfixed(326305509.0/4294967296.0,1,-nbitq), 
to_sfixed(-507545449.0/4294967296.0,1,-nbitq), 
to_sfixed(493712547.0/4294967296.0,1,-nbitq), 
to_sfixed(-297040829.0/4294967296.0,1,-nbitq), 
to_sfixed(-110816805.0/4294967296.0,1,-nbitq), 
to_sfixed(-177779755.0/4294967296.0,1,-nbitq), 
to_sfixed(-298685453.0/4294967296.0,1,-nbitq), 
to_sfixed(-445060584.0/4294967296.0,1,-nbitq), 
to_sfixed(-274769733.0/4294967296.0,1,-nbitq), 
to_sfixed(-486889571.0/4294967296.0,1,-nbitq), 
to_sfixed(199528684.0/4294967296.0,1,-nbitq), 
to_sfixed(-180311294.0/4294967296.0,1,-nbitq), 
to_sfixed(257906868.0/4294967296.0,1,-nbitq), 
to_sfixed(-103304029.0/4294967296.0,1,-nbitq), 
to_sfixed(-77204683.0/4294967296.0,1,-nbitq), 
to_sfixed(-24337945.0/4294967296.0,1,-nbitq), 
to_sfixed(408080274.0/4294967296.0,1,-nbitq), 
to_sfixed(241295155.0/4294967296.0,1,-nbitq), 
to_sfixed(-601987692.0/4294967296.0,1,-nbitq), 
to_sfixed(162558653.0/4294967296.0,1,-nbitq), 
to_sfixed(-61147205.0/4294967296.0,1,-nbitq), 
to_sfixed(-96949315.0/4294967296.0,1,-nbitq), 
to_sfixed(-194460790.0/4294967296.0,1,-nbitq), 
to_sfixed(-363649001.0/4294967296.0,1,-nbitq), 
to_sfixed(121831879.0/4294967296.0,1,-nbitq), 
to_sfixed(-25187920.0/4294967296.0,1,-nbitq), 
to_sfixed(-102598648.0/4294967296.0,1,-nbitq), 
to_sfixed(402467204.0/4294967296.0,1,-nbitq), 
to_sfixed(-279915485.0/4294967296.0,1,-nbitq), 
to_sfixed(-267299998.0/4294967296.0,1,-nbitq), 
to_sfixed(-265926556.0/4294967296.0,1,-nbitq), 
to_sfixed(22305593.0/4294967296.0,1,-nbitq), 
to_sfixed(394689384.0/4294967296.0,1,-nbitq), 
to_sfixed(-297456230.0/4294967296.0,1,-nbitq), 
to_sfixed(204595101.0/4294967296.0,1,-nbitq), 
to_sfixed(-49610319.0/4294967296.0,1,-nbitq), 
to_sfixed(-54140273.0/4294967296.0,1,-nbitq), 
to_sfixed(678512592.0/4294967296.0,1,-nbitq), 
to_sfixed(293235314.0/4294967296.0,1,-nbitq), 
to_sfixed(-111961917.0/4294967296.0,1,-nbitq), 
to_sfixed(170996302.0/4294967296.0,1,-nbitq), 
to_sfixed(84567043.0/4294967296.0,1,-nbitq), 
to_sfixed(-76086666.0/4294967296.0,1,-nbitq), 
to_sfixed(-398344339.0/4294967296.0,1,-nbitq), 
to_sfixed(381054711.0/4294967296.0,1,-nbitq), 
to_sfixed(-186498681.0/4294967296.0,1,-nbitq), 
to_sfixed(-307887419.0/4294967296.0,1,-nbitq), 
to_sfixed(-491684106.0/4294967296.0,1,-nbitq), 
to_sfixed(-431516016.0/4294967296.0,1,-nbitq), 
to_sfixed(267212596.0/4294967296.0,1,-nbitq), 
to_sfixed(-6997684.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-375304116.0/4294967296.0,1,-nbitq), 
to_sfixed(-507703815.0/4294967296.0,1,-nbitq), 
to_sfixed(520196801.0/4294967296.0,1,-nbitq), 
to_sfixed(-1158910114.0/4294967296.0,1,-nbitq), 
to_sfixed(-524679200.0/4294967296.0,1,-nbitq), 
to_sfixed(-351765062.0/4294967296.0,1,-nbitq), 
to_sfixed(245428887.0/4294967296.0,1,-nbitq), 
to_sfixed(-18600020.0/4294967296.0,1,-nbitq), 
to_sfixed(-338267297.0/4294967296.0,1,-nbitq), 
to_sfixed(-110998163.0/4294967296.0,1,-nbitq), 
to_sfixed(132783824.0/4294967296.0,1,-nbitq), 
to_sfixed(-73316268.0/4294967296.0,1,-nbitq), 
to_sfixed(747863320.0/4294967296.0,1,-nbitq), 
to_sfixed(524049633.0/4294967296.0,1,-nbitq), 
to_sfixed(272310797.0/4294967296.0,1,-nbitq), 
to_sfixed(646957245.0/4294967296.0,1,-nbitq), 
to_sfixed(57190151.0/4294967296.0,1,-nbitq), 
to_sfixed(370176497.0/4294967296.0,1,-nbitq), 
to_sfixed(-349051713.0/4294967296.0,1,-nbitq), 
to_sfixed(58138753.0/4294967296.0,1,-nbitq), 
to_sfixed(9071777.0/4294967296.0,1,-nbitq), 
to_sfixed(6240631.0/4294967296.0,1,-nbitq), 
to_sfixed(-514558914.0/4294967296.0,1,-nbitq), 
to_sfixed(98627547.0/4294967296.0,1,-nbitq), 
to_sfixed(-124989830.0/4294967296.0,1,-nbitq), 
to_sfixed(-458938903.0/4294967296.0,1,-nbitq), 
to_sfixed(287524007.0/4294967296.0,1,-nbitq), 
to_sfixed(-230439059.0/4294967296.0,1,-nbitq), 
to_sfixed(-63877506.0/4294967296.0,1,-nbitq), 
to_sfixed(511555554.0/4294967296.0,1,-nbitq), 
to_sfixed(266594329.0/4294967296.0,1,-nbitq), 
to_sfixed(432379663.0/4294967296.0,1,-nbitq), 
to_sfixed(-141832325.0/4294967296.0,1,-nbitq), 
to_sfixed(-54260146.0/4294967296.0,1,-nbitq), 
to_sfixed(-336726451.0/4294967296.0,1,-nbitq), 
to_sfixed(326088591.0/4294967296.0,1,-nbitq), 
to_sfixed(-112263338.0/4294967296.0,1,-nbitq), 
to_sfixed(155650505.0/4294967296.0,1,-nbitq), 
to_sfixed(180348176.0/4294967296.0,1,-nbitq), 
to_sfixed(-303334757.0/4294967296.0,1,-nbitq), 
to_sfixed(-529795773.0/4294967296.0,1,-nbitq), 
to_sfixed(-143993430.0/4294967296.0,1,-nbitq), 
to_sfixed(-463074020.0/4294967296.0,1,-nbitq), 
to_sfixed(-352859357.0/4294967296.0,1,-nbitq), 
to_sfixed(-542800514.0/4294967296.0,1,-nbitq), 
to_sfixed(-435616263.0/4294967296.0,1,-nbitq), 
to_sfixed(-92222803.0/4294967296.0,1,-nbitq), 
to_sfixed(-462810330.0/4294967296.0,1,-nbitq), 
to_sfixed(43456768.0/4294967296.0,1,-nbitq), 
to_sfixed(161146459.0/4294967296.0,1,-nbitq), 
to_sfixed(205947679.0/4294967296.0,1,-nbitq), 
to_sfixed(-128037914.0/4294967296.0,1,-nbitq), 
to_sfixed(-44611896.0/4294967296.0,1,-nbitq), 
to_sfixed(-151507445.0/4294967296.0,1,-nbitq), 
to_sfixed(326236708.0/4294967296.0,1,-nbitq), 
to_sfixed(-269090494.0/4294967296.0,1,-nbitq), 
to_sfixed(135081090.0/4294967296.0,1,-nbitq), 
to_sfixed(-206401986.0/4294967296.0,1,-nbitq), 
to_sfixed(93581479.0/4294967296.0,1,-nbitq), 
to_sfixed(-227876679.0/4294967296.0,1,-nbitq), 
to_sfixed(-296352584.0/4294967296.0,1,-nbitq), 
to_sfixed(104133284.0/4294967296.0,1,-nbitq), 
to_sfixed(394025860.0/4294967296.0,1,-nbitq), 
to_sfixed(-348429947.0/4294967296.0,1,-nbitq), 
to_sfixed(-300859347.0/4294967296.0,1,-nbitq), 
to_sfixed(212769989.0/4294967296.0,1,-nbitq), 
to_sfixed(57056202.0/4294967296.0,1,-nbitq), 
to_sfixed(265838575.0/4294967296.0,1,-nbitq), 
to_sfixed(96647115.0/4294967296.0,1,-nbitq), 
to_sfixed(872141762.0/4294967296.0,1,-nbitq), 
to_sfixed(689058171.0/4294967296.0,1,-nbitq), 
to_sfixed(123508625.0/4294967296.0,1,-nbitq), 
to_sfixed(-95644824.0/4294967296.0,1,-nbitq), 
to_sfixed(-280487774.0/4294967296.0,1,-nbitq), 
to_sfixed(469493320.0/4294967296.0,1,-nbitq), 
to_sfixed(61970593.0/4294967296.0,1,-nbitq), 
to_sfixed(-58166577.0/4294967296.0,1,-nbitq), 
to_sfixed(-504624366.0/4294967296.0,1,-nbitq), 
to_sfixed(95245290.0/4294967296.0,1,-nbitq), 
to_sfixed(-185815677.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(346429409.0/4294967296.0,1,-nbitq), 
to_sfixed(37965915.0/4294967296.0,1,-nbitq), 
to_sfixed(873023333.0/4294967296.0,1,-nbitq), 
to_sfixed(-1907527790.0/4294967296.0,1,-nbitq), 
to_sfixed(-1254514965.0/4294967296.0,1,-nbitq), 
to_sfixed(-113842939.0/4294967296.0,1,-nbitq), 
to_sfixed(-393238899.0/4294967296.0,1,-nbitq), 
to_sfixed(158569524.0/4294967296.0,1,-nbitq), 
to_sfixed(-435041087.0/4294967296.0,1,-nbitq), 
to_sfixed(116638741.0/4294967296.0,1,-nbitq), 
to_sfixed(-534099430.0/4294967296.0,1,-nbitq), 
to_sfixed(-676337339.0/4294967296.0,1,-nbitq), 
to_sfixed(1568052947.0/4294967296.0,1,-nbitq), 
to_sfixed(1156887438.0/4294967296.0,1,-nbitq), 
to_sfixed(127228477.0/4294967296.0,1,-nbitq), 
to_sfixed(942206762.0/4294967296.0,1,-nbitq), 
to_sfixed(-288820632.0/4294967296.0,1,-nbitq), 
to_sfixed(-313909663.0/4294967296.0,1,-nbitq), 
to_sfixed(-148272798.0/4294967296.0,1,-nbitq), 
to_sfixed(497173503.0/4294967296.0,1,-nbitq), 
to_sfixed(-407253501.0/4294967296.0,1,-nbitq), 
to_sfixed(-396175368.0/4294967296.0,1,-nbitq), 
to_sfixed(-1200981255.0/4294967296.0,1,-nbitq), 
to_sfixed(1063872812.0/4294967296.0,1,-nbitq), 
to_sfixed(-165882819.0/4294967296.0,1,-nbitq), 
to_sfixed(-759011035.0/4294967296.0,1,-nbitq), 
to_sfixed(319605381.0/4294967296.0,1,-nbitq), 
to_sfixed(283970886.0/4294967296.0,1,-nbitq), 
to_sfixed(398774389.0/4294967296.0,1,-nbitq), 
to_sfixed(1149236135.0/4294967296.0,1,-nbitq), 
to_sfixed(-168864443.0/4294967296.0,1,-nbitq), 
to_sfixed(-5753927.0/4294967296.0,1,-nbitq), 
to_sfixed(-886786502.0/4294967296.0,1,-nbitq), 
to_sfixed(779957376.0/4294967296.0,1,-nbitq), 
to_sfixed(118040007.0/4294967296.0,1,-nbitq), 
to_sfixed(464186631.0/4294967296.0,1,-nbitq), 
to_sfixed(34155041.0/4294967296.0,1,-nbitq), 
to_sfixed(-811293401.0/4294967296.0,1,-nbitq), 
to_sfixed(56330376.0/4294967296.0,1,-nbitq), 
to_sfixed(-268779754.0/4294967296.0,1,-nbitq), 
to_sfixed(-420705919.0/4294967296.0,1,-nbitq), 
to_sfixed(-514813025.0/4294967296.0,1,-nbitq), 
to_sfixed(-954019499.0/4294967296.0,1,-nbitq), 
to_sfixed(-42380540.0/4294967296.0,1,-nbitq), 
to_sfixed(-45984165.0/4294967296.0,1,-nbitq), 
to_sfixed(-343367998.0/4294967296.0,1,-nbitq), 
to_sfixed(237545839.0/4294967296.0,1,-nbitq), 
to_sfixed(297415063.0/4294967296.0,1,-nbitq), 
to_sfixed(-435662532.0/4294967296.0,1,-nbitq), 
to_sfixed(-214803181.0/4294967296.0,1,-nbitq), 
to_sfixed(239832599.0/4294967296.0,1,-nbitq), 
to_sfixed(-1096990476.0/4294967296.0,1,-nbitq), 
to_sfixed(-157331341.0/4294967296.0,1,-nbitq), 
to_sfixed(-528392738.0/4294967296.0,1,-nbitq), 
to_sfixed(404940988.0/4294967296.0,1,-nbitq), 
to_sfixed(-194721222.0/4294967296.0,1,-nbitq), 
to_sfixed(135180589.0/4294967296.0,1,-nbitq), 
to_sfixed(-908497089.0/4294967296.0,1,-nbitq), 
to_sfixed(225823053.0/4294967296.0,1,-nbitq), 
to_sfixed(50810995.0/4294967296.0,1,-nbitq), 
to_sfixed(282193516.0/4294967296.0,1,-nbitq), 
to_sfixed(-391431942.0/4294967296.0,1,-nbitq), 
to_sfixed(393150141.0/4294967296.0,1,-nbitq), 
to_sfixed(152842658.0/4294967296.0,1,-nbitq), 
to_sfixed(-212288882.0/4294967296.0,1,-nbitq), 
to_sfixed(317379182.0/4294967296.0,1,-nbitq), 
to_sfixed(216115883.0/4294967296.0,1,-nbitq), 
to_sfixed(121746056.0/4294967296.0,1,-nbitq), 
to_sfixed(453617255.0/4294967296.0,1,-nbitq), 
to_sfixed(487691183.0/4294967296.0,1,-nbitq), 
to_sfixed(996221716.0/4294967296.0,1,-nbitq), 
to_sfixed(149442264.0/4294967296.0,1,-nbitq), 
to_sfixed(167265381.0/4294967296.0,1,-nbitq), 
to_sfixed(200973047.0/4294967296.0,1,-nbitq), 
to_sfixed(527075357.0/4294967296.0,1,-nbitq), 
to_sfixed(107922389.0/4294967296.0,1,-nbitq), 
to_sfixed(-167510705.0/4294967296.0,1,-nbitq), 
to_sfixed(-404196848.0/4294967296.0,1,-nbitq), 
to_sfixed(973562354.0/4294967296.0,1,-nbitq), 
to_sfixed(321496121.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(347162397.0/4294967296.0,1,-nbitq), 
to_sfixed(392898595.0/4294967296.0,1,-nbitq), 
to_sfixed(907293814.0/4294967296.0,1,-nbitq), 
to_sfixed(-1956477397.0/4294967296.0,1,-nbitq), 
to_sfixed(-900279085.0/4294967296.0,1,-nbitq), 
to_sfixed(1185519573.0/4294967296.0,1,-nbitq), 
to_sfixed(-261891195.0/4294967296.0,1,-nbitq), 
to_sfixed(-184478530.0/4294967296.0,1,-nbitq), 
to_sfixed(-481655346.0/4294967296.0,1,-nbitq), 
to_sfixed(103886583.0/4294967296.0,1,-nbitq), 
to_sfixed(-10955564.0/4294967296.0,1,-nbitq), 
to_sfixed(-126497224.0/4294967296.0,1,-nbitq), 
to_sfixed(1045491084.0/4294967296.0,1,-nbitq), 
to_sfixed(1092157212.0/4294967296.0,1,-nbitq), 
to_sfixed(-85226205.0/4294967296.0,1,-nbitq), 
to_sfixed(1508580946.0/4294967296.0,1,-nbitq), 
to_sfixed(208179632.0/4294967296.0,1,-nbitq), 
to_sfixed(158496752.0/4294967296.0,1,-nbitq), 
to_sfixed(-1083227555.0/4294967296.0,1,-nbitq), 
to_sfixed(1188247661.0/4294967296.0,1,-nbitq), 
to_sfixed(81526560.0/4294967296.0,1,-nbitq), 
to_sfixed(-98467173.0/4294967296.0,1,-nbitq), 
to_sfixed(-1583332864.0/4294967296.0,1,-nbitq), 
to_sfixed(1169513297.0/4294967296.0,1,-nbitq), 
to_sfixed(229179328.0/4294967296.0,1,-nbitq), 
to_sfixed(-259141624.0/4294967296.0,1,-nbitq), 
to_sfixed(-196746641.0/4294967296.0,1,-nbitq), 
to_sfixed(-95342839.0/4294967296.0,1,-nbitq), 
to_sfixed(540170095.0/4294967296.0,1,-nbitq), 
to_sfixed(1047882017.0/4294967296.0,1,-nbitq), 
to_sfixed(-82847537.0/4294967296.0,1,-nbitq), 
to_sfixed(-414983787.0/4294967296.0,1,-nbitq), 
to_sfixed(-391632544.0/4294967296.0,1,-nbitq), 
to_sfixed(695895008.0/4294967296.0,1,-nbitq), 
to_sfixed(94348555.0/4294967296.0,1,-nbitq), 
to_sfixed(1002158082.0/4294967296.0,1,-nbitq), 
to_sfixed(-176915956.0/4294967296.0,1,-nbitq), 
to_sfixed(-1376591194.0/4294967296.0,1,-nbitq), 
to_sfixed(-246139819.0/4294967296.0,1,-nbitq), 
to_sfixed(-392452228.0/4294967296.0,1,-nbitq), 
to_sfixed(99622393.0/4294967296.0,1,-nbitq), 
to_sfixed(-292262718.0/4294967296.0,1,-nbitq), 
to_sfixed(190449155.0/4294967296.0,1,-nbitq), 
to_sfixed(482287263.0/4294967296.0,1,-nbitq), 
to_sfixed(-1033304927.0/4294967296.0,1,-nbitq), 
to_sfixed(25823999.0/4294967296.0,1,-nbitq), 
to_sfixed(-314375153.0/4294967296.0,1,-nbitq), 
to_sfixed(-61103803.0/4294967296.0,1,-nbitq), 
to_sfixed(287819287.0/4294967296.0,1,-nbitq), 
to_sfixed(429073912.0/4294967296.0,1,-nbitq), 
to_sfixed(-867942462.0/4294967296.0,1,-nbitq), 
to_sfixed(-1921881355.0/4294967296.0,1,-nbitq), 
to_sfixed(244485910.0/4294967296.0,1,-nbitq), 
to_sfixed(-819780829.0/4294967296.0,1,-nbitq), 
to_sfixed(-352216081.0/4294967296.0,1,-nbitq), 
to_sfixed(-1061989336.0/4294967296.0,1,-nbitq), 
to_sfixed(-343072064.0/4294967296.0,1,-nbitq), 
to_sfixed(-800890298.0/4294967296.0,1,-nbitq), 
to_sfixed(-279966161.0/4294967296.0,1,-nbitq), 
to_sfixed(182670254.0/4294967296.0,1,-nbitq), 
to_sfixed(-402079123.0/4294967296.0,1,-nbitq), 
to_sfixed(-100694534.0/4294967296.0,1,-nbitq), 
to_sfixed(607735801.0/4294967296.0,1,-nbitq), 
to_sfixed(-148631102.0/4294967296.0,1,-nbitq), 
to_sfixed(-653069.0/4294967296.0,1,-nbitq), 
to_sfixed(-84086794.0/4294967296.0,1,-nbitq), 
to_sfixed(572344995.0/4294967296.0,1,-nbitq), 
to_sfixed(1165340056.0/4294967296.0,1,-nbitq), 
to_sfixed(1489609.0/4294967296.0,1,-nbitq), 
to_sfixed(-106984450.0/4294967296.0,1,-nbitq), 
to_sfixed(633803041.0/4294967296.0,1,-nbitq), 
to_sfixed(-11457987.0/4294967296.0,1,-nbitq), 
to_sfixed(446567362.0/4294967296.0,1,-nbitq), 
to_sfixed(60784164.0/4294967296.0,1,-nbitq), 
to_sfixed(-78725297.0/4294967296.0,1,-nbitq), 
to_sfixed(64338458.0/4294967296.0,1,-nbitq), 
to_sfixed(-426814251.0/4294967296.0,1,-nbitq), 
to_sfixed(320186653.0/4294967296.0,1,-nbitq), 
to_sfixed(1137432863.0/4294967296.0,1,-nbitq), 
to_sfixed(165820164.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(159657358.0/4294967296.0,1,-nbitq), 
to_sfixed(-293184987.0/4294967296.0,1,-nbitq), 
to_sfixed(-954790759.0/4294967296.0,1,-nbitq), 
to_sfixed(-1134872217.0/4294967296.0,1,-nbitq), 
to_sfixed(-374034845.0/4294967296.0,1,-nbitq), 
to_sfixed(1976471222.0/4294967296.0,1,-nbitq), 
to_sfixed(-62955442.0/4294967296.0,1,-nbitq), 
to_sfixed(276872493.0/4294967296.0,1,-nbitq), 
to_sfixed(-476204205.0/4294967296.0,1,-nbitq), 
to_sfixed(198500831.0/4294967296.0,1,-nbitq), 
to_sfixed(-93316753.0/4294967296.0,1,-nbitq), 
to_sfixed(-482060006.0/4294967296.0,1,-nbitq), 
to_sfixed(357957078.0/4294967296.0,1,-nbitq), 
to_sfixed(950298952.0/4294967296.0,1,-nbitq), 
to_sfixed(399421171.0/4294967296.0,1,-nbitq), 
to_sfixed(871123984.0/4294967296.0,1,-nbitq), 
to_sfixed(-84171887.0/4294967296.0,1,-nbitq), 
to_sfixed(3219918.0/4294967296.0,1,-nbitq), 
to_sfixed(-1310424850.0/4294967296.0,1,-nbitq), 
to_sfixed(1118055195.0/4294967296.0,1,-nbitq), 
to_sfixed(46906921.0/4294967296.0,1,-nbitq), 
to_sfixed(-319038639.0/4294967296.0,1,-nbitq), 
to_sfixed(-518509804.0/4294967296.0,1,-nbitq), 
to_sfixed(1200790519.0/4294967296.0,1,-nbitq), 
to_sfixed(276192395.0/4294967296.0,1,-nbitq), 
to_sfixed(141071261.0/4294967296.0,1,-nbitq), 
to_sfixed(189711248.0/4294967296.0,1,-nbitq), 
to_sfixed(-294693790.0/4294967296.0,1,-nbitq), 
to_sfixed(957269524.0/4294967296.0,1,-nbitq), 
to_sfixed(645522094.0/4294967296.0,1,-nbitq), 
to_sfixed(4051924.0/4294967296.0,1,-nbitq), 
to_sfixed(58230687.0/4294967296.0,1,-nbitq), 
to_sfixed(-312538744.0/4294967296.0,1,-nbitq), 
to_sfixed(708706546.0/4294967296.0,1,-nbitq), 
to_sfixed(-2568364.0/4294967296.0,1,-nbitq), 
to_sfixed(70481672.0/4294967296.0,1,-nbitq), 
to_sfixed(-27466867.0/4294967296.0,1,-nbitq), 
to_sfixed(-229972617.0/4294967296.0,1,-nbitq), 
to_sfixed(-219710901.0/4294967296.0,1,-nbitq), 
to_sfixed(113797420.0/4294967296.0,1,-nbitq), 
to_sfixed(-257110240.0/4294967296.0,1,-nbitq), 
to_sfixed(-216035940.0/4294967296.0,1,-nbitq), 
to_sfixed(248716027.0/4294967296.0,1,-nbitq), 
to_sfixed(364586516.0/4294967296.0,1,-nbitq), 
to_sfixed(-330363247.0/4294967296.0,1,-nbitq), 
to_sfixed(187282705.0/4294967296.0,1,-nbitq), 
to_sfixed(-84375956.0/4294967296.0,1,-nbitq), 
to_sfixed(1388558067.0/4294967296.0,1,-nbitq), 
to_sfixed(63992859.0/4294967296.0,1,-nbitq), 
to_sfixed(-576467891.0/4294967296.0,1,-nbitq), 
to_sfixed(-710525215.0/4294967296.0,1,-nbitq), 
to_sfixed(-1388360900.0/4294967296.0,1,-nbitq), 
to_sfixed(52366227.0/4294967296.0,1,-nbitq), 
to_sfixed(-637781575.0/4294967296.0,1,-nbitq), 
to_sfixed(279404966.0/4294967296.0,1,-nbitq), 
to_sfixed(-627276260.0/4294967296.0,1,-nbitq), 
to_sfixed(-352769261.0/4294967296.0,1,-nbitq), 
to_sfixed(-362813300.0/4294967296.0,1,-nbitq), 
to_sfixed(79350750.0/4294967296.0,1,-nbitq), 
to_sfixed(6813596.0/4294967296.0,1,-nbitq), 
to_sfixed(221907696.0/4294967296.0,1,-nbitq), 
to_sfixed(-266992488.0/4294967296.0,1,-nbitq), 
to_sfixed(304236559.0/4294967296.0,1,-nbitq), 
to_sfixed(-128756359.0/4294967296.0,1,-nbitq), 
to_sfixed(63190239.0/4294967296.0,1,-nbitq), 
to_sfixed(-151416981.0/4294967296.0,1,-nbitq), 
to_sfixed(417845376.0/4294967296.0,1,-nbitq), 
to_sfixed(898317514.0/4294967296.0,1,-nbitq), 
to_sfixed(299794260.0/4294967296.0,1,-nbitq), 
to_sfixed(-1100907111.0/4294967296.0,1,-nbitq), 
to_sfixed(-209153792.0/4294967296.0,1,-nbitq), 
to_sfixed(-168646193.0/4294967296.0,1,-nbitq), 
to_sfixed(-194580364.0/4294967296.0,1,-nbitq), 
to_sfixed(-1873207.0/4294967296.0,1,-nbitq), 
to_sfixed(219889125.0/4294967296.0,1,-nbitq), 
to_sfixed(-201626429.0/4294967296.0,1,-nbitq), 
to_sfixed(-311007642.0/4294967296.0,1,-nbitq), 
to_sfixed(122551780.0/4294967296.0,1,-nbitq), 
to_sfixed(349069662.0/4294967296.0,1,-nbitq), 
to_sfixed(-191603981.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(13459871.0/4294967296.0,1,-nbitq), 
to_sfixed(426034671.0/4294967296.0,1,-nbitq), 
to_sfixed(-1549895428.0/4294967296.0,1,-nbitq), 
to_sfixed(-1209363282.0/4294967296.0,1,-nbitq), 
to_sfixed(276630875.0/4294967296.0,1,-nbitq), 
to_sfixed(2692776842.0/4294967296.0,1,-nbitq), 
to_sfixed(157492753.0/4294967296.0,1,-nbitq), 
to_sfixed(526757433.0/4294967296.0,1,-nbitq), 
to_sfixed(-763431197.0/4294967296.0,1,-nbitq), 
to_sfixed(92319086.0/4294967296.0,1,-nbitq), 
to_sfixed(698707515.0/4294967296.0,1,-nbitq), 
to_sfixed(-762309578.0/4294967296.0,1,-nbitq), 
to_sfixed(387660659.0/4294967296.0,1,-nbitq), 
to_sfixed(1728616695.0/4294967296.0,1,-nbitq), 
to_sfixed(-125661723.0/4294967296.0,1,-nbitq), 
to_sfixed(1048398290.0/4294967296.0,1,-nbitq), 
to_sfixed(268408282.0/4294967296.0,1,-nbitq), 
to_sfixed(-18720824.0/4294967296.0,1,-nbitq), 
to_sfixed(262507291.0/4294967296.0,1,-nbitq), 
to_sfixed(947948714.0/4294967296.0,1,-nbitq), 
to_sfixed(368073662.0/4294967296.0,1,-nbitq), 
to_sfixed(-812506595.0/4294967296.0,1,-nbitq), 
to_sfixed(-955193277.0/4294967296.0,1,-nbitq), 
to_sfixed(721369114.0/4294967296.0,1,-nbitq), 
to_sfixed(-130679408.0/4294967296.0,1,-nbitq), 
to_sfixed(-559947661.0/4294967296.0,1,-nbitq), 
to_sfixed(596721032.0/4294967296.0,1,-nbitq), 
to_sfixed(-313771076.0/4294967296.0,1,-nbitq), 
to_sfixed(556577006.0/4294967296.0,1,-nbitq), 
to_sfixed(954124468.0/4294967296.0,1,-nbitq), 
to_sfixed(267558542.0/4294967296.0,1,-nbitq), 
to_sfixed(-129858849.0/4294967296.0,1,-nbitq), 
to_sfixed(-579826950.0/4294967296.0,1,-nbitq), 
to_sfixed(-48503057.0/4294967296.0,1,-nbitq), 
to_sfixed(-174668502.0/4294967296.0,1,-nbitq), 
to_sfixed(-1205509201.0/4294967296.0,1,-nbitq), 
to_sfixed(-753556727.0/4294967296.0,1,-nbitq), 
to_sfixed(442988284.0/4294967296.0,1,-nbitq), 
to_sfixed(178993747.0/4294967296.0,1,-nbitq), 
to_sfixed(-453278424.0/4294967296.0,1,-nbitq), 
to_sfixed(196618901.0/4294967296.0,1,-nbitq), 
to_sfixed(-71478519.0/4294967296.0,1,-nbitq), 
to_sfixed(-259484097.0/4294967296.0,1,-nbitq), 
to_sfixed(-226057529.0/4294967296.0,1,-nbitq), 
to_sfixed(-619751693.0/4294967296.0,1,-nbitq), 
to_sfixed(108019354.0/4294967296.0,1,-nbitq), 
to_sfixed(244909074.0/4294967296.0,1,-nbitq), 
to_sfixed(1182985315.0/4294967296.0,1,-nbitq), 
to_sfixed(346590683.0/4294967296.0,1,-nbitq), 
to_sfixed(-284120267.0/4294967296.0,1,-nbitq), 
to_sfixed(-618118722.0/4294967296.0,1,-nbitq), 
to_sfixed(-1393865928.0/4294967296.0,1,-nbitq), 
to_sfixed(856219435.0/4294967296.0,1,-nbitq), 
to_sfixed(-768476647.0/4294967296.0,1,-nbitq), 
to_sfixed(1557105717.0/4294967296.0,1,-nbitq), 
to_sfixed(-893414762.0/4294967296.0,1,-nbitq), 
to_sfixed(-1039970641.0/4294967296.0,1,-nbitq), 
to_sfixed(46611630.0/4294967296.0,1,-nbitq), 
to_sfixed(286256764.0/4294967296.0,1,-nbitq), 
to_sfixed(201448567.0/4294967296.0,1,-nbitq), 
to_sfixed(-164570985.0/4294967296.0,1,-nbitq), 
to_sfixed(391338080.0/4294967296.0,1,-nbitq), 
to_sfixed(18002831.0/4294967296.0,1,-nbitq), 
to_sfixed(-269637486.0/4294967296.0,1,-nbitq), 
to_sfixed(-36326502.0/4294967296.0,1,-nbitq), 
to_sfixed(-186988623.0/4294967296.0,1,-nbitq), 
to_sfixed(119405247.0/4294967296.0,1,-nbitq), 
to_sfixed(965130563.0/4294967296.0,1,-nbitq), 
to_sfixed(238782991.0/4294967296.0,1,-nbitq), 
to_sfixed(-428678179.0/4294967296.0,1,-nbitq), 
to_sfixed(593443811.0/4294967296.0,1,-nbitq), 
to_sfixed(91829877.0/4294967296.0,1,-nbitq), 
to_sfixed(690612611.0/4294967296.0,1,-nbitq), 
to_sfixed(119364336.0/4294967296.0,1,-nbitq), 
to_sfixed(62771166.0/4294967296.0,1,-nbitq), 
to_sfixed(-288853984.0/4294967296.0,1,-nbitq), 
to_sfixed(542603480.0/4294967296.0,1,-nbitq), 
to_sfixed(30459754.0/4294967296.0,1,-nbitq), 
to_sfixed(267137334.0/4294967296.0,1,-nbitq), 
to_sfixed(-288479708.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-312459282.0/4294967296.0,1,-nbitq), 
to_sfixed(893744845.0/4294967296.0,1,-nbitq), 
to_sfixed(-442556394.0/4294967296.0,1,-nbitq), 
to_sfixed(-1297236035.0/4294967296.0,1,-nbitq), 
to_sfixed(-502326767.0/4294967296.0,1,-nbitq), 
to_sfixed(3485625899.0/4294967296.0,1,-nbitq), 
to_sfixed(53148204.0/4294967296.0,1,-nbitq), 
to_sfixed(1729250398.0/4294967296.0,1,-nbitq), 
to_sfixed(-1351151775.0/4294967296.0,1,-nbitq), 
to_sfixed(136940711.0/4294967296.0,1,-nbitq), 
to_sfixed(931828430.0/4294967296.0,1,-nbitq), 
to_sfixed(-757782456.0/4294967296.0,1,-nbitq), 
to_sfixed(659102838.0/4294967296.0,1,-nbitq), 
to_sfixed(2348423973.0/4294967296.0,1,-nbitq), 
to_sfixed(-47498534.0/4294967296.0,1,-nbitq), 
to_sfixed(442256115.0/4294967296.0,1,-nbitq), 
to_sfixed(112476919.0/4294967296.0,1,-nbitq), 
to_sfixed(-372364379.0/4294967296.0,1,-nbitq), 
to_sfixed(291286747.0/4294967296.0,1,-nbitq), 
to_sfixed(404985792.0/4294967296.0,1,-nbitq), 
to_sfixed(100018269.0/4294967296.0,1,-nbitq), 
to_sfixed(-377213478.0/4294967296.0,1,-nbitq), 
to_sfixed(-824973439.0/4294967296.0,1,-nbitq), 
to_sfixed(323794893.0/4294967296.0,1,-nbitq), 
to_sfixed(183312887.0/4294967296.0,1,-nbitq), 
to_sfixed(808199609.0/4294967296.0,1,-nbitq), 
to_sfixed(-126267792.0/4294967296.0,1,-nbitq), 
to_sfixed(285012320.0/4294967296.0,1,-nbitq), 
to_sfixed(1171948010.0/4294967296.0,1,-nbitq), 
to_sfixed(1102792001.0/4294967296.0,1,-nbitq), 
to_sfixed(256538046.0/4294967296.0,1,-nbitq), 
to_sfixed(42553932.0/4294967296.0,1,-nbitq), 
to_sfixed(-612735163.0/4294967296.0,1,-nbitq), 
to_sfixed(-605414866.0/4294967296.0,1,-nbitq), 
to_sfixed(-44638943.0/4294967296.0,1,-nbitq), 
to_sfixed(-42134532.0/4294967296.0,1,-nbitq), 
to_sfixed(-972454426.0/4294967296.0,1,-nbitq), 
to_sfixed(607229332.0/4294967296.0,1,-nbitq), 
to_sfixed(1135637.0/4294967296.0,1,-nbitq), 
to_sfixed(118492550.0/4294967296.0,1,-nbitq), 
to_sfixed(-268271308.0/4294967296.0,1,-nbitq), 
to_sfixed(-285277955.0/4294967296.0,1,-nbitq), 
to_sfixed(-875496207.0/4294967296.0,1,-nbitq), 
to_sfixed(84880735.0/4294967296.0,1,-nbitq), 
to_sfixed(-1117249990.0/4294967296.0,1,-nbitq), 
to_sfixed(-479862324.0/4294967296.0,1,-nbitq), 
to_sfixed(-37248858.0/4294967296.0,1,-nbitq), 
to_sfixed(1246348706.0/4294967296.0,1,-nbitq), 
to_sfixed(296944015.0/4294967296.0,1,-nbitq), 
to_sfixed(-1289150831.0/4294967296.0,1,-nbitq), 
to_sfixed(314094769.0/4294967296.0,1,-nbitq), 
to_sfixed(-1976403598.0/4294967296.0,1,-nbitq), 
to_sfixed(933179385.0/4294967296.0,1,-nbitq), 
to_sfixed(-532713921.0/4294967296.0,1,-nbitq), 
to_sfixed(1497672447.0/4294967296.0,1,-nbitq), 
to_sfixed(-1148933223.0/4294967296.0,1,-nbitq), 
to_sfixed(-504982332.0/4294967296.0,1,-nbitq), 
to_sfixed(-170192038.0/4294967296.0,1,-nbitq), 
to_sfixed(-334748877.0/4294967296.0,1,-nbitq), 
to_sfixed(-191289060.0/4294967296.0,1,-nbitq), 
to_sfixed(510397397.0/4294967296.0,1,-nbitq), 
to_sfixed(651911237.0/4294967296.0,1,-nbitq), 
to_sfixed(-772062132.0/4294967296.0,1,-nbitq), 
to_sfixed(-513359963.0/4294967296.0,1,-nbitq), 
to_sfixed(-445809054.0/4294967296.0,1,-nbitq), 
to_sfixed(-90477901.0/4294967296.0,1,-nbitq), 
to_sfixed(-2421880409.0/4294967296.0,1,-nbitq), 
to_sfixed(367510326.0/4294967296.0,1,-nbitq), 
to_sfixed(294896202.0/4294967296.0,1,-nbitq), 
to_sfixed(-837772740.0/4294967296.0,1,-nbitq), 
to_sfixed(1870680747.0/4294967296.0,1,-nbitq), 
to_sfixed(176478930.0/4294967296.0,1,-nbitq), 
to_sfixed(239541915.0/4294967296.0,1,-nbitq), 
to_sfixed(13541406.0/4294967296.0,1,-nbitq), 
to_sfixed(429430771.0/4294967296.0,1,-nbitq), 
to_sfixed(-540184316.0/4294967296.0,1,-nbitq), 
to_sfixed(-160293913.0/4294967296.0,1,-nbitq), 
to_sfixed(-214997220.0/4294967296.0,1,-nbitq), 
to_sfixed(177869663.0/4294967296.0,1,-nbitq), 
to_sfixed(-206842241.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(516125807.0/4294967296.0,1,-nbitq), 
to_sfixed(315657829.0/4294967296.0,1,-nbitq), 
to_sfixed(-1383337016.0/4294967296.0,1,-nbitq), 
to_sfixed(-1691502051.0/4294967296.0,1,-nbitq), 
to_sfixed(-345155704.0/4294967296.0,1,-nbitq), 
to_sfixed(-114946421.0/4294967296.0,1,-nbitq), 
to_sfixed(576334314.0/4294967296.0,1,-nbitq), 
to_sfixed(1223749498.0/4294967296.0,1,-nbitq), 
to_sfixed(-1048288779.0/4294967296.0,1,-nbitq), 
to_sfixed(-31501468.0/4294967296.0,1,-nbitq), 
to_sfixed(921875214.0/4294967296.0,1,-nbitq), 
to_sfixed(-1067340120.0/4294967296.0,1,-nbitq), 
to_sfixed(601154826.0/4294967296.0,1,-nbitq), 
to_sfixed(1829646722.0/4294967296.0,1,-nbitq), 
to_sfixed(-73153237.0/4294967296.0,1,-nbitq), 
to_sfixed(1018885702.0/4294967296.0,1,-nbitq), 
to_sfixed(221848120.0/4294967296.0,1,-nbitq), 
to_sfixed(168158149.0/4294967296.0,1,-nbitq), 
to_sfixed(509793985.0/4294967296.0,1,-nbitq), 
to_sfixed(831962265.0/4294967296.0,1,-nbitq), 
to_sfixed(400498592.0/4294967296.0,1,-nbitq), 
to_sfixed(-749182601.0/4294967296.0,1,-nbitq), 
to_sfixed(-692261161.0/4294967296.0,1,-nbitq), 
to_sfixed(457057417.0/4294967296.0,1,-nbitq), 
to_sfixed(120235109.0/4294967296.0,1,-nbitq), 
to_sfixed(354779742.0/4294967296.0,1,-nbitq), 
to_sfixed(-45103083.0/4294967296.0,1,-nbitq), 
to_sfixed(629900313.0/4294967296.0,1,-nbitq), 
to_sfixed(1471672606.0/4294967296.0,1,-nbitq), 
to_sfixed(1374465411.0/4294967296.0,1,-nbitq), 
to_sfixed(-150564304.0/4294967296.0,1,-nbitq), 
to_sfixed(-982997606.0/4294967296.0,1,-nbitq), 
to_sfixed(-772181623.0/4294967296.0,1,-nbitq), 
to_sfixed(-86828684.0/4294967296.0,1,-nbitq), 
to_sfixed(788900257.0/4294967296.0,1,-nbitq), 
to_sfixed(-49366696.0/4294967296.0,1,-nbitq), 
to_sfixed(137558009.0/4294967296.0,1,-nbitq), 
to_sfixed(1356717740.0/4294967296.0,1,-nbitq), 
to_sfixed(-474692441.0/4294967296.0,1,-nbitq), 
to_sfixed(-27230060.0/4294967296.0,1,-nbitq), 
to_sfixed(-866685520.0/4294967296.0,1,-nbitq), 
to_sfixed(-657700513.0/4294967296.0,1,-nbitq), 
to_sfixed(-656768203.0/4294967296.0,1,-nbitq), 
to_sfixed(-214046348.0/4294967296.0,1,-nbitq), 
to_sfixed(-1309351471.0/4294967296.0,1,-nbitq), 
to_sfixed(-226549151.0/4294967296.0,1,-nbitq), 
to_sfixed(-103861037.0/4294967296.0,1,-nbitq), 
to_sfixed(934916134.0/4294967296.0,1,-nbitq), 
to_sfixed(144710088.0/4294967296.0,1,-nbitq), 
to_sfixed(-1777870511.0/4294967296.0,1,-nbitq), 
to_sfixed(19556555.0/4294967296.0,1,-nbitq), 
to_sfixed(-1187027369.0/4294967296.0,1,-nbitq), 
to_sfixed(711258206.0/4294967296.0,1,-nbitq), 
to_sfixed(-33077582.0/4294967296.0,1,-nbitq), 
to_sfixed(1613989206.0/4294967296.0,1,-nbitq), 
to_sfixed(-1099941484.0/4294967296.0,1,-nbitq), 
to_sfixed(-231847486.0/4294967296.0,1,-nbitq), 
to_sfixed(-140858597.0/4294967296.0,1,-nbitq), 
to_sfixed(147777945.0/4294967296.0,1,-nbitq), 
to_sfixed(146890458.0/4294967296.0,1,-nbitq), 
to_sfixed(196722252.0/4294967296.0,1,-nbitq), 
to_sfixed(979827015.0/4294967296.0,1,-nbitq), 
to_sfixed(-448508723.0/4294967296.0,1,-nbitq), 
to_sfixed(-1222914606.0/4294967296.0,1,-nbitq), 
to_sfixed(19111285.0/4294967296.0,1,-nbitq), 
to_sfixed(-554527824.0/4294967296.0,1,-nbitq), 
to_sfixed(-2100091954.0/4294967296.0,1,-nbitq), 
to_sfixed(1568561254.0/4294967296.0,1,-nbitq), 
to_sfixed(-403922214.0/4294967296.0,1,-nbitq), 
to_sfixed(-194370625.0/4294967296.0,1,-nbitq), 
to_sfixed(1826275138.0/4294967296.0,1,-nbitq), 
to_sfixed(337222142.0/4294967296.0,1,-nbitq), 
to_sfixed(949479449.0/4294967296.0,1,-nbitq), 
to_sfixed(297799080.0/4294967296.0,1,-nbitq), 
to_sfixed(436310262.0/4294967296.0,1,-nbitq), 
to_sfixed(-485310754.0/4294967296.0,1,-nbitq), 
to_sfixed(-932105903.0/4294967296.0,1,-nbitq), 
to_sfixed(254906360.0/4294967296.0,1,-nbitq), 
to_sfixed(-1548507611.0/4294967296.0,1,-nbitq), 
to_sfixed(190125737.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(342889554.0/4294967296.0,1,-nbitq), 
to_sfixed(387880635.0/4294967296.0,1,-nbitq), 
to_sfixed(-2132292156.0/4294967296.0,1,-nbitq), 
to_sfixed(-1375282008.0/4294967296.0,1,-nbitq), 
to_sfixed(306420060.0/4294967296.0,1,-nbitq), 
to_sfixed(-1248129070.0/4294967296.0,1,-nbitq), 
to_sfixed(729390381.0/4294967296.0,1,-nbitq), 
to_sfixed(-838527952.0/4294967296.0,1,-nbitq), 
to_sfixed(-276912792.0/4294967296.0,1,-nbitq), 
to_sfixed(-393243907.0/4294967296.0,1,-nbitq), 
to_sfixed(277658784.0/4294967296.0,1,-nbitq), 
to_sfixed(-2052491860.0/4294967296.0,1,-nbitq), 
to_sfixed(1614169431.0/4294967296.0,1,-nbitq), 
to_sfixed(1678180850.0/4294967296.0,1,-nbitq), 
to_sfixed(233623626.0/4294967296.0,1,-nbitq), 
to_sfixed(1243044916.0/4294967296.0,1,-nbitq), 
to_sfixed(-263020916.0/4294967296.0,1,-nbitq), 
to_sfixed(-283985685.0/4294967296.0,1,-nbitq), 
to_sfixed(-548235567.0/4294967296.0,1,-nbitq), 
to_sfixed(1222067882.0/4294967296.0,1,-nbitq), 
to_sfixed(326123816.0/4294967296.0,1,-nbitq), 
to_sfixed(-1434439039.0/4294967296.0,1,-nbitq), 
to_sfixed(-1347382635.0/4294967296.0,1,-nbitq), 
to_sfixed(1098883485.0/4294967296.0,1,-nbitq), 
to_sfixed(-290030139.0/4294967296.0,1,-nbitq), 
to_sfixed(210196430.0/4294967296.0,1,-nbitq), 
to_sfixed(-176664569.0/4294967296.0,1,-nbitq), 
to_sfixed(1298441761.0/4294967296.0,1,-nbitq), 
to_sfixed(894172342.0/4294967296.0,1,-nbitq), 
to_sfixed(1080416441.0/4294967296.0,1,-nbitq), 
to_sfixed(-157480662.0/4294967296.0,1,-nbitq), 
to_sfixed(-909362522.0/4294967296.0,1,-nbitq), 
to_sfixed(-458915641.0/4294967296.0,1,-nbitq), 
to_sfixed(907436103.0/4294967296.0,1,-nbitq), 
to_sfixed(825179880.0/4294967296.0,1,-nbitq), 
to_sfixed(-131448201.0/4294967296.0,1,-nbitq), 
to_sfixed(-322233105.0/4294967296.0,1,-nbitq), 
to_sfixed(1874679477.0/4294967296.0,1,-nbitq), 
to_sfixed(110266989.0/4294967296.0,1,-nbitq), 
to_sfixed(257404367.0/4294967296.0,1,-nbitq), 
to_sfixed(-594951169.0/4294967296.0,1,-nbitq), 
to_sfixed(-911674124.0/4294967296.0,1,-nbitq), 
to_sfixed(-554341271.0/4294967296.0,1,-nbitq), 
to_sfixed(110086353.0/4294967296.0,1,-nbitq), 
to_sfixed(-468960246.0/4294967296.0,1,-nbitq), 
to_sfixed(-1995380596.0/4294967296.0,1,-nbitq), 
to_sfixed(223937735.0/4294967296.0,1,-nbitq), 
to_sfixed(337517794.0/4294967296.0,1,-nbitq), 
to_sfixed(410487826.0/4294967296.0,1,-nbitq), 
to_sfixed(-2015751108.0/4294967296.0,1,-nbitq), 
to_sfixed(-137019551.0/4294967296.0,1,-nbitq), 
to_sfixed(-1738158423.0/4294967296.0,1,-nbitq), 
to_sfixed(9166734.0/4294967296.0,1,-nbitq), 
to_sfixed(753631849.0/4294967296.0,1,-nbitq), 
to_sfixed(1603126773.0/4294967296.0,1,-nbitq), 
to_sfixed(-1152095662.0/4294967296.0,1,-nbitq), 
to_sfixed(646698236.0/4294967296.0,1,-nbitq), 
to_sfixed(-937073242.0/4294967296.0,1,-nbitq), 
to_sfixed(-39170116.0/4294967296.0,1,-nbitq), 
to_sfixed(314147152.0/4294967296.0,1,-nbitq), 
to_sfixed(274056946.0/4294967296.0,1,-nbitq), 
to_sfixed(1141172102.0/4294967296.0,1,-nbitq), 
to_sfixed(-1005673497.0/4294967296.0,1,-nbitq), 
to_sfixed(-1137454055.0/4294967296.0,1,-nbitq), 
to_sfixed(-122387518.0/4294967296.0,1,-nbitq), 
to_sfixed(-333922195.0/4294967296.0,1,-nbitq), 
to_sfixed(802762687.0/4294967296.0,1,-nbitq), 
to_sfixed(795517919.0/4294967296.0,1,-nbitq), 
to_sfixed(325416766.0/4294967296.0,1,-nbitq), 
to_sfixed(1732014212.0/4294967296.0,1,-nbitq), 
to_sfixed(2187628629.0/4294967296.0,1,-nbitq), 
to_sfixed(621942761.0/4294967296.0,1,-nbitq), 
to_sfixed(568359832.0/4294967296.0,1,-nbitq), 
to_sfixed(313686154.0/4294967296.0,1,-nbitq), 
to_sfixed(75361703.0/4294967296.0,1,-nbitq), 
to_sfixed(-418144934.0/4294967296.0,1,-nbitq), 
to_sfixed(-412392939.0/4294967296.0,1,-nbitq), 
to_sfixed(164333012.0/4294967296.0,1,-nbitq), 
to_sfixed(-2236570094.0/4294967296.0,1,-nbitq), 
to_sfixed(375304827.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(651673109.0/4294967296.0,1,-nbitq), 
to_sfixed(439535467.0/4294967296.0,1,-nbitq), 
to_sfixed(-1889185983.0/4294967296.0,1,-nbitq), 
to_sfixed(-948032016.0/4294967296.0,1,-nbitq), 
to_sfixed(1025641864.0/4294967296.0,1,-nbitq), 
to_sfixed(128407608.0/4294967296.0,1,-nbitq), 
to_sfixed(244232341.0/4294967296.0,1,-nbitq), 
to_sfixed(-1891334141.0/4294967296.0,1,-nbitq), 
to_sfixed(-400481702.0/4294967296.0,1,-nbitq), 
to_sfixed(-408109776.0/4294967296.0,1,-nbitq), 
to_sfixed(547351279.0/4294967296.0,1,-nbitq), 
to_sfixed(-2539495559.0/4294967296.0,1,-nbitq), 
to_sfixed(1098406593.0/4294967296.0,1,-nbitq), 
to_sfixed(350917105.0/4294967296.0,1,-nbitq), 
to_sfixed(286481914.0/4294967296.0,1,-nbitq), 
to_sfixed(929412722.0/4294967296.0,1,-nbitq), 
to_sfixed(312664018.0/4294967296.0,1,-nbitq), 
to_sfixed(68680426.0/4294967296.0,1,-nbitq), 
to_sfixed(12749861.0/4294967296.0,1,-nbitq), 
to_sfixed(1122152044.0/4294967296.0,1,-nbitq), 
to_sfixed(69280795.0/4294967296.0,1,-nbitq), 
to_sfixed(-1697366036.0/4294967296.0,1,-nbitq), 
to_sfixed(-491491552.0/4294967296.0,1,-nbitq), 
to_sfixed(1163040633.0/4294967296.0,1,-nbitq), 
to_sfixed(-365165220.0/4294967296.0,1,-nbitq), 
to_sfixed(391208146.0/4294967296.0,1,-nbitq), 
to_sfixed(-256949113.0/4294967296.0,1,-nbitq), 
to_sfixed(1136156691.0/4294967296.0,1,-nbitq), 
to_sfixed(-1487735433.0/4294967296.0,1,-nbitq), 
to_sfixed(913472916.0/4294967296.0,1,-nbitq), 
to_sfixed(1631228440.0/4294967296.0,1,-nbitq), 
to_sfixed(-17206841.0/4294967296.0,1,-nbitq), 
to_sfixed(-423101115.0/4294967296.0,1,-nbitq), 
to_sfixed(1225630631.0/4294967296.0,1,-nbitq), 
to_sfixed(880323395.0/4294967296.0,1,-nbitq), 
to_sfixed(635324361.0/4294967296.0,1,-nbitq), 
to_sfixed(-528574535.0/4294967296.0,1,-nbitq), 
to_sfixed(2073903442.0/4294967296.0,1,-nbitq), 
to_sfixed(-219705388.0/4294967296.0,1,-nbitq), 
to_sfixed(-37062641.0/4294967296.0,1,-nbitq), 
to_sfixed(688156410.0/4294967296.0,1,-nbitq), 
to_sfixed(-731510817.0/4294967296.0,1,-nbitq), 
to_sfixed(-840903681.0/4294967296.0,1,-nbitq), 
to_sfixed(-566936694.0/4294967296.0,1,-nbitq), 
to_sfixed(-10542980.0/4294967296.0,1,-nbitq), 
to_sfixed(-1518802296.0/4294967296.0,1,-nbitq), 
to_sfixed(-80649438.0/4294967296.0,1,-nbitq), 
to_sfixed(162293938.0/4294967296.0,1,-nbitq), 
to_sfixed(281640028.0/4294967296.0,1,-nbitq), 
to_sfixed(-1619342023.0/4294967296.0,1,-nbitq), 
to_sfixed(245697331.0/4294967296.0,1,-nbitq), 
to_sfixed(-714611947.0/4294967296.0,1,-nbitq), 
to_sfixed(-151500592.0/4294967296.0,1,-nbitq), 
to_sfixed(929911191.0/4294967296.0,1,-nbitq), 
to_sfixed(1600252731.0/4294967296.0,1,-nbitq), 
to_sfixed(-1931996474.0/4294967296.0,1,-nbitq), 
to_sfixed(-390908051.0/4294967296.0,1,-nbitq), 
to_sfixed(-1016559613.0/4294967296.0,1,-nbitq), 
to_sfixed(12493623.0/4294967296.0,1,-nbitq), 
to_sfixed(246461564.0/4294967296.0,1,-nbitq), 
to_sfixed(349048372.0/4294967296.0,1,-nbitq), 
to_sfixed(325867695.0/4294967296.0,1,-nbitq), 
to_sfixed(-897194768.0/4294967296.0,1,-nbitq), 
to_sfixed(-1269128116.0/4294967296.0,1,-nbitq), 
to_sfixed(68839533.0/4294967296.0,1,-nbitq), 
to_sfixed(-503243056.0/4294967296.0,1,-nbitq), 
to_sfixed(2531312855.0/4294967296.0,1,-nbitq), 
to_sfixed(462337796.0/4294967296.0,1,-nbitq), 
to_sfixed(-231119552.0/4294967296.0,1,-nbitq), 
to_sfixed(2865928859.0/4294967296.0,1,-nbitq), 
to_sfixed(1680109713.0/4294967296.0,1,-nbitq), 
to_sfixed(388786630.0/4294967296.0,1,-nbitq), 
to_sfixed(353855744.0/4294967296.0,1,-nbitq), 
to_sfixed(-292830364.0/4294967296.0,1,-nbitq), 
to_sfixed(-262448554.0/4294967296.0,1,-nbitq), 
to_sfixed(-1237737462.0/4294967296.0,1,-nbitq), 
to_sfixed(-1032342239.0/4294967296.0,1,-nbitq), 
to_sfixed(77221582.0/4294967296.0,1,-nbitq), 
to_sfixed(-1897158139.0/4294967296.0,1,-nbitq), 
to_sfixed(-309117673.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(393176395.0/4294967296.0,1,-nbitq), 
to_sfixed(-380065069.0/4294967296.0,1,-nbitq), 
to_sfixed(-251933031.0/4294967296.0,1,-nbitq), 
to_sfixed(-947910832.0/4294967296.0,1,-nbitq), 
to_sfixed(1780846753.0/4294967296.0,1,-nbitq), 
to_sfixed(738206855.0/4294967296.0,1,-nbitq), 
to_sfixed(23764899.0/4294967296.0,1,-nbitq), 
to_sfixed(-1310233198.0/4294967296.0,1,-nbitq), 
to_sfixed(-1976009974.0/4294967296.0,1,-nbitq), 
to_sfixed(268046746.0/4294967296.0,1,-nbitq), 
to_sfixed(179652919.0/4294967296.0,1,-nbitq), 
to_sfixed(-2933146061.0/4294967296.0,1,-nbitq), 
to_sfixed(728579379.0/4294967296.0,1,-nbitq), 
to_sfixed(-2681895.0/4294967296.0,1,-nbitq), 
to_sfixed(-406238542.0/4294967296.0,1,-nbitq), 
to_sfixed(288076761.0/4294967296.0,1,-nbitq), 
to_sfixed(-102728872.0/4294967296.0,1,-nbitq), 
to_sfixed(-244631288.0/4294967296.0,1,-nbitq), 
to_sfixed(134113649.0/4294967296.0,1,-nbitq), 
to_sfixed(347358862.0/4294967296.0,1,-nbitq), 
to_sfixed(-170553570.0/4294967296.0,1,-nbitq), 
to_sfixed(-697453458.0/4294967296.0,1,-nbitq), 
to_sfixed(605268060.0/4294967296.0,1,-nbitq), 
to_sfixed(3545706624.0/4294967296.0,1,-nbitq), 
to_sfixed(353498551.0/4294967296.0,1,-nbitq), 
to_sfixed(456707492.0/4294967296.0,1,-nbitq), 
to_sfixed(455210834.0/4294967296.0,1,-nbitq), 
to_sfixed(-268168900.0/4294967296.0,1,-nbitq), 
to_sfixed(-3009009835.0/4294967296.0,1,-nbitq), 
to_sfixed(971506554.0/4294967296.0,1,-nbitq), 
to_sfixed(2461119435.0/4294967296.0,1,-nbitq), 
to_sfixed(-689060657.0/4294967296.0,1,-nbitq), 
to_sfixed(-832524380.0/4294967296.0,1,-nbitq), 
to_sfixed(1353743967.0/4294967296.0,1,-nbitq), 
to_sfixed(-194440163.0/4294967296.0,1,-nbitq), 
to_sfixed(658071557.0/4294967296.0,1,-nbitq), 
to_sfixed(-58962989.0/4294967296.0,1,-nbitq), 
to_sfixed(1500485998.0/4294967296.0,1,-nbitq), 
to_sfixed(-236998937.0/4294967296.0,1,-nbitq), 
to_sfixed(149703192.0/4294967296.0,1,-nbitq), 
to_sfixed(1772338073.0/4294967296.0,1,-nbitq), 
to_sfixed(217084388.0/4294967296.0,1,-nbitq), 
to_sfixed(-137828068.0/4294967296.0,1,-nbitq), 
to_sfixed(-766796856.0/4294967296.0,1,-nbitq), 
to_sfixed(-803473301.0/4294967296.0,1,-nbitq), 
to_sfixed(275485126.0/4294967296.0,1,-nbitq), 
to_sfixed(127220872.0/4294967296.0,1,-nbitq), 
to_sfixed(863142480.0/4294967296.0,1,-nbitq), 
to_sfixed(82011803.0/4294967296.0,1,-nbitq), 
to_sfixed(-1483430684.0/4294967296.0,1,-nbitq), 
to_sfixed(107715247.0/4294967296.0,1,-nbitq), 
to_sfixed(-564345525.0/4294967296.0,1,-nbitq), 
to_sfixed(55373162.0/4294967296.0,1,-nbitq), 
to_sfixed(1566147150.0/4294967296.0,1,-nbitq), 
to_sfixed(1298774685.0/4294967296.0,1,-nbitq), 
to_sfixed(-2212036161.0/4294967296.0,1,-nbitq), 
to_sfixed(-365957068.0/4294967296.0,1,-nbitq), 
to_sfixed(-1297732006.0/4294967296.0,1,-nbitq), 
to_sfixed(429865879.0/4294967296.0,1,-nbitq), 
to_sfixed(219229314.0/4294967296.0,1,-nbitq), 
to_sfixed(468050464.0/4294967296.0,1,-nbitq), 
to_sfixed(260007312.0/4294967296.0,1,-nbitq), 
to_sfixed(230881015.0/4294967296.0,1,-nbitq), 
to_sfixed(-318474230.0/4294967296.0,1,-nbitq), 
to_sfixed(102324996.0/4294967296.0,1,-nbitq), 
to_sfixed(-136763473.0/4294967296.0,1,-nbitq), 
to_sfixed(1681558768.0/4294967296.0,1,-nbitq), 
to_sfixed(1021433828.0/4294967296.0,1,-nbitq), 
to_sfixed(-25435216.0/4294967296.0,1,-nbitq), 
to_sfixed(957573965.0/4294967296.0,1,-nbitq), 
to_sfixed(1101890958.0/4294967296.0,1,-nbitq), 
to_sfixed(188833184.0/4294967296.0,1,-nbitq), 
to_sfixed(-69109083.0/4294967296.0,1,-nbitq), 
to_sfixed(-7111098.0/4294967296.0,1,-nbitq), 
to_sfixed(17210746.0/4294967296.0,1,-nbitq), 
to_sfixed(-1086004920.0/4294967296.0,1,-nbitq), 
to_sfixed(-1887925826.0/4294967296.0,1,-nbitq), 
to_sfixed(-4895660.0/4294967296.0,1,-nbitq), 
to_sfixed(-1320883726.0/4294967296.0,1,-nbitq), 
to_sfixed(186226583.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(160268709.0/4294967296.0,1,-nbitq), 
to_sfixed(-373790689.0/4294967296.0,1,-nbitq), 
to_sfixed(-671430612.0/4294967296.0,1,-nbitq), 
to_sfixed(-815559655.0/4294967296.0,1,-nbitq), 
to_sfixed(1508275750.0/4294967296.0,1,-nbitq), 
to_sfixed(1520747792.0/4294967296.0,1,-nbitq), 
to_sfixed(-400890719.0/4294967296.0,1,-nbitq), 
to_sfixed(361515267.0/4294967296.0,1,-nbitq), 
to_sfixed(-1590209305.0/4294967296.0,1,-nbitq), 
to_sfixed(146160738.0/4294967296.0,1,-nbitq), 
to_sfixed(199197794.0/4294967296.0,1,-nbitq), 
to_sfixed(-1509189672.0/4294967296.0,1,-nbitq), 
to_sfixed(1345666255.0/4294967296.0,1,-nbitq), 
to_sfixed(464122576.0/4294967296.0,1,-nbitq), 
to_sfixed(-399683418.0/4294967296.0,1,-nbitq), 
to_sfixed(-503704090.0/4294967296.0,1,-nbitq), 
to_sfixed(-162697590.0/4294967296.0,1,-nbitq), 
to_sfixed(341168307.0/4294967296.0,1,-nbitq), 
to_sfixed(-1660118206.0/4294967296.0,1,-nbitq), 
to_sfixed(-88172331.0/4294967296.0,1,-nbitq), 
to_sfixed(35644752.0/4294967296.0,1,-nbitq), 
to_sfixed(-407215399.0/4294967296.0,1,-nbitq), 
to_sfixed(1789029297.0/4294967296.0,1,-nbitq), 
to_sfixed(628953839.0/4294967296.0,1,-nbitq), 
to_sfixed(251178299.0/4294967296.0,1,-nbitq), 
to_sfixed(-537581828.0/4294967296.0,1,-nbitq), 
to_sfixed(-410878627.0/4294967296.0,1,-nbitq), 
to_sfixed(-1559419859.0/4294967296.0,1,-nbitq), 
to_sfixed(-1125308028.0/4294967296.0,1,-nbitq), 
to_sfixed(1138431109.0/4294967296.0,1,-nbitq), 
to_sfixed(-444940806.0/4294967296.0,1,-nbitq), 
to_sfixed(-319934687.0/4294967296.0,1,-nbitq), 
to_sfixed(-769296952.0/4294967296.0,1,-nbitq), 
to_sfixed(1064286473.0/4294967296.0,1,-nbitq), 
to_sfixed(495501178.0/4294967296.0,1,-nbitq), 
to_sfixed(220580711.0/4294967296.0,1,-nbitq), 
to_sfixed(35405721.0/4294967296.0,1,-nbitq), 
to_sfixed(854260115.0/4294967296.0,1,-nbitq), 
to_sfixed(241068120.0/4294967296.0,1,-nbitq), 
to_sfixed(51570822.0/4294967296.0,1,-nbitq), 
to_sfixed(1670386272.0/4294967296.0,1,-nbitq), 
to_sfixed(1135170267.0/4294967296.0,1,-nbitq), 
to_sfixed(-47337336.0/4294967296.0,1,-nbitq), 
to_sfixed(-829040069.0/4294967296.0,1,-nbitq), 
to_sfixed(-1276521556.0/4294967296.0,1,-nbitq), 
to_sfixed(-1051946283.0/4294967296.0,1,-nbitq), 
to_sfixed(200188813.0/4294967296.0,1,-nbitq), 
to_sfixed(623255168.0/4294967296.0,1,-nbitq), 
to_sfixed(-22717121.0/4294967296.0,1,-nbitq), 
to_sfixed(-434849256.0/4294967296.0,1,-nbitq), 
to_sfixed(-184858501.0/4294967296.0,1,-nbitq), 
to_sfixed(-435008991.0/4294967296.0,1,-nbitq), 
to_sfixed(824285235.0/4294967296.0,1,-nbitq), 
to_sfixed(1295648083.0/4294967296.0,1,-nbitq), 
to_sfixed(-210297699.0/4294967296.0,1,-nbitq), 
to_sfixed(-867453475.0/4294967296.0,1,-nbitq), 
to_sfixed(-458054877.0/4294967296.0,1,-nbitq), 
to_sfixed(-1082675423.0/4294967296.0,1,-nbitq), 
to_sfixed(288200551.0/4294967296.0,1,-nbitq), 
to_sfixed(37394501.0/4294967296.0,1,-nbitq), 
to_sfixed(-1132089.0/4294967296.0,1,-nbitq), 
to_sfixed(-851448282.0/4294967296.0,1,-nbitq), 
to_sfixed(181896948.0/4294967296.0,1,-nbitq), 
to_sfixed(-429807930.0/4294967296.0,1,-nbitq), 
to_sfixed(-11068145.0/4294967296.0,1,-nbitq), 
to_sfixed(-303876666.0/4294967296.0,1,-nbitq), 
to_sfixed(2172346218.0/4294967296.0,1,-nbitq), 
to_sfixed(948639811.0/4294967296.0,1,-nbitq), 
to_sfixed(256906790.0/4294967296.0,1,-nbitq), 
to_sfixed(721220420.0/4294967296.0,1,-nbitq), 
to_sfixed(615394855.0/4294967296.0,1,-nbitq), 
to_sfixed(-463254411.0/4294967296.0,1,-nbitq), 
to_sfixed(-1413248045.0/4294967296.0,1,-nbitq), 
to_sfixed(-79864625.0/4294967296.0,1,-nbitq), 
to_sfixed(93351431.0/4294967296.0,1,-nbitq), 
to_sfixed(-1039495886.0/4294967296.0,1,-nbitq), 
to_sfixed(-1598368106.0/4294967296.0,1,-nbitq), 
to_sfixed(-557804363.0/4294967296.0,1,-nbitq), 
to_sfixed(-799491083.0/4294967296.0,1,-nbitq), 
to_sfixed(214263641.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(27278741.0/4294967296.0,1,-nbitq), 
to_sfixed(1214807628.0/4294967296.0,1,-nbitq), 
to_sfixed(406500436.0/4294967296.0,1,-nbitq), 
to_sfixed(-14679580.0/4294967296.0,1,-nbitq), 
to_sfixed(1118005282.0/4294967296.0,1,-nbitq), 
to_sfixed(971826026.0/4294967296.0,1,-nbitq), 
to_sfixed(83056322.0/4294967296.0,1,-nbitq), 
to_sfixed(668933958.0/4294967296.0,1,-nbitq), 
to_sfixed(-955136082.0/4294967296.0,1,-nbitq), 
to_sfixed(201320372.0/4294967296.0,1,-nbitq), 
to_sfixed(-371599345.0/4294967296.0,1,-nbitq), 
to_sfixed(-421470044.0/4294967296.0,1,-nbitq), 
to_sfixed(1070089147.0/4294967296.0,1,-nbitq), 
to_sfixed(-139044201.0/4294967296.0,1,-nbitq), 
to_sfixed(-205468144.0/4294967296.0,1,-nbitq), 
to_sfixed(-449269161.0/4294967296.0,1,-nbitq), 
to_sfixed(107239938.0/4294967296.0,1,-nbitq), 
to_sfixed(150047198.0/4294967296.0,1,-nbitq), 
to_sfixed(-1620009479.0/4294967296.0,1,-nbitq), 
to_sfixed(-984206582.0/4294967296.0,1,-nbitq), 
to_sfixed(50892940.0/4294967296.0,1,-nbitq), 
to_sfixed(996151325.0/4294967296.0,1,-nbitq), 
to_sfixed(733696088.0/4294967296.0,1,-nbitq), 
to_sfixed(-3055499145.0/4294967296.0,1,-nbitq), 
to_sfixed(-289964935.0/4294967296.0,1,-nbitq), 
to_sfixed(49514680.0/4294967296.0,1,-nbitq), 
to_sfixed(-698596948.0/4294967296.0,1,-nbitq), 
to_sfixed(-1466138697.0/4294967296.0,1,-nbitq), 
to_sfixed(304478360.0/4294967296.0,1,-nbitq), 
to_sfixed(1023049067.0/4294967296.0,1,-nbitq), 
to_sfixed(-2000293437.0/4294967296.0,1,-nbitq), 
to_sfixed(237697361.0/4294967296.0,1,-nbitq), 
to_sfixed(-221820642.0/4294967296.0,1,-nbitq), 
to_sfixed(893337518.0/4294967296.0,1,-nbitq), 
to_sfixed(1066801617.0/4294967296.0,1,-nbitq), 
to_sfixed(-916023661.0/4294967296.0,1,-nbitq), 
to_sfixed(8512655.0/4294967296.0,1,-nbitq), 
to_sfixed(-1212233427.0/4294967296.0,1,-nbitq), 
to_sfixed(51944734.0/4294967296.0,1,-nbitq), 
to_sfixed(-101857378.0/4294967296.0,1,-nbitq), 
to_sfixed(917458262.0/4294967296.0,1,-nbitq), 
to_sfixed(1751990422.0/4294967296.0,1,-nbitq), 
to_sfixed(420504760.0/4294967296.0,1,-nbitq), 
to_sfixed(-711423878.0/4294967296.0,1,-nbitq), 
to_sfixed(-1284922799.0/4294967296.0,1,-nbitq), 
to_sfixed(-503725792.0/4294967296.0,1,-nbitq), 
to_sfixed(148211578.0/4294967296.0,1,-nbitq), 
to_sfixed(750585377.0/4294967296.0,1,-nbitq), 
to_sfixed(50974097.0/4294967296.0,1,-nbitq), 
to_sfixed(47306965.0/4294967296.0,1,-nbitq), 
to_sfixed(-24431268.0/4294967296.0,1,-nbitq), 
to_sfixed(-1363007.0/4294967296.0,1,-nbitq), 
to_sfixed(2116499018.0/4294967296.0,1,-nbitq), 
to_sfixed(423417452.0/4294967296.0,1,-nbitq), 
to_sfixed(-860523622.0/4294967296.0,1,-nbitq), 
to_sfixed(-1330963685.0/4294967296.0,1,-nbitq), 
to_sfixed(-1016235149.0/4294967296.0,1,-nbitq), 
to_sfixed(157327373.0/4294967296.0,1,-nbitq), 
to_sfixed(-207032247.0/4294967296.0,1,-nbitq), 
to_sfixed(-253875550.0/4294967296.0,1,-nbitq), 
to_sfixed(-70153067.0/4294967296.0,1,-nbitq), 
to_sfixed(-1133275978.0/4294967296.0,1,-nbitq), 
to_sfixed(1152620374.0/4294967296.0,1,-nbitq), 
to_sfixed(33915348.0/4294967296.0,1,-nbitq), 
to_sfixed(-138646122.0/4294967296.0,1,-nbitq), 
to_sfixed(-292940635.0/4294967296.0,1,-nbitq), 
to_sfixed(1760226195.0/4294967296.0,1,-nbitq), 
to_sfixed(1704888702.0/4294967296.0,1,-nbitq), 
to_sfixed(108299414.0/4294967296.0,1,-nbitq), 
to_sfixed(365496983.0/4294967296.0,1,-nbitq), 
to_sfixed(361259025.0/4294967296.0,1,-nbitq), 
to_sfixed(-373516384.0/4294967296.0,1,-nbitq), 
to_sfixed(-1663021220.0/4294967296.0,1,-nbitq), 
to_sfixed(98135467.0/4294967296.0,1,-nbitq), 
to_sfixed(11231730.0/4294967296.0,1,-nbitq), 
to_sfixed(75056868.0/4294967296.0,1,-nbitq), 
to_sfixed(-1699990231.0/4294967296.0,1,-nbitq), 
to_sfixed(-720558704.0/4294967296.0,1,-nbitq), 
to_sfixed(21710564.0/4294967296.0,1,-nbitq), 
to_sfixed(294018698.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-443708998.0/4294967296.0,1,-nbitq), 
to_sfixed(1378654299.0/4294967296.0,1,-nbitq), 
to_sfixed(-542027864.0/4294967296.0,1,-nbitq), 
to_sfixed(-41277183.0/4294967296.0,1,-nbitq), 
to_sfixed(480369397.0/4294967296.0,1,-nbitq), 
to_sfixed(864449276.0/4294967296.0,1,-nbitq), 
to_sfixed(-432654883.0/4294967296.0,1,-nbitq), 
to_sfixed(331376529.0/4294967296.0,1,-nbitq), 
to_sfixed(-407154578.0/4294967296.0,1,-nbitq), 
to_sfixed(201355238.0/4294967296.0,1,-nbitq), 
to_sfixed(-202073947.0/4294967296.0,1,-nbitq), 
to_sfixed(1167147588.0/4294967296.0,1,-nbitq), 
to_sfixed(407131202.0/4294967296.0,1,-nbitq), 
to_sfixed(-639817684.0/4294967296.0,1,-nbitq), 
to_sfixed(21506145.0/4294967296.0,1,-nbitq), 
to_sfixed(-84217409.0/4294967296.0,1,-nbitq), 
to_sfixed(159589105.0/4294967296.0,1,-nbitq), 
to_sfixed(308580415.0/4294967296.0,1,-nbitq), 
to_sfixed(-1041403098.0/4294967296.0,1,-nbitq), 
to_sfixed(-954301391.0/4294967296.0,1,-nbitq), 
to_sfixed(-294825678.0/4294967296.0,1,-nbitq), 
to_sfixed(756933106.0/4294967296.0,1,-nbitq), 
to_sfixed(285330034.0/4294967296.0,1,-nbitq), 
to_sfixed(-2436285047.0/4294967296.0,1,-nbitq), 
to_sfixed(-113664247.0/4294967296.0,1,-nbitq), 
to_sfixed(314299605.0/4294967296.0,1,-nbitq), 
to_sfixed(-1203895326.0/4294967296.0,1,-nbitq), 
to_sfixed(-421249202.0/4294967296.0,1,-nbitq), 
to_sfixed(-287753372.0/4294967296.0,1,-nbitq), 
to_sfixed(1215592768.0/4294967296.0,1,-nbitq), 
to_sfixed(-1433244276.0/4294967296.0,1,-nbitq), 
to_sfixed(1802063478.0/4294967296.0,1,-nbitq), 
to_sfixed(-79352116.0/4294967296.0,1,-nbitq), 
to_sfixed(-21105117.0/4294967296.0,1,-nbitq), 
to_sfixed(-131731163.0/4294967296.0,1,-nbitq), 
to_sfixed(-544569251.0/4294967296.0,1,-nbitq), 
to_sfixed(-165597356.0/4294967296.0,1,-nbitq), 
to_sfixed(-1218943015.0/4294967296.0,1,-nbitq), 
to_sfixed(-33537275.0/4294967296.0,1,-nbitq), 
to_sfixed(118866060.0/4294967296.0,1,-nbitq), 
to_sfixed(403362539.0/4294967296.0,1,-nbitq), 
to_sfixed(1097320671.0/4294967296.0,1,-nbitq), 
to_sfixed(-538485404.0/4294967296.0,1,-nbitq), 
to_sfixed(-1741437091.0/4294967296.0,1,-nbitq), 
to_sfixed(-1086228658.0/4294967296.0,1,-nbitq), 
to_sfixed(-670024727.0/4294967296.0,1,-nbitq), 
to_sfixed(-362384219.0/4294967296.0,1,-nbitq), 
to_sfixed(691313231.0/4294967296.0,1,-nbitq), 
to_sfixed(-545214691.0/4294967296.0,1,-nbitq), 
to_sfixed(541679090.0/4294967296.0,1,-nbitq), 
to_sfixed(25311898.0/4294967296.0,1,-nbitq), 
to_sfixed(-360738068.0/4294967296.0,1,-nbitq), 
to_sfixed(1262816204.0/4294967296.0,1,-nbitq), 
to_sfixed(521409633.0/4294967296.0,1,-nbitq), 
to_sfixed(-785197497.0/4294967296.0,1,-nbitq), 
to_sfixed(-1269601055.0/4294967296.0,1,-nbitq), 
to_sfixed(-762123382.0/4294967296.0,1,-nbitq), 
to_sfixed(41736053.0/4294967296.0,1,-nbitq), 
to_sfixed(261300651.0/4294967296.0,1,-nbitq), 
to_sfixed(-53386627.0/4294967296.0,1,-nbitq), 
to_sfixed(-9051756.0/4294967296.0,1,-nbitq), 
to_sfixed(-1367336192.0/4294967296.0,1,-nbitq), 
to_sfixed(545528196.0/4294967296.0,1,-nbitq), 
to_sfixed(953315204.0/4294967296.0,1,-nbitq), 
to_sfixed(-437489300.0/4294967296.0,1,-nbitq), 
to_sfixed(152056061.0/4294967296.0,1,-nbitq), 
to_sfixed(-97523221.0/4294967296.0,1,-nbitq), 
to_sfixed(291470508.0/4294967296.0,1,-nbitq), 
to_sfixed(-290777288.0/4294967296.0,1,-nbitq), 
to_sfixed(898918186.0/4294967296.0,1,-nbitq), 
to_sfixed(539136786.0/4294967296.0,1,-nbitq), 
to_sfixed(-608442898.0/4294967296.0,1,-nbitq), 
to_sfixed(-1353524169.0/4294967296.0,1,-nbitq), 
to_sfixed(-73236258.0/4294967296.0,1,-nbitq), 
to_sfixed(255416603.0/4294967296.0,1,-nbitq), 
to_sfixed(295987241.0/4294967296.0,1,-nbitq), 
to_sfixed(-1420039033.0/4294967296.0,1,-nbitq), 
to_sfixed(-396698416.0/4294967296.0,1,-nbitq), 
to_sfixed(200623137.0/4294967296.0,1,-nbitq), 
to_sfixed(-255609212.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-489323825.0/4294967296.0,1,-nbitq), 
to_sfixed(1820606585.0/4294967296.0,1,-nbitq), 
to_sfixed(-1062662570.0/4294967296.0,1,-nbitq), 
to_sfixed(659911606.0/4294967296.0,1,-nbitq), 
to_sfixed(595634494.0/4294967296.0,1,-nbitq), 
to_sfixed(838302309.0/4294967296.0,1,-nbitq), 
to_sfixed(-19827433.0/4294967296.0,1,-nbitq), 
to_sfixed(131324919.0/4294967296.0,1,-nbitq), 
to_sfixed(-463128716.0/4294967296.0,1,-nbitq), 
to_sfixed(340712629.0/4294967296.0,1,-nbitq), 
to_sfixed(-617844132.0/4294967296.0,1,-nbitq), 
to_sfixed(1543414891.0/4294967296.0,1,-nbitq), 
to_sfixed(-567012347.0/4294967296.0,1,-nbitq), 
to_sfixed(-1678778858.0/4294967296.0,1,-nbitq), 
to_sfixed(341348108.0/4294967296.0,1,-nbitq), 
to_sfixed(104472140.0/4294967296.0,1,-nbitq), 
to_sfixed(273922679.0/4294967296.0,1,-nbitq), 
to_sfixed(-140910975.0/4294967296.0,1,-nbitq), 
to_sfixed(-890821815.0/4294967296.0,1,-nbitq), 
to_sfixed(-107872037.0/4294967296.0,1,-nbitq), 
to_sfixed(303517114.0/4294967296.0,1,-nbitq), 
to_sfixed(371630795.0/4294967296.0,1,-nbitq), 
to_sfixed(247096354.0/4294967296.0,1,-nbitq), 
to_sfixed(-1295077854.0/4294967296.0,1,-nbitq), 
to_sfixed(-217677659.0/4294967296.0,1,-nbitq), 
to_sfixed(692816875.0/4294967296.0,1,-nbitq), 
to_sfixed(-685600017.0/4294967296.0,1,-nbitq), 
to_sfixed(-354513339.0/4294967296.0,1,-nbitq), 
to_sfixed(177889945.0/4294967296.0,1,-nbitq), 
to_sfixed(1375268377.0/4294967296.0,1,-nbitq), 
to_sfixed(-538348397.0/4294967296.0,1,-nbitq), 
to_sfixed(2207498310.0/4294967296.0,1,-nbitq), 
to_sfixed(29978614.0/4294967296.0,1,-nbitq), 
to_sfixed(-69954744.0/4294967296.0,1,-nbitq), 
to_sfixed(-596299915.0/4294967296.0,1,-nbitq), 
to_sfixed(-593476271.0/4294967296.0,1,-nbitq), 
to_sfixed(-451062060.0/4294967296.0,1,-nbitq), 
to_sfixed(-983400087.0/4294967296.0,1,-nbitq), 
to_sfixed(391168759.0/4294967296.0,1,-nbitq), 
to_sfixed(201820889.0/4294967296.0,1,-nbitq), 
to_sfixed(-515453397.0/4294967296.0,1,-nbitq), 
to_sfixed(313672023.0/4294967296.0,1,-nbitq), 
to_sfixed(-439241699.0/4294967296.0,1,-nbitq), 
to_sfixed(-1181920529.0/4294967296.0,1,-nbitq), 
to_sfixed(-475410799.0/4294967296.0,1,-nbitq), 
to_sfixed(-377136719.0/4294967296.0,1,-nbitq), 
to_sfixed(-370812225.0/4294967296.0,1,-nbitq), 
to_sfixed(951064954.0/4294967296.0,1,-nbitq), 
to_sfixed(-937208490.0/4294967296.0,1,-nbitq), 
to_sfixed(572004375.0/4294967296.0,1,-nbitq), 
to_sfixed(-145508.0/4294967296.0,1,-nbitq), 
to_sfixed(-953454290.0/4294967296.0,1,-nbitq), 
to_sfixed(1219354953.0/4294967296.0,1,-nbitq), 
to_sfixed(674033191.0/4294967296.0,1,-nbitq), 
to_sfixed(-805015271.0/4294967296.0,1,-nbitq), 
to_sfixed(-851503633.0/4294967296.0,1,-nbitq), 
to_sfixed(68404748.0/4294967296.0,1,-nbitq), 
to_sfixed(-138806582.0/4294967296.0,1,-nbitq), 
to_sfixed(-140278660.0/4294967296.0,1,-nbitq), 
to_sfixed(-11787469.0/4294967296.0,1,-nbitq), 
to_sfixed(98089584.0/4294967296.0,1,-nbitq), 
to_sfixed(-1598573772.0/4294967296.0,1,-nbitq), 
to_sfixed(385525050.0/4294967296.0,1,-nbitq), 
to_sfixed(1134479529.0/4294967296.0,1,-nbitq), 
to_sfixed(-224697892.0/4294967296.0,1,-nbitq), 
to_sfixed(196619329.0/4294967296.0,1,-nbitq), 
to_sfixed(-2564147883.0/4294967296.0,1,-nbitq), 
to_sfixed(-322794098.0/4294967296.0,1,-nbitq), 
to_sfixed(97881756.0/4294967296.0,1,-nbitq), 
to_sfixed(698138808.0/4294967296.0,1,-nbitq), 
to_sfixed(68389821.0/4294967296.0,1,-nbitq), 
to_sfixed(-233660522.0/4294967296.0,1,-nbitq), 
to_sfixed(-1279621561.0/4294967296.0,1,-nbitq), 
to_sfixed(310441037.0/4294967296.0,1,-nbitq), 
to_sfixed(8326842.0/4294967296.0,1,-nbitq), 
to_sfixed(758193250.0/4294967296.0,1,-nbitq), 
to_sfixed(-1458209949.0/4294967296.0,1,-nbitq), 
to_sfixed(-22783483.0/4294967296.0,1,-nbitq), 
to_sfixed(-218256015.0/4294967296.0,1,-nbitq), 
to_sfixed(-107748205.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-520248985.0/4294967296.0,1,-nbitq), 
to_sfixed(1116512090.0/4294967296.0,1,-nbitq), 
to_sfixed(-644610235.0/4294967296.0,1,-nbitq), 
to_sfixed(355009934.0/4294967296.0,1,-nbitq), 
to_sfixed(-867576309.0/4294967296.0,1,-nbitq), 
to_sfixed(553529064.0/4294967296.0,1,-nbitq), 
to_sfixed(350599279.0/4294967296.0,1,-nbitq), 
to_sfixed(-406176415.0/4294967296.0,1,-nbitq), 
to_sfixed(-1076754417.0/4294967296.0,1,-nbitq), 
to_sfixed(-267203965.0/4294967296.0,1,-nbitq), 
to_sfixed(4089407.0/4294967296.0,1,-nbitq), 
to_sfixed(920225336.0/4294967296.0,1,-nbitq), 
to_sfixed(965412525.0/4294967296.0,1,-nbitq), 
to_sfixed(-2308069360.0/4294967296.0,1,-nbitq), 
to_sfixed(100428051.0/4294967296.0,1,-nbitq), 
to_sfixed(332754709.0/4294967296.0,1,-nbitq), 
to_sfixed(148571307.0/4294967296.0,1,-nbitq), 
to_sfixed(420315451.0/4294967296.0,1,-nbitq), 
to_sfixed(-62148210.0/4294967296.0,1,-nbitq), 
to_sfixed(-168448275.0/4294967296.0,1,-nbitq), 
to_sfixed(138015545.0/4294967296.0,1,-nbitq), 
to_sfixed(599559147.0/4294967296.0,1,-nbitq), 
to_sfixed(-349339229.0/4294967296.0,1,-nbitq), 
to_sfixed(-1648835596.0/4294967296.0,1,-nbitq), 
to_sfixed(-404076037.0/4294967296.0,1,-nbitq), 
to_sfixed(488943856.0/4294967296.0,1,-nbitq), 
to_sfixed(-768160770.0/4294967296.0,1,-nbitq), 
to_sfixed(183270345.0/4294967296.0,1,-nbitq), 
to_sfixed(-652823152.0/4294967296.0,1,-nbitq), 
to_sfixed(1300868962.0/4294967296.0,1,-nbitq), 
to_sfixed(-800322417.0/4294967296.0,1,-nbitq), 
to_sfixed(1913866007.0/4294967296.0,1,-nbitq), 
to_sfixed(-333013581.0/4294967296.0,1,-nbitq), 
to_sfixed(-227238831.0/4294967296.0,1,-nbitq), 
to_sfixed(119411513.0/4294967296.0,1,-nbitq), 
to_sfixed(-1145281945.0/4294967296.0,1,-nbitq), 
to_sfixed(-152230254.0/4294967296.0,1,-nbitq), 
to_sfixed(-665066997.0/4294967296.0,1,-nbitq), 
to_sfixed(-4442132.0/4294967296.0,1,-nbitq), 
to_sfixed(147149556.0/4294967296.0,1,-nbitq), 
to_sfixed(-1169475393.0/4294967296.0,1,-nbitq), 
to_sfixed(164006122.0/4294967296.0,1,-nbitq), 
to_sfixed(3788556.0/4294967296.0,1,-nbitq), 
to_sfixed(-522546688.0/4294967296.0,1,-nbitq), 
to_sfixed(-822783487.0/4294967296.0,1,-nbitq), 
to_sfixed(-841969742.0/4294967296.0,1,-nbitq), 
to_sfixed(-352808644.0/4294967296.0,1,-nbitq), 
to_sfixed(1007954327.0/4294967296.0,1,-nbitq), 
to_sfixed(-610000923.0/4294967296.0,1,-nbitq), 
to_sfixed(886246969.0/4294967296.0,1,-nbitq), 
to_sfixed(-156961340.0/4294967296.0,1,-nbitq), 
to_sfixed(-381294613.0/4294967296.0,1,-nbitq), 
to_sfixed(1310137009.0/4294967296.0,1,-nbitq), 
to_sfixed(383419324.0/4294967296.0,1,-nbitq), 
to_sfixed(-318773804.0/4294967296.0,1,-nbitq), 
to_sfixed(-19984276.0/4294967296.0,1,-nbitq), 
to_sfixed(497447760.0/4294967296.0,1,-nbitq), 
to_sfixed(-252197724.0/4294967296.0,1,-nbitq), 
to_sfixed(379561961.0/4294967296.0,1,-nbitq), 
to_sfixed(112908011.0/4294967296.0,1,-nbitq), 
to_sfixed(-171088020.0/4294967296.0,1,-nbitq), 
to_sfixed(667757711.0/4294967296.0,1,-nbitq), 
to_sfixed(71107558.0/4294967296.0,1,-nbitq), 
to_sfixed(1047352889.0/4294967296.0,1,-nbitq), 
to_sfixed(-126194705.0/4294967296.0,1,-nbitq), 
to_sfixed(219316710.0/4294967296.0,1,-nbitq), 
to_sfixed(-1984369260.0/4294967296.0,1,-nbitq), 
to_sfixed(167438633.0/4294967296.0,1,-nbitq), 
to_sfixed(24157245.0/4294967296.0,1,-nbitq), 
to_sfixed(636393307.0/4294967296.0,1,-nbitq), 
to_sfixed(567247566.0/4294967296.0,1,-nbitq), 
to_sfixed(-680328274.0/4294967296.0,1,-nbitq), 
to_sfixed(-499205540.0/4294967296.0,1,-nbitq), 
to_sfixed(300662206.0/4294967296.0,1,-nbitq), 
to_sfixed(-203167561.0/4294967296.0,1,-nbitq), 
to_sfixed(254782564.0/4294967296.0,1,-nbitq), 
to_sfixed(-1550427289.0/4294967296.0,1,-nbitq), 
to_sfixed(134251650.0/4294967296.0,1,-nbitq), 
to_sfixed(-511521145.0/4294967296.0,1,-nbitq), 
to_sfixed(187614615.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-461036897.0/4294967296.0,1,-nbitq), 
to_sfixed(1031178158.0/4294967296.0,1,-nbitq), 
to_sfixed(-880631878.0/4294967296.0,1,-nbitq), 
to_sfixed(-413650915.0/4294967296.0,1,-nbitq), 
to_sfixed(-1386507252.0/4294967296.0,1,-nbitq), 
to_sfixed(240302162.0/4294967296.0,1,-nbitq), 
to_sfixed(-216320822.0/4294967296.0,1,-nbitq), 
to_sfixed(-256410366.0/4294967296.0,1,-nbitq), 
to_sfixed(-940463065.0/4294967296.0,1,-nbitq), 
to_sfixed(-17420874.0/4294967296.0,1,-nbitq), 
to_sfixed(261812565.0/4294967296.0,1,-nbitq), 
to_sfixed(300227731.0/4294967296.0,1,-nbitq), 
to_sfixed(363581692.0/4294967296.0,1,-nbitq), 
to_sfixed(-1382122848.0/4294967296.0,1,-nbitq), 
to_sfixed(153736269.0/4294967296.0,1,-nbitq), 
to_sfixed(-150498313.0/4294967296.0,1,-nbitq), 
to_sfixed(-49479810.0/4294967296.0,1,-nbitq), 
to_sfixed(227105932.0/4294967296.0,1,-nbitq), 
to_sfixed(479975971.0/4294967296.0,1,-nbitq), 
to_sfixed(-83115925.0/4294967296.0,1,-nbitq), 
to_sfixed(-335877689.0/4294967296.0,1,-nbitq), 
to_sfixed(-370734151.0/4294967296.0,1,-nbitq), 
to_sfixed(-1291985210.0/4294967296.0,1,-nbitq), 
to_sfixed(-1283859294.0/4294967296.0,1,-nbitq), 
to_sfixed(252497003.0/4294967296.0,1,-nbitq), 
to_sfixed(751640450.0/4294967296.0,1,-nbitq), 
to_sfixed(-127808592.0/4294967296.0,1,-nbitq), 
to_sfixed(470473752.0/4294967296.0,1,-nbitq), 
to_sfixed(-957759147.0/4294967296.0,1,-nbitq), 
to_sfixed(1339989296.0/4294967296.0,1,-nbitq), 
to_sfixed(-484624249.0/4294967296.0,1,-nbitq), 
to_sfixed(1564779699.0/4294967296.0,1,-nbitq), 
to_sfixed(-597020285.0/4294967296.0,1,-nbitq), 
to_sfixed(-175032742.0/4294967296.0,1,-nbitq), 
to_sfixed(409380398.0/4294967296.0,1,-nbitq), 
to_sfixed(-573521744.0/4294967296.0,1,-nbitq), 
to_sfixed(-586361472.0/4294967296.0,1,-nbitq), 
to_sfixed(-677032856.0/4294967296.0,1,-nbitq), 
to_sfixed(628762466.0/4294967296.0,1,-nbitq), 
to_sfixed(558248988.0/4294967296.0,1,-nbitq), 
to_sfixed(-705327728.0/4294967296.0,1,-nbitq), 
to_sfixed(-348114408.0/4294967296.0,1,-nbitq), 
to_sfixed(-413167428.0/4294967296.0,1,-nbitq), 
to_sfixed(-436284307.0/4294967296.0,1,-nbitq), 
to_sfixed(-392311100.0/4294967296.0,1,-nbitq), 
to_sfixed(192473720.0/4294967296.0,1,-nbitq), 
to_sfixed(-247921093.0/4294967296.0,1,-nbitq), 
to_sfixed(485356705.0/4294967296.0,1,-nbitq), 
to_sfixed(-408310680.0/4294967296.0,1,-nbitq), 
to_sfixed(720382647.0/4294967296.0,1,-nbitq), 
to_sfixed(-496065305.0/4294967296.0,1,-nbitq), 
to_sfixed(-393139621.0/4294967296.0,1,-nbitq), 
to_sfixed(1370996204.0/4294967296.0,1,-nbitq), 
to_sfixed(334547320.0/4294967296.0,1,-nbitq), 
to_sfixed(-1164042798.0/4294967296.0,1,-nbitq), 
to_sfixed(476324105.0/4294967296.0,1,-nbitq), 
to_sfixed(378579794.0/4294967296.0,1,-nbitq), 
to_sfixed(-29583750.0/4294967296.0,1,-nbitq), 
to_sfixed(194384106.0/4294967296.0,1,-nbitq), 
to_sfixed(254671993.0/4294967296.0,1,-nbitq), 
to_sfixed(-274203927.0/4294967296.0,1,-nbitq), 
to_sfixed(535839593.0/4294967296.0,1,-nbitq), 
to_sfixed(17163850.0/4294967296.0,1,-nbitq), 
to_sfixed(551056492.0/4294967296.0,1,-nbitq), 
to_sfixed(-151476607.0/4294967296.0,1,-nbitq), 
to_sfixed(339725189.0/4294967296.0,1,-nbitq), 
to_sfixed(-1062418027.0/4294967296.0,1,-nbitq), 
to_sfixed(-512282114.0/4294967296.0,1,-nbitq), 
to_sfixed(359406632.0/4294967296.0,1,-nbitq), 
to_sfixed(374743835.0/4294967296.0,1,-nbitq), 
to_sfixed(423862057.0/4294967296.0,1,-nbitq), 
to_sfixed(-393889627.0/4294967296.0,1,-nbitq), 
to_sfixed(-28612203.0/4294967296.0,1,-nbitq), 
to_sfixed(40597540.0/4294967296.0,1,-nbitq), 
to_sfixed(-95900675.0/4294967296.0,1,-nbitq), 
to_sfixed(1096489484.0/4294967296.0,1,-nbitq), 
to_sfixed(-1542352843.0/4294967296.0,1,-nbitq), 
to_sfixed(78374376.0/4294967296.0,1,-nbitq), 
to_sfixed(-2219980.0/4294967296.0,1,-nbitq), 
to_sfixed(-214378532.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-171319159.0/4294967296.0,1,-nbitq), 
to_sfixed(644281144.0/4294967296.0,1,-nbitq), 
to_sfixed(-1137535758.0/4294967296.0,1,-nbitq), 
to_sfixed(621578244.0/4294967296.0,1,-nbitq), 
to_sfixed(-1550076578.0/4294967296.0,1,-nbitq), 
to_sfixed(297219170.0/4294967296.0,1,-nbitq), 
to_sfixed(-314100540.0/4294967296.0,1,-nbitq), 
to_sfixed(-226024462.0/4294967296.0,1,-nbitq), 
to_sfixed(-2221736232.0/4294967296.0,1,-nbitq), 
to_sfixed(133074917.0/4294967296.0,1,-nbitq), 
to_sfixed(-224626042.0/4294967296.0,1,-nbitq), 
to_sfixed(434627054.0/4294967296.0,1,-nbitq), 
to_sfixed(247406558.0/4294967296.0,1,-nbitq), 
to_sfixed(-880602448.0/4294967296.0,1,-nbitq), 
to_sfixed(478016622.0/4294967296.0,1,-nbitq), 
to_sfixed(-100881427.0/4294967296.0,1,-nbitq), 
to_sfixed(-13897284.0/4294967296.0,1,-nbitq), 
to_sfixed(-342456187.0/4294967296.0,1,-nbitq), 
to_sfixed(-436489935.0/4294967296.0,1,-nbitq), 
to_sfixed(-301308149.0/4294967296.0,1,-nbitq), 
to_sfixed(356236564.0/4294967296.0,1,-nbitq), 
to_sfixed(-1110427734.0/4294967296.0,1,-nbitq), 
to_sfixed(-1417947705.0/4294967296.0,1,-nbitq), 
to_sfixed(-1177633700.0/4294967296.0,1,-nbitq), 
to_sfixed(-269228551.0/4294967296.0,1,-nbitq), 
to_sfixed(918208765.0/4294967296.0,1,-nbitq), 
to_sfixed(-703190321.0/4294967296.0,1,-nbitq), 
to_sfixed(975148731.0/4294967296.0,1,-nbitq), 
to_sfixed(-502574178.0/4294967296.0,1,-nbitq), 
to_sfixed(1347469897.0/4294967296.0,1,-nbitq), 
to_sfixed(980550398.0/4294967296.0,1,-nbitq), 
to_sfixed(1507431970.0/4294967296.0,1,-nbitq), 
to_sfixed(-363752512.0/4294967296.0,1,-nbitq), 
to_sfixed(342380533.0/4294967296.0,1,-nbitq), 
to_sfixed(1035498823.0/4294967296.0,1,-nbitq), 
to_sfixed(402024767.0/4294967296.0,1,-nbitq), 
to_sfixed(-959011656.0/4294967296.0,1,-nbitq), 
to_sfixed(-119832323.0/4294967296.0,1,-nbitq), 
to_sfixed(508387291.0/4294967296.0,1,-nbitq), 
to_sfixed(484781012.0/4294967296.0,1,-nbitq), 
to_sfixed(-62145776.0/4294967296.0,1,-nbitq), 
to_sfixed(66076965.0/4294967296.0,1,-nbitq), 
to_sfixed(-1200744623.0/4294967296.0,1,-nbitq), 
to_sfixed(-1317974084.0/4294967296.0,1,-nbitq), 
to_sfixed(-598080297.0/4294967296.0,1,-nbitq), 
to_sfixed(-916255983.0/4294967296.0,1,-nbitq), 
to_sfixed(92164830.0/4294967296.0,1,-nbitq), 
to_sfixed(705953832.0/4294967296.0,1,-nbitq), 
to_sfixed(-25268703.0/4294967296.0,1,-nbitq), 
to_sfixed(841489073.0/4294967296.0,1,-nbitq), 
to_sfixed(20448472.0/4294967296.0,1,-nbitq), 
to_sfixed(-419216129.0/4294967296.0,1,-nbitq), 
to_sfixed(674651008.0/4294967296.0,1,-nbitq), 
to_sfixed(329171962.0/4294967296.0,1,-nbitq), 
to_sfixed(-519367098.0/4294967296.0,1,-nbitq), 
to_sfixed(-93213779.0/4294967296.0,1,-nbitq), 
to_sfixed(-14911899.0/4294967296.0,1,-nbitq), 
to_sfixed(58583899.0/4294967296.0,1,-nbitq), 
to_sfixed(254137490.0/4294967296.0,1,-nbitq), 
to_sfixed(-267652416.0/4294967296.0,1,-nbitq), 
to_sfixed(-261987233.0/4294967296.0,1,-nbitq), 
to_sfixed(326069420.0/4294967296.0,1,-nbitq), 
to_sfixed(303812566.0/4294967296.0,1,-nbitq), 
to_sfixed(356328547.0/4294967296.0,1,-nbitq), 
to_sfixed(366302883.0/4294967296.0,1,-nbitq), 
to_sfixed(-89244938.0/4294967296.0,1,-nbitq), 
to_sfixed(-342400215.0/4294967296.0,1,-nbitq), 
to_sfixed(-585826952.0/4294967296.0,1,-nbitq), 
to_sfixed(-331354166.0/4294967296.0,1,-nbitq), 
to_sfixed(814222460.0/4294967296.0,1,-nbitq), 
to_sfixed(423683185.0/4294967296.0,1,-nbitq), 
to_sfixed(-105337111.0/4294967296.0,1,-nbitq), 
to_sfixed(122017545.0/4294967296.0,1,-nbitq), 
to_sfixed(303220568.0/4294967296.0,1,-nbitq), 
to_sfixed(385264731.0/4294967296.0,1,-nbitq), 
to_sfixed(676047473.0/4294967296.0,1,-nbitq), 
to_sfixed(-2107680254.0/4294967296.0,1,-nbitq), 
to_sfixed(137092915.0/4294967296.0,1,-nbitq), 
to_sfixed(-90613546.0/4294967296.0,1,-nbitq), 
to_sfixed(210407981.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-303002883.0/4294967296.0,1,-nbitq), 
to_sfixed(804852615.0/4294967296.0,1,-nbitq), 
to_sfixed(-1011111172.0/4294967296.0,1,-nbitq), 
to_sfixed(-130348373.0/4294967296.0,1,-nbitq), 
to_sfixed(-1315017049.0/4294967296.0,1,-nbitq), 
to_sfixed(-487371871.0/4294967296.0,1,-nbitq), 
to_sfixed(-172312859.0/4294967296.0,1,-nbitq), 
to_sfixed(717902453.0/4294967296.0,1,-nbitq), 
to_sfixed(-1359226714.0/4294967296.0,1,-nbitq), 
to_sfixed(59560313.0/4294967296.0,1,-nbitq), 
to_sfixed(-7260917.0/4294967296.0,1,-nbitq), 
to_sfixed(-27172336.0/4294967296.0,1,-nbitq), 
to_sfixed(121541717.0/4294967296.0,1,-nbitq), 
to_sfixed(-600604252.0/4294967296.0,1,-nbitq), 
to_sfixed(-289121460.0/4294967296.0,1,-nbitq), 
to_sfixed(152155717.0/4294967296.0,1,-nbitq), 
to_sfixed(166095381.0/4294967296.0,1,-nbitq), 
to_sfixed(233321093.0/4294967296.0,1,-nbitq), 
to_sfixed(-100957635.0/4294967296.0,1,-nbitq), 
to_sfixed(-47755794.0/4294967296.0,1,-nbitq), 
to_sfixed(-358970273.0/4294967296.0,1,-nbitq), 
to_sfixed(-588853164.0/4294967296.0,1,-nbitq), 
to_sfixed(-1140270025.0/4294967296.0,1,-nbitq), 
to_sfixed(-1039965345.0/4294967296.0,1,-nbitq), 
to_sfixed(332662442.0/4294967296.0,1,-nbitq), 
to_sfixed(-367436859.0/4294967296.0,1,-nbitq), 
to_sfixed(-88603561.0/4294967296.0,1,-nbitq), 
to_sfixed(398846211.0/4294967296.0,1,-nbitq), 
to_sfixed(-97546987.0/4294967296.0,1,-nbitq), 
to_sfixed(467501105.0/4294967296.0,1,-nbitq), 
to_sfixed(724802652.0/4294967296.0,1,-nbitq), 
to_sfixed(1052794233.0/4294967296.0,1,-nbitq), 
to_sfixed(-243653556.0/4294967296.0,1,-nbitq), 
to_sfixed(923506988.0/4294967296.0,1,-nbitq), 
to_sfixed(-37056785.0/4294967296.0,1,-nbitq), 
to_sfixed(623437615.0/4294967296.0,1,-nbitq), 
to_sfixed(-478709590.0/4294967296.0,1,-nbitq), 
to_sfixed(599893334.0/4294967296.0,1,-nbitq), 
to_sfixed(213629559.0/4294967296.0,1,-nbitq), 
to_sfixed(430199819.0/4294967296.0,1,-nbitq), 
to_sfixed(-176282592.0/4294967296.0,1,-nbitq), 
to_sfixed(-139565059.0/4294967296.0,1,-nbitq), 
to_sfixed(-1286645501.0/4294967296.0,1,-nbitq), 
to_sfixed(-420252041.0/4294967296.0,1,-nbitq), 
to_sfixed(-918922471.0/4294967296.0,1,-nbitq), 
to_sfixed(-553080407.0/4294967296.0,1,-nbitq), 
to_sfixed(-392682407.0/4294967296.0,1,-nbitq), 
to_sfixed(920503739.0/4294967296.0,1,-nbitq), 
to_sfixed(212117575.0/4294967296.0,1,-nbitq), 
to_sfixed(213500337.0/4294967296.0,1,-nbitq), 
to_sfixed(504647875.0/4294967296.0,1,-nbitq), 
to_sfixed(-259522602.0/4294967296.0,1,-nbitq), 
to_sfixed(1150988646.0/4294967296.0,1,-nbitq), 
to_sfixed(171931871.0/4294967296.0,1,-nbitq), 
to_sfixed(-198309142.0/4294967296.0,1,-nbitq), 
to_sfixed(-393699780.0/4294967296.0,1,-nbitq), 
to_sfixed(863610353.0/4294967296.0,1,-nbitq), 
to_sfixed(237529989.0/4294967296.0,1,-nbitq), 
to_sfixed(-192386007.0/4294967296.0,1,-nbitq), 
to_sfixed(-341218598.0/4294967296.0,1,-nbitq), 
to_sfixed(-146723443.0/4294967296.0,1,-nbitq), 
to_sfixed(-788219694.0/4294967296.0,1,-nbitq), 
to_sfixed(46845678.0/4294967296.0,1,-nbitq), 
to_sfixed(-205036382.0/4294967296.0,1,-nbitq), 
to_sfixed(-185153760.0/4294967296.0,1,-nbitq), 
to_sfixed(397969884.0/4294967296.0,1,-nbitq), 
to_sfixed(246704929.0/4294967296.0,1,-nbitq), 
to_sfixed(-313227853.0/4294967296.0,1,-nbitq), 
to_sfixed(391295330.0/4294967296.0,1,-nbitq), 
to_sfixed(697069477.0/4294967296.0,1,-nbitq), 
to_sfixed(-222149553.0/4294967296.0,1,-nbitq), 
to_sfixed(48412691.0/4294967296.0,1,-nbitq), 
to_sfixed(349680983.0/4294967296.0,1,-nbitq), 
to_sfixed(-184815589.0/4294967296.0,1,-nbitq), 
to_sfixed(76470594.0/4294967296.0,1,-nbitq), 
to_sfixed(597194192.0/4294967296.0,1,-nbitq), 
to_sfixed(-887805595.0/4294967296.0,1,-nbitq), 
to_sfixed(-190663821.0/4294967296.0,1,-nbitq), 
to_sfixed(-419074947.0/4294967296.0,1,-nbitq), 
to_sfixed(-230121194.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(79991788.0/4294967296.0,1,-nbitq), 
to_sfixed(504698405.0/4294967296.0,1,-nbitq), 
to_sfixed(-1225168311.0/4294967296.0,1,-nbitq), 
to_sfixed(-1116602609.0/4294967296.0,1,-nbitq), 
to_sfixed(-1499970311.0/4294967296.0,1,-nbitq), 
to_sfixed(-167719152.0/4294967296.0,1,-nbitq), 
to_sfixed(-322665652.0/4294967296.0,1,-nbitq), 
to_sfixed(495759863.0/4294967296.0,1,-nbitq), 
to_sfixed(-1132814641.0/4294967296.0,1,-nbitq), 
to_sfixed(419000183.0/4294967296.0,1,-nbitq), 
to_sfixed(647174956.0/4294967296.0,1,-nbitq), 
to_sfixed(128799150.0/4294967296.0,1,-nbitq), 
to_sfixed(697658272.0/4294967296.0,1,-nbitq), 
to_sfixed(-1038023476.0/4294967296.0,1,-nbitq), 
to_sfixed(229206430.0/4294967296.0,1,-nbitq), 
to_sfixed(45990435.0/4294967296.0,1,-nbitq), 
to_sfixed(-119080933.0/4294967296.0,1,-nbitq), 
to_sfixed(-194707069.0/4294967296.0,1,-nbitq), 
to_sfixed(730896567.0/4294967296.0,1,-nbitq), 
to_sfixed(18118119.0/4294967296.0,1,-nbitq), 
to_sfixed(169495919.0/4294967296.0,1,-nbitq), 
to_sfixed(-570044414.0/4294967296.0,1,-nbitq), 
to_sfixed(-352105110.0/4294967296.0,1,-nbitq), 
to_sfixed(-1158567284.0/4294967296.0,1,-nbitq), 
to_sfixed(-62645726.0/4294967296.0,1,-nbitq), 
to_sfixed(-1288192125.0/4294967296.0,1,-nbitq), 
to_sfixed(184771863.0/4294967296.0,1,-nbitq), 
to_sfixed(435289243.0/4294967296.0,1,-nbitq), 
to_sfixed(-253377961.0/4294967296.0,1,-nbitq), 
to_sfixed(374779304.0/4294967296.0,1,-nbitq), 
to_sfixed(496880967.0/4294967296.0,1,-nbitq), 
to_sfixed(382629948.0/4294967296.0,1,-nbitq), 
to_sfixed(-379444240.0/4294967296.0,1,-nbitq), 
to_sfixed(1366173819.0/4294967296.0,1,-nbitq), 
to_sfixed(-750543380.0/4294967296.0,1,-nbitq), 
to_sfixed(179812433.0/4294967296.0,1,-nbitq), 
to_sfixed(-142931680.0/4294967296.0,1,-nbitq), 
to_sfixed(-252878658.0/4294967296.0,1,-nbitq), 
to_sfixed(-163564233.0/4294967296.0,1,-nbitq), 
to_sfixed(-175930999.0/4294967296.0,1,-nbitq), 
to_sfixed(-200896208.0/4294967296.0,1,-nbitq), 
to_sfixed(-483025412.0/4294967296.0,1,-nbitq), 
to_sfixed(-523565534.0/4294967296.0,1,-nbitq), 
to_sfixed(-389812561.0/4294967296.0,1,-nbitq), 
to_sfixed(-786085939.0/4294967296.0,1,-nbitq), 
to_sfixed(105235851.0/4294967296.0,1,-nbitq), 
to_sfixed(297915077.0/4294967296.0,1,-nbitq), 
to_sfixed(407146424.0/4294967296.0,1,-nbitq), 
to_sfixed(179100104.0/4294967296.0,1,-nbitq), 
to_sfixed(-50511313.0/4294967296.0,1,-nbitq), 
to_sfixed(138586793.0/4294967296.0,1,-nbitq), 
to_sfixed(-871037112.0/4294967296.0,1,-nbitq), 
to_sfixed(755352931.0/4294967296.0,1,-nbitq), 
to_sfixed(-532628880.0/4294967296.0,1,-nbitq), 
to_sfixed(-506038021.0/4294967296.0,1,-nbitq), 
to_sfixed(-117291556.0/4294967296.0,1,-nbitq), 
to_sfixed(809180265.0/4294967296.0,1,-nbitq), 
to_sfixed(17747060.0/4294967296.0,1,-nbitq), 
to_sfixed(-77458706.0/4294967296.0,1,-nbitq), 
to_sfixed(-242109206.0/4294967296.0,1,-nbitq), 
to_sfixed(405365933.0/4294967296.0,1,-nbitq), 
to_sfixed(-859255109.0/4294967296.0,1,-nbitq), 
to_sfixed(451062257.0/4294967296.0,1,-nbitq), 
to_sfixed(-568717569.0/4294967296.0,1,-nbitq), 
to_sfixed(153564796.0/4294967296.0,1,-nbitq), 
to_sfixed(-196423164.0/4294967296.0,1,-nbitq), 
to_sfixed(10150199.0/4294967296.0,1,-nbitq), 
to_sfixed(-90360801.0/4294967296.0,1,-nbitq), 
to_sfixed(64272992.0/4294967296.0,1,-nbitq), 
to_sfixed(576159502.0/4294967296.0,1,-nbitq), 
to_sfixed(-346635650.0/4294967296.0,1,-nbitq), 
to_sfixed(63737056.0/4294967296.0,1,-nbitq), 
to_sfixed(262962076.0/4294967296.0,1,-nbitq), 
to_sfixed(-192291759.0/4294967296.0,1,-nbitq), 
to_sfixed(-1047350.0/4294967296.0,1,-nbitq), 
to_sfixed(455116127.0/4294967296.0,1,-nbitq), 
to_sfixed(-1108855629.0/4294967296.0,1,-nbitq), 
to_sfixed(158009048.0/4294967296.0,1,-nbitq), 
to_sfixed(303166493.0/4294967296.0,1,-nbitq), 
to_sfixed(-331257090.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-337080620.0/4294967296.0,1,-nbitq), 
to_sfixed(649746531.0/4294967296.0,1,-nbitq), 
to_sfixed(-980144315.0/4294967296.0,1,-nbitq), 
to_sfixed(-912143357.0/4294967296.0,1,-nbitq), 
to_sfixed(-839820654.0/4294967296.0,1,-nbitq), 
to_sfixed(-392721259.0/4294967296.0,1,-nbitq), 
to_sfixed(-238972875.0/4294967296.0,1,-nbitq), 
to_sfixed(480602033.0/4294967296.0,1,-nbitq), 
to_sfixed(-1170877467.0/4294967296.0,1,-nbitq), 
to_sfixed(114425375.0/4294967296.0,1,-nbitq), 
to_sfixed(479925573.0/4294967296.0,1,-nbitq), 
to_sfixed(284493546.0/4294967296.0,1,-nbitq), 
to_sfixed(389964490.0/4294967296.0,1,-nbitq), 
to_sfixed(-615739038.0/4294967296.0,1,-nbitq), 
to_sfixed(-186949889.0/4294967296.0,1,-nbitq), 
to_sfixed(336576268.0/4294967296.0,1,-nbitq), 
to_sfixed(314929593.0/4294967296.0,1,-nbitq), 
to_sfixed(-358800035.0/4294967296.0,1,-nbitq), 
to_sfixed(-31674783.0/4294967296.0,1,-nbitq), 
to_sfixed(266918177.0/4294967296.0,1,-nbitq), 
to_sfixed(278161239.0/4294967296.0,1,-nbitq), 
to_sfixed(36208524.0/4294967296.0,1,-nbitq), 
to_sfixed(-384044270.0/4294967296.0,1,-nbitq), 
to_sfixed(-618719965.0/4294967296.0,1,-nbitq), 
to_sfixed(344848551.0/4294967296.0,1,-nbitq), 
to_sfixed(-923223872.0/4294967296.0,1,-nbitq), 
to_sfixed(-104426800.0/4294967296.0,1,-nbitq), 
to_sfixed(507999988.0/4294967296.0,1,-nbitq), 
to_sfixed(-141016581.0/4294967296.0,1,-nbitq), 
to_sfixed(111101535.0/4294967296.0,1,-nbitq), 
to_sfixed(-86472945.0/4294967296.0,1,-nbitq), 
to_sfixed(-66649433.0/4294967296.0,1,-nbitq), 
to_sfixed(328074950.0/4294967296.0,1,-nbitq), 
to_sfixed(250172778.0/4294967296.0,1,-nbitq), 
to_sfixed(70551646.0/4294967296.0,1,-nbitq), 
to_sfixed(205679713.0/4294967296.0,1,-nbitq), 
to_sfixed(-311199021.0/4294967296.0,1,-nbitq), 
to_sfixed(-141299920.0/4294967296.0,1,-nbitq), 
to_sfixed(-182695232.0/4294967296.0,1,-nbitq), 
to_sfixed(413677435.0/4294967296.0,1,-nbitq), 
to_sfixed(469633387.0/4294967296.0,1,-nbitq), 
to_sfixed(-812728273.0/4294967296.0,1,-nbitq), 
to_sfixed(-388647290.0/4294967296.0,1,-nbitq), 
to_sfixed(-1102204058.0/4294967296.0,1,-nbitq), 
to_sfixed(-557796021.0/4294967296.0,1,-nbitq), 
to_sfixed(-322070790.0/4294967296.0,1,-nbitq), 
to_sfixed(241906949.0/4294967296.0,1,-nbitq), 
to_sfixed(-12175535.0/4294967296.0,1,-nbitq), 
to_sfixed(109257000.0/4294967296.0,1,-nbitq), 
to_sfixed(154452769.0/4294967296.0,1,-nbitq), 
to_sfixed(382044888.0/4294967296.0,1,-nbitq), 
to_sfixed(-57525724.0/4294967296.0,1,-nbitq), 
to_sfixed(806536690.0/4294967296.0,1,-nbitq), 
to_sfixed(-704660656.0/4294967296.0,1,-nbitq), 
to_sfixed(-827497414.0/4294967296.0,1,-nbitq), 
to_sfixed(-603400548.0/4294967296.0,1,-nbitq), 
to_sfixed(1090338615.0/4294967296.0,1,-nbitq), 
to_sfixed(515177463.0/4294967296.0,1,-nbitq), 
to_sfixed(356920116.0/4294967296.0,1,-nbitq), 
to_sfixed(205685987.0/4294967296.0,1,-nbitq), 
to_sfixed(272320816.0/4294967296.0,1,-nbitq), 
to_sfixed(-967670372.0/4294967296.0,1,-nbitq), 
to_sfixed(-24785229.0/4294967296.0,1,-nbitq), 
to_sfixed(55987466.0/4294967296.0,1,-nbitq), 
to_sfixed(-224190118.0/4294967296.0,1,-nbitq), 
to_sfixed(110767826.0/4294967296.0,1,-nbitq), 
to_sfixed(-50890444.0/4294967296.0,1,-nbitq), 
to_sfixed(-591291744.0/4294967296.0,1,-nbitq), 
to_sfixed(-19246326.0/4294967296.0,1,-nbitq), 
to_sfixed(922996622.0/4294967296.0,1,-nbitq), 
to_sfixed(-506229179.0/4294967296.0,1,-nbitq), 
to_sfixed(-60292273.0/4294967296.0,1,-nbitq), 
to_sfixed(813564956.0/4294967296.0,1,-nbitq), 
to_sfixed(414481482.0/4294967296.0,1,-nbitq), 
to_sfixed(451335069.0/4294967296.0,1,-nbitq), 
to_sfixed(185896059.0/4294967296.0,1,-nbitq), 
to_sfixed(-1171667377.0/4294967296.0,1,-nbitq), 
to_sfixed(-653522493.0/4294967296.0,1,-nbitq), 
to_sfixed(71414625.0/4294967296.0,1,-nbitq), 
to_sfixed(-122664400.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(194406940.0/4294967296.0,1,-nbitq), 
to_sfixed(668450358.0/4294967296.0,1,-nbitq), 
to_sfixed(-688878469.0/4294967296.0,1,-nbitq), 
to_sfixed(-203104100.0/4294967296.0,1,-nbitq), 
to_sfixed(-791158970.0/4294967296.0,1,-nbitq), 
to_sfixed(-791346121.0/4294967296.0,1,-nbitq), 
to_sfixed(125564162.0/4294967296.0,1,-nbitq), 
to_sfixed(702064400.0/4294967296.0,1,-nbitq), 
to_sfixed(-588882497.0/4294967296.0,1,-nbitq), 
to_sfixed(329086735.0/4294967296.0,1,-nbitq), 
to_sfixed(688950133.0/4294967296.0,1,-nbitq), 
to_sfixed(119699766.0/4294967296.0,1,-nbitq), 
to_sfixed(77346388.0/4294967296.0,1,-nbitq), 
to_sfixed(-143565432.0/4294967296.0,1,-nbitq), 
to_sfixed(124367609.0/4294967296.0,1,-nbitq), 
to_sfixed(-230648090.0/4294967296.0,1,-nbitq), 
to_sfixed(272851659.0/4294967296.0,1,-nbitq), 
to_sfixed(-426321896.0/4294967296.0,1,-nbitq), 
to_sfixed(-21735711.0/4294967296.0,1,-nbitq), 
to_sfixed(-333309914.0/4294967296.0,1,-nbitq), 
to_sfixed(-157066584.0/4294967296.0,1,-nbitq), 
to_sfixed(-258862542.0/4294967296.0,1,-nbitq), 
to_sfixed(-179877619.0/4294967296.0,1,-nbitq), 
to_sfixed(-342995149.0/4294967296.0,1,-nbitq), 
to_sfixed(-130190116.0/4294967296.0,1,-nbitq), 
to_sfixed(-870330389.0/4294967296.0,1,-nbitq), 
to_sfixed(479928636.0/4294967296.0,1,-nbitq), 
to_sfixed(454584679.0/4294967296.0,1,-nbitq), 
to_sfixed(-434418221.0/4294967296.0,1,-nbitq), 
to_sfixed(573120643.0/4294967296.0,1,-nbitq), 
to_sfixed(-9697197.0/4294967296.0,1,-nbitq), 
to_sfixed(407960877.0/4294967296.0,1,-nbitq), 
to_sfixed(295074866.0/4294967296.0,1,-nbitq), 
to_sfixed(95541042.0/4294967296.0,1,-nbitq), 
to_sfixed(-764103823.0/4294967296.0,1,-nbitq), 
to_sfixed(111978240.0/4294967296.0,1,-nbitq), 
to_sfixed(-373624751.0/4294967296.0,1,-nbitq), 
to_sfixed(-74179329.0/4294967296.0,1,-nbitq), 
to_sfixed(172769841.0/4294967296.0,1,-nbitq), 
to_sfixed(-222439726.0/4294967296.0,1,-nbitq), 
to_sfixed(2866153.0/4294967296.0,1,-nbitq), 
to_sfixed(-255653131.0/4294967296.0,1,-nbitq), 
to_sfixed(-250364521.0/4294967296.0,1,-nbitq), 
to_sfixed(-1111860625.0/4294967296.0,1,-nbitq), 
to_sfixed(-229161036.0/4294967296.0,1,-nbitq), 
to_sfixed(-423526410.0/4294967296.0,1,-nbitq), 
to_sfixed(-97986820.0/4294967296.0,1,-nbitq), 
to_sfixed(-416656157.0/4294967296.0,1,-nbitq), 
to_sfixed(87513929.0/4294967296.0,1,-nbitq), 
to_sfixed(-114063126.0/4294967296.0,1,-nbitq), 
to_sfixed(-152715087.0/4294967296.0,1,-nbitq), 
to_sfixed(-123453751.0/4294967296.0,1,-nbitq), 
to_sfixed(898163559.0/4294967296.0,1,-nbitq), 
to_sfixed(73200941.0/4294967296.0,1,-nbitq), 
to_sfixed(-351067683.0/4294967296.0,1,-nbitq), 
to_sfixed(-339760886.0/4294967296.0,1,-nbitq), 
to_sfixed(426353187.0/4294967296.0,1,-nbitq), 
to_sfixed(485280788.0/4294967296.0,1,-nbitq), 
to_sfixed(-229537727.0/4294967296.0,1,-nbitq), 
to_sfixed(-46588752.0/4294967296.0,1,-nbitq), 
to_sfixed(-195738668.0/4294967296.0,1,-nbitq), 
to_sfixed(-623704294.0/4294967296.0,1,-nbitq), 
to_sfixed(-63940648.0/4294967296.0,1,-nbitq), 
to_sfixed(-219571231.0/4294967296.0,1,-nbitq), 
to_sfixed(-62942729.0/4294967296.0,1,-nbitq), 
to_sfixed(226580068.0/4294967296.0,1,-nbitq), 
to_sfixed(188613089.0/4294967296.0,1,-nbitq), 
to_sfixed(-138505345.0/4294967296.0,1,-nbitq), 
to_sfixed(-220308899.0/4294967296.0,1,-nbitq), 
to_sfixed(86502313.0/4294967296.0,1,-nbitq), 
to_sfixed(376007783.0/4294967296.0,1,-nbitq), 
to_sfixed(27526287.0/4294967296.0,1,-nbitq), 
to_sfixed(998774163.0/4294967296.0,1,-nbitq), 
to_sfixed(-126986314.0/4294967296.0,1,-nbitq), 
to_sfixed(311491924.0/4294967296.0,1,-nbitq), 
to_sfixed(-314427486.0/4294967296.0,1,-nbitq), 
to_sfixed(-478760363.0/4294967296.0,1,-nbitq), 
to_sfixed(-223686398.0/4294967296.0,1,-nbitq), 
to_sfixed(-68630847.0/4294967296.0,1,-nbitq), 
to_sfixed(-51218232.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-75590613.0/4294967296.0,1,-nbitq), 
to_sfixed(159178697.0/4294967296.0,1,-nbitq), 
to_sfixed(474958858.0/4294967296.0,1,-nbitq), 
to_sfixed(-690363668.0/4294967296.0,1,-nbitq), 
to_sfixed(-173184472.0/4294967296.0,1,-nbitq), 
to_sfixed(-285588876.0/4294967296.0,1,-nbitq), 
to_sfixed(-4103565.0/4294967296.0,1,-nbitq), 
to_sfixed(390891320.0/4294967296.0,1,-nbitq), 
to_sfixed(-543083886.0/4294967296.0,1,-nbitq), 
to_sfixed(195115339.0/4294967296.0,1,-nbitq), 
to_sfixed(489743582.0/4294967296.0,1,-nbitq), 
to_sfixed(-149170863.0/4294967296.0,1,-nbitq), 
to_sfixed(-413732506.0/4294967296.0,1,-nbitq), 
to_sfixed(65072977.0/4294967296.0,1,-nbitq), 
to_sfixed(-107312856.0/4294967296.0,1,-nbitq), 
to_sfixed(168364700.0/4294967296.0,1,-nbitq), 
to_sfixed(147027906.0/4294967296.0,1,-nbitq), 
to_sfixed(-40676812.0/4294967296.0,1,-nbitq), 
to_sfixed(307362302.0/4294967296.0,1,-nbitq), 
to_sfixed(355667926.0/4294967296.0,1,-nbitq), 
to_sfixed(266347235.0/4294967296.0,1,-nbitq), 
to_sfixed(-307307211.0/4294967296.0,1,-nbitq), 
to_sfixed(126679673.0/4294967296.0,1,-nbitq), 
to_sfixed(303464769.0/4294967296.0,1,-nbitq), 
to_sfixed(-10341151.0/4294967296.0,1,-nbitq), 
to_sfixed(-182366571.0/4294967296.0,1,-nbitq), 
to_sfixed(136358242.0/4294967296.0,1,-nbitq), 
to_sfixed(-427158966.0/4294967296.0,1,-nbitq), 
to_sfixed(380361022.0/4294967296.0,1,-nbitq), 
to_sfixed(-192874951.0/4294967296.0,1,-nbitq), 
to_sfixed(-40207885.0/4294967296.0,1,-nbitq), 
to_sfixed(289782644.0/4294967296.0,1,-nbitq), 
to_sfixed(41445207.0/4294967296.0,1,-nbitq), 
to_sfixed(-104589195.0/4294967296.0,1,-nbitq), 
to_sfixed(-401655655.0/4294967296.0,1,-nbitq), 
to_sfixed(-261886013.0/4294967296.0,1,-nbitq), 
to_sfixed(101460298.0/4294967296.0,1,-nbitq), 
to_sfixed(-309607266.0/4294967296.0,1,-nbitq), 
to_sfixed(-226898172.0/4294967296.0,1,-nbitq), 
to_sfixed(10619726.0/4294967296.0,1,-nbitq), 
to_sfixed(82151993.0/4294967296.0,1,-nbitq), 
to_sfixed(40258906.0/4294967296.0,1,-nbitq), 
to_sfixed(-517907032.0/4294967296.0,1,-nbitq), 
to_sfixed(-496339664.0/4294967296.0,1,-nbitq), 
to_sfixed(189172248.0/4294967296.0,1,-nbitq), 
to_sfixed(-488421059.0/4294967296.0,1,-nbitq), 
to_sfixed(-300067555.0/4294967296.0,1,-nbitq), 
to_sfixed(-343209621.0/4294967296.0,1,-nbitq), 
to_sfixed(-403651139.0/4294967296.0,1,-nbitq), 
to_sfixed(-268364615.0/4294967296.0,1,-nbitq), 
to_sfixed(13193406.0/4294967296.0,1,-nbitq), 
to_sfixed(458852122.0/4294967296.0,1,-nbitq), 
to_sfixed(-40927509.0/4294967296.0,1,-nbitq), 
to_sfixed(-153344243.0/4294967296.0,1,-nbitq), 
to_sfixed(-155825870.0/4294967296.0,1,-nbitq), 
to_sfixed(-272134920.0/4294967296.0,1,-nbitq), 
to_sfixed(279427355.0/4294967296.0,1,-nbitq), 
to_sfixed(-73724605.0/4294967296.0,1,-nbitq), 
to_sfixed(262009552.0/4294967296.0,1,-nbitq), 
to_sfixed(191810608.0/4294967296.0,1,-nbitq), 
to_sfixed(274835578.0/4294967296.0,1,-nbitq), 
to_sfixed(189753352.0/4294967296.0,1,-nbitq), 
to_sfixed(287888974.0/4294967296.0,1,-nbitq), 
to_sfixed(120191554.0/4294967296.0,1,-nbitq), 
to_sfixed(10560483.0/4294967296.0,1,-nbitq), 
to_sfixed(-5736739.0/4294967296.0,1,-nbitq), 
to_sfixed(820486391.0/4294967296.0,1,-nbitq), 
to_sfixed(-204725676.0/4294967296.0,1,-nbitq), 
to_sfixed(-229835197.0/4294967296.0,1,-nbitq), 
to_sfixed(549581886.0/4294967296.0,1,-nbitq), 
to_sfixed(-127638579.0/4294967296.0,1,-nbitq), 
to_sfixed(-127171272.0/4294967296.0,1,-nbitq), 
to_sfixed(482573433.0/4294967296.0,1,-nbitq), 
to_sfixed(359321759.0/4294967296.0,1,-nbitq), 
to_sfixed(168471349.0/4294967296.0,1,-nbitq), 
to_sfixed(-157380666.0/4294967296.0,1,-nbitq), 
to_sfixed(-64391589.0/4294967296.0,1,-nbitq), 
to_sfixed(-427982156.0/4294967296.0,1,-nbitq), 
to_sfixed(-168054431.0/4294967296.0,1,-nbitq), 
to_sfixed(-103536261.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(81218944.0/4294967296.0,1,-nbitq), 
to_sfixed(-424671325.0/4294967296.0,1,-nbitq), 
to_sfixed(-264307416.0/4294967296.0,1,-nbitq), 
to_sfixed(-340365344.0/4294967296.0,1,-nbitq), 
to_sfixed(-64054846.0/4294967296.0,1,-nbitq), 
to_sfixed(-457221890.0/4294967296.0,1,-nbitq), 
to_sfixed(-329695737.0/4294967296.0,1,-nbitq), 
to_sfixed(8593489.0/4294967296.0,1,-nbitq), 
to_sfixed(-187739589.0/4294967296.0,1,-nbitq), 
to_sfixed(143581404.0/4294967296.0,1,-nbitq), 
to_sfixed(254968210.0/4294967296.0,1,-nbitq), 
to_sfixed(84128526.0/4294967296.0,1,-nbitq), 
to_sfixed(34423602.0/4294967296.0,1,-nbitq), 
to_sfixed(284310917.0/4294967296.0,1,-nbitq), 
to_sfixed(33684837.0/4294967296.0,1,-nbitq), 
to_sfixed(-94559076.0/4294967296.0,1,-nbitq), 
to_sfixed(-140488111.0/4294967296.0,1,-nbitq), 
to_sfixed(134786075.0/4294967296.0,1,-nbitq), 
to_sfixed(-80666503.0/4294967296.0,1,-nbitq), 
to_sfixed(-215498976.0/4294967296.0,1,-nbitq), 
to_sfixed(-269842738.0/4294967296.0,1,-nbitq), 
to_sfixed(-58755015.0/4294967296.0,1,-nbitq), 
to_sfixed(161139927.0/4294967296.0,1,-nbitq), 
to_sfixed(-65540055.0/4294967296.0,1,-nbitq), 
to_sfixed(197679143.0/4294967296.0,1,-nbitq), 
to_sfixed(-363247000.0/4294967296.0,1,-nbitq), 
to_sfixed(-128219131.0/4294967296.0,1,-nbitq), 
to_sfixed(118206416.0/4294967296.0,1,-nbitq), 
to_sfixed(26903343.0/4294967296.0,1,-nbitq), 
to_sfixed(252324695.0/4294967296.0,1,-nbitq), 
to_sfixed(-241664628.0/4294967296.0,1,-nbitq), 
to_sfixed(-36145913.0/4294967296.0,1,-nbitq), 
to_sfixed(-192380612.0/4294967296.0,1,-nbitq), 
to_sfixed(-462511620.0/4294967296.0,1,-nbitq), 
to_sfixed(-550501035.0/4294967296.0,1,-nbitq), 
to_sfixed(38534620.0/4294967296.0,1,-nbitq), 
to_sfixed(-498679403.0/4294967296.0,1,-nbitq), 
to_sfixed(83872885.0/4294967296.0,1,-nbitq), 
to_sfixed(224060728.0/4294967296.0,1,-nbitq), 
to_sfixed(102296210.0/4294967296.0,1,-nbitq), 
to_sfixed(446399099.0/4294967296.0,1,-nbitq), 
to_sfixed(-207364990.0/4294967296.0,1,-nbitq), 
to_sfixed(-46819089.0/4294967296.0,1,-nbitq), 
to_sfixed(-412370605.0/4294967296.0,1,-nbitq), 
to_sfixed(-127031174.0/4294967296.0,1,-nbitq), 
to_sfixed(-149233397.0/4294967296.0,1,-nbitq), 
to_sfixed(-390508444.0/4294967296.0,1,-nbitq), 
to_sfixed(9129594.0/4294967296.0,1,-nbitq), 
to_sfixed(-378291551.0/4294967296.0,1,-nbitq), 
to_sfixed(131097263.0/4294967296.0,1,-nbitq), 
to_sfixed(198374603.0/4294967296.0,1,-nbitq), 
to_sfixed(-295477151.0/4294967296.0,1,-nbitq), 
to_sfixed(216527047.0/4294967296.0,1,-nbitq), 
to_sfixed(74711258.0/4294967296.0,1,-nbitq), 
to_sfixed(446974931.0/4294967296.0,1,-nbitq), 
to_sfixed(221140310.0/4294967296.0,1,-nbitq), 
to_sfixed(535992221.0/4294967296.0,1,-nbitq), 
to_sfixed(-292715535.0/4294967296.0,1,-nbitq), 
to_sfixed(7639014.0/4294967296.0,1,-nbitq), 
to_sfixed(42019037.0/4294967296.0,1,-nbitq), 
to_sfixed(-123055790.0/4294967296.0,1,-nbitq), 
to_sfixed(38199522.0/4294967296.0,1,-nbitq), 
to_sfixed(-114768568.0/4294967296.0,1,-nbitq), 
to_sfixed(-180510627.0/4294967296.0,1,-nbitq), 
to_sfixed(-157002765.0/4294967296.0,1,-nbitq), 
to_sfixed(-100279692.0/4294967296.0,1,-nbitq), 
to_sfixed(844171496.0/4294967296.0,1,-nbitq), 
to_sfixed(182968718.0/4294967296.0,1,-nbitq), 
to_sfixed(-199148971.0/4294967296.0,1,-nbitq), 
to_sfixed(-16287859.0/4294967296.0,1,-nbitq), 
to_sfixed(-433871798.0/4294967296.0,1,-nbitq), 
to_sfixed(-334343628.0/4294967296.0,1,-nbitq), 
to_sfixed(-187682172.0/4294967296.0,1,-nbitq), 
to_sfixed(-7841747.0/4294967296.0,1,-nbitq), 
to_sfixed(95331385.0/4294967296.0,1,-nbitq), 
to_sfixed(-67925292.0/4294967296.0,1,-nbitq), 
to_sfixed(-205033555.0/4294967296.0,1,-nbitq), 
to_sfixed(-378885348.0/4294967296.0,1,-nbitq), 
to_sfixed(342211631.0/4294967296.0,1,-nbitq), 
to_sfixed(246084276.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-373819852.0/4294967296.0,1,-nbitq), 
to_sfixed(121259243.0/4294967296.0,1,-nbitq), 
to_sfixed(507867596.0/4294967296.0,1,-nbitq), 
to_sfixed(-528064168.0/4294967296.0,1,-nbitq), 
to_sfixed(-199302116.0/4294967296.0,1,-nbitq), 
to_sfixed(255194691.0/4294967296.0,1,-nbitq), 
to_sfixed(-280535694.0/4294967296.0,1,-nbitq), 
to_sfixed(-173666659.0/4294967296.0,1,-nbitq), 
to_sfixed(263922999.0/4294967296.0,1,-nbitq), 
to_sfixed(-18503443.0/4294967296.0,1,-nbitq), 
to_sfixed(-352794268.0/4294967296.0,1,-nbitq), 
to_sfixed(-262070450.0/4294967296.0,1,-nbitq), 
to_sfixed(105793212.0/4294967296.0,1,-nbitq), 
to_sfixed(460711978.0/4294967296.0,1,-nbitq), 
to_sfixed(-114965650.0/4294967296.0,1,-nbitq), 
to_sfixed(-321285643.0/4294967296.0,1,-nbitq), 
to_sfixed(255022082.0/4294967296.0,1,-nbitq), 
to_sfixed(-37029421.0/4294967296.0,1,-nbitq), 
to_sfixed(-108763994.0/4294967296.0,1,-nbitq), 
to_sfixed(35720032.0/4294967296.0,1,-nbitq), 
to_sfixed(-7109728.0/4294967296.0,1,-nbitq), 
to_sfixed(-336265599.0/4294967296.0,1,-nbitq), 
to_sfixed(485288300.0/4294967296.0,1,-nbitq), 
to_sfixed(-28470425.0/4294967296.0,1,-nbitq), 
to_sfixed(131930105.0/4294967296.0,1,-nbitq), 
to_sfixed(420929154.0/4294967296.0,1,-nbitq), 
to_sfixed(-78142387.0/4294967296.0,1,-nbitq), 
to_sfixed(-644491467.0/4294967296.0,1,-nbitq), 
to_sfixed(338372771.0/4294967296.0,1,-nbitq), 
to_sfixed(-327286233.0/4294967296.0,1,-nbitq), 
to_sfixed(-505299344.0/4294967296.0,1,-nbitq), 
to_sfixed(-231204492.0/4294967296.0,1,-nbitq), 
to_sfixed(29102256.0/4294967296.0,1,-nbitq), 
to_sfixed(-271553656.0/4294967296.0,1,-nbitq), 
to_sfixed(-37787679.0/4294967296.0,1,-nbitq), 
to_sfixed(-297451603.0/4294967296.0,1,-nbitq), 
to_sfixed(-22146508.0/4294967296.0,1,-nbitq), 
to_sfixed(288119553.0/4294967296.0,1,-nbitq), 
to_sfixed(-202871199.0/4294967296.0,1,-nbitq), 
to_sfixed(-84100659.0/4294967296.0,1,-nbitq), 
to_sfixed(129928850.0/4294967296.0,1,-nbitq), 
to_sfixed(-121176971.0/4294967296.0,1,-nbitq), 
to_sfixed(293545163.0/4294967296.0,1,-nbitq), 
to_sfixed(-12195671.0/4294967296.0,1,-nbitq), 
to_sfixed(-188974254.0/4294967296.0,1,-nbitq), 
to_sfixed(-69859649.0/4294967296.0,1,-nbitq), 
to_sfixed(50491115.0/4294967296.0,1,-nbitq), 
to_sfixed(165306054.0/4294967296.0,1,-nbitq), 
to_sfixed(-76372265.0/4294967296.0,1,-nbitq), 
to_sfixed(76403246.0/4294967296.0,1,-nbitq), 
to_sfixed(186996053.0/4294967296.0,1,-nbitq), 
to_sfixed(24376986.0/4294967296.0,1,-nbitq), 
to_sfixed(229146233.0/4294967296.0,1,-nbitq), 
to_sfixed(137349543.0/4294967296.0,1,-nbitq), 
to_sfixed(-62674669.0/4294967296.0,1,-nbitq), 
to_sfixed(390229.0/4294967296.0,1,-nbitq), 
to_sfixed(427143377.0/4294967296.0,1,-nbitq), 
to_sfixed(-126654514.0/4294967296.0,1,-nbitq), 
to_sfixed(-330542806.0/4294967296.0,1,-nbitq), 
to_sfixed(346720158.0/4294967296.0,1,-nbitq), 
to_sfixed(327873767.0/4294967296.0,1,-nbitq), 
to_sfixed(-3666501.0/4294967296.0,1,-nbitq), 
to_sfixed(-447856032.0/4294967296.0,1,-nbitq), 
to_sfixed(-3588519.0/4294967296.0,1,-nbitq), 
to_sfixed(156874703.0/4294967296.0,1,-nbitq), 
to_sfixed(-278794641.0/4294967296.0,1,-nbitq), 
to_sfixed(756357404.0/4294967296.0,1,-nbitq), 
to_sfixed(266313518.0/4294967296.0,1,-nbitq), 
to_sfixed(263775595.0/4294967296.0,1,-nbitq), 
to_sfixed(537177547.0/4294967296.0,1,-nbitq), 
to_sfixed(155986187.0/4294967296.0,1,-nbitq), 
to_sfixed(-350576375.0/4294967296.0,1,-nbitq), 
to_sfixed(268660454.0/4294967296.0,1,-nbitq), 
to_sfixed(-4378396.0/4294967296.0,1,-nbitq), 
to_sfixed(157312244.0/4294967296.0,1,-nbitq), 
to_sfixed(-132354406.0/4294967296.0,1,-nbitq), 
to_sfixed(52947935.0/4294967296.0,1,-nbitq), 
to_sfixed(-292521105.0/4294967296.0,1,-nbitq), 
to_sfixed(-240084641.0/4294967296.0,1,-nbitq), 
to_sfixed(355948944.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(282666197.0/4294967296.0,1,-nbitq), 
to_sfixed(296300954.0/4294967296.0,1,-nbitq), 
to_sfixed(403287120.0/4294967296.0,1,-nbitq), 
to_sfixed(-520795001.0/4294967296.0,1,-nbitq), 
to_sfixed(405246633.0/4294967296.0,1,-nbitq), 
to_sfixed(-247060144.0/4294967296.0,1,-nbitq), 
to_sfixed(411497569.0/4294967296.0,1,-nbitq), 
to_sfixed(183734659.0/4294967296.0,1,-nbitq), 
to_sfixed(-168527409.0/4294967296.0,1,-nbitq), 
to_sfixed(-343758792.0/4294967296.0,1,-nbitq), 
to_sfixed(-109241896.0/4294967296.0,1,-nbitq), 
to_sfixed(2175680.0/4294967296.0,1,-nbitq), 
to_sfixed(529158123.0/4294967296.0,1,-nbitq), 
to_sfixed(14906735.0/4294967296.0,1,-nbitq), 
to_sfixed(-271109155.0/4294967296.0,1,-nbitq), 
to_sfixed(-138228084.0/4294967296.0,1,-nbitq), 
to_sfixed(-223073398.0/4294967296.0,1,-nbitq), 
to_sfixed(272778942.0/4294967296.0,1,-nbitq), 
to_sfixed(278769972.0/4294967296.0,1,-nbitq), 
to_sfixed(-78119618.0/4294967296.0,1,-nbitq), 
to_sfixed(-327621119.0/4294967296.0,1,-nbitq), 
to_sfixed(58428726.0/4294967296.0,1,-nbitq), 
to_sfixed(154290496.0/4294967296.0,1,-nbitq), 
to_sfixed(270482011.0/4294967296.0,1,-nbitq), 
to_sfixed(-100798407.0/4294967296.0,1,-nbitq), 
to_sfixed(460400764.0/4294967296.0,1,-nbitq), 
to_sfixed(-185927439.0/4294967296.0,1,-nbitq), 
to_sfixed(-396766353.0/4294967296.0,1,-nbitq), 
to_sfixed(-130378230.0/4294967296.0,1,-nbitq), 
to_sfixed(88688281.0/4294967296.0,1,-nbitq), 
to_sfixed(4400990.0/4294967296.0,1,-nbitq), 
to_sfixed(-327755363.0/4294967296.0,1,-nbitq), 
to_sfixed(-161506267.0/4294967296.0,1,-nbitq), 
to_sfixed(95010635.0/4294967296.0,1,-nbitq), 
to_sfixed(330514911.0/4294967296.0,1,-nbitq), 
to_sfixed(63207729.0/4294967296.0,1,-nbitq), 
to_sfixed(-266618240.0/4294967296.0,1,-nbitq), 
to_sfixed(-62752042.0/4294967296.0,1,-nbitq), 
to_sfixed(-474416031.0/4294967296.0,1,-nbitq), 
to_sfixed(220795661.0/4294967296.0,1,-nbitq), 
to_sfixed(9503456.0/4294967296.0,1,-nbitq), 
to_sfixed(67408531.0/4294967296.0,1,-nbitq), 
to_sfixed(135671902.0/4294967296.0,1,-nbitq), 
to_sfixed(87086328.0/4294967296.0,1,-nbitq), 
to_sfixed(149387677.0/4294967296.0,1,-nbitq), 
to_sfixed(-426885136.0/4294967296.0,1,-nbitq), 
to_sfixed(-18077450.0/4294967296.0,1,-nbitq), 
to_sfixed(-282942009.0/4294967296.0,1,-nbitq), 
to_sfixed(257891960.0/4294967296.0,1,-nbitq), 
to_sfixed(-195712586.0/4294967296.0,1,-nbitq), 
to_sfixed(55661421.0/4294967296.0,1,-nbitq), 
to_sfixed(-198557237.0/4294967296.0,1,-nbitq), 
to_sfixed(-139367604.0/4294967296.0,1,-nbitq), 
to_sfixed(-23220695.0/4294967296.0,1,-nbitq), 
to_sfixed(53954092.0/4294967296.0,1,-nbitq), 
to_sfixed(296519011.0/4294967296.0,1,-nbitq), 
to_sfixed(-2504885.0/4294967296.0,1,-nbitq), 
to_sfixed(268269168.0/4294967296.0,1,-nbitq), 
to_sfixed(373157018.0/4294967296.0,1,-nbitq), 
to_sfixed(386970451.0/4294967296.0,1,-nbitq), 
to_sfixed(-191438075.0/4294967296.0,1,-nbitq), 
to_sfixed(-49843959.0/4294967296.0,1,-nbitq), 
to_sfixed(-228622951.0/4294967296.0,1,-nbitq), 
to_sfixed(-238197945.0/4294967296.0,1,-nbitq), 
to_sfixed(-427495472.0/4294967296.0,1,-nbitq), 
to_sfixed(-323601433.0/4294967296.0,1,-nbitq), 
to_sfixed(293242456.0/4294967296.0,1,-nbitq), 
to_sfixed(129431004.0/4294967296.0,1,-nbitq), 
to_sfixed(-256652065.0/4294967296.0,1,-nbitq), 
to_sfixed(4989587.0/4294967296.0,1,-nbitq), 
to_sfixed(337237712.0/4294967296.0,1,-nbitq), 
to_sfixed(223369312.0/4294967296.0,1,-nbitq), 
to_sfixed(-208993066.0/4294967296.0,1,-nbitq), 
to_sfixed(-340139285.0/4294967296.0,1,-nbitq), 
to_sfixed(-9861337.0/4294967296.0,1,-nbitq), 
to_sfixed(122842683.0/4294967296.0,1,-nbitq), 
to_sfixed(-510068151.0/4294967296.0,1,-nbitq), 
to_sfixed(-361036263.0/4294967296.0,1,-nbitq), 
to_sfixed(-347079986.0/4294967296.0,1,-nbitq), 
to_sfixed(-87019711.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-224965574.0/4294967296.0,1,-nbitq), 
to_sfixed(130242147.0/4294967296.0,1,-nbitq), 
to_sfixed(353835474.0/4294967296.0,1,-nbitq), 
to_sfixed(-569781394.0/4294967296.0,1,-nbitq), 
to_sfixed(226427779.0/4294967296.0,1,-nbitq), 
to_sfixed(-411495420.0/4294967296.0,1,-nbitq), 
to_sfixed(-195488554.0/4294967296.0,1,-nbitq), 
to_sfixed(481125861.0/4294967296.0,1,-nbitq), 
to_sfixed(-262521236.0/4294967296.0,1,-nbitq), 
to_sfixed(-305848616.0/4294967296.0,1,-nbitq), 
to_sfixed(44089175.0/4294967296.0,1,-nbitq), 
to_sfixed(-327359641.0/4294967296.0,1,-nbitq), 
to_sfixed(248482688.0/4294967296.0,1,-nbitq), 
to_sfixed(468854637.0/4294967296.0,1,-nbitq), 
to_sfixed(335914120.0/4294967296.0,1,-nbitq), 
to_sfixed(-175123190.0/4294967296.0,1,-nbitq), 
to_sfixed(-401346521.0/4294967296.0,1,-nbitq), 
to_sfixed(248194188.0/4294967296.0,1,-nbitq), 
to_sfixed(162762718.0/4294967296.0,1,-nbitq), 
to_sfixed(-94276391.0/4294967296.0,1,-nbitq), 
to_sfixed(367808040.0/4294967296.0,1,-nbitq), 
to_sfixed(-59947658.0/4294967296.0,1,-nbitq), 
to_sfixed(129601937.0/4294967296.0,1,-nbitq), 
to_sfixed(-94397686.0/4294967296.0,1,-nbitq), 
to_sfixed(275729398.0/4294967296.0,1,-nbitq), 
to_sfixed(555804866.0/4294967296.0,1,-nbitq), 
to_sfixed(-215105359.0/4294967296.0,1,-nbitq), 
to_sfixed(33851848.0/4294967296.0,1,-nbitq), 
to_sfixed(382048422.0/4294967296.0,1,-nbitq), 
to_sfixed(-115175533.0/4294967296.0,1,-nbitq), 
to_sfixed(-229925641.0/4294967296.0,1,-nbitq), 
to_sfixed(-207382583.0/4294967296.0,1,-nbitq), 
to_sfixed(197743130.0/4294967296.0,1,-nbitq), 
to_sfixed(-64500164.0/4294967296.0,1,-nbitq), 
to_sfixed(355767252.0/4294967296.0,1,-nbitq), 
to_sfixed(-165880223.0/4294967296.0,1,-nbitq), 
to_sfixed(-91111389.0/4294967296.0,1,-nbitq), 
to_sfixed(-73336023.0/4294967296.0,1,-nbitq), 
to_sfixed(279199699.0/4294967296.0,1,-nbitq), 
to_sfixed(114035453.0/4294967296.0,1,-nbitq), 
to_sfixed(-68075603.0/4294967296.0,1,-nbitq), 
to_sfixed(-497466423.0/4294967296.0,1,-nbitq), 
to_sfixed(-93362028.0/4294967296.0,1,-nbitq), 
to_sfixed(-92327486.0/4294967296.0,1,-nbitq), 
to_sfixed(-304340253.0/4294967296.0,1,-nbitq), 
to_sfixed(305359822.0/4294967296.0,1,-nbitq), 
to_sfixed(17937592.0/4294967296.0,1,-nbitq), 
to_sfixed(-87146779.0/4294967296.0,1,-nbitq), 
to_sfixed(-80775180.0/4294967296.0,1,-nbitq), 
to_sfixed(-39151990.0/4294967296.0,1,-nbitq), 
to_sfixed(-397159028.0/4294967296.0,1,-nbitq), 
to_sfixed(-37694530.0/4294967296.0,1,-nbitq), 
to_sfixed(-644971054.0/4294967296.0,1,-nbitq), 
to_sfixed(242086571.0/4294967296.0,1,-nbitq), 
to_sfixed(13988531.0/4294967296.0,1,-nbitq), 
to_sfixed(-76734580.0/4294967296.0,1,-nbitq), 
to_sfixed(313973671.0/4294967296.0,1,-nbitq), 
to_sfixed(-571284243.0/4294967296.0,1,-nbitq), 
to_sfixed(-56514000.0/4294967296.0,1,-nbitq), 
to_sfixed(368459410.0/4294967296.0,1,-nbitq), 
to_sfixed(-32543612.0/4294967296.0,1,-nbitq), 
to_sfixed(471828348.0/4294967296.0,1,-nbitq), 
to_sfixed(207768077.0/4294967296.0,1,-nbitq), 
to_sfixed(8611463.0/4294967296.0,1,-nbitq), 
to_sfixed(-424800341.0/4294967296.0,1,-nbitq), 
to_sfixed(-187094785.0/4294967296.0,1,-nbitq), 
to_sfixed(508300773.0/4294967296.0,1,-nbitq), 
to_sfixed(388983572.0/4294967296.0,1,-nbitq), 
to_sfixed(-285599405.0/4294967296.0,1,-nbitq), 
to_sfixed(6205230.0/4294967296.0,1,-nbitq), 
to_sfixed(454185281.0/4294967296.0,1,-nbitq), 
to_sfixed(-102362077.0/4294967296.0,1,-nbitq), 
to_sfixed(226191529.0/4294967296.0,1,-nbitq), 
to_sfixed(436983985.0/4294967296.0,1,-nbitq), 
to_sfixed(-29654126.0/4294967296.0,1,-nbitq), 
to_sfixed(-304194808.0/4294967296.0,1,-nbitq), 
to_sfixed(-591438267.0/4294967296.0,1,-nbitq), 
to_sfixed(56764395.0/4294967296.0,1,-nbitq), 
to_sfixed(285458879.0/4294967296.0,1,-nbitq), 
to_sfixed(335212193.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(73568806.0/4294967296.0,1,-nbitq), 
to_sfixed(154051559.0/4294967296.0,1,-nbitq), 
to_sfixed(731434917.0/4294967296.0,1,-nbitq), 
to_sfixed(-424219613.0/4294967296.0,1,-nbitq), 
to_sfixed(110009598.0/4294967296.0,1,-nbitq), 
to_sfixed(-343585773.0/4294967296.0,1,-nbitq), 
to_sfixed(172985427.0/4294967296.0,1,-nbitq), 
to_sfixed(-80088705.0/4294967296.0,1,-nbitq), 
to_sfixed(-984486978.0/4294967296.0,1,-nbitq), 
to_sfixed(276378462.0/4294967296.0,1,-nbitq), 
to_sfixed(-123384776.0/4294967296.0,1,-nbitq), 
to_sfixed(119307657.0/4294967296.0,1,-nbitq), 
to_sfixed(956308483.0/4294967296.0,1,-nbitq), 
to_sfixed(821557025.0/4294967296.0,1,-nbitq), 
to_sfixed(-137910712.0/4294967296.0,1,-nbitq), 
to_sfixed(519240207.0/4294967296.0,1,-nbitq), 
to_sfixed(313420417.0/4294967296.0,1,-nbitq), 
to_sfixed(-257495972.0/4294967296.0,1,-nbitq), 
to_sfixed(184626342.0/4294967296.0,1,-nbitq), 
to_sfixed(419863138.0/4294967296.0,1,-nbitq), 
to_sfixed(103663226.0/4294967296.0,1,-nbitq), 
to_sfixed(-87534915.0/4294967296.0,1,-nbitq), 
to_sfixed(-232367887.0/4294967296.0,1,-nbitq), 
to_sfixed(604315551.0/4294967296.0,1,-nbitq), 
to_sfixed(-73308159.0/4294967296.0,1,-nbitq), 
to_sfixed(314981857.0/4294967296.0,1,-nbitq), 
to_sfixed(356333318.0/4294967296.0,1,-nbitq), 
to_sfixed(-294387945.0/4294967296.0,1,-nbitq), 
to_sfixed(-160103365.0/4294967296.0,1,-nbitq), 
to_sfixed(314580774.0/4294967296.0,1,-nbitq), 
to_sfixed(-128465771.0/4294967296.0,1,-nbitq), 
to_sfixed(465036710.0/4294967296.0,1,-nbitq), 
to_sfixed(-282710908.0/4294967296.0,1,-nbitq), 
to_sfixed(13100479.0/4294967296.0,1,-nbitq), 
to_sfixed(-166100078.0/4294967296.0,1,-nbitq), 
to_sfixed(-35811706.0/4294967296.0,1,-nbitq), 
to_sfixed(27470855.0/4294967296.0,1,-nbitq), 
to_sfixed(-530550345.0/4294967296.0,1,-nbitq), 
to_sfixed(-228092917.0/4294967296.0,1,-nbitq), 
to_sfixed(53511230.0/4294967296.0,1,-nbitq), 
to_sfixed(146739372.0/4294967296.0,1,-nbitq), 
to_sfixed(-245474189.0/4294967296.0,1,-nbitq), 
to_sfixed(-189133288.0/4294967296.0,1,-nbitq), 
to_sfixed(-225614025.0/4294967296.0,1,-nbitq), 
to_sfixed(231938268.0/4294967296.0,1,-nbitq), 
to_sfixed(-322791009.0/4294967296.0,1,-nbitq), 
to_sfixed(-356477203.0/4294967296.0,1,-nbitq), 
to_sfixed(20326561.0/4294967296.0,1,-nbitq), 
to_sfixed(-191643810.0/4294967296.0,1,-nbitq), 
to_sfixed(209150293.0/4294967296.0,1,-nbitq), 
to_sfixed(-243591539.0/4294967296.0,1,-nbitq), 
to_sfixed(-57098525.0/4294967296.0,1,-nbitq), 
to_sfixed(116472976.0/4294967296.0,1,-nbitq), 
to_sfixed(84073973.0/4294967296.0,1,-nbitq), 
to_sfixed(798707576.0/4294967296.0,1,-nbitq), 
to_sfixed(84155458.0/4294967296.0,1,-nbitq), 
to_sfixed(168556360.0/4294967296.0,1,-nbitq), 
to_sfixed(-351192968.0/4294967296.0,1,-nbitq), 
to_sfixed(-216162306.0/4294967296.0,1,-nbitq), 
to_sfixed(-265445275.0/4294967296.0,1,-nbitq), 
to_sfixed(123619463.0/4294967296.0,1,-nbitq), 
to_sfixed(229065699.0/4294967296.0,1,-nbitq), 
to_sfixed(-328109145.0/4294967296.0,1,-nbitq), 
to_sfixed(348126958.0/4294967296.0,1,-nbitq), 
to_sfixed(184631834.0/4294967296.0,1,-nbitq), 
to_sfixed(-156695246.0/4294967296.0,1,-nbitq), 
to_sfixed(36356303.0/4294967296.0,1,-nbitq), 
to_sfixed(2063894.0/4294967296.0,1,-nbitq), 
to_sfixed(-244302674.0/4294967296.0,1,-nbitq), 
to_sfixed(326948303.0/4294967296.0,1,-nbitq), 
to_sfixed(435129193.0/4294967296.0,1,-nbitq), 
to_sfixed(218415499.0/4294967296.0,1,-nbitq), 
to_sfixed(-128314321.0/4294967296.0,1,-nbitq), 
to_sfixed(429887132.0/4294967296.0,1,-nbitq), 
to_sfixed(484096979.0/4294967296.0,1,-nbitq), 
to_sfixed(-291379277.0/4294967296.0,1,-nbitq), 
to_sfixed(-39392759.0/4294967296.0,1,-nbitq), 
to_sfixed(-405612749.0/4294967296.0,1,-nbitq), 
to_sfixed(-16708136.0/4294967296.0,1,-nbitq), 
to_sfixed(-367407341.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-193247142.0/4294967296.0,1,-nbitq), 
to_sfixed(-385318545.0/4294967296.0,1,-nbitq), 
to_sfixed(1000650130.0/4294967296.0,1,-nbitq), 
to_sfixed(-1102812485.0/4294967296.0,1,-nbitq), 
to_sfixed(-1037086865.0/4294967296.0,1,-nbitq), 
to_sfixed(-154224948.0/4294967296.0,1,-nbitq), 
to_sfixed(323977381.0/4294967296.0,1,-nbitq), 
to_sfixed(-659657901.0/4294967296.0,1,-nbitq), 
to_sfixed(-1355689619.0/4294967296.0,1,-nbitq), 
to_sfixed(-15106814.0/4294967296.0,1,-nbitq), 
to_sfixed(-62210637.0/4294967296.0,1,-nbitq), 
to_sfixed(30944727.0/4294967296.0,1,-nbitq), 
to_sfixed(1534020136.0/4294967296.0,1,-nbitq), 
to_sfixed(1086297647.0/4294967296.0,1,-nbitq), 
to_sfixed(57954341.0/4294967296.0,1,-nbitq), 
to_sfixed(914580298.0/4294967296.0,1,-nbitq), 
to_sfixed(-48494750.0/4294967296.0,1,-nbitq), 
to_sfixed(381244780.0/4294967296.0,1,-nbitq), 
to_sfixed(-513244706.0/4294967296.0,1,-nbitq), 
to_sfixed(771354900.0/4294967296.0,1,-nbitq), 
to_sfixed(-103728308.0/4294967296.0,1,-nbitq), 
to_sfixed(-457325299.0/4294967296.0,1,-nbitq), 
to_sfixed(-618689741.0/4294967296.0,1,-nbitq), 
to_sfixed(1419404142.0/4294967296.0,1,-nbitq), 
to_sfixed(321563396.0/4294967296.0,1,-nbitq), 
to_sfixed(279612421.0/4294967296.0,1,-nbitq), 
to_sfixed(-174199417.0/4294967296.0,1,-nbitq), 
to_sfixed(-422034266.0/4294967296.0,1,-nbitq), 
to_sfixed(-78886244.0/4294967296.0,1,-nbitq), 
to_sfixed(527805162.0/4294967296.0,1,-nbitq), 
to_sfixed(-154960835.0/4294967296.0,1,-nbitq), 
to_sfixed(211289757.0/4294967296.0,1,-nbitq), 
to_sfixed(-895561010.0/4294967296.0,1,-nbitq), 
to_sfixed(468830723.0/4294967296.0,1,-nbitq), 
to_sfixed(-86272472.0/4294967296.0,1,-nbitq), 
to_sfixed(956050605.0/4294967296.0,1,-nbitq), 
to_sfixed(302537261.0/4294967296.0,1,-nbitq), 
to_sfixed(-699233827.0/4294967296.0,1,-nbitq), 
to_sfixed(-510456358.0/4294967296.0,1,-nbitq), 
to_sfixed(68133764.0/4294967296.0,1,-nbitq), 
to_sfixed(328142782.0/4294967296.0,1,-nbitq), 
to_sfixed(-858136377.0/4294967296.0,1,-nbitq), 
to_sfixed(-22648586.0/4294967296.0,1,-nbitq), 
to_sfixed(-120135607.0/4294967296.0,1,-nbitq), 
to_sfixed(-365761891.0/4294967296.0,1,-nbitq), 
to_sfixed(-545604966.0/4294967296.0,1,-nbitq), 
to_sfixed(216197963.0/4294967296.0,1,-nbitq), 
to_sfixed(-66882029.0/4294967296.0,1,-nbitq), 
to_sfixed(327182249.0/4294967296.0,1,-nbitq), 
to_sfixed(-39579212.0/4294967296.0,1,-nbitq), 
to_sfixed(33502229.0/4294967296.0,1,-nbitq), 
to_sfixed(-1237915891.0/4294967296.0,1,-nbitq), 
to_sfixed(642775731.0/4294967296.0,1,-nbitq), 
to_sfixed(-911759599.0/4294967296.0,1,-nbitq), 
to_sfixed(612241019.0/4294967296.0,1,-nbitq), 
to_sfixed(-244571253.0/4294967296.0,1,-nbitq), 
to_sfixed(378010064.0/4294967296.0,1,-nbitq), 
to_sfixed(-939504491.0/4294967296.0,1,-nbitq), 
to_sfixed(365820776.0/4294967296.0,1,-nbitq), 
to_sfixed(8174758.0/4294967296.0,1,-nbitq), 
to_sfixed(153170118.0/4294967296.0,1,-nbitq), 
to_sfixed(-420104282.0/4294967296.0,1,-nbitq), 
to_sfixed(-281520994.0/4294967296.0,1,-nbitq), 
to_sfixed(568155789.0/4294967296.0,1,-nbitq), 
to_sfixed(40028546.0/4294967296.0,1,-nbitq), 
to_sfixed(-361087946.0/4294967296.0,1,-nbitq), 
to_sfixed(362894356.0/4294967296.0,1,-nbitq), 
to_sfixed(386497595.0/4294967296.0,1,-nbitq), 
to_sfixed(455593712.0/4294967296.0,1,-nbitq), 
to_sfixed(354289587.0/4294967296.0,1,-nbitq), 
to_sfixed(604348221.0/4294967296.0,1,-nbitq), 
to_sfixed(-333176943.0/4294967296.0,1,-nbitq), 
to_sfixed(-175068490.0/4294967296.0,1,-nbitq), 
to_sfixed(428925338.0/4294967296.0,1,-nbitq), 
to_sfixed(-155065627.0/4294967296.0,1,-nbitq), 
to_sfixed(-15956618.0/4294967296.0,1,-nbitq), 
to_sfixed(41083409.0/4294967296.0,1,-nbitq), 
to_sfixed(62306861.0/4294967296.0,1,-nbitq), 
to_sfixed(990428990.0/4294967296.0,1,-nbitq), 
to_sfixed(-314369607.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-55610011.0/4294967296.0,1,-nbitq), 
to_sfixed(-1187922901.0/4294967296.0,1,-nbitq), 
to_sfixed(510131414.0/4294967296.0,1,-nbitq), 
to_sfixed(-1125079561.0/4294967296.0,1,-nbitq), 
to_sfixed(-958997819.0/4294967296.0,1,-nbitq), 
to_sfixed(558636004.0/4294967296.0,1,-nbitq), 
to_sfixed(-163107322.0/4294967296.0,1,-nbitq), 
to_sfixed(-109613397.0/4294967296.0,1,-nbitq), 
to_sfixed(-1103127736.0/4294967296.0,1,-nbitq), 
to_sfixed(129188450.0/4294967296.0,1,-nbitq), 
to_sfixed(364585870.0/4294967296.0,1,-nbitq), 
to_sfixed(-249378481.0/4294967296.0,1,-nbitq), 
to_sfixed(1798493551.0/4294967296.0,1,-nbitq), 
to_sfixed(1145847692.0/4294967296.0,1,-nbitq), 
to_sfixed(380728020.0/4294967296.0,1,-nbitq), 
to_sfixed(554688080.0/4294967296.0,1,-nbitq), 
to_sfixed(10910958.0/4294967296.0,1,-nbitq), 
to_sfixed(-192060767.0/4294967296.0,1,-nbitq), 
to_sfixed(-1658637818.0/4294967296.0,1,-nbitq), 
to_sfixed(643222195.0/4294967296.0,1,-nbitq), 
to_sfixed(302934089.0/4294967296.0,1,-nbitq), 
to_sfixed(-406063356.0/4294967296.0,1,-nbitq), 
to_sfixed(-722898341.0/4294967296.0,1,-nbitq), 
to_sfixed(1064191356.0/4294967296.0,1,-nbitq), 
to_sfixed(75403306.0/4294967296.0,1,-nbitq), 
to_sfixed(564187451.0/4294967296.0,1,-nbitq), 
to_sfixed(-477551242.0/4294967296.0,1,-nbitq), 
to_sfixed(-477010904.0/4294967296.0,1,-nbitq), 
to_sfixed(115892445.0/4294967296.0,1,-nbitq), 
to_sfixed(588957552.0/4294967296.0,1,-nbitq), 
to_sfixed(-158843270.0/4294967296.0,1,-nbitq), 
to_sfixed(219555570.0/4294967296.0,1,-nbitq), 
to_sfixed(-365696149.0/4294967296.0,1,-nbitq), 
to_sfixed(484420286.0/4294967296.0,1,-nbitq), 
to_sfixed(181361177.0/4294967296.0,1,-nbitq), 
to_sfixed(1276380041.0/4294967296.0,1,-nbitq), 
to_sfixed(75972724.0/4294967296.0,1,-nbitq), 
to_sfixed(-1188594578.0/4294967296.0,1,-nbitq), 
to_sfixed(-531085274.0/4294967296.0,1,-nbitq), 
to_sfixed(-337323224.0/4294967296.0,1,-nbitq), 
to_sfixed(99546806.0/4294967296.0,1,-nbitq), 
to_sfixed(-928430881.0/4294967296.0,1,-nbitq), 
to_sfixed(-323642146.0/4294967296.0,1,-nbitq), 
to_sfixed(-206213781.0/4294967296.0,1,-nbitq), 
to_sfixed(-192597906.0/4294967296.0,1,-nbitq), 
to_sfixed(17035789.0/4294967296.0,1,-nbitq), 
to_sfixed(48709321.0/4294967296.0,1,-nbitq), 
to_sfixed(67599814.0/4294967296.0,1,-nbitq), 
to_sfixed(-397888167.0/4294967296.0,1,-nbitq), 
to_sfixed(243090946.0/4294967296.0,1,-nbitq), 
to_sfixed(-372540176.0/4294967296.0,1,-nbitq), 
to_sfixed(-1461527920.0/4294967296.0,1,-nbitq), 
to_sfixed(1005241200.0/4294967296.0,1,-nbitq), 
to_sfixed(-793112457.0/4294967296.0,1,-nbitq), 
to_sfixed(-81481712.0/4294967296.0,1,-nbitq), 
to_sfixed(-272974021.0/4294967296.0,1,-nbitq), 
to_sfixed(-119830177.0/4294967296.0,1,-nbitq), 
to_sfixed(-770748452.0/4294967296.0,1,-nbitq), 
to_sfixed(-361167450.0/4294967296.0,1,-nbitq), 
to_sfixed(191296535.0/4294967296.0,1,-nbitq), 
to_sfixed(-154857931.0/4294967296.0,1,-nbitq), 
to_sfixed(-607175572.0/4294967296.0,1,-nbitq), 
to_sfixed(-122111832.0/4294967296.0,1,-nbitq), 
to_sfixed(-41029671.0/4294967296.0,1,-nbitq), 
to_sfixed(-25543961.0/4294967296.0,1,-nbitq), 
to_sfixed(-110313930.0/4294967296.0,1,-nbitq), 
to_sfixed(-29823619.0/4294967296.0,1,-nbitq), 
to_sfixed(943515200.0/4294967296.0,1,-nbitq), 
to_sfixed(397397258.0/4294967296.0,1,-nbitq), 
to_sfixed(-533730687.0/4294967296.0,1,-nbitq), 
to_sfixed(645965103.0/4294967296.0,1,-nbitq), 
to_sfixed(-415342470.0/4294967296.0,1,-nbitq), 
to_sfixed(-228676616.0/4294967296.0,1,-nbitq), 
to_sfixed(-88528436.0/4294967296.0,1,-nbitq), 
to_sfixed(-206386559.0/4294967296.0,1,-nbitq), 
to_sfixed(333116859.0/4294967296.0,1,-nbitq), 
to_sfixed(287876493.0/4294967296.0,1,-nbitq), 
to_sfixed(54498460.0/4294967296.0,1,-nbitq), 
to_sfixed(695459744.0/4294967296.0,1,-nbitq), 
to_sfixed(2276348.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(582628502.0/4294967296.0,1,-nbitq), 
to_sfixed(-629638703.0/4294967296.0,1,-nbitq), 
to_sfixed(-372230963.0/4294967296.0,1,-nbitq), 
to_sfixed(-1314835543.0/4294967296.0,1,-nbitq), 
to_sfixed(-679048923.0/4294967296.0,1,-nbitq), 
to_sfixed(959481068.0/4294967296.0,1,-nbitq), 
to_sfixed(83122511.0/4294967296.0,1,-nbitq), 
to_sfixed(585257533.0/4294967296.0,1,-nbitq), 
to_sfixed(-603958975.0/4294967296.0,1,-nbitq), 
to_sfixed(254757468.0/4294967296.0,1,-nbitq), 
to_sfixed(-53575989.0/4294967296.0,1,-nbitq), 
to_sfixed(691690562.0/4294967296.0,1,-nbitq), 
to_sfixed(960280737.0/4294967296.0,1,-nbitq), 
to_sfixed(947304930.0/4294967296.0,1,-nbitq), 
to_sfixed(419994155.0/4294967296.0,1,-nbitq), 
to_sfixed(515070618.0/4294967296.0,1,-nbitq), 
to_sfixed(6793244.0/4294967296.0,1,-nbitq), 
to_sfixed(-90992990.0/4294967296.0,1,-nbitq), 
to_sfixed(-1087593966.0/4294967296.0,1,-nbitq), 
to_sfixed(885617473.0/4294967296.0,1,-nbitq), 
to_sfixed(85685162.0/4294967296.0,1,-nbitq), 
to_sfixed(-429887358.0/4294967296.0,1,-nbitq), 
to_sfixed(-1228263558.0/4294967296.0,1,-nbitq), 
to_sfixed(1113260584.0/4294967296.0,1,-nbitq), 
to_sfixed(-162438933.0/4294967296.0,1,-nbitq), 
to_sfixed(299560031.0/4294967296.0,1,-nbitq), 
to_sfixed(92684408.0/4294967296.0,1,-nbitq), 
to_sfixed(-230893972.0/4294967296.0,1,-nbitq), 
to_sfixed(576736671.0/4294967296.0,1,-nbitq), 
to_sfixed(702722058.0/4294967296.0,1,-nbitq), 
to_sfixed(-444257290.0/4294967296.0,1,-nbitq), 
to_sfixed(457358832.0/4294967296.0,1,-nbitq), 
to_sfixed(-301897253.0/4294967296.0,1,-nbitq), 
to_sfixed(976967689.0/4294967296.0,1,-nbitq), 
to_sfixed(-679757368.0/4294967296.0,1,-nbitq), 
to_sfixed(-291282840.0/4294967296.0,1,-nbitq), 
to_sfixed(-446863334.0/4294967296.0,1,-nbitq), 
to_sfixed(-393263169.0/4294967296.0,1,-nbitq), 
to_sfixed(299476943.0/4294967296.0,1,-nbitq), 
to_sfixed(-436433448.0/4294967296.0,1,-nbitq), 
to_sfixed(124142911.0/4294967296.0,1,-nbitq), 
to_sfixed(-811471966.0/4294967296.0,1,-nbitq), 
to_sfixed(619539246.0/4294967296.0,1,-nbitq), 
to_sfixed(870972142.0/4294967296.0,1,-nbitq), 
to_sfixed(-434068586.0/4294967296.0,1,-nbitq), 
to_sfixed(-191130756.0/4294967296.0,1,-nbitq), 
to_sfixed(-240411058.0/4294967296.0,1,-nbitq), 
to_sfixed(983902646.0/4294967296.0,1,-nbitq), 
to_sfixed(-252010324.0/4294967296.0,1,-nbitq), 
to_sfixed(564803562.0/4294967296.0,1,-nbitq), 
to_sfixed(-853935918.0/4294967296.0,1,-nbitq), 
to_sfixed(-743257304.0/4294967296.0,1,-nbitq), 
to_sfixed(141928042.0/4294967296.0,1,-nbitq), 
to_sfixed(-1605468458.0/4294967296.0,1,-nbitq), 
to_sfixed(-496150725.0/4294967296.0,1,-nbitq), 
to_sfixed(-516032566.0/4294967296.0,1,-nbitq), 
to_sfixed(-680555211.0/4294967296.0,1,-nbitq), 
to_sfixed(-485308814.0/4294967296.0,1,-nbitq), 
to_sfixed(21860277.0/4294967296.0,1,-nbitq), 
to_sfixed(178804066.0/4294967296.0,1,-nbitq), 
to_sfixed(87496234.0/4294967296.0,1,-nbitq), 
to_sfixed(-217515361.0/4294967296.0,1,-nbitq), 
to_sfixed(-576332733.0/4294967296.0,1,-nbitq), 
to_sfixed(-842512016.0/4294967296.0,1,-nbitq), 
to_sfixed(165068967.0/4294967296.0,1,-nbitq), 
to_sfixed(93929719.0/4294967296.0,1,-nbitq), 
to_sfixed(129591136.0/4294967296.0,1,-nbitq), 
to_sfixed(1679715613.0/4294967296.0,1,-nbitq), 
to_sfixed(331009374.0/4294967296.0,1,-nbitq), 
to_sfixed(-624038904.0/4294967296.0,1,-nbitq), 
to_sfixed(401282610.0/4294967296.0,1,-nbitq), 
to_sfixed(-503547493.0/4294967296.0,1,-nbitq), 
to_sfixed(447237153.0/4294967296.0,1,-nbitq), 
to_sfixed(-202147699.0/4294967296.0,1,-nbitq), 
to_sfixed(143414238.0/4294967296.0,1,-nbitq), 
to_sfixed(482378683.0/4294967296.0,1,-nbitq), 
to_sfixed(390707657.0/4294967296.0,1,-nbitq), 
to_sfixed(167749655.0/4294967296.0,1,-nbitq), 
to_sfixed(1111002825.0/4294967296.0,1,-nbitq), 
to_sfixed(-421718747.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-364469057.0/4294967296.0,1,-nbitq), 
to_sfixed(-1236235630.0/4294967296.0,1,-nbitq), 
to_sfixed(-1374370107.0/4294967296.0,1,-nbitq), 
to_sfixed(-1287045519.0/4294967296.0,1,-nbitq), 
to_sfixed(-583947351.0/4294967296.0,1,-nbitq), 
to_sfixed(2605506463.0/4294967296.0,1,-nbitq), 
to_sfixed(-330755065.0/4294967296.0,1,-nbitq), 
to_sfixed(53174977.0/4294967296.0,1,-nbitq), 
to_sfixed(-182611205.0/4294967296.0,1,-nbitq), 
to_sfixed(-245119071.0/4294967296.0,1,-nbitq), 
to_sfixed(-447221598.0/4294967296.0,1,-nbitq), 
to_sfixed(-107569472.0/4294967296.0,1,-nbitq), 
to_sfixed(464736594.0/4294967296.0,1,-nbitq), 
to_sfixed(1280611695.0/4294967296.0,1,-nbitq), 
to_sfixed(-74510893.0/4294967296.0,1,-nbitq), 
to_sfixed(604950861.0/4294967296.0,1,-nbitq), 
to_sfixed(-118940212.0/4294967296.0,1,-nbitq), 
to_sfixed(57519350.0/4294967296.0,1,-nbitq), 
to_sfixed(-21312760.0/4294967296.0,1,-nbitq), 
to_sfixed(420604916.0/4294967296.0,1,-nbitq), 
to_sfixed(-281483509.0/4294967296.0,1,-nbitq), 
to_sfixed(-987241072.0/4294967296.0,1,-nbitq), 
to_sfixed(-883109247.0/4294967296.0,1,-nbitq), 
to_sfixed(536141442.0/4294967296.0,1,-nbitq), 
to_sfixed(-97503172.0/4294967296.0,1,-nbitq), 
to_sfixed(235297835.0/4294967296.0,1,-nbitq), 
to_sfixed(-110708796.0/4294967296.0,1,-nbitq), 
to_sfixed(-598925606.0/4294967296.0,1,-nbitq), 
to_sfixed(918720226.0/4294967296.0,1,-nbitq), 
to_sfixed(794416880.0/4294967296.0,1,-nbitq), 
to_sfixed(-159707878.0/4294967296.0,1,-nbitq), 
to_sfixed(73863767.0/4294967296.0,1,-nbitq), 
to_sfixed(16070698.0/4294967296.0,1,-nbitq), 
to_sfixed(5225566.0/4294967296.0,1,-nbitq), 
to_sfixed(-665468264.0/4294967296.0,1,-nbitq), 
to_sfixed(-855388229.0/4294967296.0,1,-nbitq), 
to_sfixed(-329849905.0/4294967296.0,1,-nbitq), 
to_sfixed(5977385.0/4294967296.0,1,-nbitq), 
to_sfixed(-145170581.0/4294967296.0,1,-nbitq), 
to_sfixed(8697661.0/4294967296.0,1,-nbitq), 
to_sfixed(-243028192.0/4294967296.0,1,-nbitq), 
to_sfixed(-392100253.0/4294967296.0,1,-nbitq), 
to_sfixed(570763353.0/4294967296.0,1,-nbitq), 
to_sfixed(1035841894.0/4294967296.0,1,-nbitq), 
to_sfixed(-720930548.0/4294967296.0,1,-nbitq), 
to_sfixed(-1184565359.0/4294967296.0,1,-nbitq), 
to_sfixed(280866204.0/4294967296.0,1,-nbitq), 
to_sfixed(1030859716.0/4294967296.0,1,-nbitq), 
to_sfixed(-142826685.0/4294967296.0,1,-nbitq), 
to_sfixed(721476211.0/4294967296.0,1,-nbitq), 
to_sfixed(-420764899.0/4294967296.0,1,-nbitq), 
to_sfixed(-1250453869.0/4294967296.0,1,-nbitq), 
to_sfixed(775521250.0/4294967296.0,1,-nbitq), 
to_sfixed(-1313211176.0/4294967296.0,1,-nbitq), 
to_sfixed(840726339.0/4294967296.0,1,-nbitq), 
to_sfixed(-575890619.0/4294967296.0,1,-nbitq), 
to_sfixed(-635548802.0/4294967296.0,1,-nbitq), 
to_sfixed(-78312451.0/4294967296.0,1,-nbitq), 
to_sfixed(-36679025.0/4294967296.0,1,-nbitq), 
to_sfixed(83867597.0/4294967296.0,1,-nbitq), 
to_sfixed(23456987.0/4294967296.0,1,-nbitq), 
to_sfixed(827232285.0/4294967296.0,1,-nbitq), 
to_sfixed(-116092719.0/4294967296.0,1,-nbitq), 
to_sfixed(-899249680.0/4294967296.0,1,-nbitq), 
to_sfixed(-167497375.0/4294967296.0,1,-nbitq), 
to_sfixed(-12421237.0/4294967296.0,1,-nbitq), 
to_sfixed(121469863.0/4294967296.0,1,-nbitq), 
to_sfixed(990482078.0/4294967296.0,1,-nbitq), 
to_sfixed(280796758.0/4294967296.0,1,-nbitq), 
to_sfixed(-413681605.0/4294967296.0,1,-nbitq), 
to_sfixed(1424770210.0/4294967296.0,1,-nbitq), 
to_sfixed(-209120573.0/4294967296.0,1,-nbitq), 
to_sfixed(743867001.0/4294967296.0,1,-nbitq), 
to_sfixed(280723159.0/4294967296.0,1,-nbitq), 
to_sfixed(316778555.0/4294967296.0,1,-nbitq), 
to_sfixed(-127867739.0/4294967296.0,1,-nbitq), 
to_sfixed(1195104436.0/4294967296.0,1,-nbitq), 
to_sfixed(-60505056.0/4294967296.0,1,-nbitq), 
to_sfixed(1356657344.0/4294967296.0,1,-nbitq), 
to_sfixed(365502697.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(177894462.0/4294967296.0,1,-nbitq), 
to_sfixed(-340738619.0/4294967296.0,1,-nbitq), 
to_sfixed(-2159982910.0/4294967296.0,1,-nbitq), 
to_sfixed(-1056029873.0/4294967296.0,1,-nbitq), 
to_sfixed(-581903143.0/4294967296.0,1,-nbitq), 
to_sfixed(2706675658.0/4294967296.0,1,-nbitq), 
to_sfixed(401192755.0/4294967296.0,1,-nbitq), 
to_sfixed(651376754.0/4294967296.0,1,-nbitq), 
to_sfixed(-1211099680.0/4294967296.0,1,-nbitq), 
to_sfixed(-296308863.0/4294967296.0,1,-nbitq), 
to_sfixed(1068244473.0/4294967296.0,1,-nbitq), 
to_sfixed(234696962.0/4294967296.0,1,-nbitq), 
to_sfixed(657571890.0/4294967296.0,1,-nbitq), 
to_sfixed(1501452084.0/4294967296.0,1,-nbitq), 
to_sfixed(-184816683.0/4294967296.0,1,-nbitq), 
to_sfixed(934627794.0/4294967296.0,1,-nbitq), 
to_sfixed(-87438443.0/4294967296.0,1,-nbitq), 
to_sfixed(33073385.0/4294967296.0,1,-nbitq), 
to_sfixed(215891556.0/4294967296.0,1,-nbitq), 
to_sfixed(139500792.0/4294967296.0,1,-nbitq), 
to_sfixed(-150287317.0/4294967296.0,1,-nbitq), 
to_sfixed(-538371699.0/4294967296.0,1,-nbitq), 
to_sfixed(-1162777304.0/4294967296.0,1,-nbitq), 
to_sfixed(714912437.0/4294967296.0,1,-nbitq), 
to_sfixed(458066417.0/4294967296.0,1,-nbitq), 
to_sfixed(841422156.0/4294967296.0,1,-nbitq), 
to_sfixed(-313762066.0/4294967296.0,1,-nbitq), 
to_sfixed(-40289598.0/4294967296.0,1,-nbitq), 
to_sfixed(812433250.0/4294967296.0,1,-nbitq), 
to_sfixed(907342072.0/4294967296.0,1,-nbitq), 
to_sfixed(690081351.0/4294967296.0,1,-nbitq), 
to_sfixed(-309944971.0/4294967296.0,1,-nbitq), 
to_sfixed(-179295413.0/4294967296.0,1,-nbitq), 
to_sfixed(-805609863.0/4294967296.0,1,-nbitq), 
to_sfixed(-59066544.0/4294967296.0,1,-nbitq), 
to_sfixed(201773500.0/4294967296.0,1,-nbitq), 
to_sfixed(-664704291.0/4294967296.0,1,-nbitq), 
to_sfixed(953008345.0/4294967296.0,1,-nbitq), 
to_sfixed(-259673281.0/4294967296.0,1,-nbitq), 
to_sfixed(-307785169.0/4294967296.0,1,-nbitq), 
to_sfixed(-621249818.0/4294967296.0,1,-nbitq), 
to_sfixed(-904723879.0/4294967296.0,1,-nbitq), 
to_sfixed(121178348.0/4294967296.0,1,-nbitq), 
to_sfixed(-37430812.0/4294967296.0,1,-nbitq), 
to_sfixed(-1298335520.0/4294967296.0,1,-nbitq), 
to_sfixed(24118314.0/4294967296.0,1,-nbitq), 
to_sfixed(-310143296.0/4294967296.0,1,-nbitq), 
to_sfixed(714260321.0/4294967296.0,1,-nbitq), 
to_sfixed(105389999.0/4294967296.0,1,-nbitq), 
to_sfixed(667249465.0/4294967296.0,1,-nbitq), 
to_sfixed(-614123627.0/4294967296.0,1,-nbitq), 
to_sfixed(-1458343942.0/4294967296.0,1,-nbitq), 
to_sfixed(-44495448.0/4294967296.0,1,-nbitq), 
to_sfixed(-1798147796.0/4294967296.0,1,-nbitq), 
to_sfixed(1383193431.0/4294967296.0,1,-nbitq), 
to_sfixed(-826587755.0/4294967296.0,1,-nbitq), 
to_sfixed(-307515892.0/4294967296.0,1,-nbitq), 
to_sfixed(706893759.0/4294967296.0,1,-nbitq), 
to_sfixed(-241179156.0/4294967296.0,1,-nbitq), 
to_sfixed(-192477336.0/4294967296.0,1,-nbitq), 
to_sfixed(514242523.0/4294967296.0,1,-nbitq), 
to_sfixed(605458555.0/4294967296.0,1,-nbitq), 
to_sfixed(-581661744.0/4294967296.0,1,-nbitq), 
to_sfixed(-730157086.0/4294967296.0,1,-nbitq), 
to_sfixed(-75656801.0/4294967296.0,1,-nbitq), 
to_sfixed(-571971122.0/4294967296.0,1,-nbitq), 
to_sfixed(-828664138.0/4294967296.0,1,-nbitq), 
to_sfixed(1394020803.0/4294967296.0,1,-nbitq), 
to_sfixed(-140067333.0/4294967296.0,1,-nbitq), 
to_sfixed(-1390832722.0/4294967296.0,1,-nbitq), 
to_sfixed(1235802676.0/4294967296.0,1,-nbitq), 
to_sfixed(-45979898.0/4294967296.0,1,-nbitq), 
to_sfixed(680232764.0/4294967296.0,1,-nbitq), 
to_sfixed(-79758099.0/4294967296.0,1,-nbitq), 
to_sfixed(-113706099.0/4294967296.0,1,-nbitq), 
to_sfixed(-1093756757.0/4294967296.0,1,-nbitq), 
to_sfixed(1399062751.0/4294967296.0,1,-nbitq), 
to_sfixed(-140015681.0/4294967296.0,1,-nbitq), 
to_sfixed(1379799481.0/4294967296.0,1,-nbitq), 
to_sfixed(345517177.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(621203006.0/4294967296.0,1,-nbitq), 
to_sfixed(-1381957285.0/4294967296.0,1,-nbitq), 
to_sfixed(-3062578246.0/4294967296.0,1,-nbitq), 
to_sfixed(-1380792006.0/4294967296.0,1,-nbitq), 
to_sfixed(-828542571.0/4294967296.0,1,-nbitq), 
to_sfixed(328350461.0/4294967296.0,1,-nbitq), 
to_sfixed(323583783.0/4294967296.0,1,-nbitq), 
to_sfixed(698859144.0/4294967296.0,1,-nbitq), 
to_sfixed(-987024019.0/4294967296.0,1,-nbitq), 
to_sfixed(185102999.0/4294967296.0,1,-nbitq), 
to_sfixed(1482959657.0/4294967296.0,1,-nbitq), 
to_sfixed(13793160.0/4294967296.0,1,-nbitq), 
to_sfixed(-25342091.0/4294967296.0,1,-nbitq), 
to_sfixed(1106001523.0/4294967296.0,1,-nbitq), 
to_sfixed(385586508.0/4294967296.0,1,-nbitq), 
to_sfixed(849553750.0/4294967296.0,1,-nbitq), 
to_sfixed(284401235.0/4294967296.0,1,-nbitq), 
to_sfixed(383252559.0/4294967296.0,1,-nbitq), 
to_sfixed(-329533958.0/4294967296.0,1,-nbitq), 
to_sfixed(779122162.0/4294967296.0,1,-nbitq), 
to_sfixed(-377663775.0/4294967296.0,1,-nbitq), 
to_sfixed(-1935515746.0/4294967296.0,1,-nbitq), 
to_sfixed(-1009696690.0/4294967296.0,1,-nbitq), 
to_sfixed(222637595.0/4294967296.0,1,-nbitq), 
to_sfixed(-192370103.0/4294967296.0,1,-nbitq), 
to_sfixed(1192234518.0/4294967296.0,1,-nbitq), 
to_sfixed(207913048.0/4294967296.0,1,-nbitq), 
to_sfixed(295903229.0/4294967296.0,1,-nbitq), 
to_sfixed(1101651634.0/4294967296.0,1,-nbitq), 
to_sfixed(1137966041.0/4294967296.0,1,-nbitq), 
to_sfixed(-112461710.0/4294967296.0,1,-nbitq), 
to_sfixed(-1017445230.0/4294967296.0,1,-nbitq), 
to_sfixed(-73341887.0/4294967296.0,1,-nbitq), 
to_sfixed(-393365345.0/4294967296.0,1,-nbitq), 
to_sfixed(158813885.0/4294967296.0,1,-nbitq), 
to_sfixed(-884436867.0/4294967296.0,1,-nbitq), 
to_sfixed(-683061249.0/4294967296.0,1,-nbitq), 
to_sfixed(1528055773.0/4294967296.0,1,-nbitq), 
to_sfixed(-285945788.0/4294967296.0,1,-nbitq), 
to_sfixed(90329185.0/4294967296.0,1,-nbitq), 
to_sfixed(-1036464818.0/4294967296.0,1,-nbitq), 
to_sfixed(-911467421.0/4294967296.0,1,-nbitq), 
to_sfixed(-80836195.0/4294967296.0,1,-nbitq), 
to_sfixed(-401502464.0/4294967296.0,1,-nbitq), 
to_sfixed(-1493649262.0/4294967296.0,1,-nbitq), 
to_sfixed(132522869.0/4294967296.0,1,-nbitq), 
to_sfixed(-348800284.0/4294967296.0,1,-nbitq), 
to_sfixed(811877281.0/4294967296.0,1,-nbitq), 
to_sfixed(102191973.0/4294967296.0,1,-nbitq), 
to_sfixed(874256519.0/4294967296.0,1,-nbitq), 
to_sfixed(-81748721.0/4294967296.0,1,-nbitq), 
to_sfixed(-1377248740.0/4294967296.0,1,-nbitq), 
to_sfixed(544938045.0/4294967296.0,1,-nbitq), 
to_sfixed(-1323282598.0/4294967296.0,1,-nbitq), 
to_sfixed(666435691.0/4294967296.0,1,-nbitq), 
to_sfixed(-655598264.0/4294967296.0,1,-nbitq), 
to_sfixed(-399594232.0/4294967296.0,1,-nbitq), 
to_sfixed(955825473.0/4294967296.0,1,-nbitq), 
to_sfixed(10548643.0/4294967296.0,1,-nbitq), 
to_sfixed(-86411640.0/4294967296.0,1,-nbitq), 
to_sfixed(307720858.0/4294967296.0,1,-nbitq), 
to_sfixed(1085632276.0/4294967296.0,1,-nbitq), 
to_sfixed(-1017797384.0/4294967296.0,1,-nbitq), 
to_sfixed(-1246229673.0/4294967296.0,1,-nbitq), 
to_sfixed(-199906005.0/4294967296.0,1,-nbitq), 
to_sfixed(-319293022.0/4294967296.0,1,-nbitq), 
to_sfixed(-37802512.0/4294967296.0,1,-nbitq), 
to_sfixed(1599545183.0/4294967296.0,1,-nbitq), 
to_sfixed(15127695.0/4294967296.0,1,-nbitq), 
to_sfixed(-310156711.0/4294967296.0,1,-nbitq), 
to_sfixed(716285036.0/4294967296.0,1,-nbitq), 
to_sfixed(28989845.0/4294967296.0,1,-nbitq), 
to_sfixed(612912201.0/4294967296.0,1,-nbitq), 
to_sfixed(313666113.0/4294967296.0,1,-nbitq), 
to_sfixed(137271706.0/4294967296.0,1,-nbitq), 
to_sfixed(-1388513535.0/4294967296.0,1,-nbitq), 
to_sfixed(561431768.0/4294967296.0,1,-nbitq), 
to_sfixed(209457446.0/4294967296.0,1,-nbitq), 
to_sfixed(839410000.0/4294967296.0,1,-nbitq), 
to_sfixed(-173766266.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(741592783.0/4294967296.0,1,-nbitq), 
to_sfixed(-1210164814.0/4294967296.0,1,-nbitq), 
to_sfixed(-3186443972.0/4294967296.0,1,-nbitq), 
to_sfixed(-1265415945.0/4294967296.0,1,-nbitq), 
to_sfixed(32372000.0/4294967296.0,1,-nbitq), 
to_sfixed(-155547871.0/4294967296.0,1,-nbitq), 
to_sfixed(270208146.0/4294967296.0,1,-nbitq), 
to_sfixed(-2139273484.0/4294967296.0,1,-nbitq), 
to_sfixed(-790751114.0/4294967296.0,1,-nbitq), 
to_sfixed(-57933957.0/4294967296.0,1,-nbitq), 
to_sfixed(1656890517.0/4294967296.0,1,-nbitq), 
to_sfixed(-385593141.0/4294967296.0,1,-nbitq), 
to_sfixed(784398707.0/4294967296.0,1,-nbitq), 
to_sfixed(369003570.0/4294967296.0,1,-nbitq), 
to_sfixed(389906805.0/4294967296.0,1,-nbitq), 
to_sfixed(1030496107.0/4294967296.0,1,-nbitq), 
to_sfixed(73414925.0/4294967296.0,1,-nbitq), 
to_sfixed(9978139.0/4294967296.0,1,-nbitq), 
to_sfixed(-1284770546.0/4294967296.0,1,-nbitq), 
to_sfixed(-79513175.0/4294967296.0,1,-nbitq), 
to_sfixed(335555274.0/4294967296.0,1,-nbitq), 
to_sfixed(-1601250209.0/4294967296.0,1,-nbitq), 
to_sfixed(-945778826.0/4294967296.0,1,-nbitq), 
to_sfixed(911875720.0/4294967296.0,1,-nbitq), 
to_sfixed(-226707805.0/4294967296.0,1,-nbitq), 
to_sfixed(1837367128.0/4294967296.0,1,-nbitq), 
to_sfixed(-15997217.0/4294967296.0,1,-nbitq), 
to_sfixed(1396967205.0/4294967296.0,1,-nbitq), 
to_sfixed(824302318.0/4294967296.0,1,-nbitq), 
to_sfixed(753644806.0/4294967296.0,1,-nbitq), 
to_sfixed(632505328.0/4294967296.0,1,-nbitq), 
to_sfixed(-1440298747.0/4294967296.0,1,-nbitq), 
to_sfixed(135784813.0/4294967296.0,1,-nbitq), 
to_sfixed(373118248.0/4294967296.0,1,-nbitq), 
to_sfixed(518711512.0/4294967296.0,1,-nbitq), 
to_sfixed(-837412337.0/4294967296.0,1,-nbitq), 
to_sfixed(-674193380.0/4294967296.0,1,-nbitq), 
to_sfixed(2091970699.0/4294967296.0,1,-nbitq), 
to_sfixed(-306753698.0/4294967296.0,1,-nbitq), 
to_sfixed(-49975030.0/4294967296.0,1,-nbitq), 
to_sfixed(-437303821.0/4294967296.0,1,-nbitq), 
to_sfixed(-701817376.0/4294967296.0,1,-nbitq), 
to_sfixed(-678900695.0/4294967296.0,1,-nbitq), 
to_sfixed(102302060.0/4294967296.0,1,-nbitq), 
to_sfixed(-549264298.0/4294967296.0,1,-nbitq), 
to_sfixed(-609400736.0/4294967296.0,1,-nbitq), 
to_sfixed(-353466173.0/4294967296.0,1,-nbitq), 
to_sfixed(206073553.0/4294967296.0,1,-nbitq), 
to_sfixed(224634316.0/4294967296.0,1,-nbitq), 
to_sfixed(912984981.0/4294967296.0,1,-nbitq), 
to_sfixed(-266029385.0/4294967296.0,1,-nbitq), 
to_sfixed(-652373985.0/4294967296.0,1,-nbitq), 
to_sfixed(-41362493.0/4294967296.0,1,-nbitq), 
to_sfixed(-105887191.0/4294967296.0,1,-nbitq), 
to_sfixed(426403020.0/4294967296.0,1,-nbitq), 
to_sfixed(-68240692.0/4294967296.0,1,-nbitq), 
to_sfixed(281667330.0/4294967296.0,1,-nbitq), 
to_sfixed(381731140.0/4294967296.0,1,-nbitq), 
to_sfixed(-169496980.0/4294967296.0,1,-nbitq), 
to_sfixed(252636892.0/4294967296.0,1,-nbitq), 
to_sfixed(-45730801.0/4294967296.0,1,-nbitq), 
to_sfixed(894944796.0/4294967296.0,1,-nbitq), 
to_sfixed(-916689611.0/4294967296.0,1,-nbitq), 
to_sfixed(-952832690.0/4294967296.0,1,-nbitq), 
to_sfixed(-255723637.0/4294967296.0,1,-nbitq), 
to_sfixed(-303391614.0/4294967296.0,1,-nbitq), 
to_sfixed(416334257.0/4294967296.0,1,-nbitq), 
to_sfixed(1543438212.0/4294967296.0,1,-nbitq), 
to_sfixed(308434143.0/4294967296.0,1,-nbitq), 
to_sfixed(1477601213.0/4294967296.0,1,-nbitq), 
to_sfixed(1400891541.0/4294967296.0,1,-nbitq), 
to_sfixed(52735695.0/4294967296.0,1,-nbitq), 
to_sfixed(900398011.0/4294967296.0,1,-nbitq), 
to_sfixed(230260853.0/4294967296.0,1,-nbitq), 
to_sfixed(-206733635.0/4294967296.0,1,-nbitq), 
to_sfixed(-2453181430.0/4294967296.0,1,-nbitq), 
to_sfixed(14301833.0/4294967296.0,1,-nbitq), 
to_sfixed(-332155203.0/4294967296.0,1,-nbitq), 
to_sfixed(-403742981.0/4294967296.0,1,-nbitq), 
to_sfixed(326483162.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(36058713.0/4294967296.0,1,-nbitq), 
to_sfixed(-346449119.0/4294967296.0,1,-nbitq), 
to_sfixed(-1011716042.0/4294967296.0,1,-nbitq), 
to_sfixed(-1035710083.0/4294967296.0,1,-nbitq), 
to_sfixed(426677771.0/4294967296.0,1,-nbitq), 
to_sfixed(355481353.0/4294967296.0,1,-nbitq), 
to_sfixed(609283999.0/4294967296.0,1,-nbitq), 
to_sfixed(-2522443841.0/4294967296.0,1,-nbitq), 
to_sfixed(-809391003.0/4294967296.0,1,-nbitq), 
to_sfixed(261632047.0/4294967296.0,1,-nbitq), 
to_sfixed(1211191973.0/4294967296.0,1,-nbitq), 
to_sfixed(-1864973385.0/4294967296.0,1,-nbitq), 
to_sfixed(261741905.0/4294967296.0,1,-nbitq), 
to_sfixed(-212315129.0/4294967296.0,1,-nbitq), 
to_sfixed(195323978.0/4294967296.0,1,-nbitq), 
to_sfixed(453025705.0/4294967296.0,1,-nbitq), 
to_sfixed(-275274639.0/4294967296.0,1,-nbitq), 
to_sfixed(-9329271.0/4294967296.0,1,-nbitq), 
to_sfixed(102406610.0/4294967296.0,1,-nbitq), 
to_sfixed(464174223.0/4294967296.0,1,-nbitq), 
to_sfixed(181472430.0/4294967296.0,1,-nbitq), 
to_sfixed(-736456899.0/4294967296.0,1,-nbitq), 
to_sfixed(-969674383.0/4294967296.0,1,-nbitq), 
to_sfixed(1515601674.0/4294967296.0,1,-nbitq), 
to_sfixed(291428653.0/4294967296.0,1,-nbitq), 
to_sfixed(938551793.0/4294967296.0,1,-nbitq), 
to_sfixed(751831677.0/4294967296.0,1,-nbitq), 
to_sfixed(1284913718.0/4294967296.0,1,-nbitq), 
to_sfixed(-2200702832.0/4294967296.0,1,-nbitq), 
to_sfixed(786500505.0/4294967296.0,1,-nbitq), 
to_sfixed(1625352789.0/4294967296.0,1,-nbitq), 
to_sfixed(-1482368309.0/4294967296.0,1,-nbitq), 
to_sfixed(724379323.0/4294967296.0,1,-nbitq), 
to_sfixed(127242547.0/4294967296.0,1,-nbitq), 
to_sfixed(-428261043.0/4294967296.0,1,-nbitq), 
to_sfixed(-1003359480.0/4294967296.0,1,-nbitq), 
to_sfixed(-291358580.0/4294967296.0,1,-nbitq), 
to_sfixed(1541860988.0/4294967296.0,1,-nbitq), 
to_sfixed(66407043.0/4294967296.0,1,-nbitq), 
to_sfixed(641763812.0/4294967296.0,1,-nbitq), 
to_sfixed(1602780077.0/4294967296.0,1,-nbitq), 
to_sfixed(-897277552.0/4294967296.0,1,-nbitq), 
to_sfixed(-645102914.0/4294967296.0,1,-nbitq), 
to_sfixed(-614858913.0/4294967296.0,1,-nbitq), 
to_sfixed(-134171049.0/4294967296.0,1,-nbitq), 
to_sfixed(-753333658.0/4294967296.0,1,-nbitq), 
to_sfixed(-381464122.0/4294967296.0,1,-nbitq), 
to_sfixed(-453360195.0/4294967296.0,1,-nbitq), 
to_sfixed(51288423.0/4294967296.0,1,-nbitq), 
to_sfixed(870485489.0/4294967296.0,1,-nbitq), 
to_sfixed(655066148.0/4294967296.0,1,-nbitq), 
to_sfixed(-1443328370.0/4294967296.0,1,-nbitq), 
to_sfixed(-485778650.0/4294967296.0,1,-nbitq), 
to_sfixed(696689526.0/4294967296.0,1,-nbitq), 
to_sfixed(285235441.0/4294967296.0,1,-nbitq), 
to_sfixed(-1394693060.0/4294967296.0,1,-nbitq), 
to_sfixed(6999112.0/4294967296.0,1,-nbitq), 
to_sfixed(163063059.0/4294967296.0,1,-nbitq), 
to_sfixed(-233634320.0/4294967296.0,1,-nbitq), 
to_sfixed(-146231892.0/4294967296.0,1,-nbitq), 
to_sfixed(-159505809.0/4294967296.0,1,-nbitq), 
to_sfixed(981946890.0/4294967296.0,1,-nbitq), 
to_sfixed(702690093.0/4294967296.0,1,-nbitq), 
to_sfixed(131484090.0/4294967296.0,1,-nbitq), 
to_sfixed(-289696359.0/4294967296.0,1,-nbitq), 
to_sfixed(-412448397.0/4294967296.0,1,-nbitq), 
to_sfixed(1407940872.0/4294967296.0,1,-nbitq), 
to_sfixed(1618918663.0/4294967296.0,1,-nbitq), 
to_sfixed(27645143.0/4294967296.0,1,-nbitq), 
to_sfixed(1851638691.0/4294967296.0,1,-nbitq), 
to_sfixed(777365084.0/4294967296.0,1,-nbitq), 
to_sfixed(204698825.0/4294967296.0,1,-nbitq), 
to_sfixed(625507024.0/4294967296.0,1,-nbitq), 
to_sfixed(184781012.0/4294967296.0,1,-nbitq), 
to_sfixed(-151945302.0/4294967296.0,1,-nbitq), 
to_sfixed(-2254075843.0/4294967296.0,1,-nbitq), 
to_sfixed(-482771921.0/4294967296.0,1,-nbitq), 
to_sfixed(-18321890.0/4294967296.0,1,-nbitq), 
to_sfixed(-1526206384.0/4294967296.0,1,-nbitq), 
to_sfixed(124679815.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(104105713.0/4294967296.0,1,-nbitq), 
to_sfixed(575226084.0/4294967296.0,1,-nbitq), 
to_sfixed(342902136.0/4294967296.0,1,-nbitq), 
to_sfixed(-686026226.0/4294967296.0,1,-nbitq), 
to_sfixed(504455804.0/4294967296.0,1,-nbitq), 
to_sfixed(-787071915.0/4294967296.0,1,-nbitq), 
to_sfixed(324601540.0/4294967296.0,1,-nbitq), 
to_sfixed(-1082858786.0/4294967296.0,1,-nbitq), 
to_sfixed(-445641856.0/4294967296.0,1,-nbitq), 
to_sfixed(341640133.0/4294967296.0,1,-nbitq), 
to_sfixed(1047034432.0/4294967296.0,1,-nbitq), 
to_sfixed(-1770742460.0/4294967296.0,1,-nbitq), 
to_sfixed(498173430.0/4294967296.0,1,-nbitq), 
to_sfixed(-497566494.0/4294967296.0,1,-nbitq), 
to_sfixed(82927410.0/4294967296.0,1,-nbitq), 
to_sfixed(1946344558.0/4294967296.0,1,-nbitq), 
to_sfixed(-178375672.0/4294967296.0,1,-nbitq), 
to_sfixed(76702057.0/4294967296.0,1,-nbitq), 
to_sfixed(-22000438.0/4294967296.0,1,-nbitq), 
to_sfixed(824654234.0/4294967296.0,1,-nbitq), 
to_sfixed(-3032691.0/4294967296.0,1,-nbitq), 
to_sfixed(-508502376.0/4294967296.0,1,-nbitq), 
to_sfixed(637063819.0/4294967296.0,1,-nbitq), 
to_sfixed(3388194479.0/4294967296.0,1,-nbitq), 
to_sfixed(300641529.0/4294967296.0,1,-nbitq), 
to_sfixed(426659390.0/4294967296.0,1,-nbitq), 
to_sfixed(479394173.0/4294967296.0,1,-nbitq), 
to_sfixed(-215095589.0/4294967296.0,1,-nbitq), 
to_sfixed(-3331570430.0/4294967296.0,1,-nbitq), 
to_sfixed(-249831141.0/4294967296.0,1,-nbitq), 
to_sfixed(1646442488.0/4294967296.0,1,-nbitq), 
to_sfixed(-262342485.0/4294967296.0,1,-nbitq), 
to_sfixed(-152831881.0/4294967296.0,1,-nbitq), 
to_sfixed(770551759.0/4294967296.0,1,-nbitq), 
to_sfixed(-50118590.0/4294967296.0,1,-nbitq), 
to_sfixed(-333170834.0/4294967296.0,1,-nbitq), 
to_sfixed(-20840542.0/4294967296.0,1,-nbitq), 
to_sfixed(1090827432.0/4294967296.0,1,-nbitq), 
to_sfixed(-90185861.0/4294967296.0,1,-nbitq), 
to_sfixed(541394817.0/4294967296.0,1,-nbitq), 
to_sfixed(2296030357.0/4294967296.0,1,-nbitq), 
to_sfixed(486929899.0/4294967296.0,1,-nbitq), 
to_sfixed(-965211178.0/4294967296.0,1,-nbitq), 
to_sfixed(-542687092.0/4294967296.0,1,-nbitq), 
to_sfixed(-582960747.0/4294967296.0,1,-nbitq), 
to_sfixed(735305.0/4294967296.0,1,-nbitq), 
to_sfixed(57878242.0/4294967296.0,1,-nbitq), 
to_sfixed(1067427231.0/4294967296.0,1,-nbitq), 
to_sfixed(269949025.0/4294967296.0,1,-nbitq), 
to_sfixed(26566029.0/4294967296.0,1,-nbitq), 
to_sfixed(474820394.0/4294967296.0,1,-nbitq), 
to_sfixed(-1716193689.0/4294967296.0,1,-nbitq), 
to_sfixed(-273391715.0/4294967296.0,1,-nbitq), 
to_sfixed(1432796570.0/4294967296.0,1,-nbitq), 
to_sfixed(978538743.0/4294967296.0,1,-nbitq), 
to_sfixed(-1663225951.0/4294967296.0,1,-nbitq), 
to_sfixed(-1117122474.0/4294967296.0,1,-nbitq), 
to_sfixed(-547583209.0/4294967296.0,1,-nbitq), 
to_sfixed(-141374993.0/4294967296.0,1,-nbitq), 
to_sfixed(-221201245.0/4294967296.0,1,-nbitq), 
to_sfixed(-352515395.0/4294967296.0,1,-nbitq), 
to_sfixed(111425189.0/4294967296.0,1,-nbitq), 
to_sfixed(1450737317.0/4294967296.0,1,-nbitq), 
to_sfixed(-48037406.0/4294967296.0,1,-nbitq), 
to_sfixed(74444438.0/4294967296.0,1,-nbitq), 
to_sfixed(119918439.0/4294967296.0,1,-nbitq), 
to_sfixed(61797285.0/4294967296.0,1,-nbitq), 
to_sfixed(1170251020.0/4294967296.0,1,-nbitq), 
to_sfixed(-79902305.0/4294967296.0,1,-nbitq), 
to_sfixed(834793559.0/4294967296.0,1,-nbitq), 
to_sfixed(996780438.0/4294967296.0,1,-nbitq), 
to_sfixed(-404457186.0/4294967296.0,1,-nbitq), 
to_sfixed(-587104914.0/4294967296.0,1,-nbitq), 
to_sfixed(194422143.0/4294967296.0,1,-nbitq), 
to_sfixed(-426375184.0/4294967296.0,1,-nbitq), 
to_sfixed(-1431378889.0/4294967296.0,1,-nbitq), 
to_sfixed(-631305315.0/4294967296.0,1,-nbitq), 
to_sfixed(-1203693836.0/4294967296.0,1,-nbitq), 
to_sfixed(-1403189623.0/4294967296.0,1,-nbitq), 
to_sfixed(269921331.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(374228754.0/4294967296.0,1,-nbitq), 
to_sfixed(1584269275.0/4294967296.0,1,-nbitq), 
to_sfixed(-1555645866.0/4294967296.0,1,-nbitq), 
to_sfixed(-612558808.0/4294967296.0,1,-nbitq), 
to_sfixed(3881713.0/4294967296.0,1,-nbitq), 
to_sfixed(-621713832.0/4294967296.0,1,-nbitq), 
to_sfixed(-343537788.0/4294967296.0,1,-nbitq), 
to_sfixed(907305043.0/4294967296.0,1,-nbitq), 
to_sfixed(-566340970.0/4294967296.0,1,-nbitq), 
to_sfixed(135078824.0/4294967296.0,1,-nbitq), 
to_sfixed(376379947.0/4294967296.0,1,-nbitq), 
to_sfixed(-3429507298.0/4294967296.0,1,-nbitq), 
to_sfixed(1230626885.0/4294967296.0,1,-nbitq), 
to_sfixed(-437093535.0/4294967296.0,1,-nbitq), 
to_sfixed(-108807347.0/4294967296.0,1,-nbitq), 
to_sfixed(1307476125.0/4294967296.0,1,-nbitq), 
to_sfixed(132955290.0/4294967296.0,1,-nbitq), 
to_sfixed(-266840144.0/4294967296.0,1,-nbitq), 
to_sfixed(-879292030.0/4294967296.0,1,-nbitq), 
to_sfixed(711342882.0/4294967296.0,1,-nbitq), 
to_sfixed(117922105.0/4294967296.0,1,-nbitq), 
to_sfixed(-388797275.0/4294967296.0,1,-nbitq), 
to_sfixed(760454350.0/4294967296.0,1,-nbitq), 
to_sfixed(-963612228.0/4294967296.0,1,-nbitq), 
to_sfixed(277915246.0/4294967296.0,1,-nbitq), 
to_sfixed(-64267668.0/4294967296.0,1,-nbitq), 
to_sfixed(-108468352.0/4294967296.0,1,-nbitq), 
to_sfixed(-1313456470.0/4294967296.0,1,-nbitq), 
to_sfixed(-1728560936.0/4294967296.0,1,-nbitq), 
to_sfixed(435681398.0/4294967296.0,1,-nbitq), 
to_sfixed(-364065429.0/4294967296.0,1,-nbitq), 
to_sfixed(690652703.0/4294967296.0,1,-nbitq), 
to_sfixed(211100746.0/4294967296.0,1,-nbitq), 
to_sfixed(667143679.0/4294967296.0,1,-nbitq), 
to_sfixed(741294722.0/4294967296.0,1,-nbitq), 
to_sfixed(-149372322.0/4294967296.0,1,-nbitq), 
to_sfixed(-130302954.0/4294967296.0,1,-nbitq), 
to_sfixed(756532168.0/4294967296.0,1,-nbitq), 
to_sfixed(-368291604.0/4294967296.0,1,-nbitq), 
to_sfixed(403934805.0/4294967296.0,1,-nbitq), 
to_sfixed(1555724281.0/4294967296.0,1,-nbitq), 
to_sfixed(811381338.0/4294967296.0,1,-nbitq), 
to_sfixed(-115322763.0/4294967296.0,1,-nbitq), 
to_sfixed(-166368082.0/4294967296.0,1,-nbitq), 
to_sfixed(-362820023.0/4294967296.0,1,-nbitq), 
to_sfixed(-33032556.0/4294967296.0,1,-nbitq), 
to_sfixed(231156573.0/4294967296.0,1,-nbitq), 
to_sfixed(441407286.0/4294967296.0,1,-nbitq), 
to_sfixed(-13108396.0/4294967296.0,1,-nbitq), 
to_sfixed(763152042.0/4294967296.0,1,-nbitq), 
to_sfixed(418988854.0/4294967296.0,1,-nbitq), 
to_sfixed(-729525666.0/4294967296.0,1,-nbitq), 
to_sfixed(1431111554.0/4294967296.0,1,-nbitq), 
to_sfixed(1379418947.0/4294967296.0,1,-nbitq), 
to_sfixed(410377452.0/4294967296.0,1,-nbitq), 
to_sfixed(-1068609120.0/4294967296.0,1,-nbitq), 
to_sfixed(-385093021.0/4294967296.0,1,-nbitq), 
to_sfixed(5732651.0/4294967296.0,1,-nbitq), 
to_sfixed(-24145128.0/4294967296.0,1,-nbitq), 
to_sfixed(190331385.0/4294967296.0,1,-nbitq), 
to_sfixed(-127334654.0/4294967296.0,1,-nbitq), 
to_sfixed(-1049240209.0/4294967296.0,1,-nbitq), 
to_sfixed(686901371.0/4294967296.0,1,-nbitq), 
to_sfixed(292133463.0/4294967296.0,1,-nbitq), 
to_sfixed(-379394109.0/4294967296.0,1,-nbitq), 
to_sfixed(-51827766.0/4294967296.0,1,-nbitq), 
to_sfixed(1507757036.0/4294967296.0,1,-nbitq), 
to_sfixed(1247991469.0/4294967296.0,1,-nbitq), 
to_sfixed(-158476941.0/4294967296.0,1,-nbitq), 
to_sfixed(326378245.0/4294967296.0,1,-nbitq), 
to_sfixed(1574415292.0/4294967296.0,1,-nbitq), 
to_sfixed(139913896.0/4294967296.0,1,-nbitq), 
to_sfixed(-963465931.0/4294967296.0,1,-nbitq), 
to_sfixed(153756891.0/4294967296.0,1,-nbitq), 
to_sfixed(-512745043.0/4294967296.0,1,-nbitq), 
to_sfixed(-815336342.0/4294967296.0,1,-nbitq), 
to_sfixed(-850525235.0/4294967296.0,1,-nbitq), 
to_sfixed(-855541162.0/4294967296.0,1,-nbitq), 
to_sfixed(-581166168.0/4294967296.0,1,-nbitq), 
to_sfixed(109451664.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(75619949.0/4294967296.0,1,-nbitq), 
to_sfixed(2103862275.0/4294967296.0,1,-nbitq), 
to_sfixed(-521480760.0/4294967296.0,1,-nbitq), 
to_sfixed(-798729066.0/4294967296.0,1,-nbitq), 
to_sfixed(262043377.0/4294967296.0,1,-nbitq), 
to_sfixed(790795402.0/4294967296.0,1,-nbitq), 
to_sfixed(-121038586.0/4294967296.0,1,-nbitq), 
to_sfixed(594616524.0/4294967296.0,1,-nbitq), 
to_sfixed(-475946016.0/4294967296.0,1,-nbitq), 
to_sfixed(-100610760.0/4294967296.0,1,-nbitq), 
to_sfixed(-765741827.0/4294967296.0,1,-nbitq), 
to_sfixed(-2069590427.0/4294967296.0,1,-nbitq), 
to_sfixed(-279564407.0/4294967296.0,1,-nbitq), 
to_sfixed(-259225622.0/4294967296.0,1,-nbitq), 
to_sfixed(289585094.0/4294967296.0,1,-nbitq), 
to_sfixed(913155570.0/4294967296.0,1,-nbitq), 
to_sfixed(295901542.0/4294967296.0,1,-nbitq), 
to_sfixed(-301898848.0/4294967296.0,1,-nbitq), 
to_sfixed(-162467570.0/4294967296.0,1,-nbitq), 
to_sfixed(437792759.0/4294967296.0,1,-nbitq), 
to_sfixed(-164228169.0/4294967296.0,1,-nbitq), 
to_sfixed(786745564.0/4294967296.0,1,-nbitq), 
to_sfixed(278694719.0/4294967296.0,1,-nbitq), 
to_sfixed(-4222323294.0/4294967296.0,1,-nbitq), 
to_sfixed(328001854.0/4294967296.0,1,-nbitq), 
to_sfixed(-341967037.0/4294967296.0,1,-nbitq), 
to_sfixed(-721835915.0/4294967296.0,1,-nbitq), 
to_sfixed(-405861347.0/4294967296.0,1,-nbitq), 
to_sfixed(121021690.0/4294967296.0,1,-nbitq), 
to_sfixed(1124563278.0/4294967296.0,1,-nbitq), 
to_sfixed(-1220641153.0/4294967296.0,1,-nbitq), 
to_sfixed(1391366998.0/4294967296.0,1,-nbitq), 
to_sfixed(561440134.0/4294967296.0,1,-nbitq), 
to_sfixed(1055385217.0/4294967296.0,1,-nbitq), 
to_sfixed(1155948519.0/4294967296.0,1,-nbitq), 
to_sfixed(-458633496.0/4294967296.0,1,-nbitq), 
to_sfixed(508178165.0/4294967296.0,1,-nbitq), 
to_sfixed(-68185379.0/4294967296.0,1,-nbitq), 
to_sfixed(146140486.0/4294967296.0,1,-nbitq), 
to_sfixed(-129374428.0/4294967296.0,1,-nbitq), 
to_sfixed(262941072.0/4294967296.0,1,-nbitq), 
to_sfixed(1176041380.0/4294967296.0,1,-nbitq), 
to_sfixed(553249608.0/4294967296.0,1,-nbitq), 
to_sfixed(-320055583.0/4294967296.0,1,-nbitq), 
to_sfixed(-1733596777.0/4294967296.0,1,-nbitq), 
to_sfixed(-190054820.0/4294967296.0,1,-nbitq), 
to_sfixed(228914126.0/4294967296.0,1,-nbitq), 
to_sfixed(1170008919.0/4294967296.0,1,-nbitq), 
to_sfixed(246530931.0/4294967296.0,1,-nbitq), 
to_sfixed(512604678.0/4294967296.0,1,-nbitq), 
to_sfixed(357452493.0/4294967296.0,1,-nbitq), 
to_sfixed(418653611.0/4294967296.0,1,-nbitq), 
to_sfixed(1217145085.0/4294967296.0,1,-nbitq), 
to_sfixed(1616622288.0/4294967296.0,1,-nbitq), 
to_sfixed(-364297682.0/4294967296.0,1,-nbitq), 
to_sfixed(-1883660122.0/4294967296.0,1,-nbitq), 
to_sfixed(-1332135598.0/4294967296.0,1,-nbitq), 
to_sfixed(1034555118.0/4294967296.0,1,-nbitq), 
to_sfixed(-133636810.0/4294967296.0,1,-nbitq), 
to_sfixed(365413810.0/4294967296.0,1,-nbitq), 
to_sfixed(292142697.0/4294967296.0,1,-nbitq), 
to_sfixed(-628953291.0/4294967296.0,1,-nbitq), 
to_sfixed(361430480.0/4294967296.0,1,-nbitq), 
to_sfixed(241668688.0/4294967296.0,1,-nbitq), 
to_sfixed(-293691690.0/4294967296.0,1,-nbitq), 
to_sfixed(64686992.0/4294967296.0,1,-nbitq), 
to_sfixed(1162933888.0/4294967296.0,1,-nbitq), 
to_sfixed(697742143.0/4294967296.0,1,-nbitq), 
to_sfixed(-181031.0/4294967296.0,1,-nbitq), 
to_sfixed(-22688828.0/4294967296.0,1,-nbitq), 
to_sfixed(1378383949.0/4294967296.0,1,-nbitq), 
to_sfixed(-498530648.0/4294967296.0,1,-nbitq), 
to_sfixed(-1082257034.0/4294967296.0,1,-nbitq), 
to_sfixed(-185860474.0/4294967296.0,1,-nbitq), 
to_sfixed(-112173300.0/4294967296.0,1,-nbitq), 
to_sfixed(-495960771.0/4294967296.0,1,-nbitq), 
to_sfixed(-868888247.0/4294967296.0,1,-nbitq), 
to_sfixed(-40857679.0/4294967296.0,1,-nbitq), 
to_sfixed(-419673890.0/4294967296.0,1,-nbitq), 
to_sfixed(215128670.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(304534447.0/4294967296.0,1,-nbitq), 
to_sfixed(2599898453.0/4294967296.0,1,-nbitq), 
to_sfixed(-1023618458.0/4294967296.0,1,-nbitq), 
to_sfixed(-68046310.0/4294967296.0,1,-nbitq), 
to_sfixed(438185048.0/4294967296.0,1,-nbitq), 
to_sfixed(287520075.0/4294967296.0,1,-nbitq), 
to_sfixed(-387387695.0/4294967296.0,1,-nbitq), 
to_sfixed(477995888.0/4294967296.0,1,-nbitq), 
to_sfixed(-314867380.0/4294967296.0,1,-nbitq), 
to_sfixed(-253758378.0/4294967296.0,1,-nbitq), 
to_sfixed(-1955480927.0/4294967296.0,1,-nbitq), 
to_sfixed(-1674563343.0/4294967296.0,1,-nbitq), 
to_sfixed(-736104067.0/4294967296.0,1,-nbitq), 
to_sfixed(29352958.0/4294967296.0,1,-nbitq), 
to_sfixed(-137712572.0/4294967296.0,1,-nbitq), 
to_sfixed(103009635.0/4294967296.0,1,-nbitq), 
to_sfixed(46770221.0/4294967296.0,1,-nbitq), 
to_sfixed(68246175.0/4294967296.0,1,-nbitq), 
to_sfixed(-536842171.0/4294967296.0,1,-nbitq), 
to_sfixed(139594408.0/4294967296.0,1,-nbitq), 
to_sfixed(123990214.0/4294967296.0,1,-nbitq), 
to_sfixed(-294766137.0/4294967296.0,1,-nbitq), 
to_sfixed(256385422.0/4294967296.0,1,-nbitq), 
to_sfixed(-2408708296.0/4294967296.0,1,-nbitq), 
to_sfixed(188659639.0/4294967296.0,1,-nbitq), 
to_sfixed(-233198064.0/4294967296.0,1,-nbitq), 
to_sfixed(-757455878.0/4294967296.0,1,-nbitq), 
to_sfixed(-192628565.0/4294967296.0,1,-nbitq), 
to_sfixed(325858044.0/4294967296.0,1,-nbitq), 
to_sfixed(2102957550.0/4294967296.0,1,-nbitq), 
to_sfixed(-1798720166.0/4294967296.0,1,-nbitq), 
to_sfixed(1593380755.0/4294967296.0,1,-nbitq), 
to_sfixed(542044766.0/4294967296.0,1,-nbitq), 
to_sfixed(450845970.0/4294967296.0,1,-nbitq), 
to_sfixed(387592150.0/4294967296.0,1,-nbitq), 
to_sfixed(-719227008.0/4294967296.0,1,-nbitq), 
to_sfixed(60233291.0/4294967296.0,1,-nbitq), 
to_sfixed(-256859621.0/4294967296.0,1,-nbitq), 
to_sfixed(-257250551.0/4294967296.0,1,-nbitq), 
to_sfixed(-70455259.0/4294967296.0,1,-nbitq), 
to_sfixed(-699126769.0/4294967296.0,1,-nbitq), 
to_sfixed(327187910.0/4294967296.0,1,-nbitq), 
to_sfixed(-183323505.0/4294967296.0,1,-nbitq), 
to_sfixed(-1144294769.0/4294967296.0,1,-nbitq), 
to_sfixed(-1314838908.0/4294967296.0,1,-nbitq), 
to_sfixed(-58751312.0/4294967296.0,1,-nbitq), 
to_sfixed(-324637213.0/4294967296.0,1,-nbitq), 
to_sfixed(1245899987.0/4294967296.0,1,-nbitq), 
to_sfixed(268258587.0/4294967296.0,1,-nbitq), 
to_sfixed(939383287.0/4294967296.0,1,-nbitq), 
to_sfixed(-275691491.0/4294967296.0,1,-nbitq), 
to_sfixed(-128658360.0/4294967296.0,1,-nbitq), 
to_sfixed(1435997929.0/4294967296.0,1,-nbitq), 
to_sfixed(1240905088.0/4294967296.0,1,-nbitq), 
to_sfixed(-362142872.0/4294967296.0,1,-nbitq), 
to_sfixed(-1174989691.0/4294967296.0,1,-nbitq), 
to_sfixed(-662523195.0/4294967296.0,1,-nbitq), 
to_sfixed(481605170.0/4294967296.0,1,-nbitq), 
to_sfixed(361386245.0/4294967296.0,1,-nbitq), 
to_sfixed(367198254.0/4294967296.0,1,-nbitq), 
to_sfixed(-210185203.0/4294967296.0,1,-nbitq), 
to_sfixed(-492748255.0/4294967296.0,1,-nbitq), 
to_sfixed(112873944.0/4294967296.0,1,-nbitq), 
to_sfixed(1208586741.0/4294967296.0,1,-nbitq), 
to_sfixed(-316609293.0/4294967296.0,1,-nbitq), 
to_sfixed(90858664.0/4294967296.0,1,-nbitq), 
to_sfixed(482565704.0/4294967296.0,1,-nbitq), 
to_sfixed(-176884224.0/4294967296.0,1,-nbitq), 
to_sfixed(349638861.0/4294967296.0,1,-nbitq), 
to_sfixed(633824574.0/4294967296.0,1,-nbitq), 
to_sfixed(699299914.0/4294967296.0,1,-nbitq), 
to_sfixed(-100509305.0/4294967296.0,1,-nbitq), 
to_sfixed(-966103035.0/4294967296.0,1,-nbitq), 
to_sfixed(-17618755.0/4294967296.0,1,-nbitq), 
to_sfixed(-237045130.0/4294967296.0,1,-nbitq), 
to_sfixed(-795075561.0/4294967296.0,1,-nbitq), 
to_sfixed(-895723015.0/4294967296.0,1,-nbitq), 
to_sfixed(-238134857.0/4294967296.0,1,-nbitq), 
to_sfixed(-35329992.0/4294967296.0,1,-nbitq), 
to_sfixed(-226032790.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-443411963.0/4294967296.0,1,-nbitq), 
to_sfixed(2172653375.0/4294967296.0,1,-nbitq), 
to_sfixed(-1495892332.0/4294967296.0,1,-nbitq), 
to_sfixed(419991333.0/4294967296.0,1,-nbitq), 
to_sfixed(1109045725.0/4294967296.0,1,-nbitq), 
to_sfixed(136843797.0/4294967296.0,1,-nbitq), 
to_sfixed(104282488.0/4294967296.0,1,-nbitq), 
to_sfixed(-209686874.0/4294967296.0,1,-nbitq), 
to_sfixed(-401437184.0/4294967296.0,1,-nbitq), 
to_sfixed(-337810479.0/4294967296.0,1,-nbitq), 
to_sfixed(-1115969719.0/4294967296.0,1,-nbitq), 
to_sfixed(366590371.0/4294967296.0,1,-nbitq), 
to_sfixed(-124903841.0/4294967296.0,1,-nbitq), 
to_sfixed(-259085550.0/4294967296.0,1,-nbitq), 
to_sfixed(-71024573.0/4294967296.0,1,-nbitq), 
to_sfixed(644342303.0/4294967296.0,1,-nbitq), 
to_sfixed(46333823.0/4294967296.0,1,-nbitq), 
to_sfixed(-50890084.0/4294967296.0,1,-nbitq), 
to_sfixed(27234925.0/4294967296.0,1,-nbitq), 
to_sfixed(-362128062.0/4294967296.0,1,-nbitq), 
to_sfixed(-222135954.0/4294967296.0,1,-nbitq), 
to_sfixed(-545901731.0/4294967296.0,1,-nbitq), 
to_sfixed(898136670.0/4294967296.0,1,-nbitq), 
to_sfixed(-1446080983.0/4294967296.0,1,-nbitq), 
to_sfixed(-43804637.0/4294967296.0,1,-nbitq), 
to_sfixed(-622507179.0/4294967296.0,1,-nbitq), 
to_sfixed(-200147346.0/4294967296.0,1,-nbitq), 
to_sfixed(-524082247.0/4294967296.0,1,-nbitq), 
to_sfixed(-219793351.0/4294967296.0,1,-nbitq), 
to_sfixed(1065935991.0/4294967296.0,1,-nbitq), 
to_sfixed(-1075827467.0/4294967296.0,1,-nbitq), 
to_sfixed(1362149332.0/4294967296.0,1,-nbitq), 
to_sfixed(81165908.0/4294967296.0,1,-nbitq), 
to_sfixed(-133154119.0/4294967296.0,1,-nbitq), 
to_sfixed(506129511.0/4294967296.0,1,-nbitq), 
to_sfixed(-708113029.0/4294967296.0,1,-nbitq), 
to_sfixed(-217160831.0/4294967296.0,1,-nbitq), 
to_sfixed(49268553.0/4294967296.0,1,-nbitq), 
to_sfixed(31944794.0/4294967296.0,1,-nbitq), 
to_sfixed(-443695964.0/4294967296.0,1,-nbitq), 
to_sfixed(-1119967582.0/4294967296.0,1,-nbitq), 
to_sfixed(-290666626.0/4294967296.0,1,-nbitq), 
to_sfixed(-322758118.0/4294967296.0,1,-nbitq), 
to_sfixed(-451600617.0/4294967296.0,1,-nbitq), 
to_sfixed(-639882202.0/4294967296.0,1,-nbitq), 
to_sfixed(-487200485.0/4294967296.0,1,-nbitq), 
to_sfixed(-255605821.0/4294967296.0,1,-nbitq), 
to_sfixed(1443841765.0/4294967296.0,1,-nbitq), 
to_sfixed(221253605.0/4294967296.0,1,-nbitq), 
to_sfixed(806011979.0/4294967296.0,1,-nbitq), 
to_sfixed(-30152959.0/4294967296.0,1,-nbitq), 
to_sfixed(-285798150.0/4294967296.0,1,-nbitq), 
to_sfixed(1106409965.0/4294967296.0,1,-nbitq), 
to_sfixed(-57396505.0/4294967296.0,1,-nbitq), 
to_sfixed(-286610364.0/4294967296.0,1,-nbitq), 
to_sfixed(-492833288.0/4294967296.0,1,-nbitq), 
to_sfixed(-392679066.0/4294967296.0,1,-nbitq), 
to_sfixed(-241733931.0/4294967296.0,1,-nbitq), 
to_sfixed(-38809610.0/4294967296.0,1,-nbitq), 
to_sfixed(264354641.0/4294967296.0,1,-nbitq), 
to_sfixed(326515807.0/4294967296.0,1,-nbitq), 
to_sfixed(-243748664.0/4294967296.0,1,-nbitq), 
to_sfixed(-470577503.0/4294967296.0,1,-nbitq), 
to_sfixed(1155110426.0/4294967296.0,1,-nbitq), 
to_sfixed(-113207450.0/4294967296.0,1,-nbitq), 
to_sfixed(55632449.0/4294967296.0,1,-nbitq), 
to_sfixed(-1940676144.0/4294967296.0,1,-nbitq), 
to_sfixed(-281553303.0/4294967296.0,1,-nbitq), 
to_sfixed(-164172255.0/4294967296.0,1,-nbitq), 
to_sfixed(-439641026.0/4294967296.0,1,-nbitq), 
to_sfixed(-160141189.0/4294967296.0,1,-nbitq), 
to_sfixed(15496082.0/4294967296.0,1,-nbitq), 
to_sfixed(-1692675421.0/4294967296.0,1,-nbitq), 
to_sfixed(223474020.0/4294967296.0,1,-nbitq), 
to_sfixed(-223273872.0/4294967296.0,1,-nbitq), 
to_sfixed(-86494098.0/4294967296.0,1,-nbitq), 
to_sfixed(-1821627846.0/4294967296.0,1,-nbitq), 
to_sfixed(276851228.0/4294967296.0,1,-nbitq), 
to_sfixed(-11532838.0/4294967296.0,1,-nbitq), 
to_sfixed(-234850441.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-441576498.0/4294967296.0,1,-nbitq), 
to_sfixed(1677724388.0/4294967296.0,1,-nbitq), 
to_sfixed(-996726084.0/4294967296.0,1,-nbitq), 
to_sfixed(-26279152.0/4294967296.0,1,-nbitq), 
to_sfixed(432306366.0/4294967296.0,1,-nbitq), 
to_sfixed(-536180283.0/4294967296.0,1,-nbitq), 
to_sfixed(68008336.0/4294967296.0,1,-nbitq), 
to_sfixed(-621211839.0/4294967296.0,1,-nbitq), 
to_sfixed(-991084174.0/4294967296.0,1,-nbitq), 
to_sfixed(241847674.0/4294967296.0,1,-nbitq), 
to_sfixed(25758565.0/4294967296.0,1,-nbitq), 
to_sfixed(744315059.0/4294967296.0,1,-nbitq), 
to_sfixed(579898786.0/4294967296.0,1,-nbitq), 
to_sfixed(-1481755812.0/4294967296.0,1,-nbitq), 
to_sfixed(546342080.0/4294967296.0,1,-nbitq), 
to_sfixed(204623256.0/4294967296.0,1,-nbitq), 
to_sfixed(-114308999.0/4294967296.0,1,-nbitq), 
to_sfixed(-133892794.0/4294967296.0,1,-nbitq), 
to_sfixed(629545938.0/4294967296.0,1,-nbitq), 
to_sfixed(218746704.0/4294967296.0,1,-nbitq), 
to_sfixed(-422936667.0/4294967296.0,1,-nbitq), 
to_sfixed(249260238.0/4294967296.0,1,-nbitq), 
to_sfixed(176457374.0/4294967296.0,1,-nbitq), 
to_sfixed(-1392222124.0/4294967296.0,1,-nbitq), 
to_sfixed(19133541.0/4294967296.0,1,-nbitq), 
to_sfixed(557561147.0/4294967296.0,1,-nbitq), 
to_sfixed(-936064372.0/4294967296.0,1,-nbitq), 
to_sfixed(-157801130.0/4294967296.0,1,-nbitq), 
to_sfixed(-520967836.0/4294967296.0,1,-nbitq), 
to_sfixed(661521982.0/4294967296.0,1,-nbitq), 
to_sfixed(-1476999201.0/4294967296.0,1,-nbitq), 
to_sfixed(1361533381.0/4294967296.0,1,-nbitq), 
to_sfixed(-572767162.0/4294967296.0,1,-nbitq), 
to_sfixed(-34050590.0/4294967296.0,1,-nbitq), 
to_sfixed(336946016.0/4294967296.0,1,-nbitq), 
to_sfixed(-1263545454.0/4294967296.0,1,-nbitq), 
to_sfixed(-529510818.0/4294967296.0,1,-nbitq), 
to_sfixed(-80790582.0/4294967296.0,1,-nbitq), 
to_sfixed(-78675160.0/4294967296.0,1,-nbitq), 
to_sfixed(33065766.0/4294967296.0,1,-nbitq), 
to_sfixed(-645116968.0/4294967296.0,1,-nbitq), 
to_sfixed(179263179.0/4294967296.0,1,-nbitq), 
to_sfixed(-444123639.0/4294967296.0,1,-nbitq), 
to_sfixed(25321048.0/4294967296.0,1,-nbitq), 
to_sfixed(-801016898.0/4294967296.0,1,-nbitq), 
to_sfixed(-177405177.0/4294967296.0,1,-nbitq), 
to_sfixed(117976316.0/4294967296.0,1,-nbitq), 
to_sfixed(1490842811.0/4294967296.0,1,-nbitq), 
to_sfixed(-776937129.0/4294967296.0,1,-nbitq), 
to_sfixed(504953803.0/4294967296.0,1,-nbitq), 
to_sfixed(-231254020.0/4294967296.0,1,-nbitq), 
to_sfixed(-1066383365.0/4294967296.0,1,-nbitq), 
to_sfixed(493446101.0/4294967296.0,1,-nbitq), 
to_sfixed(-439225357.0/4294967296.0,1,-nbitq), 
to_sfixed(-1218487502.0/4294967296.0,1,-nbitq), 
to_sfixed(378744079.0/4294967296.0,1,-nbitq), 
to_sfixed(-127738424.0/4294967296.0,1,-nbitq), 
to_sfixed(-176566330.0/4294967296.0,1,-nbitq), 
to_sfixed(-256264623.0/4294967296.0,1,-nbitq), 
to_sfixed(-309057860.0/4294967296.0,1,-nbitq), 
to_sfixed(-371787208.0/4294967296.0,1,-nbitq), 
to_sfixed(70980622.0/4294967296.0,1,-nbitq), 
to_sfixed(203911587.0/4294967296.0,1,-nbitq), 
to_sfixed(686302492.0/4294967296.0,1,-nbitq), 
to_sfixed(-466403250.0/4294967296.0,1,-nbitq), 
to_sfixed(-253280433.0/4294967296.0,1,-nbitq), 
to_sfixed(-1501910577.0/4294967296.0,1,-nbitq), 
to_sfixed(-331370527.0/4294967296.0,1,-nbitq), 
to_sfixed(314952443.0/4294967296.0,1,-nbitq), 
to_sfixed(-474183149.0/4294967296.0,1,-nbitq), 
to_sfixed(-78584170.0/4294967296.0,1,-nbitq), 
to_sfixed(-69657237.0/4294967296.0,1,-nbitq), 
to_sfixed(-670565727.0/4294967296.0,1,-nbitq), 
to_sfixed(-62114956.0/4294967296.0,1,-nbitq), 
to_sfixed(410489520.0/4294967296.0,1,-nbitq), 
to_sfixed(1104603535.0/4294967296.0,1,-nbitq), 
to_sfixed(-1870812862.0/4294967296.0,1,-nbitq), 
to_sfixed(92313260.0/4294967296.0,1,-nbitq), 
to_sfixed(-371221939.0/4294967296.0,1,-nbitq), 
to_sfixed(-349829517.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(179554715.0/4294967296.0,1,-nbitq), 
to_sfixed(1293288057.0/4294967296.0,1,-nbitq), 
to_sfixed(-1228871702.0/4294967296.0,1,-nbitq), 
to_sfixed(-128054892.0/4294967296.0,1,-nbitq), 
to_sfixed(-332859652.0/4294967296.0,1,-nbitq), 
to_sfixed(-7829687.0/4294967296.0,1,-nbitq), 
to_sfixed(-374793443.0/4294967296.0,1,-nbitq), 
to_sfixed(-5108902.0/4294967296.0,1,-nbitq), 
to_sfixed(-957530833.0/4294967296.0,1,-nbitq), 
to_sfixed(265589790.0/4294967296.0,1,-nbitq), 
to_sfixed(-227004358.0/4294967296.0,1,-nbitq), 
to_sfixed(1084757032.0/4294967296.0,1,-nbitq), 
to_sfixed(311803258.0/4294967296.0,1,-nbitq), 
to_sfixed(-1741112785.0/4294967296.0,1,-nbitq), 
to_sfixed(42774085.0/4294967296.0,1,-nbitq), 
to_sfixed(183200223.0/4294967296.0,1,-nbitq), 
to_sfixed(75776120.0/4294967296.0,1,-nbitq), 
to_sfixed(-99927215.0/4294967296.0,1,-nbitq), 
to_sfixed(285948564.0/4294967296.0,1,-nbitq), 
to_sfixed(-477480949.0/4294967296.0,1,-nbitq), 
to_sfixed(288599040.0/4294967296.0,1,-nbitq), 
to_sfixed(732817232.0/4294967296.0,1,-nbitq), 
to_sfixed(-723935650.0/4294967296.0,1,-nbitq), 
to_sfixed(-876005380.0/4294967296.0,1,-nbitq), 
to_sfixed(27229369.0/4294967296.0,1,-nbitq), 
to_sfixed(474148998.0/4294967296.0,1,-nbitq), 
to_sfixed(-751391363.0/4294967296.0,1,-nbitq), 
to_sfixed(692069643.0/4294967296.0,1,-nbitq), 
to_sfixed(-815468260.0/4294967296.0,1,-nbitq), 
to_sfixed(821829324.0/4294967296.0,1,-nbitq), 
to_sfixed(-756991093.0/4294967296.0,1,-nbitq), 
to_sfixed(1510780636.0/4294967296.0,1,-nbitq), 
to_sfixed(-58427872.0/4294967296.0,1,-nbitq), 
to_sfixed(211175600.0/4294967296.0,1,-nbitq), 
to_sfixed(149712513.0/4294967296.0,1,-nbitq), 
to_sfixed(-513223266.0/4294967296.0,1,-nbitq), 
to_sfixed(-224105473.0/4294967296.0,1,-nbitq), 
to_sfixed(-506484231.0/4294967296.0,1,-nbitq), 
to_sfixed(540807619.0/4294967296.0,1,-nbitq), 
to_sfixed(-159655576.0/4294967296.0,1,-nbitq), 
to_sfixed(-149099699.0/4294967296.0,1,-nbitq), 
to_sfixed(691319056.0/4294967296.0,1,-nbitq), 
to_sfixed(-794970933.0/4294967296.0,1,-nbitq), 
to_sfixed(-647188159.0/4294967296.0,1,-nbitq), 
to_sfixed(-542266260.0/4294967296.0,1,-nbitq), 
to_sfixed(693396971.0/4294967296.0,1,-nbitq), 
to_sfixed(180933396.0/4294967296.0,1,-nbitq), 
to_sfixed(859052670.0/4294967296.0,1,-nbitq), 
to_sfixed(-648312647.0/4294967296.0,1,-nbitq), 
to_sfixed(864481123.0/4294967296.0,1,-nbitq), 
to_sfixed(83772497.0/4294967296.0,1,-nbitq), 
to_sfixed(-373379124.0/4294967296.0,1,-nbitq), 
to_sfixed(674917497.0/4294967296.0,1,-nbitq), 
to_sfixed(-397172923.0/4294967296.0,1,-nbitq), 
to_sfixed(-938600760.0/4294967296.0,1,-nbitq), 
to_sfixed(288656279.0/4294967296.0,1,-nbitq), 
to_sfixed(430633078.0/4294967296.0,1,-nbitq), 
to_sfixed(264899766.0/4294967296.0,1,-nbitq), 
to_sfixed(78875119.0/4294967296.0,1,-nbitq), 
to_sfixed(35621702.0/4294967296.0,1,-nbitq), 
to_sfixed(-512028882.0/4294967296.0,1,-nbitq), 
to_sfixed(277188827.0/4294967296.0,1,-nbitq), 
to_sfixed(163797093.0/4294967296.0,1,-nbitq), 
to_sfixed(30536568.0/4294967296.0,1,-nbitq), 
to_sfixed(-110330860.0/4294967296.0,1,-nbitq), 
to_sfixed(-418860257.0/4294967296.0,1,-nbitq), 
to_sfixed(-1107052636.0/4294967296.0,1,-nbitq), 
to_sfixed(-267867068.0/4294967296.0,1,-nbitq), 
to_sfixed(80006311.0/4294967296.0,1,-nbitq), 
to_sfixed(349738165.0/4294967296.0,1,-nbitq), 
to_sfixed(163637182.0/4294967296.0,1,-nbitq), 
to_sfixed(162645589.0/4294967296.0,1,-nbitq), 
to_sfixed(-445174538.0/4294967296.0,1,-nbitq), 
to_sfixed(-352490774.0/4294967296.0,1,-nbitq), 
to_sfixed(-76529525.0/4294967296.0,1,-nbitq), 
to_sfixed(1127684334.0/4294967296.0,1,-nbitq), 
to_sfixed(-1192766033.0/4294967296.0,1,-nbitq), 
to_sfixed(179957229.0/4294967296.0,1,-nbitq), 
to_sfixed(-503053602.0/4294967296.0,1,-nbitq), 
to_sfixed(180327730.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-524559252.0/4294967296.0,1,-nbitq), 
to_sfixed(688907114.0/4294967296.0,1,-nbitq), 
to_sfixed(-1027117248.0/4294967296.0,1,-nbitq), 
to_sfixed(-348352914.0/4294967296.0,1,-nbitq), 
to_sfixed(-991612949.0/4294967296.0,1,-nbitq), 
to_sfixed(-711157599.0/4294967296.0,1,-nbitq), 
to_sfixed(-382041071.0/4294967296.0,1,-nbitq), 
to_sfixed(415124853.0/4294967296.0,1,-nbitq), 
to_sfixed(-1908081307.0/4294967296.0,1,-nbitq), 
to_sfixed(-68039336.0/4294967296.0,1,-nbitq), 
to_sfixed(-619921171.0/4294967296.0,1,-nbitq), 
to_sfixed(382268737.0/4294967296.0,1,-nbitq), 
to_sfixed(-576001335.0/4294967296.0,1,-nbitq), 
to_sfixed(-1027241862.0/4294967296.0,1,-nbitq), 
to_sfixed(317099577.0/4294967296.0,1,-nbitq), 
to_sfixed(348810117.0/4294967296.0,1,-nbitq), 
to_sfixed(-362069854.0/4294967296.0,1,-nbitq), 
to_sfixed(-11942694.0/4294967296.0,1,-nbitq), 
to_sfixed(240117673.0/4294967296.0,1,-nbitq), 
to_sfixed(-507646081.0/4294967296.0,1,-nbitq), 
to_sfixed(-334742700.0/4294967296.0,1,-nbitq), 
to_sfixed(-262356028.0/4294967296.0,1,-nbitq), 
to_sfixed(-770612314.0/4294967296.0,1,-nbitq), 
to_sfixed(-310925610.0/4294967296.0,1,-nbitq), 
to_sfixed(29055391.0/4294967296.0,1,-nbitq), 
to_sfixed(355903264.0/4294967296.0,1,-nbitq), 
to_sfixed(-519521696.0/4294967296.0,1,-nbitq), 
to_sfixed(901838775.0/4294967296.0,1,-nbitq), 
to_sfixed(-703402799.0/4294967296.0,1,-nbitq), 
to_sfixed(-474474069.0/4294967296.0,1,-nbitq), 
to_sfixed(151883259.0/4294967296.0,1,-nbitq), 
to_sfixed(454805480.0/4294967296.0,1,-nbitq), 
to_sfixed(69048217.0/4294967296.0,1,-nbitq), 
to_sfixed(222271257.0/4294967296.0,1,-nbitq), 
to_sfixed(147856308.0/4294967296.0,1,-nbitq), 
to_sfixed(588340759.0/4294967296.0,1,-nbitq), 
to_sfixed(-467450592.0/4294967296.0,1,-nbitq), 
to_sfixed(-109238738.0/4294967296.0,1,-nbitq), 
to_sfixed(30746155.0/4294967296.0,1,-nbitq), 
to_sfixed(-34630492.0/4294967296.0,1,-nbitq), 
to_sfixed(-296834806.0/4294967296.0,1,-nbitq), 
to_sfixed(270357708.0/4294967296.0,1,-nbitq), 
to_sfixed(-517117904.0/4294967296.0,1,-nbitq), 
to_sfixed(-1032201919.0/4294967296.0,1,-nbitq), 
to_sfixed(-829889807.0/4294967296.0,1,-nbitq), 
to_sfixed(-554036779.0/4294967296.0,1,-nbitq), 
to_sfixed(192819863.0/4294967296.0,1,-nbitq), 
to_sfixed(313134405.0/4294967296.0,1,-nbitq), 
to_sfixed(-474419574.0/4294967296.0,1,-nbitq), 
to_sfixed(1020425682.0/4294967296.0,1,-nbitq), 
to_sfixed(-304127247.0/4294967296.0,1,-nbitq), 
to_sfixed(-165138513.0/4294967296.0,1,-nbitq), 
to_sfixed(189662623.0/4294967296.0,1,-nbitq), 
to_sfixed(-127828866.0/4294967296.0,1,-nbitq), 
to_sfixed(-845960750.0/4294967296.0,1,-nbitq), 
to_sfixed(-76909802.0/4294967296.0,1,-nbitq), 
to_sfixed(298602921.0/4294967296.0,1,-nbitq), 
to_sfixed(-421897264.0/4294967296.0,1,-nbitq), 
to_sfixed(163151682.0/4294967296.0,1,-nbitq), 
to_sfixed(303739607.0/4294967296.0,1,-nbitq), 
to_sfixed(-206957192.0/4294967296.0,1,-nbitq), 
to_sfixed(48064101.0/4294967296.0,1,-nbitq), 
to_sfixed(410336071.0/4294967296.0,1,-nbitq), 
to_sfixed(-646142973.0/4294967296.0,1,-nbitq), 
to_sfixed(86548254.0/4294967296.0,1,-nbitq), 
to_sfixed(-210927763.0/4294967296.0,1,-nbitq), 
to_sfixed(-361104766.0/4294967296.0,1,-nbitq), 
to_sfixed(-535631888.0/4294967296.0,1,-nbitq), 
to_sfixed(101344258.0/4294967296.0,1,-nbitq), 
to_sfixed(675519649.0/4294967296.0,1,-nbitq), 
to_sfixed(-843485878.0/4294967296.0,1,-nbitq), 
to_sfixed(367499381.0/4294967296.0,1,-nbitq), 
to_sfixed(224070791.0/4294967296.0,1,-nbitq), 
to_sfixed(-323368404.0/4294967296.0,1,-nbitq), 
to_sfixed(-165197245.0/4294967296.0,1,-nbitq), 
to_sfixed(1074598118.0/4294967296.0,1,-nbitq), 
to_sfixed(-2051610607.0/4294967296.0,1,-nbitq), 
to_sfixed(264743779.0/4294967296.0,1,-nbitq), 
to_sfixed(146417601.0/4294967296.0,1,-nbitq), 
to_sfixed(-384382916.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-167113823.0/4294967296.0,1,-nbitq), 
to_sfixed(839354001.0/4294967296.0,1,-nbitq), 
to_sfixed(-1562711643.0/4294967296.0,1,-nbitq), 
to_sfixed(-1286265668.0/4294967296.0,1,-nbitq), 
to_sfixed(-1454710140.0/4294967296.0,1,-nbitq), 
to_sfixed(-399086643.0/4294967296.0,1,-nbitq), 
to_sfixed(162876806.0/4294967296.0,1,-nbitq), 
to_sfixed(896678477.0/4294967296.0,1,-nbitq), 
to_sfixed(-1236334326.0/4294967296.0,1,-nbitq), 
to_sfixed(-270973098.0/4294967296.0,1,-nbitq), 
to_sfixed(-966165.0/4294967296.0,1,-nbitq), 
to_sfixed(64375102.0/4294967296.0,1,-nbitq), 
to_sfixed(-168272986.0/4294967296.0,1,-nbitq), 
to_sfixed(-927039991.0/4294967296.0,1,-nbitq), 
to_sfixed(186030514.0/4294967296.0,1,-nbitq), 
to_sfixed(-109987196.0/4294967296.0,1,-nbitq), 
to_sfixed(356721321.0/4294967296.0,1,-nbitq), 
to_sfixed(231468744.0/4294967296.0,1,-nbitq), 
to_sfixed(638216064.0/4294967296.0,1,-nbitq), 
to_sfixed(248649792.0/4294967296.0,1,-nbitq), 
to_sfixed(-198257603.0/4294967296.0,1,-nbitq), 
to_sfixed(-823014012.0/4294967296.0,1,-nbitq), 
to_sfixed(-829814634.0/4294967296.0,1,-nbitq), 
to_sfixed(-966608193.0/4294967296.0,1,-nbitq), 
to_sfixed(-311653642.0/4294967296.0,1,-nbitq), 
to_sfixed(-136444302.0/4294967296.0,1,-nbitq), 
to_sfixed(90728200.0/4294967296.0,1,-nbitq), 
to_sfixed(827461546.0/4294967296.0,1,-nbitq), 
to_sfixed(-206322630.0/4294967296.0,1,-nbitq), 
to_sfixed(-545547807.0/4294967296.0,1,-nbitq), 
to_sfixed(513379903.0/4294967296.0,1,-nbitq), 
to_sfixed(877804162.0/4294967296.0,1,-nbitq), 
to_sfixed(-404894270.0/4294967296.0,1,-nbitq), 
to_sfixed(1125274143.0/4294967296.0,1,-nbitq), 
to_sfixed(-282607092.0/4294967296.0,1,-nbitq), 
to_sfixed(485850191.0/4294967296.0,1,-nbitq), 
to_sfixed(-772387461.0/4294967296.0,1,-nbitq), 
to_sfixed(163914332.0/4294967296.0,1,-nbitq), 
to_sfixed(-8870917.0/4294967296.0,1,-nbitq), 
to_sfixed(-250643620.0/4294967296.0,1,-nbitq), 
to_sfixed(9602137.0/4294967296.0,1,-nbitq), 
to_sfixed(132765175.0/4294967296.0,1,-nbitq), 
to_sfixed(-604039722.0/4294967296.0,1,-nbitq), 
to_sfixed(-1078728627.0/4294967296.0,1,-nbitq), 
to_sfixed(-1172877551.0/4294967296.0,1,-nbitq), 
to_sfixed(-833106719.0/4294967296.0,1,-nbitq), 
to_sfixed(-434322292.0/4294967296.0,1,-nbitq), 
to_sfixed(570966345.0/4294967296.0,1,-nbitq), 
to_sfixed(-238131092.0/4294967296.0,1,-nbitq), 
to_sfixed(645467526.0/4294967296.0,1,-nbitq), 
to_sfixed(-136607134.0/4294967296.0,1,-nbitq), 
to_sfixed(-236963505.0/4294967296.0,1,-nbitq), 
to_sfixed(187660628.0/4294967296.0,1,-nbitq), 
to_sfixed(371772122.0/4294967296.0,1,-nbitq), 
to_sfixed(20542901.0/4294967296.0,1,-nbitq), 
to_sfixed(-307762149.0/4294967296.0,1,-nbitq), 
to_sfixed(994706948.0/4294967296.0,1,-nbitq), 
to_sfixed(-148833271.0/4294967296.0,1,-nbitq), 
to_sfixed(-17392901.0/4294967296.0,1,-nbitq), 
to_sfixed(19552459.0/4294967296.0,1,-nbitq), 
to_sfixed(-337730506.0/4294967296.0,1,-nbitq), 
to_sfixed(-915234049.0/4294967296.0,1,-nbitq), 
to_sfixed(320397996.0/4294967296.0,1,-nbitq), 
to_sfixed(-877466207.0/4294967296.0,1,-nbitq), 
to_sfixed(193494365.0/4294967296.0,1,-nbitq), 
to_sfixed(100367304.0/4294967296.0,1,-nbitq), 
to_sfixed(727987083.0/4294967296.0,1,-nbitq), 
to_sfixed(-333143441.0/4294967296.0,1,-nbitq), 
to_sfixed(324181253.0/4294967296.0,1,-nbitq), 
to_sfixed(982511426.0/4294967296.0,1,-nbitq), 
to_sfixed(-656188353.0/4294967296.0,1,-nbitq), 
to_sfixed(85862214.0/4294967296.0,1,-nbitq), 
to_sfixed(635730529.0/4294967296.0,1,-nbitq), 
to_sfixed(256913738.0/4294967296.0,1,-nbitq), 
to_sfixed(391038547.0/4294967296.0,1,-nbitq), 
to_sfixed(656271468.0/4294967296.0,1,-nbitq), 
to_sfixed(-806223509.0/4294967296.0,1,-nbitq), 
to_sfixed(246208935.0/4294967296.0,1,-nbitq), 
to_sfixed(-455157928.0/4294967296.0,1,-nbitq), 
to_sfixed(17074835.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-242236807.0/4294967296.0,1,-nbitq), 
to_sfixed(1162833247.0/4294967296.0,1,-nbitq), 
to_sfixed(-1298376823.0/4294967296.0,1,-nbitq), 
to_sfixed(-1884516791.0/4294967296.0,1,-nbitq), 
to_sfixed(-664082352.0/4294967296.0,1,-nbitq), 
to_sfixed(-847885039.0/4294967296.0,1,-nbitq), 
to_sfixed(-376922870.0/4294967296.0,1,-nbitq), 
to_sfixed(810944013.0/4294967296.0,1,-nbitq), 
to_sfixed(-913600071.0/4294967296.0,1,-nbitq), 
to_sfixed(-97043287.0/4294967296.0,1,-nbitq), 
to_sfixed(848253982.0/4294967296.0,1,-nbitq), 
to_sfixed(-104210787.0/4294967296.0,1,-nbitq), 
to_sfixed(362591954.0/4294967296.0,1,-nbitq), 
to_sfixed(-997969897.0/4294967296.0,1,-nbitq), 
to_sfixed(-96576189.0/4294967296.0,1,-nbitq), 
to_sfixed(7547402.0/4294967296.0,1,-nbitq), 
to_sfixed(376518260.0/4294967296.0,1,-nbitq), 
to_sfixed(-361708369.0/4294967296.0,1,-nbitq), 
to_sfixed(386865252.0/4294967296.0,1,-nbitq), 
to_sfixed(-108321319.0/4294967296.0,1,-nbitq), 
to_sfixed(30706187.0/4294967296.0,1,-nbitq), 
to_sfixed(-100082488.0/4294967296.0,1,-nbitq), 
to_sfixed(-5774929.0/4294967296.0,1,-nbitq), 
to_sfixed(-1334553511.0/4294967296.0,1,-nbitq), 
to_sfixed(-240852491.0/4294967296.0,1,-nbitq), 
to_sfixed(-887465942.0/4294967296.0,1,-nbitq), 
to_sfixed(140205183.0/4294967296.0,1,-nbitq), 
to_sfixed(576604228.0/4294967296.0,1,-nbitq), 
to_sfixed(69589660.0/4294967296.0,1,-nbitq), 
to_sfixed(314163704.0/4294967296.0,1,-nbitq), 
to_sfixed(488657822.0/4294967296.0,1,-nbitq), 
to_sfixed(891658916.0/4294967296.0,1,-nbitq), 
to_sfixed(-559958855.0/4294967296.0,1,-nbitq), 
to_sfixed(1007991786.0/4294967296.0,1,-nbitq), 
to_sfixed(-372155920.0/4294967296.0,1,-nbitq), 
to_sfixed(3569143.0/4294967296.0,1,-nbitq), 
to_sfixed(-399224508.0/4294967296.0,1,-nbitq), 
to_sfixed(-566534736.0/4294967296.0,1,-nbitq), 
to_sfixed(207069902.0/4294967296.0,1,-nbitq), 
to_sfixed(280883290.0/4294967296.0,1,-nbitq), 
to_sfixed(-200042926.0/4294967296.0,1,-nbitq), 
to_sfixed(-223313019.0/4294967296.0,1,-nbitq), 
to_sfixed(-736476145.0/4294967296.0,1,-nbitq), 
to_sfixed(-1025674205.0/4294967296.0,1,-nbitq), 
to_sfixed(-557733292.0/4294967296.0,1,-nbitq), 
to_sfixed(-271213462.0/4294967296.0,1,-nbitq), 
to_sfixed(99347511.0/4294967296.0,1,-nbitq), 
to_sfixed(198628114.0/4294967296.0,1,-nbitq), 
to_sfixed(-228465007.0/4294967296.0,1,-nbitq), 
to_sfixed(407700727.0/4294967296.0,1,-nbitq), 
to_sfixed(-126290114.0/4294967296.0,1,-nbitq), 
to_sfixed(-783184694.0/4294967296.0,1,-nbitq), 
to_sfixed(418575125.0/4294967296.0,1,-nbitq), 
to_sfixed(-806362568.0/4294967296.0,1,-nbitq), 
to_sfixed(-540735903.0/4294967296.0,1,-nbitq), 
to_sfixed(264518712.0/4294967296.0,1,-nbitq), 
to_sfixed(753925178.0/4294967296.0,1,-nbitq), 
to_sfixed(-204913724.0/4294967296.0,1,-nbitq), 
to_sfixed(-390433436.0/4294967296.0,1,-nbitq), 
to_sfixed(-31566914.0/4294967296.0,1,-nbitq), 
to_sfixed(-372303969.0/4294967296.0,1,-nbitq), 
to_sfixed(-764369921.0/4294967296.0,1,-nbitq), 
to_sfixed(54223424.0/4294967296.0,1,-nbitq), 
to_sfixed(-424660158.0/4294967296.0,1,-nbitq), 
to_sfixed(-283923346.0/4294967296.0,1,-nbitq), 
to_sfixed(-74423209.0/4294967296.0,1,-nbitq), 
to_sfixed(-168363048.0/4294967296.0,1,-nbitq), 
to_sfixed(1426276.0/4294967296.0,1,-nbitq), 
to_sfixed(357871806.0/4294967296.0,1,-nbitq), 
to_sfixed(970867277.0/4294967296.0,1,-nbitq), 
to_sfixed(-305252876.0/4294967296.0,1,-nbitq), 
to_sfixed(200933603.0/4294967296.0,1,-nbitq), 
to_sfixed(701689247.0/4294967296.0,1,-nbitq), 
to_sfixed(68935217.0/4294967296.0,1,-nbitq), 
to_sfixed(233811268.0/4294967296.0,1,-nbitq), 
to_sfixed(575807532.0/4294967296.0,1,-nbitq), 
to_sfixed(-786829336.0/4294967296.0,1,-nbitq), 
to_sfixed(470483271.0/4294967296.0,1,-nbitq), 
to_sfixed(-253427708.0/4294967296.0,1,-nbitq), 
to_sfixed(157261471.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-405408676.0/4294967296.0,1,-nbitq), 
to_sfixed(1144221329.0/4294967296.0,1,-nbitq), 
to_sfixed(-842494323.0/4294967296.0,1,-nbitq), 
to_sfixed(-779229619.0/4294967296.0,1,-nbitq), 
to_sfixed(-821902028.0/4294967296.0,1,-nbitq), 
to_sfixed(-260746337.0/4294967296.0,1,-nbitq), 
to_sfixed(57006430.0/4294967296.0,1,-nbitq), 
to_sfixed(891645299.0/4294967296.0,1,-nbitq), 
to_sfixed(-716388549.0/4294967296.0,1,-nbitq), 
to_sfixed(-16981210.0/4294967296.0,1,-nbitq), 
to_sfixed(398078362.0/4294967296.0,1,-nbitq), 
to_sfixed(162380523.0/4294967296.0,1,-nbitq), 
to_sfixed(29340264.0/4294967296.0,1,-nbitq), 
to_sfixed(-429585121.0/4294967296.0,1,-nbitq), 
to_sfixed(-325663378.0/4294967296.0,1,-nbitq), 
to_sfixed(-206871107.0/4294967296.0,1,-nbitq), 
to_sfixed(-11689383.0/4294967296.0,1,-nbitq), 
to_sfixed(-65363925.0/4294967296.0,1,-nbitq), 
to_sfixed(263743613.0/4294967296.0,1,-nbitq), 
to_sfixed(131530274.0/4294967296.0,1,-nbitq), 
to_sfixed(-36240409.0/4294967296.0,1,-nbitq), 
to_sfixed(38471212.0/4294967296.0,1,-nbitq), 
to_sfixed(179229816.0/4294967296.0,1,-nbitq), 
to_sfixed(-420110682.0/4294967296.0,1,-nbitq), 
to_sfixed(318247352.0/4294967296.0,1,-nbitq), 
to_sfixed(284563928.0/4294967296.0,1,-nbitq), 
to_sfixed(-166380759.0/4294967296.0,1,-nbitq), 
to_sfixed(488682710.0/4294967296.0,1,-nbitq), 
to_sfixed(212140398.0/4294967296.0,1,-nbitq), 
to_sfixed(-23913258.0/4294967296.0,1,-nbitq), 
to_sfixed(-354404311.0/4294967296.0,1,-nbitq), 
to_sfixed(167759663.0/4294967296.0,1,-nbitq), 
to_sfixed(67340878.0/4294967296.0,1,-nbitq), 
to_sfixed(611856034.0/4294967296.0,1,-nbitq), 
to_sfixed(-405719506.0/4294967296.0,1,-nbitq), 
to_sfixed(47725443.0/4294967296.0,1,-nbitq), 
to_sfixed(-506690479.0/4294967296.0,1,-nbitq), 
to_sfixed(-287444721.0/4294967296.0,1,-nbitq), 
to_sfixed(92149357.0/4294967296.0,1,-nbitq), 
to_sfixed(268836838.0/4294967296.0,1,-nbitq), 
to_sfixed(560688557.0/4294967296.0,1,-nbitq), 
to_sfixed(-380876549.0/4294967296.0,1,-nbitq), 
to_sfixed(-823858182.0/4294967296.0,1,-nbitq), 
to_sfixed(-484048785.0/4294967296.0,1,-nbitq), 
to_sfixed(-561708824.0/4294967296.0,1,-nbitq), 
to_sfixed(-869922631.0/4294967296.0,1,-nbitq), 
to_sfixed(-41510270.0/4294967296.0,1,-nbitq), 
to_sfixed(607223412.0/4294967296.0,1,-nbitq), 
to_sfixed(-187778986.0/4294967296.0,1,-nbitq), 
to_sfixed(315888877.0/4294967296.0,1,-nbitq), 
to_sfixed(298499627.0/4294967296.0,1,-nbitq), 
to_sfixed(-627456953.0/4294967296.0,1,-nbitq), 
to_sfixed(369625339.0/4294967296.0,1,-nbitq), 
to_sfixed(-438470893.0/4294967296.0,1,-nbitq), 
to_sfixed(-317445724.0/4294967296.0,1,-nbitq), 
to_sfixed(194027608.0/4294967296.0,1,-nbitq), 
to_sfixed(681919452.0/4294967296.0,1,-nbitq), 
to_sfixed(150592223.0/4294967296.0,1,-nbitq), 
to_sfixed(-36782116.0/4294967296.0,1,-nbitq), 
to_sfixed(217783636.0/4294967296.0,1,-nbitq), 
to_sfixed(85722029.0/4294967296.0,1,-nbitq), 
to_sfixed(-441392284.0/4294967296.0,1,-nbitq), 
to_sfixed(202519931.0/4294967296.0,1,-nbitq), 
to_sfixed(-569107001.0/4294967296.0,1,-nbitq), 
to_sfixed(-291222740.0/4294967296.0,1,-nbitq), 
to_sfixed(-289646259.0/4294967296.0,1,-nbitq), 
to_sfixed(94408227.0/4294967296.0,1,-nbitq), 
to_sfixed(-152969322.0/4294967296.0,1,-nbitq), 
to_sfixed(252099964.0/4294967296.0,1,-nbitq), 
to_sfixed(1005318690.0/4294967296.0,1,-nbitq), 
to_sfixed(-285638661.0/4294967296.0,1,-nbitq), 
to_sfixed(-56175270.0/4294967296.0,1,-nbitq), 
to_sfixed(227217615.0/4294967296.0,1,-nbitq), 
to_sfixed(-357971019.0/4294967296.0,1,-nbitq), 
to_sfixed(435932816.0/4294967296.0,1,-nbitq), 
to_sfixed(-243337010.0/4294967296.0,1,-nbitq), 
to_sfixed(-834315086.0/4294967296.0,1,-nbitq), 
to_sfixed(-724671641.0/4294967296.0,1,-nbitq), 
to_sfixed(-163971217.0/4294967296.0,1,-nbitq), 
to_sfixed(177387617.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(172370866.0/4294967296.0,1,-nbitq), 
to_sfixed(929443980.0/4294967296.0,1,-nbitq), 
to_sfixed(-555015588.0/4294967296.0,1,-nbitq), 
to_sfixed(-38843881.0/4294967296.0,1,-nbitq), 
to_sfixed(-619892175.0/4294967296.0,1,-nbitq), 
to_sfixed(-226182060.0/4294967296.0,1,-nbitq), 
to_sfixed(-332594858.0/4294967296.0,1,-nbitq), 
to_sfixed(388687924.0/4294967296.0,1,-nbitq), 
to_sfixed(-321758881.0/4294967296.0,1,-nbitq), 
to_sfixed(-341665966.0/4294967296.0,1,-nbitq), 
to_sfixed(308011074.0/4294967296.0,1,-nbitq), 
to_sfixed(86459202.0/4294967296.0,1,-nbitq), 
to_sfixed(-21889377.0/4294967296.0,1,-nbitq), 
to_sfixed(-227230608.0/4294967296.0,1,-nbitq), 
to_sfixed(-220012613.0/4294967296.0,1,-nbitq), 
to_sfixed(-262232975.0/4294967296.0,1,-nbitq), 
to_sfixed(-183705906.0/4294967296.0,1,-nbitq), 
to_sfixed(75175347.0/4294967296.0,1,-nbitq), 
to_sfixed(-21641868.0/4294967296.0,1,-nbitq), 
to_sfixed(-229999566.0/4294967296.0,1,-nbitq), 
to_sfixed(187472594.0/4294967296.0,1,-nbitq), 
to_sfixed(-428589847.0/4294967296.0,1,-nbitq), 
to_sfixed(-604593109.0/4294967296.0,1,-nbitq), 
to_sfixed(-409042947.0/4294967296.0,1,-nbitq), 
to_sfixed(-67741735.0/4294967296.0,1,-nbitq), 
to_sfixed(-264872631.0/4294967296.0,1,-nbitq), 
to_sfixed(20494564.0/4294967296.0,1,-nbitq), 
to_sfixed(428630965.0/4294967296.0,1,-nbitq), 
to_sfixed(-201533291.0/4294967296.0,1,-nbitq), 
to_sfixed(-125601977.0/4294967296.0,1,-nbitq), 
to_sfixed(-35324896.0/4294967296.0,1,-nbitq), 
to_sfixed(13918913.0/4294967296.0,1,-nbitq), 
to_sfixed(497544835.0/4294967296.0,1,-nbitq), 
to_sfixed(-64230917.0/4294967296.0,1,-nbitq), 
to_sfixed(-376535393.0/4294967296.0,1,-nbitq), 
to_sfixed(17531421.0/4294967296.0,1,-nbitq), 
to_sfixed(-345000584.0/4294967296.0,1,-nbitq), 
to_sfixed(-363047603.0/4294967296.0,1,-nbitq), 
to_sfixed(270448749.0/4294967296.0,1,-nbitq), 
to_sfixed(-115710169.0/4294967296.0,1,-nbitq), 
to_sfixed(-143176909.0/4294967296.0,1,-nbitq), 
to_sfixed(-486538843.0/4294967296.0,1,-nbitq), 
to_sfixed(-77588793.0/4294967296.0,1,-nbitq), 
to_sfixed(-1126416289.0/4294967296.0,1,-nbitq), 
to_sfixed(4931924.0/4294967296.0,1,-nbitq), 
to_sfixed(-916891697.0/4294967296.0,1,-nbitq), 
to_sfixed(-438045765.0/4294967296.0,1,-nbitq), 
to_sfixed(281075758.0/4294967296.0,1,-nbitq), 
to_sfixed(-390401852.0/4294967296.0,1,-nbitq), 
to_sfixed(116131038.0/4294967296.0,1,-nbitq), 
to_sfixed(54015013.0/4294967296.0,1,-nbitq), 
to_sfixed(352421355.0/4294967296.0,1,-nbitq), 
to_sfixed(10398733.0/4294967296.0,1,-nbitq), 
to_sfixed(15265997.0/4294967296.0,1,-nbitq), 
to_sfixed(-43250883.0/4294967296.0,1,-nbitq), 
to_sfixed(-121766216.0/4294967296.0,1,-nbitq), 
to_sfixed(-284302457.0/4294967296.0,1,-nbitq), 
to_sfixed(340353393.0/4294967296.0,1,-nbitq), 
to_sfixed(29273470.0/4294967296.0,1,-nbitq), 
to_sfixed(160708083.0/4294967296.0,1,-nbitq), 
to_sfixed(208405801.0/4294967296.0,1,-nbitq), 
to_sfixed(-312555019.0/4294967296.0,1,-nbitq), 
to_sfixed(-80941417.0/4294967296.0,1,-nbitq), 
to_sfixed(-90306964.0/4294967296.0,1,-nbitq), 
to_sfixed(-97941420.0/4294967296.0,1,-nbitq), 
to_sfixed(-368633605.0/4294967296.0,1,-nbitq), 
to_sfixed(313536273.0/4294967296.0,1,-nbitq), 
to_sfixed(-362794157.0/4294967296.0,1,-nbitq), 
to_sfixed(-95627599.0/4294967296.0,1,-nbitq), 
to_sfixed(17339604.0/4294967296.0,1,-nbitq), 
to_sfixed(-104012890.0/4294967296.0,1,-nbitq), 
to_sfixed(-334670040.0/4294967296.0,1,-nbitq), 
to_sfixed(493127027.0/4294967296.0,1,-nbitq), 
to_sfixed(261917974.0/4294967296.0,1,-nbitq), 
to_sfixed(33545205.0/4294967296.0,1,-nbitq), 
to_sfixed(-301531564.0/4294967296.0,1,-nbitq), 
to_sfixed(-348175794.0/4294967296.0,1,-nbitq), 
to_sfixed(-288298879.0/4294967296.0,1,-nbitq), 
to_sfixed(36169664.0/4294967296.0,1,-nbitq), 
to_sfixed(-218224831.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-82555042.0/4294967296.0,1,-nbitq), 
to_sfixed(63558955.0/4294967296.0,1,-nbitq), 
to_sfixed(-143425538.0/4294967296.0,1,-nbitq), 
to_sfixed(-245530302.0/4294967296.0,1,-nbitq), 
to_sfixed(-294230740.0/4294967296.0,1,-nbitq), 
to_sfixed(-457459165.0/4294967296.0,1,-nbitq), 
to_sfixed(-83608731.0/4294967296.0,1,-nbitq), 
to_sfixed(279731229.0/4294967296.0,1,-nbitq), 
to_sfixed(-658197847.0/4294967296.0,1,-nbitq), 
to_sfixed(271537869.0/4294967296.0,1,-nbitq), 
to_sfixed(457667188.0/4294967296.0,1,-nbitq), 
to_sfixed(43440579.0/4294967296.0,1,-nbitq), 
to_sfixed(53069542.0/4294967296.0,1,-nbitq), 
to_sfixed(-259210449.0/4294967296.0,1,-nbitq), 
to_sfixed(149122756.0/4294967296.0,1,-nbitq), 
to_sfixed(334968534.0/4294967296.0,1,-nbitq), 
to_sfixed(72955140.0/4294967296.0,1,-nbitq), 
to_sfixed(-298515217.0/4294967296.0,1,-nbitq), 
to_sfixed(482534932.0/4294967296.0,1,-nbitq), 
to_sfixed(-375685319.0/4294967296.0,1,-nbitq), 
to_sfixed(-191854365.0/4294967296.0,1,-nbitq), 
to_sfixed(-352806964.0/4294967296.0,1,-nbitq), 
to_sfixed(-243952278.0/4294967296.0,1,-nbitq), 
to_sfixed(96178567.0/4294967296.0,1,-nbitq), 
to_sfixed(245518810.0/4294967296.0,1,-nbitq), 
to_sfixed(-263202298.0/4294967296.0,1,-nbitq), 
to_sfixed(377981547.0/4294967296.0,1,-nbitq), 
to_sfixed(-49951322.0/4294967296.0,1,-nbitq), 
to_sfixed(611435637.0/4294967296.0,1,-nbitq), 
to_sfixed(-51584688.0/4294967296.0,1,-nbitq), 
to_sfixed(-374591523.0/4294967296.0,1,-nbitq), 
to_sfixed(-10015801.0/4294967296.0,1,-nbitq), 
to_sfixed(-3256661.0/4294967296.0,1,-nbitq), 
to_sfixed(182754892.0/4294967296.0,1,-nbitq), 
to_sfixed(-146733604.0/4294967296.0,1,-nbitq), 
to_sfixed(-618023604.0/4294967296.0,1,-nbitq), 
to_sfixed(-107880444.0/4294967296.0,1,-nbitq), 
to_sfixed(49341880.0/4294967296.0,1,-nbitq), 
to_sfixed(-314067264.0/4294967296.0,1,-nbitq), 
to_sfixed(120131814.0/4294967296.0,1,-nbitq), 
to_sfixed(375043636.0/4294967296.0,1,-nbitq), 
to_sfixed(301466206.0/4294967296.0,1,-nbitq), 
to_sfixed(-506140077.0/4294967296.0,1,-nbitq), 
to_sfixed(-290362168.0/4294967296.0,1,-nbitq), 
to_sfixed(330858145.0/4294967296.0,1,-nbitq), 
to_sfixed(-107438501.0/4294967296.0,1,-nbitq), 
to_sfixed(79858814.0/4294967296.0,1,-nbitq), 
to_sfixed(-301448003.0/4294967296.0,1,-nbitq), 
to_sfixed(76683763.0/4294967296.0,1,-nbitq), 
to_sfixed(138468107.0/4294967296.0,1,-nbitq), 
to_sfixed(292237575.0/4294967296.0,1,-nbitq), 
to_sfixed(-131645856.0/4294967296.0,1,-nbitq), 
to_sfixed(5731464.0/4294967296.0,1,-nbitq), 
to_sfixed(273581710.0/4294967296.0,1,-nbitq), 
to_sfixed(-226795794.0/4294967296.0,1,-nbitq), 
to_sfixed(-238653320.0/4294967296.0,1,-nbitq), 
to_sfixed(10656997.0/4294967296.0,1,-nbitq), 
to_sfixed(16228826.0/4294967296.0,1,-nbitq), 
to_sfixed(85277313.0/4294967296.0,1,-nbitq), 
to_sfixed(-106222719.0/4294967296.0,1,-nbitq), 
to_sfixed(-45714789.0/4294967296.0,1,-nbitq), 
to_sfixed(-155779415.0/4294967296.0,1,-nbitq), 
to_sfixed(346185666.0/4294967296.0,1,-nbitq), 
to_sfixed(-312773237.0/4294967296.0,1,-nbitq), 
to_sfixed(-72854158.0/4294967296.0,1,-nbitq), 
to_sfixed(142257399.0/4294967296.0,1,-nbitq), 
to_sfixed(204461181.0/4294967296.0,1,-nbitq), 
to_sfixed(254250577.0/4294967296.0,1,-nbitq), 
to_sfixed(128273097.0/4294967296.0,1,-nbitq), 
to_sfixed(627691042.0/4294967296.0,1,-nbitq), 
to_sfixed(133067182.0/4294967296.0,1,-nbitq), 
to_sfixed(-109686528.0/4294967296.0,1,-nbitq), 
to_sfixed(353143637.0/4294967296.0,1,-nbitq), 
to_sfixed(47844481.0/4294967296.0,1,-nbitq), 
to_sfixed(-16824801.0/4294967296.0,1,-nbitq), 
to_sfixed(-396744524.0/4294967296.0,1,-nbitq), 
to_sfixed(-422505119.0/4294967296.0,1,-nbitq), 
to_sfixed(-574016863.0/4294967296.0,1,-nbitq), 
to_sfixed(-280347291.0/4294967296.0,1,-nbitq), 
to_sfixed(333107770.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-169358979.0/4294967296.0,1,-nbitq), 
to_sfixed(-138671706.0/4294967296.0,1,-nbitq), 
to_sfixed(-312373337.0/4294967296.0,1,-nbitq), 
to_sfixed(25143962.0/4294967296.0,1,-nbitq), 
to_sfixed(-349300476.0/4294967296.0,1,-nbitq), 
to_sfixed(-173522167.0/4294967296.0,1,-nbitq), 
to_sfixed(-116314603.0/4294967296.0,1,-nbitq), 
to_sfixed(-62216418.0/4294967296.0,1,-nbitq), 
to_sfixed(-121483936.0/4294967296.0,1,-nbitq), 
to_sfixed(-356749580.0/4294967296.0,1,-nbitq), 
to_sfixed(202286041.0/4294967296.0,1,-nbitq), 
to_sfixed(-278751449.0/4294967296.0,1,-nbitq), 
to_sfixed(-1800061.0/4294967296.0,1,-nbitq), 
to_sfixed(-413878350.0/4294967296.0,1,-nbitq), 
to_sfixed(-397302576.0/4294967296.0,1,-nbitq), 
to_sfixed(278557710.0/4294967296.0,1,-nbitq), 
to_sfixed(-97504594.0/4294967296.0,1,-nbitq), 
to_sfixed(151447653.0/4294967296.0,1,-nbitq), 
to_sfixed(318328565.0/4294967296.0,1,-nbitq), 
to_sfixed(-346619154.0/4294967296.0,1,-nbitq), 
to_sfixed(287039666.0/4294967296.0,1,-nbitq), 
to_sfixed(235739724.0/4294967296.0,1,-nbitq), 
to_sfixed(-321059613.0/4294967296.0,1,-nbitq), 
to_sfixed(202849577.0/4294967296.0,1,-nbitq), 
to_sfixed(-95178483.0/4294967296.0,1,-nbitq), 
to_sfixed(-347520357.0/4294967296.0,1,-nbitq), 
to_sfixed(100206471.0/4294967296.0,1,-nbitq), 
to_sfixed(92744684.0/4294967296.0,1,-nbitq), 
to_sfixed(7838359.0/4294967296.0,1,-nbitq), 
to_sfixed(202505382.0/4294967296.0,1,-nbitq), 
to_sfixed(-4153790.0/4294967296.0,1,-nbitq), 
to_sfixed(-108124504.0/4294967296.0,1,-nbitq), 
to_sfixed(120261499.0/4294967296.0,1,-nbitq), 
to_sfixed(-469671763.0/4294967296.0,1,-nbitq), 
to_sfixed(-497889809.0/4294967296.0,1,-nbitq), 
to_sfixed(-93168531.0/4294967296.0,1,-nbitq), 
to_sfixed(-3039424.0/4294967296.0,1,-nbitq), 
to_sfixed(240023530.0/4294967296.0,1,-nbitq), 
to_sfixed(224724834.0/4294967296.0,1,-nbitq), 
to_sfixed(436313577.0/4294967296.0,1,-nbitq), 
to_sfixed(381925355.0/4294967296.0,1,-nbitq), 
to_sfixed(-70621969.0/4294967296.0,1,-nbitq), 
to_sfixed(-242505196.0/4294967296.0,1,-nbitq), 
to_sfixed(-269314347.0/4294967296.0,1,-nbitq), 
to_sfixed(169882793.0/4294967296.0,1,-nbitq), 
to_sfixed(-406653280.0/4294967296.0,1,-nbitq), 
to_sfixed(44750821.0/4294967296.0,1,-nbitq), 
to_sfixed(-210573436.0/4294967296.0,1,-nbitq), 
to_sfixed(312896302.0/4294967296.0,1,-nbitq), 
to_sfixed(261111593.0/4294967296.0,1,-nbitq), 
to_sfixed(387341928.0/4294967296.0,1,-nbitq), 
to_sfixed(312575178.0/4294967296.0,1,-nbitq), 
to_sfixed(193132685.0/4294967296.0,1,-nbitq), 
to_sfixed(-107784732.0/4294967296.0,1,-nbitq), 
to_sfixed(-177209456.0/4294967296.0,1,-nbitq), 
to_sfixed(371244656.0/4294967296.0,1,-nbitq), 
to_sfixed(-150441715.0/4294967296.0,1,-nbitq), 
to_sfixed(-392107106.0/4294967296.0,1,-nbitq), 
to_sfixed(402896614.0/4294967296.0,1,-nbitq), 
to_sfixed(64506551.0/4294967296.0,1,-nbitq), 
to_sfixed(105723902.0/4294967296.0,1,-nbitq), 
to_sfixed(-262164100.0/4294967296.0,1,-nbitq), 
to_sfixed(-260388410.0/4294967296.0,1,-nbitq), 
to_sfixed(66941453.0/4294967296.0,1,-nbitq), 
to_sfixed(-230682051.0/4294967296.0,1,-nbitq), 
to_sfixed(-168641428.0/4294967296.0,1,-nbitq), 
to_sfixed(840655434.0/4294967296.0,1,-nbitq), 
to_sfixed(48859685.0/4294967296.0,1,-nbitq), 
to_sfixed(-300131298.0/4294967296.0,1,-nbitq), 
to_sfixed(198883953.0/4294967296.0,1,-nbitq), 
to_sfixed(-502874666.0/4294967296.0,1,-nbitq), 
to_sfixed(-92063824.0/4294967296.0,1,-nbitq), 
to_sfixed(195624291.0/4294967296.0,1,-nbitq), 
to_sfixed(-57409103.0/4294967296.0,1,-nbitq), 
to_sfixed(-40504387.0/4294967296.0,1,-nbitq), 
to_sfixed(-294726185.0/4294967296.0,1,-nbitq), 
to_sfixed(-398415283.0/4294967296.0,1,-nbitq), 
to_sfixed(-251165278.0/4294967296.0,1,-nbitq), 
to_sfixed(-235603054.0/4294967296.0,1,-nbitq), 
to_sfixed(245977713.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(148154829.0/4294967296.0,1,-nbitq), 
to_sfixed(-352840489.0/4294967296.0,1,-nbitq), 
to_sfixed(29458581.0/4294967296.0,1,-nbitq), 
to_sfixed(226616398.0/4294967296.0,1,-nbitq), 
to_sfixed(-78279113.0/4294967296.0,1,-nbitq), 
to_sfixed(73058682.0/4294967296.0,1,-nbitq), 
to_sfixed(-139849220.0/4294967296.0,1,-nbitq), 
to_sfixed(133398977.0/4294967296.0,1,-nbitq), 
to_sfixed(-205792622.0/4294967296.0,1,-nbitq), 
to_sfixed(109782341.0/4294967296.0,1,-nbitq), 
to_sfixed(459039010.0/4294967296.0,1,-nbitq), 
to_sfixed(74739777.0/4294967296.0,1,-nbitq), 
to_sfixed(174644411.0/4294967296.0,1,-nbitq), 
to_sfixed(-368585690.0/4294967296.0,1,-nbitq), 
to_sfixed(-54739190.0/4294967296.0,1,-nbitq), 
to_sfixed(165151505.0/4294967296.0,1,-nbitq), 
to_sfixed(152935701.0/4294967296.0,1,-nbitq), 
to_sfixed(261073239.0/4294967296.0,1,-nbitq), 
to_sfixed(36512997.0/4294967296.0,1,-nbitq), 
to_sfixed(-291012703.0/4294967296.0,1,-nbitq), 
to_sfixed(44858152.0/4294967296.0,1,-nbitq), 
to_sfixed(147756541.0/4294967296.0,1,-nbitq), 
to_sfixed(172389708.0/4294967296.0,1,-nbitq), 
to_sfixed(-46469391.0/4294967296.0,1,-nbitq), 
to_sfixed(284087483.0/4294967296.0,1,-nbitq), 
to_sfixed(-264324378.0/4294967296.0,1,-nbitq), 
to_sfixed(-93542355.0/4294967296.0,1,-nbitq), 
to_sfixed(-627722246.0/4294967296.0,1,-nbitq), 
to_sfixed(216355131.0/4294967296.0,1,-nbitq), 
to_sfixed(-414319522.0/4294967296.0,1,-nbitq), 
to_sfixed(-380411707.0/4294967296.0,1,-nbitq), 
to_sfixed(228257051.0/4294967296.0,1,-nbitq), 
to_sfixed(207219032.0/4294967296.0,1,-nbitq), 
to_sfixed(-84597807.0/4294967296.0,1,-nbitq), 
to_sfixed(-302580408.0/4294967296.0,1,-nbitq), 
to_sfixed(112662975.0/4294967296.0,1,-nbitq), 
to_sfixed(306059230.0/4294967296.0,1,-nbitq), 
to_sfixed(334146998.0/4294967296.0,1,-nbitq), 
to_sfixed(319566724.0/4294967296.0,1,-nbitq), 
to_sfixed(302633085.0/4294967296.0,1,-nbitq), 
to_sfixed(-41322983.0/4294967296.0,1,-nbitq), 
to_sfixed(-209730629.0/4294967296.0,1,-nbitq), 
to_sfixed(-292938879.0/4294967296.0,1,-nbitq), 
to_sfixed(242564556.0/4294967296.0,1,-nbitq), 
to_sfixed(82099723.0/4294967296.0,1,-nbitq), 
to_sfixed(-233709106.0/4294967296.0,1,-nbitq), 
to_sfixed(234698238.0/4294967296.0,1,-nbitq), 
to_sfixed(-441587009.0/4294967296.0,1,-nbitq), 
to_sfixed(217658326.0/4294967296.0,1,-nbitq), 
to_sfixed(281147465.0/4294967296.0,1,-nbitq), 
to_sfixed(16172479.0/4294967296.0,1,-nbitq), 
to_sfixed(409243624.0/4294967296.0,1,-nbitq), 
to_sfixed(-123909324.0/4294967296.0,1,-nbitq), 
to_sfixed(-189994339.0/4294967296.0,1,-nbitq), 
to_sfixed(257845081.0/4294967296.0,1,-nbitq), 
to_sfixed(-4248593.0/4294967296.0,1,-nbitq), 
to_sfixed(429985691.0/4294967296.0,1,-nbitq), 
to_sfixed(57771254.0/4294967296.0,1,-nbitq), 
to_sfixed(-13944949.0/4294967296.0,1,-nbitq), 
to_sfixed(-351398848.0/4294967296.0,1,-nbitq), 
to_sfixed(25085954.0/4294967296.0,1,-nbitq), 
to_sfixed(103255094.0/4294967296.0,1,-nbitq), 
to_sfixed(-187464916.0/4294967296.0,1,-nbitq), 
to_sfixed(212612641.0/4294967296.0,1,-nbitq), 
to_sfixed(191838302.0/4294967296.0,1,-nbitq), 
to_sfixed(306603546.0/4294967296.0,1,-nbitq), 
to_sfixed(333496290.0/4294967296.0,1,-nbitq), 
to_sfixed(120371202.0/4294967296.0,1,-nbitq), 
to_sfixed(244892429.0/4294967296.0,1,-nbitq), 
to_sfixed(358382819.0/4294967296.0,1,-nbitq), 
to_sfixed(-238834873.0/4294967296.0,1,-nbitq), 
to_sfixed(-239860651.0/4294967296.0,1,-nbitq), 
to_sfixed(323883068.0/4294967296.0,1,-nbitq), 
to_sfixed(182443768.0/4294967296.0,1,-nbitq), 
to_sfixed(126589503.0/4294967296.0,1,-nbitq), 
to_sfixed(112011726.0/4294967296.0,1,-nbitq), 
to_sfixed(247257384.0/4294967296.0,1,-nbitq), 
to_sfixed(-99480803.0/4294967296.0,1,-nbitq), 
to_sfixed(-503671059.0/4294967296.0,1,-nbitq), 
to_sfixed(73002824.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-370059547.0/4294967296.0,1,-nbitq), 
to_sfixed(-24871842.0/4294967296.0,1,-nbitq), 
to_sfixed(-178276423.0/4294967296.0,1,-nbitq), 
to_sfixed(690730506.0/4294967296.0,1,-nbitq), 
to_sfixed(713923471.0/4294967296.0,1,-nbitq), 
to_sfixed(283810084.0/4294967296.0,1,-nbitq), 
to_sfixed(-260048535.0/4294967296.0,1,-nbitq), 
to_sfixed(-481896471.0/4294967296.0,1,-nbitq), 
to_sfixed(49546837.0/4294967296.0,1,-nbitq), 
to_sfixed(-137438171.0/4294967296.0,1,-nbitq), 
to_sfixed(-450990245.0/4294967296.0,1,-nbitq), 
to_sfixed(95907357.0/4294967296.0,1,-nbitq), 
to_sfixed(-582225286.0/4294967296.0,1,-nbitq), 
to_sfixed(1247225.0/4294967296.0,1,-nbitq), 
to_sfixed(-66249866.0/4294967296.0,1,-nbitq), 
to_sfixed(228814147.0/4294967296.0,1,-nbitq), 
to_sfixed(-202321696.0/4294967296.0,1,-nbitq), 
to_sfixed(250317884.0/4294967296.0,1,-nbitq), 
to_sfixed(144058376.0/4294967296.0,1,-nbitq), 
to_sfixed(-98631492.0/4294967296.0,1,-nbitq), 
to_sfixed(379421348.0/4294967296.0,1,-nbitq), 
to_sfixed(-722349.0/4294967296.0,1,-nbitq), 
to_sfixed(-111699767.0/4294967296.0,1,-nbitq), 
to_sfixed(340030039.0/4294967296.0,1,-nbitq), 
to_sfixed(-331800743.0/4294967296.0,1,-nbitq), 
to_sfixed(-71686252.0/4294967296.0,1,-nbitq), 
to_sfixed(360646230.0/4294967296.0,1,-nbitq), 
to_sfixed(-561988870.0/4294967296.0,1,-nbitq), 
to_sfixed(189414350.0/4294967296.0,1,-nbitq), 
to_sfixed(205535680.0/4294967296.0,1,-nbitq), 
to_sfixed(-650976331.0/4294967296.0,1,-nbitq), 
to_sfixed(-625126974.0/4294967296.0,1,-nbitq), 
to_sfixed(467409305.0/4294967296.0,1,-nbitq), 
to_sfixed(12998823.0/4294967296.0,1,-nbitq), 
to_sfixed(39348297.0/4294967296.0,1,-nbitq), 
to_sfixed(-499838553.0/4294967296.0,1,-nbitq), 
to_sfixed(-317618370.0/4294967296.0,1,-nbitq), 
to_sfixed(261901370.0/4294967296.0,1,-nbitq), 
to_sfixed(281256412.0/4294967296.0,1,-nbitq), 
to_sfixed(206180523.0/4294967296.0,1,-nbitq), 
to_sfixed(16827637.0/4294967296.0,1,-nbitq), 
to_sfixed(337003758.0/4294967296.0,1,-nbitq), 
to_sfixed(688998803.0/4294967296.0,1,-nbitq), 
to_sfixed(71206259.0/4294967296.0,1,-nbitq), 
to_sfixed(4921222.0/4294967296.0,1,-nbitq), 
to_sfixed(106888826.0/4294967296.0,1,-nbitq), 
to_sfixed(232911692.0/4294967296.0,1,-nbitq), 
to_sfixed(-509797104.0/4294967296.0,1,-nbitq), 
to_sfixed(-63290920.0/4294967296.0,1,-nbitq), 
to_sfixed(-10344857.0/4294967296.0,1,-nbitq), 
to_sfixed(418262760.0/4294967296.0,1,-nbitq), 
to_sfixed(495727745.0/4294967296.0,1,-nbitq), 
to_sfixed(-392965742.0/4294967296.0,1,-nbitq), 
to_sfixed(653223695.0/4294967296.0,1,-nbitq), 
to_sfixed(195765399.0/4294967296.0,1,-nbitq), 
to_sfixed(178608878.0/4294967296.0,1,-nbitq), 
to_sfixed(-84639055.0/4294967296.0,1,-nbitq), 
to_sfixed(-403452339.0/4294967296.0,1,-nbitq), 
to_sfixed(271284182.0/4294967296.0,1,-nbitq), 
to_sfixed(-81497710.0/4294967296.0,1,-nbitq), 
to_sfixed(-528690.0/4294967296.0,1,-nbitq), 
to_sfixed(519908121.0/4294967296.0,1,-nbitq), 
to_sfixed(314458366.0/4294967296.0,1,-nbitq), 
to_sfixed(236032581.0/4294967296.0,1,-nbitq), 
to_sfixed(219802166.0/4294967296.0,1,-nbitq), 
to_sfixed(-387420007.0/4294967296.0,1,-nbitq), 
to_sfixed(313265241.0/4294967296.0,1,-nbitq), 
to_sfixed(231007301.0/4294967296.0,1,-nbitq), 
to_sfixed(386860497.0/4294967296.0,1,-nbitq), 
to_sfixed(263611419.0/4294967296.0,1,-nbitq), 
to_sfixed(-321159773.0/4294967296.0,1,-nbitq), 
to_sfixed(373850664.0/4294967296.0,1,-nbitq), 
to_sfixed(-292038091.0/4294967296.0,1,-nbitq), 
to_sfixed(283704582.0/4294967296.0,1,-nbitq), 
to_sfixed(-155442860.0/4294967296.0,1,-nbitq), 
to_sfixed(60343586.0/4294967296.0,1,-nbitq), 
to_sfixed(-67513011.0/4294967296.0,1,-nbitq), 
to_sfixed(42023154.0/4294967296.0,1,-nbitq), 
to_sfixed(120197736.0/4294967296.0,1,-nbitq), 
to_sfixed(175231147.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(29765318.0/4294967296.0,1,-nbitq), 
to_sfixed(-409200457.0/4294967296.0,1,-nbitq), 
to_sfixed(-133776033.0/4294967296.0,1,-nbitq), 
to_sfixed(267241382.0/4294967296.0,1,-nbitq), 
to_sfixed(759959905.0/4294967296.0,1,-nbitq), 
to_sfixed(-254880853.0/4294967296.0,1,-nbitq), 
to_sfixed(170871968.0/4294967296.0,1,-nbitq), 
to_sfixed(39662299.0/4294967296.0,1,-nbitq), 
to_sfixed(227079458.0/4294967296.0,1,-nbitq), 
to_sfixed(-245014773.0/4294967296.0,1,-nbitq), 
to_sfixed(-31121717.0/4294967296.0,1,-nbitq), 
to_sfixed(272818816.0/4294967296.0,1,-nbitq), 
to_sfixed(-191659248.0/4294967296.0,1,-nbitq), 
to_sfixed(109439518.0/4294967296.0,1,-nbitq), 
to_sfixed(-19128792.0/4294967296.0,1,-nbitq), 
to_sfixed(115929095.0/4294967296.0,1,-nbitq), 
to_sfixed(-364936016.0/4294967296.0,1,-nbitq), 
to_sfixed(-5858296.0/4294967296.0,1,-nbitq), 
to_sfixed(-207850468.0/4294967296.0,1,-nbitq), 
to_sfixed(155272089.0/4294967296.0,1,-nbitq), 
to_sfixed(-349640938.0/4294967296.0,1,-nbitq), 
to_sfixed(-23211471.0/4294967296.0,1,-nbitq), 
to_sfixed(346236608.0/4294967296.0,1,-nbitq), 
to_sfixed(108075307.0/4294967296.0,1,-nbitq), 
to_sfixed(26533684.0/4294967296.0,1,-nbitq), 
to_sfixed(279931285.0/4294967296.0,1,-nbitq), 
to_sfixed(46970645.0/4294967296.0,1,-nbitq), 
to_sfixed(-451863613.0/4294967296.0,1,-nbitq), 
to_sfixed(500981992.0/4294967296.0,1,-nbitq), 
to_sfixed(-56001991.0/4294967296.0,1,-nbitq), 
to_sfixed(90769621.0/4294967296.0,1,-nbitq), 
to_sfixed(-103019666.0/4294967296.0,1,-nbitq), 
to_sfixed(87652435.0/4294967296.0,1,-nbitq), 
to_sfixed(-381984886.0/4294967296.0,1,-nbitq), 
to_sfixed(-29173131.0/4294967296.0,1,-nbitq), 
to_sfixed(-666398052.0/4294967296.0,1,-nbitq), 
to_sfixed(-58043650.0/4294967296.0,1,-nbitq), 
to_sfixed(468806989.0/4294967296.0,1,-nbitq), 
to_sfixed(-273330334.0/4294967296.0,1,-nbitq), 
to_sfixed(33352568.0/4294967296.0,1,-nbitq), 
to_sfixed(244927264.0/4294967296.0,1,-nbitq), 
to_sfixed(-11935313.0/4294967296.0,1,-nbitq), 
to_sfixed(-98074895.0/4294967296.0,1,-nbitq), 
to_sfixed(534980554.0/4294967296.0,1,-nbitq), 
to_sfixed(248781095.0/4294967296.0,1,-nbitq), 
to_sfixed(361132978.0/4294967296.0,1,-nbitq), 
to_sfixed(-338542984.0/4294967296.0,1,-nbitq), 
to_sfixed(-18359522.0/4294967296.0,1,-nbitq), 
to_sfixed(-111577993.0/4294967296.0,1,-nbitq), 
to_sfixed(-323690324.0/4294967296.0,1,-nbitq), 
to_sfixed(-82582013.0/4294967296.0,1,-nbitq), 
to_sfixed(295894753.0/4294967296.0,1,-nbitq), 
to_sfixed(-278341547.0/4294967296.0,1,-nbitq), 
to_sfixed(505254610.0/4294967296.0,1,-nbitq), 
to_sfixed(516908148.0/4294967296.0,1,-nbitq), 
to_sfixed(-264462912.0/4294967296.0,1,-nbitq), 
to_sfixed(-135367397.0/4294967296.0,1,-nbitq), 
to_sfixed(-286717885.0/4294967296.0,1,-nbitq), 
to_sfixed(383486731.0/4294967296.0,1,-nbitq), 
to_sfixed(-99692142.0/4294967296.0,1,-nbitq), 
to_sfixed(-413853071.0/4294967296.0,1,-nbitq), 
to_sfixed(683517099.0/4294967296.0,1,-nbitq), 
to_sfixed(-33041458.0/4294967296.0,1,-nbitq), 
to_sfixed(440589874.0/4294967296.0,1,-nbitq), 
to_sfixed(-101098809.0/4294967296.0,1,-nbitq), 
to_sfixed(-92886544.0/4294967296.0,1,-nbitq), 
to_sfixed(262840104.0/4294967296.0,1,-nbitq), 
to_sfixed(257491123.0/4294967296.0,1,-nbitq), 
to_sfixed(380235076.0/4294967296.0,1,-nbitq), 
to_sfixed(219470147.0/4294967296.0,1,-nbitq), 
to_sfixed(-122062363.0/4294967296.0,1,-nbitq), 
to_sfixed(-295203820.0/4294967296.0,1,-nbitq), 
to_sfixed(-125463216.0/4294967296.0,1,-nbitq), 
to_sfixed(269777933.0/4294967296.0,1,-nbitq), 
to_sfixed(-132895269.0/4294967296.0,1,-nbitq), 
to_sfixed(223782132.0/4294967296.0,1,-nbitq), 
to_sfixed(-139389780.0/4294967296.0,1,-nbitq), 
to_sfixed(303925280.0/4294967296.0,1,-nbitq), 
to_sfixed(43764657.0/4294967296.0,1,-nbitq), 
to_sfixed(-63284711.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(204348990.0/4294967296.0,1,-nbitq), 
to_sfixed(-436629953.0/4294967296.0,1,-nbitq), 
to_sfixed(-1333665.0/4294967296.0,1,-nbitq), 
to_sfixed(109138235.0/4294967296.0,1,-nbitq), 
to_sfixed(204519822.0/4294967296.0,1,-nbitq), 
to_sfixed(-1571767.0/4294967296.0,1,-nbitq), 
to_sfixed(186735483.0/4294967296.0,1,-nbitq), 
to_sfixed(-257432585.0/4294967296.0,1,-nbitq), 
to_sfixed(-303407001.0/4294967296.0,1,-nbitq), 
to_sfixed(-257265452.0/4294967296.0,1,-nbitq), 
to_sfixed(-319300398.0/4294967296.0,1,-nbitq), 
to_sfixed(-352136587.0/4294967296.0,1,-nbitq), 
to_sfixed(623505160.0/4294967296.0,1,-nbitq), 
to_sfixed(719437556.0/4294967296.0,1,-nbitq), 
to_sfixed(132766058.0/4294967296.0,1,-nbitq), 
to_sfixed(245858939.0/4294967296.0,1,-nbitq), 
to_sfixed(77201925.0/4294967296.0,1,-nbitq), 
to_sfixed(-201923841.0/4294967296.0,1,-nbitq), 
to_sfixed(195552174.0/4294967296.0,1,-nbitq), 
to_sfixed(443615674.0/4294967296.0,1,-nbitq), 
to_sfixed(-244243058.0/4294967296.0,1,-nbitq), 
to_sfixed(63440154.0/4294967296.0,1,-nbitq), 
to_sfixed(-212047392.0/4294967296.0,1,-nbitq), 
to_sfixed(118241372.0/4294967296.0,1,-nbitq), 
to_sfixed(-148201130.0/4294967296.0,1,-nbitq), 
to_sfixed(531540114.0/4294967296.0,1,-nbitq), 
to_sfixed(-279109555.0/4294967296.0,1,-nbitq), 
to_sfixed(74014336.0/4294967296.0,1,-nbitq), 
to_sfixed(23318632.0/4294967296.0,1,-nbitq), 
to_sfixed(38987550.0/4294967296.0,1,-nbitq), 
to_sfixed(262661965.0/4294967296.0,1,-nbitq), 
to_sfixed(259415963.0/4294967296.0,1,-nbitq), 
to_sfixed(-164389291.0/4294967296.0,1,-nbitq), 
to_sfixed(44812749.0/4294967296.0,1,-nbitq), 
to_sfixed(-155523748.0/4294967296.0,1,-nbitq), 
to_sfixed(126693125.0/4294967296.0,1,-nbitq), 
to_sfixed(-366178076.0/4294967296.0,1,-nbitq), 
to_sfixed(-154630554.0/4294967296.0,1,-nbitq), 
to_sfixed(33450957.0/4294967296.0,1,-nbitq), 
to_sfixed(173074431.0/4294967296.0,1,-nbitq), 
to_sfixed(-370332108.0/4294967296.0,1,-nbitq), 
to_sfixed(249402404.0/4294967296.0,1,-nbitq), 
to_sfixed(300841319.0/4294967296.0,1,-nbitq), 
to_sfixed(-21585140.0/4294967296.0,1,-nbitq), 
to_sfixed(-352011003.0/4294967296.0,1,-nbitq), 
to_sfixed(386494819.0/4294967296.0,1,-nbitq), 
to_sfixed(58037767.0/4294967296.0,1,-nbitq), 
to_sfixed(-377760980.0/4294967296.0,1,-nbitq), 
to_sfixed(-110520308.0/4294967296.0,1,-nbitq), 
to_sfixed(-492242668.0/4294967296.0,1,-nbitq), 
to_sfixed(40821276.0/4294967296.0,1,-nbitq), 
to_sfixed(298703114.0/4294967296.0,1,-nbitq), 
to_sfixed(-42732751.0/4294967296.0,1,-nbitq), 
to_sfixed(610607455.0/4294967296.0,1,-nbitq), 
to_sfixed(261859016.0/4294967296.0,1,-nbitq), 
to_sfixed(208457300.0/4294967296.0,1,-nbitq), 
to_sfixed(85079921.0/4294967296.0,1,-nbitq), 
to_sfixed(-203052875.0/4294967296.0,1,-nbitq), 
to_sfixed(304601173.0/4294967296.0,1,-nbitq), 
to_sfixed(63608521.0/4294967296.0,1,-nbitq), 
to_sfixed(-176381125.0/4294967296.0,1,-nbitq), 
to_sfixed(479329270.0/4294967296.0,1,-nbitq), 
to_sfixed(52840800.0/4294967296.0,1,-nbitq), 
to_sfixed(142119897.0/4294967296.0,1,-nbitq), 
to_sfixed(-147328574.0/4294967296.0,1,-nbitq), 
to_sfixed(254240679.0/4294967296.0,1,-nbitq), 
to_sfixed(308424470.0/4294967296.0,1,-nbitq), 
to_sfixed(-58419160.0/4294967296.0,1,-nbitq), 
to_sfixed(441894166.0/4294967296.0,1,-nbitq), 
to_sfixed(187830963.0/4294967296.0,1,-nbitq), 
to_sfixed(498698516.0/4294967296.0,1,-nbitq), 
to_sfixed(-347351841.0/4294967296.0,1,-nbitq), 
to_sfixed(-451465899.0/4294967296.0,1,-nbitq), 
to_sfixed(371629395.0/4294967296.0,1,-nbitq), 
to_sfixed(289207806.0/4294967296.0,1,-nbitq), 
to_sfixed(157416101.0/4294967296.0,1,-nbitq), 
to_sfixed(-271807819.0/4294967296.0,1,-nbitq), 
to_sfixed(-54982847.0/4294967296.0,1,-nbitq), 
to_sfixed(164894458.0/4294967296.0,1,-nbitq), 
to_sfixed(152724247.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-213875606.0/4294967296.0,1,-nbitq), 
to_sfixed(174484972.0/4294967296.0,1,-nbitq), 
to_sfixed(797764943.0/4294967296.0,1,-nbitq), 
to_sfixed(-345932946.0/4294967296.0,1,-nbitq), 
to_sfixed(67474616.0/4294967296.0,1,-nbitq), 
to_sfixed(-298789226.0/4294967296.0,1,-nbitq), 
to_sfixed(-193063711.0/4294967296.0,1,-nbitq), 
to_sfixed(-606653602.0/4294967296.0,1,-nbitq), 
to_sfixed(-1078557835.0/4294967296.0,1,-nbitq), 
to_sfixed(304682392.0/4294967296.0,1,-nbitq), 
to_sfixed(55284124.0/4294967296.0,1,-nbitq), 
to_sfixed(-101410311.0/4294967296.0,1,-nbitq), 
to_sfixed(465812564.0/4294967296.0,1,-nbitq), 
to_sfixed(1034384614.0/4294967296.0,1,-nbitq), 
to_sfixed(392227147.0/4294967296.0,1,-nbitq), 
to_sfixed(55675223.0/4294967296.0,1,-nbitq), 
to_sfixed(-158577616.0/4294967296.0,1,-nbitq), 
to_sfixed(-117898608.0/4294967296.0,1,-nbitq), 
to_sfixed(-453898846.0/4294967296.0,1,-nbitq), 
to_sfixed(312224481.0/4294967296.0,1,-nbitq), 
to_sfixed(-278539739.0/4294967296.0,1,-nbitq), 
to_sfixed(-529281276.0/4294967296.0,1,-nbitq), 
to_sfixed(-425508877.0/4294967296.0,1,-nbitq), 
to_sfixed(642046045.0/4294967296.0,1,-nbitq), 
to_sfixed(161745385.0/4294967296.0,1,-nbitq), 
to_sfixed(822740208.0/4294967296.0,1,-nbitq), 
to_sfixed(180748094.0/4294967296.0,1,-nbitq), 
to_sfixed(-274393158.0/4294967296.0,1,-nbitq), 
to_sfixed(83353317.0/4294967296.0,1,-nbitq), 
to_sfixed(362580084.0/4294967296.0,1,-nbitq), 
to_sfixed(-171197565.0/4294967296.0,1,-nbitq), 
to_sfixed(-154172846.0/4294967296.0,1,-nbitq), 
to_sfixed(-287633071.0/4294967296.0,1,-nbitq), 
to_sfixed(-349450332.0/4294967296.0,1,-nbitq), 
to_sfixed(238227216.0/4294967296.0,1,-nbitq), 
to_sfixed(-218479730.0/4294967296.0,1,-nbitq), 
to_sfixed(-250478790.0/4294967296.0,1,-nbitq), 
to_sfixed(39323916.0/4294967296.0,1,-nbitq), 
to_sfixed(-274008987.0/4294967296.0,1,-nbitq), 
to_sfixed(8783441.0/4294967296.0,1,-nbitq), 
to_sfixed(-141528088.0/4294967296.0,1,-nbitq), 
to_sfixed(-224410833.0/4294967296.0,1,-nbitq), 
to_sfixed(77022360.0/4294967296.0,1,-nbitq), 
to_sfixed(177923836.0/4294967296.0,1,-nbitq), 
to_sfixed(25983952.0/4294967296.0,1,-nbitq), 
to_sfixed(174474498.0/4294967296.0,1,-nbitq), 
to_sfixed(188550255.0/4294967296.0,1,-nbitq), 
to_sfixed(-231682232.0/4294967296.0,1,-nbitq), 
to_sfixed(-55934643.0/4294967296.0,1,-nbitq), 
to_sfixed(-215079447.0/4294967296.0,1,-nbitq), 
to_sfixed(-182494588.0/4294967296.0,1,-nbitq), 
to_sfixed(-36976420.0/4294967296.0,1,-nbitq), 
to_sfixed(-206775437.0/4294967296.0,1,-nbitq), 
to_sfixed(235355902.0/4294967296.0,1,-nbitq), 
to_sfixed(752316326.0/4294967296.0,1,-nbitq), 
to_sfixed(-639896496.0/4294967296.0,1,-nbitq), 
to_sfixed(56209997.0/4294967296.0,1,-nbitq), 
to_sfixed(-476823134.0/4294967296.0,1,-nbitq), 
to_sfixed(188252389.0/4294967296.0,1,-nbitq), 
to_sfixed(337008071.0/4294967296.0,1,-nbitq), 
to_sfixed(291757377.0/4294967296.0,1,-nbitq), 
to_sfixed(473579805.0/4294967296.0,1,-nbitq), 
to_sfixed(36307143.0/4294967296.0,1,-nbitq), 
to_sfixed(780350738.0/4294967296.0,1,-nbitq), 
to_sfixed(108565349.0/4294967296.0,1,-nbitq), 
to_sfixed(-365276380.0/4294967296.0,1,-nbitq), 
to_sfixed(124054187.0/4294967296.0,1,-nbitq), 
to_sfixed(427338491.0/4294967296.0,1,-nbitq), 
to_sfixed(-111667436.0/4294967296.0,1,-nbitq), 
to_sfixed(-269111877.0/4294967296.0,1,-nbitq), 
to_sfixed(477785384.0/4294967296.0,1,-nbitq), 
to_sfixed(311896301.0/4294967296.0,1,-nbitq), 
to_sfixed(-447865009.0/4294967296.0,1,-nbitq), 
to_sfixed(-348760734.0/4294967296.0,1,-nbitq), 
to_sfixed(-205686783.0/4294967296.0,1,-nbitq), 
to_sfixed(586371844.0/4294967296.0,1,-nbitq), 
to_sfixed(-362468685.0/4294967296.0,1,-nbitq), 
to_sfixed(121000150.0/4294967296.0,1,-nbitq), 
to_sfixed(-255843050.0/4294967296.0,1,-nbitq), 
to_sfixed(102995114.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(305399766.0/4294967296.0,1,-nbitq), 
to_sfixed(29456424.0/4294967296.0,1,-nbitq), 
to_sfixed(1198034828.0/4294967296.0,1,-nbitq), 
to_sfixed(-998286581.0/4294967296.0,1,-nbitq), 
to_sfixed(-90621219.0/4294967296.0,1,-nbitq), 
to_sfixed(-255545773.0/4294967296.0,1,-nbitq), 
to_sfixed(-84469474.0/4294967296.0,1,-nbitq), 
to_sfixed(85396544.0/4294967296.0,1,-nbitq), 
to_sfixed(-986680236.0/4294967296.0,1,-nbitq), 
to_sfixed(336460612.0/4294967296.0,1,-nbitq), 
to_sfixed(-407770419.0/4294967296.0,1,-nbitq), 
to_sfixed(-260588926.0/4294967296.0,1,-nbitq), 
to_sfixed(987484476.0/4294967296.0,1,-nbitq), 
to_sfixed(1309123233.0/4294967296.0,1,-nbitq), 
to_sfixed(-67803661.0/4294967296.0,1,-nbitq), 
to_sfixed(-45857239.0/4294967296.0,1,-nbitq), 
to_sfixed(-203231706.0/4294967296.0,1,-nbitq), 
to_sfixed(-298595556.0/4294967296.0,1,-nbitq), 
to_sfixed(-519994087.0/4294967296.0,1,-nbitq), 
to_sfixed(627039257.0/4294967296.0,1,-nbitq), 
to_sfixed(80595388.0/4294967296.0,1,-nbitq), 
to_sfixed(-146989456.0/4294967296.0,1,-nbitq), 
to_sfixed(-10282566.0/4294967296.0,1,-nbitq), 
to_sfixed(695188177.0/4294967296.0,1,-nbitq), 
to_sfixed(388745871.0/4294967296.0,1,-nbitq), 
to_sfixed(376858201.0/4294967296.0,1,-nbitq), 
to_sfixed(-433278106.0/4294967296.0,1,-nbitq), 
to_sfixed(111533258.0/4294967296.0,1,-nbitq), 
to_sfixed(255563541.0/4294967296.0,1,-nbitq), 
to_sfixed(106866578.0/4294967296.0,1,-nbitq), 
to_sfixed(212109176.0/4294967296.0,1,-nbitq), 
to_sfixed(-102929309.0/4294967296.0,1,-nbitq), 
to_sfixed(-578853361.0/4294967296.0,1,-nbitq), 
to_sfixed(56000835.0/4294967296.0,1,-nbitq), 
to_sfixed(-174737957.0/4294967296.0,1,-nbitq), 
to_sfixed(184351088.0/4294967296.0,1,-nbitq), 
to_sfixed(-53662126.0/4294967296.0,1,-nbitq), 
to_sfixed(-474346502.0/4294967296.0,1,-nbitq), 
to_sfixed(-57115058.0/4294967296.0,1,-nbitq), 
to_sfixed(-110261970.0/4294967296.0,1,-nbitq), 
to_sfixed(-261255097.0/4294967296.0,1,-nbitq), 
to_sfixed(9008902.0/4294967296.0,1,-nbitq), 
to_sfixed(-421983159.0/4294967296.0,1,-nbitq), 
to_sfixed(512914183.0/4294967296.0,1,-nbitq), 
to_sfixed(88434660.0/4294967296.0,1,-nbitq), 
to_sfixed(-127381469.0/4294967296.0,1,-nbitq), 
to_sfixed(-305635951.0/4294967296.0,1,-nbitq), 
to_sfixed(-144786355.0/4294967296.0,1,-nbitq), 
to_sfixed(-169317213.0/4294967296.0,1,-nbitq), 
to_sfixed(-197369130.0/4294967296.0,1,-nbitq), 
to_sfixed(65492225.0/4294967296.0,1,-nbitq), 
to_sfixed(-247801293.0/4294967296.0,1,-nbitq), 
to_sfixed(265294974.0/4294967296.0,1,-nbitq), 
to_sfixed(-559756948.0/4294967296.0,1,-nbitq), 
to_sfixed(399448273.0/4294967296.0,1,-nbitq), 
to_sfixed(61864923.0/4294967296.0,1,-nbitq), 
to_sfixed(396809383.0/4294967296.0,1,-nbitq), 
to_sfixed(-820127371.0/4294967296.0,1,-nbitq), 
to_sfixed(41178264.0/4294967296.0,1,-nbitq), 
to_sfixed(-172659314.0/4294967296.0,1,-nbitq), 
to_sfixed(-168616427.0/4294967296.0,1,-nbitq), 
to_sfixed(-139722198.0/4294967296.0,1,-nbitq), 
to_sfixed(-289657984.0/4294967296.0,1,-nbitq), 
to_sfixed(-33121133.0/4294967296.0,1,-nbitq), 
to_sfixed(-308771827.0/4294967296.0,1,-nbitq), 
to_sfixed(-106244670.0/4294967296.0,1,-nbitq), 
to_sfixed(190698726.0/4294967296.0,1,-nbitq), 
to_sfixed(888224007.0/4294967296.0,1,-nbitq), 
to_sfixed(130774833.0/4294967296.0,1,-nbitq), 
to_sfixed(-571228421.0/4294967296.0,1,-nbitq), 
to_sfixed(300627015.0/4294967296.0,1,-nbitq), 
to_sfixed(14140409.0/4294967296.0,1,-nbitq), 
to_sfixed(-312966580.0/4294967296.0,1,-nbitq), 
to_sfixed(14393235.0/4294967296.0,1,-nbitq), 
to_sfixed(85503241.0/4294967296.0,1,-nbitq), 
to_sfixed(670564984.0/4294967296.0,1,-nbitq), 
to_sfixed(321777896.0/4294967296.0,1,-nbitq), 
to_sfixed(-484687410.0/4294967296.0,1,-nbitq), 
to_sfixed(720913202.0/4294967296.0,1,-nbitq), 
to_sfixed(342797649.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(131325052.0/4294967296.0,1,-nbitq), 
to_sfixed(-469362763.0/4294967296.0,1,-nbitq), 
to_sfixed(272234432.0/4294967296.0,1,-nbitq), 
to_sfixed(-918578552.0/4294967296.0,1,-nbitq), 
to_sfixed(-479242715.0/4294967296.0,1,-nbitq), 
to_sfixed(-9610466.0/4294967296.0,1,-nbitq), 
to_sfixed(397287539.0/4294967296.0,1,-nbitq), 
to_sfixed(116884228.0/4294967296.0,1,-nbitq), 
to_sfixed(-917289548.0/4294967296.0,1,-nbitq), 
to_sfixed(-166738559.0/4294967296.0,1,-nbitq), 
to_sfixed(265494257.0/4294967296.0,1,-nbitq), 
to_sfixed(9095553.0/4294967296.0,1,-nbitq), 
to_sfixed(1560591868.0/4294967296.0,1,-nbitq), 
to_sfixed(1216765942.0/4294967296.0,1,-nbitq), 
to_sfixed(307935825.0/4294967296.0,1,-nbitq), 
to_sfixed(524437680.0/4294967296.0,1,-nbitq), 
to_sfixed(98833277.0/4294967296.0,1,-nbitq), 
to_sfixed(115545852.0/4294967296.0,1,-nbitq), 
to_sfixed(-940043307.0/4294967296.0,1,-nbitq), 
to_sfixed(369801043.0/4294967296.0,1,-nbitq), 
to_sfixed(210481506.0/4294967296.0,1,-nbitq), 
to_sfixed(-50100754.0/4294967296.0,1,-nbitq), 
to_sfixed(-42628490.0/4294967296.0,1,-nbitq), 
to_sfixed(1108344854.0/4294967296.0,1,-nbitq), 
to_sfixed(407452058.0/4294967296.0,1,-nbitq), 
to_sfixed(921166705.0/4294967296.0,1,-nbitq), 
to_sfixed(-412471825.0/4294967296.0,1,-nbitq), 
to_sfixed(-166016447.0/4294967296.0,1,-nbitq), 
to_sfixed(249243941.0/4294967296.0,1,-nbitq), 
to_sfixed(592859891.0/4294967296.0,1,-nbitq), 
to_sfixed(-451188478.0/4294967296.0,1,-nbitq), 
to_sfixed(938832850.0/4294967296.0,1,-nbitq), 
to_sfixed(-422559021.0/4294967296.0,1,-nbitq), 
to_sfixed(124128769.0/4294967296.0,1,-nbitq), 
to_sfixed(-290729875.0/4294967296.0,1,-nbitq), 
to_sfixed(745185987.0/4294967296.0,1,-nbitq), 
to_sfixed(12070623.0/4294967296.0,1,-nbitq), 
to_sfixed(-1372309603.0/4294967296.0,1,-nbitq), 
to_sfixed(-32412811.0/4294967296.0,1,-nbitq), 
to_sfixed(529982099.0/4294967296.0,1,-nbitq), 
to_sfixed(18963390.0/4294967296.0,1,-nbitq), 
to_sfixed(-149296304.0/4294967296.0,1,-nbitq), 
to_sfixed(-215291502.0/4294967296.0,1,-nbitq), 
to_sfixed(48697986.0/4294967296.0,1,-nbitq), 
to_sfixed(-337727789.0/4294967296.0,1,-nbitq), 
to_sfixed(391525107.0/4294967296.0,1,-nbitq), 
to_sfixed(-25189318.0/4294967296.0,1,-nbitq), 
to_sfixed(258612715.0/4294967296.0,1,-nbitq), 
to_sfixed(178162732.0/4294967296.0,1,-nbitq), 
to_sfixed(-83621371.0/4294967296.0,1,-nbitq), 
to_sfixed(-1040396.0/4294967296.0,1,-nbitq), 
to_sfixed(-716219513.0/4294967296.0,1,-nbitq), 
to_sfixed(1091089404.0/4294967296.0,1,-nbitq), 
to_sfixed(-640950973.0/4294967296.0,1,-nbitq), 
to_sfixed(37451298.0/4294967296.0,1,-nbitq), 
to_sfixed(-298707721.0/4294967296.0,1,-nbitq), 
to_sfixed(107264167.0/4294967296.0,1,-nbitq), 
to_sfixed(-272084427.0/4294967296.0,1,-nbitq), 
to_sfixed(-340171113.0/4294967296.0,1,-nbitq), 
to_sfixed(356306106.0/4294967296.0,1,-nbitq), 
to_sfixed(201020521.0/4294967296.0,1,-nbitq), 
to_sfixed(-574627572.0/4294967296.0,1,-nbitq), 
to_sfixed(-509570822.0/4294967296.0,1,-nbitq), 
to_sfixed(-107069404.0/4294967296.0,1,-nbitq), 
to_sfixed(78807550.0/4294967296.0,1,-nbitq), 
to_sfixed(220175484.0/4294967296.0,1,-nbitq), 
to_sfixed(275384396.0/4294967296.0,1,-nbitq), 
to_sfixed(672349971.0/4294967296.0,1,-nbitq), 
to_sfixed(286098316.0/4294967296.0,1,-nbitq), 
to_sfixed(-312897508.0/4294967296.0,1,-nbitq), 
to_sfixed(691195995.0/4294967296.0,1,-nbitq), 
to_sfixed(63040713.0/4294967296.0,1,-nbitq), 
to_sfixed(195540432.0/4294967296.0,1,-nbitq), 
to_sfixed(-15164172.0/4294967296.0,1,-nbitq), 
to_sfixed(-231322726.0/4294967296.0,1,-nbitq), 
to_sfixed(911828787.0/4294967296.0,1,-nbitq), 
to_sfixed(400364725.0/4294967296.0,1,-nbitq), 
to_sfixed(-489301450.0/4294967296.0,1,-nbitq), 
to_sfixed(772903275.0/4294967296.0,1,-nbitq), 
to_sfixed(-106428862.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(457598091.0/4294967296.0,1,-nbitq), 
to_sfixed(73499954.0/4294967296.0,1,-nbitq), 
to_sfixed(-368773849.0/4294967296.0,1,-nbitq), 
to_sfixed(-865247791.0/4294967296.0,1,-nbitq), 
to_sfixed(-440518947.0/4294967296.0,1,-nbitq), 
to_sfixed(871938334.0/4294967296.0,1,-nbitq), 
to_sfixed(-36713434.0/4294967296.0,1,-nbitq), 
to_sfixed(-288286452.0/4294967296.0,1,-nbitq), 
to_sfixed(-842103945.0/4294967296.0,1,-nbitq), 
to_sfixed(-233051751.0/4294967296.0,1,-nbitq), 
to_sfixed(165462141.0/4294967296.0,1,-nbitq), 
to_sfixed(-63896321.0/4294967296.0,1,-nbitq), 
to_sfixed(1867714215.0/4294967296.0,1,-nbitq), 
to_sfixed(1249333268.0/4294967296.0,1,-nbitq), 
to_sfixed(-192944320.0/4294967296.0,1,-nbitq), 
to_sfixed(-87269546.0/4294967296.0,1,-nbitq), 
to_sfixed(150729834.0/4294967296.0,1,-nbitq), 
to_sfixed(483659731.0/4294967296.0,1,-nbitq), 
to_sfixed(-986938736.0/4294967296.0,1,-nbitq), 
to_sfixed(502504087.0/4294967296.0,1,-nbitq), 
to_sfixed(-198609671.0/4294967296.0,1,-nbitq), 
to_sfixed(-1128322707.0/4294967296.0,1,-nbitq), 
to_sfixed(-675173844.0/4294967296.0,1,-nbitq), 
to_sfixed(207824358.0/4294967296.0,1,-nbitq), 
to_sfixed(-155505340.0/4294967296.0,1,-nbitq), 
to_sfixed(838022541.0/4294967296.0,1,-nbitq), 
to_sfixed(-121540939.0/4294967296.0,1,-nbitq), 
to_sfixed(32660243.0/4294967296.0,1,-nbitq), 
to_sfixed(859073121.0/4294967296.0,1,-nbitq), 
to_sfixed(281006091.0/4294967296.0,1,-nbitq), 
to_sfixed(-8942991.0/4294967296.0,1,-nbitq), 
to_sfixed(694827666.0/4294967296.0,1,-nbitq), 
to_sfixed(7855511.0/4294967296.0,1,-nbitq), 
to_sfixed(978552204.0/4294967296.0,1,-nbitq), 
to_sfixed(-8341337.0/4294967296.0,1,-nbitq), 
to_sfixed(172132587.0/4294967296.0,1,-nbitq), 
to_sfixed(-678551346.0/4294967296.0,1,-nbitq), 
to_sfixed(-1144286399.0/4294967296.0,1,-nbitq), 
to_sfixed(109754603.0/4294967296.0,1,-nbitq), 
to_sfixed(-380991311.0/4294967296.0,1,-nbitq), 
to_sfixed(338462066.0/4294967296.0,1,-nbitq), 
to_sfixed(-752737574.0/4294967296.0,1,-nbitq), 
to_sfixed(222196597.0/4294967296.0,1,-nbitq), 
to_sfixed(29084732.0/4294967296.0,1,-nbitq), 
to_sfixed(-535137306.0/4294967296.0,1,-nbitq), 
to_sfixed(707224528.0/4294967296.0,1,-nbitq), 
to_sfixed(-388741995.0/4294967296.0,1,-nbitq), 
to_sfixed(-407020209.0/4294967296.0,1,-nbitq), 
to_sfixed(-184208394.0/4294967296.0,1,-nbitq), 
to_sfixed(809729211.0/4294967296.0,1,-nbitq), 
to_sfixed(-677918073.0/4294967296.0,1,-nbitq), 
to_sfixed(-285588099.0/4294967296.0,1,-nbitq), 
to_sfixed(562260321.0/4294967296.0,1,-nbitq), 
to_sfixed(-534545645.0/4294967296.0,1,-nbitq), 
to_sfixed(717443202.0/4294967296.0,1,-nbitq), 
to_sfixed(704137181.0/4294967296.0,1,-nbitq), 
to_sfixed(62862605.0/4294967296.0,1,-nbitq), 
to_sfixed(102818695.0/4294967296.0,1,-nbitq), 
to_sfixed(333338152.0/4294967296.0,1,-nbitq), 
to_sfixed(256294050.0/4294967296.0,1,-nbitq), 
to_sfixed(-310056880.0/4294967296.0,1,-nbitq), 
to_sfixed(-424025144.0/4294967296.0,1,-nbitq), 
to_sfixed(-1334376432.0/4294967296.0,1,-nbitq), 
to_sfixed(-242709314.0/4294967296.0,1,-nbitq), 
to_sfixed(-425611865.0/4294967296.0,1,-nbitq), 
to_sfixed(210706652.0/4294967296.0,1,-nbitq), 
to_sfixed(479878667.0/4294967296.0,1,-nbitq), 
to_sfixed(1253683407.0/4294967296.0,1,-nbitq), 
to_sfixed(369883791.0/4294967296.0,1,-nbitq), 
to_sfixed(-229700163.0/4294967296.0,1,-nbitq), 
to_sfixed(278833987.0/4294967296.0,1,-nbitq), 
to_sfixed(89375273.0/4294967296.0,1,-nbitq), 
to_sfixed(142038482.0/4294967296.0,1,-nbitq), 
to_sfixed(166979693.0/4294967296.0,1,-nbitq), 
to_sfixed(-162144999.0/4294967296.0,1,-nbitq), 
to_sfixed(655758181.0/4294967296.0,1,-nbitq), 
to_sfixed(125763080.0/4294967296.0,1,-nbitq), 
to_sfixed(-361433306.0/4294967296.0,1,-nbitq), 
to_sfixed(860415838.0/4294967296.0,1,-nbitq), 
to_sfixed(95041494.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(424249889.0/4294967296.0,1,-nbitq), 
to_sfixed(-515204146.0/4294967296.0,1,-nbitq), 
to_sfixed(-1665226167.0/4294967296.0,1,-nbitq), 
to_sfixed(-887488990.0/4294967296.0,1,-nbitq), 
to_sfixed(184946830.0/4294967296.0,1,-nbitq), 
to_sfixed(2303612908.0/4294967296.0,1,-nbitq), 
to_sfixed(420619113.0/4294967296.0,1,-nbitq), 
to_sfixed(620522834.0/4294967296.0,1,-nbitq), 
to_sfixed(86512246.0/4294967296.0,1,-nbitq), 
to_sfixed(199752158.0/4294967296.0,1,-nbitq), 
to_sfixed(-333904253.0/4294967296.0,1,-nbitq), 
to_sfixed(666568780.0/4294967296.0,1,-nbitq), 
to_sfixed(1150066827.0/4294967296.0,1,-nbitq), 
to_sfixed(905704941.0/4294967296.0,1,-nbitq), 
to_sfixed(80296659.0/4294967296.0,1,-nbitq), 
to_sfixed(520030334.0/4294967296.0,1,-nbitq), 
to_sfixed(149976128.0/4294967296.0,1,-nbitq), 
to_sfixed(319753139.0/4294967296.0,1,-nbitq), 
to_sfixed(-406561364.0/4294967296.0,1,-nbitq), 
to_sfixed(653837242.0/4294967296.0,1,-nbitq), 
to_sfixed(-225046725.0/4294967296.0,1,-nbitq), 
to_sfixed(-1282537319.0/4294967296.0,1,-nbitq), 
to_sfixed(-1032161018.0/4294967296.0,1,-nbitq), 
to_sfixed(336279388.0/4294967296.0,1,-nbitq), 
to_sfixed(-40201733.0/4294967296.0,1,-nbitq), 
to_sfixed(530026076.0/4294967296.0,1,-nbitq), 
to_sfixed(220616650.0/4294967296.0,1,-nbitq), 
to_sfixed(-512832833.0/4294967296.0,1,-nbitq), 
to_sfixed(781601320.0/4294967296.0,1,-nbitq), 
to_sfixed(940430398.0/4294967296.0,1,-nbitq), 
to_sfixed(-478938271.0/4294967296.0,1,-nbitq), 
to_sfixed(528295167.0/4294967296.0,1,-nbitq), 
to_sfixed(-135774342.0/4294967296.0,1,-nbitq), 
to_sfixed(570011314.0/4294967296.0,1,-nbitq), 
to_sfixed(-196727815.0/4294967296.0,1,-nbitq), 
to_sfixed(-213781297.0/4294967296.0,1,-nbitq), 
to_sfixed(-126655862.0/4294967296.0,1,-nbitq), 
to_sfixed(613346946.0/4294967296.0,1,-nbitq), 
to_sfixed(169310353.0/4294967296.0,1,-nbitq), 
to_sfixed(-23960742.0/4294967296.0,1,-nbitq), 
to_sfixed(-221832493.0/4294967296.0,1,-nbitq), 
to_sfixed(-350197066.0/4294967296.0,1,-nbitq), 
to_sfixed(-18489943.0/4294967296.0,1,-nbitq), 
to_sfixed(-239465614.0/4294967296.0,1,-nbitq), 
to_sfixed(-739685265.0/4294967296.0,1,-nbitq), 
to_sfixed(43717133.0/4294967296.0,1,-nbitq), 
to_sfixed(223809487.0/4294967296.0,1,-nbitq), 
to_sfixed(317656765.0/4294967296.0,1,-nbitq), 
to_sfixed(198449740.0/4294967296.0,1,-nbitq), 
to_sfixed(883959206.0/4294967296.0,1,-nbitq), 
to_sfixed(8483698.0/4294967296.0,1,-nbitq), 
to_sfixed(-694978762.0/4294967296.0,1,-nbitq), 
to_sfixed(1187329390.0/4294967296.0,1,-nbitq), 
to_sfixed(-1193019271.0/4294967296.0,1,-nbitq), 
to_sfixed(1157311852.0/4294967296.0,1,-nbitq), 
to_sfixed(400184310.0/4294967296.0,1,-nbitq), 
to_sfixed(41622977.0/4294967296.0,1,-nbitq), 
to_sfixed(744292029.0/4294967296.0,1,-nbitq), 
to_sfixed(-169416925.0/4294967296.0,1,-nbitq), 
to_sfixed(354574755.0/4294967296.0,1,-nbitq), 
to_sfixed(122022643.0/4294967296.0,1,-nbitq), 
to_sfixed(294699179.0/4294967296.0,1,-nbitq), 
to_sfixed(-969622672.0/4294967296.0,1,-nbitq), 
to_sfixed(-904030563.0/4294967296.0,1,-nbitq), 
to_sfixed(170855573.0/4294967296.0,1,-nbitq), 
to_sfixed(-594013418.0/4294967296.0,1,-nbitq), 
to_sfixed(56837691.0/4294967296.0,1,-nbitq), 
to_sfixed(1335877510.0/4294967296.0,1,-nbitq), 
to_sfixed(393393574.0/4294967296.0,1,-nbitq), 
to_sfixed(-841729395.0/4294967296.0,1,-nbitq), 
to_sfixed(1077389816.0/4294967296.0,1,-nbitq), 
to_sfixed(-612742117.0/4294967296.0,1,-nbitq), 
to_sfixed(81580567.0/4294967296.0,1,-nbitq), 
to_sfixed(-228043466.0/4294967296.0,1,-nbitq), 
to_sfixed(-273879358.0/4294967296.0,1,-nbitq), 
to_sfixed(190082275.0/4294967296.0,1,-nbitq), 
to_sfixed(633845108.0/4294967296.0,1,-nbitq), 
to_sfixed(-718742427.0/4294967296.0,1,-nbitq), 
to_sfixed(1610431615.0/4294967296.0,1,-nbitq), 
to_sfixed(-118505528.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(289094244.0/4294967296.0,1,-nbitq), 
to_sfixed(-602157797.0/4294967296.0,1,-nbitq), 
to_sfixed(-2434281443.0/4294967296.0,1,-nbitq), 
to_sfixed(-960800194.0/4294967296.0,1,-nbitq), 
to_sfixed(109759172.0/4294967296.0,1,-nbitq), 
to_sfixed(2209570405.0/4294967296.0,1,-nbitq), 
to_sfixed(259758897.0/4294967296.0,1,-nbitq), 
to_sfixed(736086268.0/4294967296.0,1,-nbitq), 
to_sfixed(-59020795.0/4294967296.0,1,-nbitq), 
to_sfixed(111201047.0/4294967296.0,1,-nbitq), 
to_sfixed(-36161587.0/4294967296.0,1,-nbitq), 
to_sfixed(564008041.0/4294967296.0,1,-nbitq), 
to_sfixed(621302779.0/4294967296.0,1,-nbitq), 
to_sfixed(1082370918.0/4294967296.0,1,-nbitq), 
to_sfixed(-252944116.0/4294967296.0,1,-nbitq), 
to_sfixed(678605184.0/4294967296.0,1,-nbitq), 
to_sfixed(1982570.0/4294967296.0,1,-nbitq), 
to_sfixed(-185906724.0/4294967296.0,1,-nbitq), 
to_sfixed(450982809.0/4294967296.0,1,-nbitq), 
to_sfixed(-79227376.0/4294967296.0,1,-nbitq), 
to_sfixed(-364890563.0/4294967296.0,1,-nbitq), 
to_sfixed(-1205451958.0/4294967296.0,1,-nbitq), 
to_sfixed(-840840846.0/4294967296.0,1,-nbitq), 
to_sfixed(351259121.0/4294967296.0,1,-nbitq), 
to_sfixed(-277214924.0/4294967296.0,1,-nbitq), 
to_sfixed(451006270.0/4294967296.0,1,-nbitq), 
to_sfixed(-319673803.0/4294967296.0,1,-nbitq), 
to_sfixed(-13596403.0/4294967296.0,1,-nbitq), 
to_sfixed(-274069189.0/4294967296.0,1,-nbitq), 
to_sfixed(329816672.0/4294967296.0,1,-nbitq), 
to_sfixed(-247460744.0/4294967296.0,1,-nbitq), 
to_sfixed(-277656736.0/4294967296.0,1,-nbitq), 
to_sfixed(14476252.0/4294967296.0,1,-nbitq), 
to_sfixed(581622433.0/4294967296.0,1,-nbitq), 
to_sfixed(-460708498.0/4294967296.0,1,-nbitq), 
to_sfixed(-327034870.0/4294967296.0,1,-nbitq), 
to_sfixed(25406359.0/4294967296.0,1,-nbitq), 
to_sfixed(387743870.0/4294967296.0,1,-nbitq), 
to_sfixed(76889815.0/4294967296.0,1,-nbitq), 
to_sfixed(-104604624.0/4294967296.0,1,-nbitq), 
to_sfixed(-110322763.0/4294967296.0,1,-nbitq), 
to_sfixed(-544607139.0/4294967296.0,1,-nbitq), 
to_sfixed(887552604.0/4294967296.0,1,-nbitq), 
to_sfixed(517379107.0/4294967296.0,1,-nbitq), 
to_sfixed(-332896963.0/4294967296.0,1,-nbitq), 
to_sfixed(465051458.0/4294967296.0,1,-nbitq), 
to_sfixed(310346384.0/4294967296.0,1,-nbitq), 
to_sfixed(-162753041.0/4294967296.0,1,-nbitq), 
to_sfixed(421343244.0/4294967296.0,1,-nbitq), 
to_sfixed(1066488741.0/4294967296.0,1,-nbitq), 
to_sfixed(-341907168.0/4294967296.0,1,-nbitq), 
to_sfixed(-481320926.0/4294967296.0,1,-nbitq), 
to_sfixed(77142148.0/4294967296.0,1,-nbitq), 
to_sfixed(-1089073860.0/4294967296.0,1,-nbitq), 
to_sfixed(461126577.0/4294967296.0,1,-nbitq), 
to_sfixed(-505934771.0/4294967296.0,1,-nbitq), 
to_sfixed(-67130661.0/4294967296.0,1,-nbitq), 
to_sfixed(823612894.0/4294967296.0,1,-nbitq), 
to_sfixed(76736196.0/4294967296.0,1,-nbitq), 
to_sfixed(258799368.0/4294967296.0,1,-nbitq), 
to_sfixed(394770030.0/4294967296.0,1,-nbitq), 
to_sfixed(64369708.0/4294967296.0,1,-nbitq), 
to_sfixed(-1677599171.0/4294967296.0,1,-nbitq), 
to_sfixed(-1103187992.0/4294967296.0,1,-nbitq), 
to_sfixed(-194724131.0/4294967296.0,1,-nbitq), 
to_sfixed(-216162885.0/4294967296.0,1,-nbitq), 
to_sfixed(-1020332587.0/4294967296.0,1,-nbitq), 
to_sfixed(827152981.0/4294967296.0,1,-nbitq), 
to_sfixed(238246217.0/4294967296.0,1,-nbitq), 
to_sfixed(-1306064863.0/4294967296.0,1,-nbitq), 
to_sfixed(850644693.0/4294967296.0,1,-nbitq), 
to_sfixed(-891932787.0/4294967296.0,1,-nbitq), 
to_sfixed(609598978.0/4294967296.0,1,-nbitq), 
to_sfixed(-91470709.0/4294967296.0,1,-nbitq), 
to_sfixed(102700578.0/4294967296.0,1,-nbitq), 
to_sfixed(-461822922.0/4294967296.0,1,-nbitq), 
to_sfixed(1056539539.0/4294967296.0,1,-nbitq), 
to_sfixed(-134969502.0/4294967296.0,1,-nbitq), 
to_sfixed(1884822238.0/4294967296.0,1,-nbitq), 
to_sfixed(-57417275.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(239892576.0/4294967296.0,1,-nbitq), 
to_sfixed(-1003451507.0/4294967296.0,1,-nbitq), 
to_sfixed(-3256398814.0/4294967296.0,1,-nbitq), 
to_sfixed(-281548131.0/4294967296.0,1,-nbitq), 
to_sfixed(263562771.0/4294967296.0,1,-nbitq), 
to_sfixed(1177513176.0/4294967296.0,1,-nbitq), 
to_sfixed(-219309834.0/4294967296.0,1,-nbitq), 
to_sfixed(1620008071.0/4294967296.0,1,-nbitq), 
to_sfixed(-451537642.0/4294967296.0,1,-nbitq), 
to_sfixed(-108711307.0/4294967296.0,1,-nbitq), 
to_sfixed(732501071.0/4294967296.0,1,-nbitq), 
to_sfixed(324563440.0/4294967296.0,1,-nbitq), 
to_sfixed(989310093.0/4294967296.0,1,-nbitq), 
to_sfixed(840118216.0/4294967296.0,1,-nbitq), 
to_sfixed(30302376.0/4294967296.0,1,-nbitq), 
to_sfixed(1004477171.0/4294967296.0,1,-nbitq), 
to_sfixed(303605161.0/4294967296.0,1,-nbitq), 
to_sfixed(431697573.0/4294967296.0,1,-nbitq), 
to_sfixed(-660284546.0/4294967296.0,1,-nbitq), 
to_sfixed(425398648.0/4294967296.0,1,-nbitq), 
to_sfixed(113709675.0/4294967296.0,1,-nbitq), 
to_sfixed(-1592472760.0/4294967296.0,1,-nbitq), 
to_sfixed(-795733934.0/4294967296.0,1,-nbitq), 
to_sfixed(1185438513.0/4294967296.0,1,-nbitq), 
to_sfixed(-149642259.0/4294967296.0,1,-nbitq), 
to_sfixed(726776148.0/4294967296.0,1,-nbitq), 
to_sfixed(153741979.0/4294967296.0,1,-nbitq), 
to_sfixed(801266443.0/4294967296.0,1,-nbitq), 
to_sfixed(663026325.0/4294967296.0,1,-nbitq), 
to_sfixed(591491830.0/4294967296.0,1,-nbitq), 
to_sfixed(377851567.0/4294967296.0,1,-nbitq), 
to_sfixed(175751908.0/4294967296.0,1,-nbitq), 
to_sfixed(501399573.0/4294967296.0,1,-nbitq), 
to_sfixed(-626180652.0/4294967296.0,1,-nbitq), 
to_sfixed(-402533864.0/4294967296.0,1,-nbitq), 
to_sfixed(-833014831.0/4294967296.0,1,-nbitq), 
to_sfixed(-295236095.0/4294967296.0,1,-nbitq), 
to_sfixed(628590468.0/4294967296.0,1,-nbitq), 
to_sfixed(-140869404.0/4294967296.0,1,-nbitq), 
to_sfixed(-282773334.0/4294967296.0,1,-nbitq), 
to_sfixed(-212492374.0/4294967296.0,1,-nbitq), 
to_sfixed(-918855831.0/4294967296.0,1,-nbitq), 
to_sfixed(424151711.0/4294967296.0,1,-nbitq), 
to_sfixed(134694146.0/4294967296.0,1,-nbitq), 
to_sfixed(-745824149.0/4294967296.0,1,-nbitq), 
to_sfixed(192974775.0/4294967296.0,1,-nbitq), 
to_sfixed(339213881.0/4294967296.0,1,-nbitq), 
to_sfixed(142992943.0/4294967296.0,1,-nbitq), 
to_sfixed(37514752.0/4294967296.0,1,-nbitq), 
to_sfixed(603740109.0/4294967296.0,1,-nbitq), 
to_sfixed(-599375586.0/4294967296.0,1,-nbitq), 
to_sfixed(-864677669.0/4294967296.0,1,-nbitq), 
to_sfixed(426145.0/4294967296.0,1,-nbitq), 
to_sfixed(-115401285.0/4294967296.0,1,-nbitq), 
to_sfixed(170827204.0/4294967296.0,1,-nbitq), 
to_sfixed(-815319287.0/4294967296.0,1,-nbitq), 
to_sfixed(-131616592.0/4294967296.0,1,-nbitq), 
to_sfixed(558502305.0/4294967296.0,1,-nbitq), 
to_sfixed(-29095818.0/4294967296.0,1,-nbitq), 
to_sfixed(-234346991.0/4294967296.0,1,-nbitq), 
to_sfixed(-156100259.0/4294967296.0,1,-nbitq), 
to_sfixed(283050634.0/4294967296.0,1,-nbitq), 
to_sfixed(-1357470713.0/4294967296.0,1,-nbitq), 
to_sfixed(-176249643.0/4294967296.0,1,-nbitq), 
to_sfixed(-384559122.0/4294967296.0,1,-nbitq), 
to_sfixed(178729361.0/4294967296.0,1,-nbitq), 
to_sfixed(-1039476402.0/4294967296.0,1,-nbitq), 
to_sfixed(432207566.0/4294967296.0,1,-nbitq), 
to_sfixed(10029275.0/4294967296.0,1,-nbitq), 
to_sfixed(-655276021.0/4294967296.0,1,-nbitq), 
to_sfixed(1688165686.0/4294967296.0,1,-nbitq), 
to_sfixed(-253876699.0/4294967296.0,1,-nbitq), 
to_sfixed(716247563.0/4294967296.0,1,-nbitq), 
to_sfixed(-7035487.0/4294967296.0,1,-nbitq), 
to_sfixed(-188315171.0/4294967296.0,1,-nbitq), 
to_sfixed(453597743.0/4294967296.0,1,-nbitq), 
to_sfixed(596266840.0/4294967296.0,1,-nbitq), 
to_sfixed(-434091261.0/4294967296.0,1,-nbitq), 
to_sfixed(1750996421.0/4294967296.0,1,-nbitq), 
to_sfixed(-138431844.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(744112618.0/4294967296.0,1,-nbitq), 
to_sfixed(-1049125602.0/4294967296.0,1,-nbitq), 
to_sfixed(-1409313924.0/4294967296.0,1,-nbitq), 
to_sfixed(-427104495.0/4294967296.0,1,-nbitq), 
to_sfixed(587237197.0/4294967296.0,1,-nbitq), 
to_sfixed(-103281718.0/4294967296.0,1,-nbitq), 
to_sfixed(104092810.0/4294967296.0,1,-nbitq), 
to_sfixed(-1427768296.0/4294967296.0,1,-nbitq), 
to_sfixed(-622232447.0/4294967296.0,1,-nbitq), 
to_sfixed(-198611461.0/4294967296.0,1,-nbitq), 
to_sfixed(593294567.0/4294967296.0,1,-nbitq), 
to_sfixed(-1229856029.0/4294967296.0,1,-nbitq), 
to_sfixed(741647936.0/4294967296.0,1,-nbitq), 
to_sfixed(-1039974171.0/4294967296.0,1,-nbitq), 
to_sfixed(-291336683.0/4294967296.0,1,-nbitq), 
to_sfixed(1091554646.0/4294967296.0,1,-nbitq), 
to_sfixed(-202610245.0/4294967296.0,1,-nbitq), 
to_sfixed(191869424.0/4294967296.0,1,-nbitq), 
to_sfixed(-1321227151.0/4294967296.0,1,-nbitq), 
to_sfixed(-638838211.0/4294967296.0,1,-nbitq), 
to_sfixed(-375530857.0/4294967296.0,1,-nbitq), 
to_sfixed(-1007933837.0/4294967296.0,1,-nbitq), 
to_sfixed(-557776015.0/4294967296.0,1,-nbitq), 
to_sfixed(1483765811.0/4294967296.0,1,-nbitq), 
to_sfixed(-308632101.0/4294967296.0,1,-nbitq), 
to_sfixed(1599624287.0/4294967296.0,1,-nbitq), 
to_sfixed(-90844105.0/4294967296.0,1,-nbitq), 
to_sfixed(1143252590.0/4294967296.0,1,-nbitq), 
to_sfixed(930912002.0/4294967296.0,1,-nbitq), 
to_sfixed(797187673.0/4294967296.0,1,-nbitq), 
to_sfixed(381974162.0/4294967296.0,1,-nbitq), 
to_sfixed(-48371924.0/4294967296.0,1,-nbitq), 
to_sfixed(303767904.0/4294967296.0,1,-nbitq), 
to_sfixed(-607000728.0/4294967296.0,1,-nbitq), 
to_sfixed(-24444849.0/4294967296.0,1,-nbitq), 
to_sfixed(-1567861576.0/4294967296.0,1,-nbitq), 
to_sfixed(-383573666.0/4294967296.0,1,-nbitq), 
to_sfixed(322315455.0/4294967296.0,1,-nbitq), 
to_sfixed(-297520057.0/4294967296.0,1,-nbitq), 
to_sfixed(-13403230.0/4294967296.0,1,-nbitq), 
to_sfixed(-221709535.0/4294967296.0,1,-nbitq), 
to_sfixed(-891151210.0/4294967296.0,1,-nbitq), 
to_sfixed(445721191.0/4294967296.0,1,-nbitq), 
to_sfixed(781969958.0/4294967296.0,1,-nbitq), 
to_sfixed(-952636435.0/4294967296.0,1,-nbitq), 
to_sfixed(30605475.0/4294967296.0,1,-nbitq), 
to_sfixed(-81831332.0/4294967296.0,1,-nbitq), 
to_sfixed(-195503131.0/4294967296.0,1,-nbitq), 
to_sfixed(-83800111.0/4294967296.0,1,-nbitq), 
to_sfixed(1894453675.0/4294967296.0,1,-nbitq), 
to_sfixed(-618342843.0/4294967296.0,1,-nbitq), 
to_sfixed(-1111876179.0/4294967296.0,1,-nbitq), 
to_sfixed(-399519173.0/4294967296.0,1,-nbitq), 
to_sfixed(206791754.0/4294967296.0,1,-nbitq), 
to_sfixed(-273848657.0/4294967296.0,1,-nbitq), 
to_sfixed(-1009809842.0/4294967296.0,1,-nbitq), 
to_sfixed(48666039.0/4294967296.0,1,-nbitq), 
to_sfixed(899023418.0/4294967296.0,1,-nbitq), 
to_sfixed(241742226.0/4294967296.0,1,-nbitq), 
to_sfixed(-277744519.0/4294967296.0,1,-nbitq), 
to_sfixed(-113039471.0/4294967296.0,1,-nbitq), 
to_sfixed(1111591685.0/4294967296.0,1,-nbitq), 
to_sfixed(-104948915.0/4294967296.0,1,-nbitq), 
to_sfixed(392352454.0/4294967296.0,1,-nbitq), 
to_sfixed(-822166.0/4294967296.0,1,-nbitq), 
to_sfixed(-132607098.0/4294967296.0,1,-nbitq), 
to_sfixed(-392847834.0/4294967296.0,1,-nbitq), 
to_sfixed(1892136619.0/4294967296.0,1,-nbitq), 
to_sfixed(-98013591.0/4294967296.0,1,-nbitq), 
to_sfixed(-174540796.0/4294967296.0,1,-nbitq), 
to_sfixed(1118370046.0/4294967296.0,1,-nbitq), 
to_sfixed(-707632079.0/4294967296.0,1,-nbitq), 
to_sfixed(413175634.0/4294967296.0,1,-nbitq), 
to_sfixed(172994358.0/4294967296.0,1,-nbitq), 
to_sfixed(252868594.0/4294967296.0,1,-nbitq), 
to_sfixed(554018784.0/4294967296.0,1,-nbitq), 
to_sfixed(166423730.0/4294967296.0,1,-nbitq), 
to_sfixed(-11896040.0/4294967296.0,1,-nbitq), 
to_sfixed(1366212165.0/4294967296.0,1,-nbitq), 
to_sfixed(212844321.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-31824001.0/4294967296.0,1,-nbitq), 
to_sfixed(-427269059.0/4294967296.0,1,-nbitq), 
to_sfixed(873631086.0/4294967296.0,1,-nbitq), 
to_sfixed(57271024.0/4294967296.0,1,-nbitq), 
to_sfixed(387911489.0/4294967296.0,1,-nbitq), 
to_sfixed(346942926.0/4294967296.0,1,-nbitq), 
to_sfixed(-96103832.0/4294967296.0,1,-nbitq), 
to_sfixed(-2275902923.0/4294967296.0,1,-nbitq), 
to_sfixed(456262686.0/4294967296.0,1,-nbitq), 
to_sfixed(-196019877.0/4294967296.0,1,-nbitq), 
to_sfixed(817684305.0/4294967296.0,1,-nbitq), 
to_sfixed(-602950762.0/4294967296.0,1,-nbitq), 
to_sfixed(827437149.0/4294967296.0,1,-nbitq), 
to_sfixed(-906784996.0/4294967296.0,1,-nbitq), 
to_sfixed(139334282.0/4294967296.0,1,-nbitq), 
to_sfixed(1742020325.0/4294967296.0,1,-nbitq), 
to_sfixed(-98675380.0/4294967296.0,1,-nbitq), 
to_sfixed(-231843244.0/4294967296.0,1,-nbitq), 
to_sfixed(-170173529.0/4294967296.0,1,-nbitq), 
to_sfixed(-552811750.0/4294967296.0,1,-nbitq), 
to_sfixed(48539795.0/4294967296.0,1,-nbitq), 
to_sfixed(-658105970.0/4294967296.0,1,-nbitq), 
to_sfixed(-214335340.0/4294967296.0,1,-nbitq), 
to_sfixed(2457748065.0/4294967296.0,1,-nbitq), 
to_sfixed(223349418.0/4294967296.0,1,-nbitq), 
to_sfixed(717335103.0/4294967296.0,1,-nbitq), 
to_sfixed(455152739.0/4294967296.0,1,-nbitq), 
to_sfixed(613200915.0/4294967296.0,1,-nbitq), 
to_sfixed(-1475481857.0/4294967296.0,1,-nbitq), 
to_sfixed(518421281.0/4294967296.0,1,-nbitq), 
to_sfixed(995081042.0/4294967296.0,1,-nbitq), 
to_sfixed(-111174663.0/4294967296.0,1,-nbitq), 
to_sfixed(444757947.0/4294967296.0,1,-nbitq), 
to_sfixed(-271295304.0/4294967296.0,1,-nbitq), 
to_sfixed(-905743060.0/4294967296.0,1,-nbitq), 
to_sfixed(-1289716690.0/4294967296.0,1,-nbitq), 
to_sfixed(-282916573.0/4294967296.0,1,-nbitq), 
to_sfixed(656286514.0/4294967296.0,1,-nbitq), 
to_sfixed(367371115.0/4294967296.0,1,-nbitq), 
to_sfixed(374003917.0/4294967296.0,1,-nbitq), 
to_sfixed(1360373220.0/4294967296.0,1,-nbitq), 
to_sfixed(-4899698.0/4294967296.0,1,-nbitq), 
to_sfixed(421626798.0/4294967296.0,1,-nbitq), 
to_sfixed(168551274.0/4294967296.0,1,-nbitq), 
to_sfixed(-111595880.0/4294967296.0,1,-nbitq), 
to_sfixed(-741911749.0/4294967296.0,1,-nbitq), 
to_sfixed(17493632.0/4294967296.0,1,-nbitq), 
to_sfixed(-198407978.0/4294967296.0,1,-nbitq), 
to_sfixed(-58567897.0/4294967296.0,1,-nbitq), 
to_sfixed(1298448804.0/4294967296.0,1,-nbitq), 
to_sfixed(454966522.0/4294967296.0,1,-nbitq), 
to_sfixed(-1006656247.0/4294967296.0,1,-nbitq), 
to_sfixed(-371435890.0/4294967296.0,1,-nbitq), 
to_sfixed(-78240217.0/4294967296.0,1,-nbitq), 
to_sfixed(219942124.0/4294967296.0,1,-nbitq), 
to_sfixed(-1026059738.0/4294967296.0,1,-nbitq), 
to_sfixed(41295796.0/4294967296.0,1,-nbitq), 
to_sfixed(246719622.0/4294967296.0,1,-nbitq), 
to_sfixed(13226260.0/4294967296.0,1,-nbitq), 
to_sfixed(-130587601.0/4294967296.0,1,-nbitq), 
to_sfixed(-252994249.0/4294967296.0,1,-nbitq), 
to_sfixed(432051893.0/4294967296.0,1,-nbitq), 
to_sfixed(1201373622.0/4294967296.0,1,-nbitq), 
to_sfixed(1169156427.0/4294967296.0,1,-nbitq), 
to_sfixed(78180318.0/4294967296.0,1,-nbitq), 
to_sfixed(136193352.0/4294967296.0,1,-nbitq), 
to_sfixed(618174366.0/4294967296.0,1,-nbitq), 
to_sfixed(2130175121.0/4294967296.0,1,-nbitq), 
to_sfixed(-376898281.0/4294967296.0,1,-nbitq), 
to_sfixed(1283618353.0/4294967296.0,1,-nbitq), 
to_sfixed(605935361.0/4294967296.0,1,-nbitq), 
to_sfixed(-251789384.0/4294967296.0,1,-nbitq), 
to_sfixed(589973850.0/4294967296.0,1,-nbitq), 
to_sfixed(89265424.0/4294967296.0,1,-nbitq), 
to_sfixed(222004892.0/4294967296.0,1,-nbitq), 
to_sfixed(-240994791.0/4294967296.0,1,-nbitq), 
to_sfixed(833017323.0/4294967296.0,1,-nbitq), 
to_sfixed(71482725.0/4294967296.0,1,-nbitq), 
to_sfixed(848912125.0/4294967296.0,1,-nbitq), 
to_sfixed(185745338.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(252632306.0/4294967296.0,1,-nbitq), 
to_sfixed(592217935.0/4294967296.0,1,-nbitq), 
to_sfixed(390728441.0/4294967296.0,1,-nbitq), 
to_sfixed(451719339.0/4294967296.0,1,-nbitq), 
to_sfixed(337152774.0/4294967296.0,1,-nbitq), 
to_sfixed(-193388526.0/4294967296.0,1,-nbitq), 
to_sfixed(130386192.0/4294967296.0,1,-nbitq), 
to_sfixed(-483519286.0/4294967296.0,1,-nbitq), 
to_sfixed(737788076.0/4294967296.0,1,-nbitq), 
to_sfixed(-285497966.0/4294967296.0,1,-nbitq), 
to_sfixed(1040056931.0/4294967296.0,1,-nbitq), 
to_sfixed(-1003529569.0/4294967296.0,1,-nbitq), 
to_sfixed(1055149035.0/4294967296.0,1,-nbitq), 
to_sfixed(485860714.0/4294967296.0,1,-nbitq), 
to_sfixed(-233651336.0/4294967296.0,1,-nbitq), 
to_sfixed(2300306740.0/4294967296.0,1,-nbitq), 
to_sfixed(229918937.0/4294967296.0,1,-nbitq), 
to_sfixed(347136259.0/4294967296.0,1,-nbitq), 
to_sfixed(-65726933.0/4294967296.0,1,-nbitq), 
to_sfixed(259069004.0/4294967296.0,1,-nbitq), 
to_sfixed(-376208482.0/4294967296.0,1,-nbitq), 
to_sfixed(35726754.0/4294967296.0,1,-nbitq), 
to_sfixed(718383596.0/4294967296.0,1,-nbitq), 
to_sfixed(2362198676.0/4294967296.0,1,-nbitq), 
to_sfixed(147758757.0/4294967296.0,1,-nbitq), 
to_sfixed(243787369.0/4294967296.0,1,-nbitq), 
to_sfixed(372624798.0/4294967296.0,1,-nbitq), 
to_sfixed(-203604768.0/4294967296.0,1,-nbitq), 
to_sfixed(-2275499758.0/4294967296.0,1,-nbitq), 
to_sfixed(545885908.0/4294967296.0,1,-nbitq), 
to_sfixed(771797142.0/4294967296.0,1,-nbitq), 
to_sfixed(1092215106.0/4294967296.0,1,-nbitq), 
to_sfixed(-323131195.0/4294967296.0,1,-nbitq), 
to_sfixed(-35078203.0/4294967296.0,1,-nbitq), 
to_sfixed(-809308752.0/4294967296.0,1,-nbitq), 
to_sfixed(180650940.0/4294967296.0,1,-nbitq), 
to_sfixed(137449974.0/4294967296.0,1,-nbitq), 
to_sfixed(1129676316.0/4294967296.0,1,-nbitq), 
to_sfixed(92876717.0/4294967296.0,1,-nbitq), 
to_sfixed(-15019837.0/4294967296.0,1,-nbitq), 
to_sfixed(2033977764.0/4294967296.0,1,-nbitq), 
to_sfixed(395315998.0/4294967296.0,1,-nbitq), 
to_sfixed(-528271490.0/4294967296.0,1,-nbitq), 
to_sfixed(-1134939181.0/4294967296.0,1,-nbitq), 
to_sfixed(157645286.0/4294967296.0,1,-nbitq), 
to_sfixed(-834660301.0/4294967296.0,1,-nbitq), 
to_sfixed(-442368446.0/4294967296.0,1,-nbitq), 
to_sfixed(656213673.0/4294967296.0,1,-nbitq), 
to_sfixed(-189639095.0/4294967296.0,1,-nbitq), 
to_sfixed(273608375.0/4294967296.0,1,-nbitq), 
to_sfixed(294803631.0/4294967296.0,1,-nbitq), 
to_sfixed(-1742845756.0/4294967296.0,1,-nbitq), 
to_sfixed(-329115411.0/4294967296.0,1,-nbitq), 
to_sfixed(-1086709316.0/4294967296.0,1,-nbitq), 
to_sfixed(374974523.0/4294967296.0,1,-nbitq), 
to_sfixed(-1177185710.0/4294967296.0,1,-nbitq), 
to_sfixed(-1143030457.0/4294967296.0,1,-nbitq), 
to_sfixed(387121728.0/4294967296.0,1,-nbitq), 
to_sfixed(-252581528.0/4294967296.0,1,-nbitq), 
to_sfixed(-107744743.0/4294967296.0,1,-nbitq), 
to_sfixed(-38178694.0/4294967296.0,1,-nbitq), 
to_sfixed(-231307204.0/4294967296.0,1,-nbitq), 
to_sfixed(963651378.0/4294967296.0,1,-nbitq), 
to_sfixed(307988987.0/4294967296.0,1,-nbitq), 
to_sfixed(-217362338.0/4294967296.0,1,-nbitq), 
to_sfixed(504222311.0/4294967296.0,1,-nbitq), 
to_sfixed(1308245695.0/4294967296.0,1,-nbitq), 
to_sfixed(1877485454.0/4294967296.0,1,-nbitq), 
to_sfixed(-41522418.0/4294967296.0,1,-nbitq), 
to_sfixed(1612877482.0/4294967296.0,1,-nbitq), 
to_sfixed(757023286.0/4294967296.0,1,-nbitq), 
to_sfixed(257550671.0/4294967296.0,1,-nbitq), 
to_sfixed(104284033.0/4294967296.0,1,-nbitq), 
to_sfixed(106046887.0/4294967296.0,1,-nbitq), 
to_sfixed(94855546.0/4294967296.0,1,-nbitq), 
to_sfixed(-1169407105.0/4294967296.0,1,-nbitq), 
to_sfixed(1025658837.0/4294967296.0,1,-nbitq), 
to_sfixed(-603357575.0/4294967296.0,1,-nbitq), 
to_sfixed(-480723217.0/4294967296.0,1,-nbitq), 
to_sfixed(369066445.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(459516033.0/4294967296.0,1,-nbitq), 
to_sfixed(1366512861.0/4294967296.0,1,-nbitq), 
to_sfixed(167232715.0/4294967296.0,1,-nbitq), 
to_sfixed(280411225.0/4294967296.0,1,-nbitq), 
to_sfixed(-452700460.0/4294967296.0,1,-nbitq), 
to_sfixed(-701789562.0/4294967296.0,1,-nbitq), 
to_sfixed(-59459676.0/4294967296.0,1,-nbitq), 
to_sfixed(1414128252.0/4294967296.0,1,-nbitq), 
to_sfixed(-659511055.0/4294967296.0,1,-nbitq), 
to_sfixed(-49632195.0/4294967296.0,1,-nbitq), 
to_sfixed(234263502.0/4294967296.0,1,-nbitq), 
to_sfixed(-1986701604.0/4294967296.0,1,-nbitq), 
to_sfixed(359767899.0/4294967296.0,1,-nbitq), 
to_sfixed(-194964813.0/4294967296.0,1,-nbitq), 
to_sfixed(-269479492.0/4294967296.0,1,-nbitq), 
to_sfixed(2417416264.0/4294967296.0,1,-nbitq), 
to_sfixed(-352655210.0/4294967296.0,1,-nbitq), 
to_sfixed(11214562.0/4294967296.0,1,-nbitq), 
to_sfixed(-654628473.0/4294967296.0,1,-nbitq), 
to_sfixed(1238706229.0/4294967296.0,1,-nbitq), 
to_sfixed(-10234883.0/4294967296.0,1,-nbitq), 
to_sfixed(490323744.0/4294967296.0,1,-nbitq), 
to_sfixed(939725585.0/4294967296.0,1,-nbitq), 
to_sfixed(-2299421929.0/4294967296.0,1,-nbitq), 
to_sfixed(-295300196.0/4294967296.0,1,-nbitq), 
to_sfixed(-11123133.0/4294967296.0,1,-nbitq), 
to_sfixed(14099196.0/4294967296.0,1,-nbitq), 
to_sfixed(-1458412812.0/4294967296.0,1,-nbitq), 
to_sfixed(-1252087243.0/4294967296.0,1,-nbitq), 
to_sfixed(97305309.0/4294967296.0,1,-nbitq), 
to_sfixed(-600487002.0/4294967296.0,1,-nbitq), 
to_sfixed(1758311277.0/4294967296.0,1,-nbitq), 
to_sfixed(-178443089.0/4294967296.0,1,-nbitq), 
to_sfixed(418598440.0/4294967296.0,1,-nbitq), 
to_sfixed(-18218318.0/4294967296.0,1,-nbitq), 
to_sfixed(-390943237.0/4294967296.0,1,-nbitq), 
to_sfixed(403973370.0/4294967296.0,1,-nbitq), 
to_sfixed(1612630181.0/4294967296.0,1,-nbitq), 
to_sfixed(-166486853.0/4294967296.0,1,-nbitq), 
to_sfixed(391738824.0/4294967296.0,1,-nbitq), 
to_sfixed(1124569741.0/4294967296.0,1,-nbitq), 
to_sfixed(920240455.0/4294967296.0,1,-nbitq), 
to_sfixed(-23110282.0/4294967296.0,1,-nbitq), 
to_sfixed(-471303702.0/4294967296.0,1,-nbitq), 
to_sfixed(-49988934.0/4294967296.0,1,-nbitq), 
to_sfixed(549775658.0/4294967296.0,1,-nbitq), 
to_sfixed(-376061857.0/4294967296.0,1,-nbitq), 
to_sfixed(821004544.0/4294967296.0,1,-nbitq), 
to_sfixed(388859334.0/4294967296.0,1,-nbitq), 
to_sfixed(-625302264.0/4294967296.0,1,-nbitq), 
to_sfixed(217991344.0/4294967296.0,1,-nbitq), 
to_sfixed(-1357313891.0/4294967296.0,1,-nbitq), 
to_sfixed(-830862464.0/4294967296.0,1,-nbitq), 
to_sfixed(-723132644.0/4294967296.0,1,-nbitq), 
to_sfixed(712302793.0/4294967296.0,1,-nbitq), 
to_sfixed(-1836818276.0/4294967296.0,1,-nbitq), 
to_sfixed(-909055554.0/4294967296.0,1,-nbitq), 
to_sfixed(998901573.0/4294967296.0,1,-nbitq), 
to_sfixed(4612486.0/4294967296.0,1,-nbitq), 
to_sfixed(-380264266.0/4294967296.0,1,-nbitq), 
to_sfixed(72360050.0/4294967296.0,1,-nbitq), 
to_sfixed(98843800.0/4294967296.0,1,-nbitq), 
to_sfixed(292864604.0/4294967296.0,1,-nbitq), 
to_sfixed(558885222.0/4294967296.0,1,-nbitq), 
to_sfixed(-117458862.0/4294967296.0,1,-nbitq), 
to_sfixed(237769049.0/4294967296.0,1,-nbitq), 
to_sfixed(537529885.0/4294967296.0,1,-nbitq), 
to_sfixed(1286416958.0/4294967296.0,1,-nbitq), 
to_sfixed(37895910.0/4294967296.0,1,-nbitq), 
to_sfixed(448995025.0/4294967296.0,1,-nbitq), 
to_sfixed(1151543668.0/4294967296.0,1,-nbitq), 
to_sfixed(-133741371.0/4294967296.0,1,-nbitq), 
to_sfixed(-350444968.0/4294967296.0,1,-nbitq), 
to_sfixed(430026148.0/4294967296.0,1,-nbitq), 
to_sfixed(-326088420.0/4294967296.0,1,-nbitq), 
to_sfixed(-811886423.0/4294967296.0,1,-nbitq), 
to_sfixed(-152309514.0/4294967296.0,1,-nbitq), 
to_sfixed(-172004958.0/4294967296.0,1,-nbitq), 
to_sfixed(-910713011.0/4294967296.0,1,-nbitq), 
to_sfixed(48414285.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(556970026.0/4294967296.0,1,-nbitq), 
to_sfixed(1689608687.0/4294967296.0,1,-nbitq), 
to_sfixed(-220250990.0/4294967296.0,1,-nbitq), 
to_sfixed(338859655.0/4294967296.0,1,-nbitq), 
to_sfixed(-697375738.0/4294967296.0,1,-nbitq), 
to_sfixed(87300450.0/4294967296.0,1,-nbitq), 
to_sfixed(-84371488.0/4294967296.0,1,-nbitq), 
to_sfixed(1196140914.0/4294967296.0,1,-nbitq), 
to_sfixed(-484550021.0/4294967296.0,1,-nbitq), 
to_sfixed(241973814.0/4294967296.0,1,-nbitq), 
to_sfixed(-581717648.0/4294967296.0,1,-nbitq), 
to_sfixed(-2271746602.0/4294967296.0,1,-nbitq), 
to_sfixed(23303941.0/4294967296.0,1,-nbitq), 
to_sfixed(704279950.0/4294967296.0,1,-nbitq), 
to_sfixed(259064916.0/4294967296.0,1,-nbitq), 
to_sfixed(1238149959.0/4294967296.0,1,-nbitq), 
to_sfixed(-259632326.0/4294967296.0,1,-nbitq), 
to_sfixed(359625466.0/4294967296.0,1,-nbitq), 
to_sfixed(-354986510.0/4294967296.0,1,-nbitq), 
to_sfixed(856615272.0/4294967296.0,1,-nbitq), 
to_sfixed(-13062226.0/4294967296.0,1,-nbitq), 
to_sfixed(236356851.0/4294967296.0,1,-nbitq), 
to_sfixed(74733873.0/4294967296.0,1,-nbitq), 
to_sfixed(-3070422651.0/4294967296.0,1,-nbitq), 
to_sfixed(282944037.0/4294967296.0,1,-nbitq), 
to_sfixed(-1141871529.0/4294967296.0,1,-nbitq), 
to_sfixed(-769255493.0/4294967296.0,1,-nbitq), 
to_sfixed(-907210045.0/4294967296.0,1,-nbitq), 
to_sfixed(-105492284.0/4294967296.0,1,-nbitq), 
to_sfixed(474854194.0/4294967296.0,1,-nbitq), 
to_sfixed(-1852321041.0/4294967296.0,1,-nbitq), 
to_sfixed(1145290042.0/4294967296.0,1,-nbitq), 
to_sfixed(511811746.0/4294967296.0,1,-nbitq), 
to_sfixed(826328501.0/4294967296.0,1,-nbitq), 
to_sfixed(782927616.0/4294967296.0,1,-nbitq), 
to_sfixed(-423252249.0/4294967296.0,1,-nbitq), 
to_sfixed(53507500.0/4294967296.0,1,-nbitq), 
to_sfixed(210672354.0/4294967296.0,1,-nbitq), 
to_sfixed(295245025.0/4294967296.0,1,-nbitq), 
to_sfixed(103845887.0/4294967296.0,1,-nbitq), 
to_sfixed(-363473287.0/4294967296.0,1,-nbitq), 
to_sfixed(1088360758.0/4294967296.0,1,-nbitq), 
to_sfixed(-131324143.0/4294967296.0,1,-nbitq), 
to_sfixed(-662193909.0/4294967296.0,1,-nbitq), 
to_sfixed(-908882944.0/4294967296.0,1,-nbitq), 
to_sfixed(-325669468.0/4294967296.0,1,-nbitq), 
to_sfixed(309187517.0/4294967296.0,1,-nbitq), 
to_sfixed(1326384145.0/4294967296.0,1,-nbitq), 
to_sfixed(235738096.0/4294967296.0,1,-nbitq), 
to_sfixed(-416278466.0/4294967296.0,1,-nbitq), 
to_sfixed(-48359793.0/4294967296.0,1,-nbitq), 
to_sfixed(-282645412.0/4294967296.0,1,-nbitq), 
to_sfixed(564332664.0/4294967296.0,1,-nbitq), 
to_sfixed(-836012799.0/4294967296.0,1,-nbitq), 
to_sfixed(-330276463.0/4294967296.0,1,-nbitq), 
to_sfixed(-1472342058.0/4294967296.0,1,-nbitq), 
to_sfixed(-1286010241.0/4294967296.0,1,-nbitq), 
to_sfixed(1637432473.0/4294967296.0,1,-nbitq), 
to_sfixed(55862511.0/4294967296.0,1,-nbitq), 
to_sfixed(-342189617.0/4294967296.0,1,-nbitq), 
to_sfixed(-92357026.0/4294967296.0,1,-nbitq), 
to_sfixed(141364576.0/4294967296.0,1,-nbitq), 
to_sfixed(165669324.0/4294967296.0,1,-nbitq), 
to_sfixed(560951003.0/4294967296.0,1,-nbitq), 
to_sfixed(-127531947.0/4294967296.0,1,-nbitq), 
to_sfixed(-59901545.0/4294967296.0,1,-nbitq), 
to_sfixed(1285288618.0/4294967296.0,1,-nbitq), 
to_sfixed(-333836570.0/4294967296.0,1,-nbitq), 
to_sfixed(-118049153.0/4294967296.0,1,-nbitq), 
to_sfixed(2499081.0/4294967296.0,1,-nbitq), 
to_sfixed(-85419793.0/4294967296.0,1,-nbitq), 
to_sfixed(315343046.0/4294967296.0,1,-nbitq), 
to_sfixed(-700775194.0/4294967296.0,1,-nbitq), 
to_sfixed(97081601.0/4294967296.0,1,-nbitq), 
to_sfixed(100319806.0/4294967296.0,1,-nbitq), 
to_sfixed(-713915973.0/4294967296.0,1,-nbitq), 
to_sfixed(-484222878.0/4294967296.0,1,-nbitq), 
to_sfixed(-207153458.0/4294967296.0,1,-nbitq), 
to_sfixed(-947431560.0/4294967296.0,1,-nbitq), 
to_sfixed(-241212819.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(341433916.0/4294967296.0,1,-nbitq), 
to_sfixed(2375383429.0/4294967296.0,1,-nbitq), 
to_sfixed(-444555268.0/4294967296.0,1,-nbitq), 
to_sfixed(-422095950.0/4294967296.0,1,-nbitq), 
to_sfixed(148889244.0/4294967296.0,1,-nbitq), 
to_sfixed(1155286653.0/4294967296.0,1,-nbitq), 
to_sfixed(-242320361.0/4294967296.0,1,-nbitq), 
to_sfixed(173683942.0/4294967296.0,1,-nbitq), 
to_sfixed(-864105752.0/4294967296.0,1,-nbitq), 
to_sfixed(-178145546.0/4294967296.0,1,-nbitq), 
to_sfixed(-1365854661.0/4294967296.0,1,-nbitq), 
to_sfixed(-1773046946.0/4294967296.0,1,-nbitq), 
to_sfixed(-190138039.0/4294967296.0,1,-nbitq), 
to_sfixed(291805393.0/4294967296.0,1,-nbitq), 
to_sfixed(-157878688.0/4294967296.0,1,-nbitq), 
to_sfixed(1070393560.0/4294967296.0,1,-nbitq), 
to_sfixed(-47533339.0/4294967296.0,1,-nbitq), 
to_sfixed(297750572.0/4294967296.0,1,-nbitq), 
to_sfixed(468122099.0/4294967296.0,1,-nbitq), 
to_sfixed(470739728.0/4294967296.0,1,-nbitq), 
to_sfixed(179907700.0/4294967296.0,1,-nbitq), 
to_sfixed(404592403.0/4294967296.0,1,-nbitq), 
to_sfixed(628465439.0/4294967296.0,1,-nbitq), 
to_sfixed(-1070812763.0/4294967296.0,1,-nbitq), 
to_sfixed(-109916711.0/4294967296.0,1,-nbitq), 
to_sfixed(-1409985501.0/4294967296.0,1,-nbitq), 
to_sfixed(-342145627.0/4294967296.0,1,-nbitq), 
to_sfixed(-1190274263.0/4294967296.0,1,-nbitq), 
to_sfixed(283733267.0/4294967296.0,1,-nbitq), 
to_sfixed(262768554.0/4294967296.0,1,-nbitq), 
to_sfixed(-765931161.0/4294967296.0,1,-nbitq), 
to_sfixed(846397040.0/4294967296.0,1,-nbitq), 
to_sfixed(-161625728.0/4294967296.0,1,-nbitq), 
to_sfixed(453844230.0/4294967296.0,1,-nbitq), 
to_sfixed(-59166827.0/4294967296.0,1,-nbitq), 
to_sfixed(-66468508.0/4294967296.0,1,-nbitq), 
to_sfixed(-488894594.0/4294967296.0,1,-nbitq), 
to_sfixed(-107519143.0/4294967296.0,1,-nbitq), 
to_sfixed(-83951190.0/4294967296.0,1,-nbitq), 
to_sfixed(-419626471.0/4294967296.0,1,-nbitq), 
to_sfixed(-734817383.0/4294967296.0,1,-nbitq), 
to_sfixed(532781776.0/4294967296.0,1,-nbitq), 
to_sfixed(15042753.0/4294967296.0,1,-nbitq), 
to_sfixed(250373968.0/4294967296.0,1,-nbitq), 
to_sfixed(-1394186785.0/4294967296.0,1,-nbitq), 
to_sfixed(543900916.0/4294967296.0,1,-nbitq), 
to_sfixed(-129151886.0/4294967296.0,1,-nbitq), 
to_sfixed(1372289100.0/4294967296.0,1,-nbitq), 
to_sfixed(413148795.0/4294967296.0,1,-nbitq), 
to_sfixed(-16443052.0/4294967296.0,1,-nbitq), 
to_sfixed(-206290614.0/4294967296.0,1,-nbitq), 
to_sfixed(438019799.0/4294967296.0,1,-nbitq), 
to_sfixed(767984965.0/4294967296.0,1,-nbitq), 
to_sfixed(-576541016.0/4294967296.0,1,-nbitq), 
to_sfixed(-324472596.0/4294967296.0,1,-nbitq), 
to_sfixed(-1210122032.0/4294967296.0,1,-nbitq), 
to_sfixed(-905008597.0/4294967296.0,1,-nbitq), 
to_sfixed(1326430395.0/4294967296.0,1,-nbitq), 
to_sfixed(-150771676.0/4294967296.0,1,-nbitq), 
to_sfixed(98822191.0/4294967296.0,1,-nbitq), 
to_sfixed(-44792306.0/4294967296.0,1,-nbitq), 
to_sfixed(324852528.0/4294967296.0,1,-nbitq), 
to_sfixed(-548161284.0/4294967296.0,1,-nbitq), 
to_sfixed(344947090.0/4294967296.0,1,-nbitq), 
to_sfixed(148621717.0/4294967296.0,1,-nbitq), 
to_sfixed(-234595523.0/4294967296.0,1,-nbitq), 
to_sfixed(-206218117.0/4294967296.0,1,-nbitq), 
to_sfixed(-892688282.0/4294967296.0,1,-nbitq), 
to_sfixed(62170390.0/4294967296.0,1,-nbitq), 
to_sfixed(-374213862.0/4294967296.0,1,-nbitq), 
to_sfixed(-510873822.0/4294967296.0,1,-nbitq), 
to_sfixed(419823544.0/4294967296.0,1,-nbitq), 
to_sfixed(-722190330.0/4294967296.0,1,-nbitq), 
to_sfixed(312798670.0/4294967296.0,1,-nbitq), 
to_sfixed(225198408.0/4294967296.0,1,-nbitq), 
to_sfixed(-821305177.0/4294967296.0,1,-nbitq), 
to_sfixed(-591763196.0/4294967296.0,1,-nbitq), 
to_sfixed(16021618.0/4294967296.0,1,-nbitq), 
to_sfixed(-586728678.0/4294967296.0,1,-nbitq), 
to_sfixed(-436743.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-136688930.0/4294967296.0,1,-nbitq), 
to_sfixed(2256401281.0/4294967296.0,1,-nbitq), 
to_sfixed(-1138108617.0/4294967296.0,1,-nbitq), 
to_sfixed(-310275918.0/4294967296.0,1,-nbitq), 
to_sfixed(454760254.0/4294967296.0,1,-nbitq), 
to_sfixed(-70208157.0/4294967296.0,1,-nbitq), 
to_sfixed(-226107864.0/4294967296.0,1,-nbitq), 
to_sfixed(29670988.0/4294967296.0,1,-nbitq), 
to_sfixed(-955232233.0/4294967296.0,1,-nbitq), 
to_sfixed(103173056.0/4294967296.0,1,-nbitq), 
to_sfixed(-825678963.0/4294967296.0,1,-nbitq), 
to_sfixed(-786179825.0/4294967296.0,1,-nbitq), 
to_sfixed(605407343.0/4294967296.0,1,-nbitq), 
to_sfixed(949876313.0/4294967296.0,1,-nbitq), 
to_sfixed(242666819.0/4294967296.0,1,-nbitq), 
to_sfixed(67276154.0/4294967296.0,1,-nbitq), 
to_sfixed(-108928334.0/4294967296.0,1,-nbitq), 
to_sfixed(-177810806.0/4294967296.0,1,-nbitq), 
to_sfixed(658628965.0/4294967296.0,1,-nbitq), 
to_sfixed(23579239.0/4294967296.0,1,-nbitq), 
to_sfixed(-326740542.0/4294967296.0,1,-nbitq), 
to_sfixed(-873919147.0/4294967296.0,1,-nbitq), 
to_sfixed(945206446.0/4294967296.0,1,-nbitq), 
to_sfixed(-20801755.0/4294967296.0,1,-nbitq), 
to_sfixed(131890726.0/4294967296.0,1,-nbitq), 
to_sfixed(-349341466.0/4294967296.0,1,-nbitq), 
to_sfixed(66247676.0/4294967296.0,1,-nbitq), 
to_sfixed(-802383699.0/4294967296.0,1,-nbitq), 
to_sfixed(654084755.0/4294967296.0,1,-nbitq), 
to_sfixed(-233937359.0/4294967296.0,1,-nbitq), 
to_sfixed(-590000120.0/4294967296.0,1,-nbitq), 
to_sfixed(790652684.0/4294967296.0,1,-nbitq), 
to_sfixed(162884942.0/4294967296.0,1,-nbitq), 
to_sfixed(1067447437.0/4294967296.0,1,-nbitq), 
to_sfixed(-199483796.0/4294967296.0,1,-nbitq), 
to_sfixed(-332313039.0/4294967296.0,1,-nbitq), 
to_sfixed(-607763264.0/4294967296.0,1,-nbitq), 
to_sfixed(229014291.0/4294967296.0,1,-nbitq), 
to_sfixed(-482491216.0/4294967296.0,1,-nbitq), 
to_sfixed(-55683829.0/4294967296.0,1,-nbitq), 
to_sfixed(-827694960.0/4294967296.0,1,-nbitq), 
to_sfixed(362397341.0/4294967296.0,1,-nbitq), 
to_sfixed(-536553488.0/4294967296.0,1,-nbitq), 
to_sfixed(-261658155.0/4294967296.0,1,-nbitq), 
to_sfixed(-457531486.0/4294967296.0,1,-nbitq), 
to_sfixed(387225984.0/4294967296.0,1,-nbitq), 
to_sfixed(-255170514.0/4294967296.0,1,-nbitq), 
to_sfixed(1463662591.0/4294967296.0,1,-nbitq), 
to_sfixed(505684729.0/4294967296.0,1,-nbitq), 
to_sfixed(644490814.0/4294967296.0,1,-nbitq), 
to_sfixed(-351984567.0/4294967296.0,1,-nbitq), 
to_sfixed(-568226000.0/4294967296.0,1,-nbitq), 
to_sfixed(301217714.0/4294967296.0,1,-nbitq), 
to_sfixed(-1169994995.0/4294967296.0,1,-nbitq), 
to_sfixed(273314851.0/4294967296.0,1,-nbitq), 
to_sfixed(-1085417329.0/4294967296.0,1,-nbitq), 
to_sfixed(-289548860.0/4294967296.0,1,-nbitq), 
to_sfixed(-35416197.0/4294967296.0,1,-nbitq), 
to_sfixed(-50874462.0/4294967296.0,1,-nbitq), 
to_sfixed(158242703.0/4294967296.0,1,-nbitq), 
to_sfixed(357892792.0/4294967296.0,1,-nbitq), 
to_sfixed(548945650.0/4294967296.0,1,-nbitq), 
to_sfixed(-556591497.0/4294967296.0,1,-nbitq), 
to_sfixed(347454505.0/4294967296.0,1,-nbitq), 
to_sfixed(165293135.0/4294967296.0,1,-nbitq), 
to_sfixed(-511145595.0/4294967296.0,1,-nbitq), 
to_sfixed(-1401708837.0/4294967296.0,1,-nbitq), 
to_sfixed(-368515723.0/4294967296.0,1,-nbitq), 
to_sfixed(-55183766.0/4294967296.0,1,-nbitq), 
to_sfixed(-132027875.0/4294967296.0,1,-nbitq), 
to_sfixed(-388910416.0/4294967296.0,1,-nbitq), 
to_sfixed(-223066691.0/4294967296.0,1,-nbitq), 
to_sfixed(-1493976299.0/4294967296.0,1,-nbitq), 
to_sfixed(-152384322.0/4294967296.0,1,-nbitq), 
to_sfixed(-181322916.0/4294967296.0,1,-nbitq), 
to_sfixed(84080960.0/4294967296.0,1,-nbitq), 
to_sfixed(-226824060.0/4294967296.0,1,-nbitq), 
to_sfixed(149241253.0/4294967296.0,1,-nbitq), 
to_sfixed(-116051875.0/4294967296.0,1,-nbitq), 
to_sfixed(216478607.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(200995399.0/4294967296.0,1,-nbitq), 
to_sfixed(1569357949.0/4294967296.0,1,-nbitq), 
to_sfixed(-393469805.0/4294967296.0,1,-nbitq), 
to_sfixed(-699831710.0/4294967296.0,1,-nbitq), 
to_sfixed(120467136.0/4294967296.0,1,-nbitq), 
to_sfixed(139874262.0/4294967296.0,1,-nbitq), 
to_sfixed(-327211238.0/4294967296.0,1,-nbitq), 
to_sfixed(-397880814.0/4294967296.0,1,-nbitq), 
to_sfixed(-883079606.0/4294967296.0,1,-nbitq), 
to_sfixed(230924142.0/4294967296.0,1,-nbitq), 
to_sfixed(-1036144172.0/4294967296.0,1,-nbitq), 
to_sfixed(-49164995.0/4294967296.0,1,-nbitq), 
to_sfixed(97462100.0/4294967296.0,1,-nbitq), 
to_sfixed(-16804637.0/4294967296.0,1,-nbitq), 
to_sfixed(-279467936.0/4294967296.0,1,-nbitq), 
to_sfixed(-131796431.0/4294967296.0,1,-nbitq), 
to_sfixed(66801950.0/4294967296.0,1,-nbitq), 
to_sfixed(442341189.0/4294967296.0,1,-nbitq), 
to_sfixed(441955488.0/4294967296.0,1,-nbitq), 
to_sfixed(-79703285.0/4294967296.0,1,-nbitq), 
to_sfixed(173109268.0/4294967296.0,1,-nbitq), 
to_sfixed(-557643781.0/4294967296.0,1,-nbitq), 
to_sfixed(367933276.0/4294967296.0,1,-nbitq), 
to_sfixed(-204015434.0/4294967296.0,1,-nbitq), 
to_sfixed(340072876.0/4294967296.0,1,-nbitq), 
to_sfixed(-309112228.0/4294967296.0,1,-nbitq), 
to_sfixed(-758687762.0/4294967296.0,1,-nbitq), 
to_sfixed(-5896691.0/4294967296.0,1,-nbitq), 
to_sfixed(97267725.0/4294967296.0,1,-nbitq), 
to_sfixed(-315625521.0/4294967296.0,1,-nbitq), 
to_sfixed(-1311411015.0/4294967296.0,1,-nbitq), 
to_sfixed(460979922.0/4294967296.0,1,-nbitq), 
to_sfixed(500172392.0/4294967296.0,1,-nbitq), 
to_sfixed(213079265.0/4294967296.0,1,-nbitq), 
to_sfixed(71757761.0/4294967296.0,1,-nbitq), 
to_sfixed(-645935590.0/4294967296.0,1,-nbitq), 
to_sfixed(-36447498.0/4294967296.0,1,-nbitq), 
to_sfixed(301988852.0/4294967296.0,1,-nbitq), 
to_sfixed(300038722.0/4294967296.0,1,-nbitq), 
to_sfixed(-150341753.0/4294967296.0,1,-nbitq), 
to_sfixed(-642866247.0/4294967296.0,1,-nbitq), 
to_sfixed(942423235.0/4294967296.0,1,-nbitq), 
to_sfixed(-290770674.0/4294967296.0,1,-nbitq), 
to_sfixed(-82137888.0/4294967296.0,1,-nbitq), 
to_sfixed(-722007781.0/4294967296.0,1,-nbitq), 
to_sfixed(940800997.0/4294967296.0,1,-nbitq), 
to_sfixed(61605002.0/4294967296.0,1,-nbitq), 
to_sfixed(698027530.0/4294967296.0,1,-nbitq), 
to_sfixed(184363037.0/4294967296.0,1,-nbitq), 
to_sfixed(102107872.0/4294967296.0,1,-nbitq), 
to_sfixed(20408289.0/4294967296.0,1,-nbitq), 
to_sfixed(-543371509.0/4294967296.0,1,-nbitq), 
to_sfixed(-224881914.0/4294967296.0,1,-nbitq), 
to_sfixed(-1001880315.0/4294967296.0,1,-nbitq), 
to_sfixed(-420702297.0/4294967296.0,1,-nbitq), 
to_sfixed(-834755479.0/4294967296.0,1,-nbitq), 
to_sfixed(491083448.0/4294967296.0,1,-nbitq), 
to_sfixed(213323285.0/4294967296.0,1,-nbitq), 
to_sfixed(-36573071.0/4294967296.0,1,-nbitq), 
to_sfixed(-54664834.0/4294967296.0,1,-nbitq), 
to_sfixed(20546169.0/4294967296.0,1,-nbitq), 
to_sfixed(726798392.0/4294967296.0,1,-nbitq), 
to_sfixed(-115952625.0/4294967296.0,1,-nbitq), 
to_sfixed(-833246660.0/4294967296.0,1,-nbitq), 
to_sfixed(384873676.0/4294967296.0,1,-nbitq), 
to_sfixed(-398152992.0/4294967296.0,1,-nbitq), 
to_sfixed(-1267940492.0/4294967296.0,1,-nbitq), 
to_sfixed(-998310059.0/4294967296.0,1,-nbitq), 
to_sfixed(283531774.0/4294967296.0,1,-nbitq), 
to_sfixed(-1119223193.0/4294967296.0,1,-nbitq), 
to_sfixed(-156510739.0/4294967296.0,1,-nbitq), 
to_sfixed(-339074197.0/4294967296.0,1,-nbitq), 
to_sfixed(-1168910541.0/4294967296.0,1,-nbitq), 
to_sfixed(230406888.0/4294967296.0,1,-nbitq), 
to_sfixed(129118510.0/4294967296.0,1,-nbitq), 
to_sfixed(1470784783.0/4294967296.0,1,-nbitq), 
to_sfixed(-177973725.0/4294967296.0,1,-nbitq), 
to_sfixed(22354581.0/4294967296.0,1,-nbitq), 
to_sfixed(-40341705.0/4294967296.0,1,-nbitq), 
to_sfixed(-397117536.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(121058661.0/4294967296.0,1,-nbitq), 
to_sfixed(817903185.0/4294967296.0,1,-nbitq), 
to_sfixed(-1294727871.0/4294967296.0,1,-nbitq), 
to_sfixed(-837073140.0/4294967296.0,1,-nbitq), 
to_sfixed(232321718.0/4294967296.0,1,-nbitq), 
to_sfixed(-628442825.0/4294967296.0,1,-nbitq), 
to_sfixed(169238595.0/4294967296.0,1,-nbitq), 
to_sfixed(-94438738.0/4294967296.0,1,-nbitq), 
to_sfixed(-383305912.0/4294967296.0,1,-nbitq), 
to_sfixed(-314449479.0/4294967296.0,1,-nbitq), 
to_sfixed(-703635136.0/4294967296.0,1,-nbitq), 
to_sfixed(-45699257.0/4294967296.0,1,-nbitq), 
to_sfixed(-265308452.0/4294967296.0,1,-nbitq), 
to_sfixed(-692737661.0/4294967296.0,1,-nbitq), 
to_sfixed(-209984242.0/4294967296.0,1,-nbitq), 
to_sfixed(-134052198.0/4294967296.0,1,-nbitq), 
to_sfixed(118483307.0/4294967296.0,1,-nbitq), 
to_sfixed(19364354.0/4294967296.0,1,-nbitq), 
to_sfixed(373211022.0/4294967296.0,1,-nbitq), 
to_sfixed(-373142290.0/4294967296.0,1,-nbitq), 
to_sfixed(-380330089.0/4294967296.0,1,-nbitq), 
to_sfixed(-561516227.0/4294967296.0,1,-nbitq), 
to_sfixed(88274988.0/4294967296.0,1,-nbitq), 
to_sfixed(-287109521.0/4294967296.0,1,-nbitq), 
to_sfixed(357906854.0/4294967296.0,1,-nbitq), 
to_sfixed(-476329118.0/4294967296.0,1,-nbitq), 
to_sfixed(-49552525.0/4294967296.0,1,-nbitq), 
to_sfixed(413214432.0/4294967296.0,1,-nbitq), 
to_sfixed(-521612781.0/4294967296.0,1,-nbitq), 
to_sfixed(-292043953.0/4294967296.0,1,-nbitq), 
to_sfixed(-1163249903.0/4294967296.0,1,-nbitq), 
to_sfixed(838076959.0/4294967296.0,1,-nbitq), 
to_sfixed(-26978298.0/4294967296.0,1,-nbitq), 
to_sfixed(351223774.0/4294967296.0,1,-nbitq), 
to_sfixed(339277112.0/4294967296.0,1,-nbitq), 
to_sfixed(-68257856.0/4294967296.0,1,-nbitq), 
to_sfixed(120728145.0/4294967296.0,1,-nbitq), 
to_sfixed(220769381.0/4294967296.0,1,-nbitq), 
to_sfixed(325732601.0/4294967296.0,1,-nbitq), 
to_sfixed(-41133342.0/4294967296.0,1,-nbitq), 
to_sfixed(-171755666.0/4294967296.0,1,-nbitq), 
to_sfixed(663375938.0/4294967296.0,1,-nbitq), 
to_sfixed(-958162963.0/4294967296.0,1,-nbitq), 
to_sfixed(-1330896126.0/4294967296.0,1,-nbitq), 
to_sfixed(-654880322.0/4294967296.0,1,-nbitq), 
to_sfixed(-63105790.0/4294967296.0,1,-nbitq), 
to_sfixed(-318732161.0/4294967296.0,1,-nbitq), 
to_sfixed(695748458.0/4294967296.0,1,-nbitq), 
to_sfixed(237580741.0/4294967296.0,1,-nbitq), 
to_sfixed(723967026.0/4294967296.0,1,-nbitq), 
to_sfixed(537574812.0/4294967296.0,1,-nbitq), 
to_sfixed(-144480954.0/4294967296.0,1,-nbitq), 
to_sfixed(-171190595.0/4294967296.0,1,-nbitq), 
to_sfixed(-443027787.0/4294967296.0,1,-nbitq), 
to_sfixed(-1295182157.0/4294967296.0,1,-nbitq), 
to_sfixed(-202989189.0/4294967296.0,1,-nbitq), 
to_sfixed(566496558.0/4294967296.0,1,-nbitq), 
to_sfixed(173684638.0/4294967296.0,1,-nbitq), 
to_sfixed(161436434.0/4294967296.0,1,-nbitq), 
to_sfixed(-274287124.0/4294967296.0,1,-nbitq), 
to_sfixed(50880260.0/4294967296.0,1,-nbitq), 
to_sfixed(480337419.0/4294967296.0,1,-nbitq), 
to_sfixed(-133251611.0/4294967296.0,1,-nbitq), 
to_sfixed(-963185203.0/4294967296.0,1,-nbitq), 
to_sfixed(-207085458.0/4294967296.0,1,-nbitq), 
to_sfixed(-138500849.0/4294967296.0,1,-nbitq), 
to_sfixed(-1174250642.0/4294967296.0,1,-nbitq), 
to_sfixed(-850108377.0/4294967296.0,1,-nbitq), 
to_sfixed(193105843.0/4294967296.0,1,-nbitq), 
to_sfixed(102880663.0/4294967296.0,1,-nbitq), 
to_sfixed(-341457748.0/4294967296.0,1,-nbitq), 
to_sfixed(137789533.0/4294967296.0,1,-nbitq), 
to_sfixed(-174299354.0/4294967296.0,1,-nbitq), 
to_sfixed(-263908286.0/4294967296.0,1,-nbitq), 
to_sfixed(322915280.0/4294967296.0,1,-nbitq), 
to_sfixed(1305115767.0/4294967296.0,1,-nbitq), 
to_sfixed(-733991796.0/4294967296.0,1,-nbitq), 
to_sfixed(480246715.0/4294967296.0,1,-nbitq), 
to_sfixed(123480458.0/4294967296.0,1,-nbitq), 
to_sfixed(94065460.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-413721510.0/4294967296.0,1,-nbitq), 
to_sfixed(805215098.0/4294967296.0,1,-nbitq), 
to_sfixed(-1736330543.0/4294967296.0,1,-nbitq), 
to_sfixed(-1399792264.0/4294967296.0,1,-nbitq), 
to_sfixed(-17549519.0/4294967296.0,1,-nbitq), 
to_sfixed(-186805525.0/4294967296.0,1,-nbitq), 
to_sfixed(-310410369.0/4294967296.0,1,-nbitq), 
to_sfixed(-1837296.0/4294967296.0,1,-nbitq), 
to_sfixed(-1060392258.0/4294967296.0,1,-nbitq), 
to_sfixed(-123545009.0/4294967296.0,1,-nbitq), 
to_sfixed(-181445180.0/4294967296.0,1,-nbitq), 
to_sfixed(1163039014.0/4294967296.0,1,-nbitq), 
to_sfixed(297785764.0/4294967296.0,1,-nbitq), 
to_sfixed(-977469939.0/4294967296.0,1,-nbitq), 
to_sfixed(87498953.0/4294967296.0,1,-nbitq), 
to_sfixed(-201383988.0/4294967296.0,1,-nbitq), 
to_sfixed(-112908189.0/4294967296.0,1,-nbitq), 
to_sfixed(63023370.0/4294967296.0,1,-nbitq), 
to_sfixed(430628317.0/4294967296.0,1,-nbitq), 
to_sfixed(82187208.0/4294967296.0,1,-nbitq), 
to_sfixed(216834708.0/4294967296.0,1,-nbitq), 
to_sfixed(-21907840.0/4294967296.0,1,-nbitq), 
to_sfixed(-322799263.0/4294967296.0,1,-nbitq), 
to_sfixed(-190951133.0/4294967296.0,1,-nbitq), 
to_sfixed(366004053.0/4294967296.0,1,-nbitq), 
to_sfixed(497334213.0/4294967296.0,1,-nbitq), 
to_sfixed(-119793070.0/4294967296.0,1,-nbitq), 
to_sfixed(899179139.0/4294967296.0,1,-nbitq), 
to_sfixed(-174743140.0/4294967296.0,1,-nbitq), 
to_sfixed(-812320696.0/4294967296.0,1,-nbitq), 
to_sfixed(737235935.0/4294967296.0,1,-nbitq), 
to_sfixed(914824271.0/4294967296.0,1,-nbitq), 
to_sfixed(-699417.0/4294967296.0,1,-nbitq), 
to_sfixed(349660027.0/4294967296.0,1,-nbitq), 
to_sfixed(485521603.0/4294967296.0,1,-nbitq), 
to_sfixed(451597033.0/4294967296.0,1,-nbitq), 
to_sfixed(-75185718.0/4294967296.0,1,-nbitq), 
to_sfixed(106088234.0/4294967296.0,1,-nbitq), 
to_sfixed(-76353019.0/4294967296.0,1,-nbitq), 
to_sfixed(11369193.0/4294967296.0,1,-nbitq), 
to_sfixed(68365036.0/4294967296.0,1,-nbitq), 
to_sfixed(258469494.0/4294967296.0,1,-nbitq), 
to_sfixed(-869346112.0/4294967296.0,1,-nbitq), 
to_sfixed(-708911628.0/4294967296.0,1,-nbitq), 
to_sfixed(-29969744.0/4294967296.0,1,-nbitq), 
to_sfixed(-507345063.0/4294967296.0,1,-nbitq), 
to_sfixed(-109033748.0/4294967296.0,1,-nbitq), 
to_sfixed(758462638.0/4294967296.0,1,-nbitq), 
to_sfixed(51451840.0/4294967296.0,1,-nbitq), 
to_sfixed(128274271.0/4294967296.0,1,-nbitq), 
to_sfixed(-226805728.0/4294967296.0,1,-nbitq), 
to_sfixed(137900892.0/4294967296.0,1,-nbitq), 
to_sfixed(-261456001.0/4294967296.0,1,-nbitq), 
to_sfixed(635485918.0/4294967296.0,1,-nbitq), 
to_sfixed(-839663073.0/4294967296.0,1,-nbitq), 
to_sfixed(505027786.0/4294967296.0,1,-nbitq), 
to_sfixed(457784194.0/4294967296.0,1,-nbitq), 
to_sfixed(6544513.0/4294967296.0,1,-nbitq), 
to_sfixed(-343621108.0/4294967296.0,1,-nbitq), 
to_sfixed(-48999602.0/4294967296.0,1,-nbitq), 
to_sfixed(-26697262.0/4294967296.0,1,-nbitq), 
to_sfixed(-398786880.0/4294967296.0,1,-nbitq), 
to_sfixed(-77157933.0/4294967296.0,1,-nbitq), 
to_sfixed(-1137465461.0/4294967296.0,1,-nbitq), 
to_sfixed(330063197.0/4294967296.0,1,-nbitq), 
to_sfixed(-33588201.0/4294967296.0,1,-nbitq), 
to_sfixed(-232209058.0/4294967296.0,1,-nbitq), 
to_sfixed(-357571104.0/4294967296.0,1,-nbitq), 
to_sfixed(-281210786.0/4294967296.0,1,-nbitq), 
to_sfixed(874526566.0/4294967296.0,1,-nbitq), 
to_sfixed(-15911933.0/4294967296.0,1,-nbitq), 
to_sfixed(395908811.0/4294967296.0,1,-nbitq), 
to_sfixed(-301115702.0/4294967296.0,1,-nbitq), 
to_sfixed(80275497.0/4294967296.0,1,-nbitq), 
to_sfixed(362465125.0/4294967296.0,1,-nbitq), 
to_sfixed(741809968.0/4294967296.0,1,-nbitq), 
to_sfixed(-1481377368.0/4294967296.0,1,-nbitq), 
to_sfixed(-262865294.0/4294967296.0,1,-nbitq), 
to_sfixed(-400988576.0/4294967296.0,1,-nbitq), 
to_sfixed(23973713.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-471848511.0/4294967296.0,1,-nbitq), 
to_sfixed(1218623495.0/4294967296.0,1,-nbitq), 
to_sfixed(-1816109772.0/4294967296.0,1,-nbitq), 
to_sfixed(-1892316191.0/4294967296.0,1,-nbitq), 
to_sfixed(-466419106.0/4294967296.0,1,-nbitq), 
to_sfixed(-373660608.0/4294967296.0,1,-nbitq), 
to_sfixed(-341813653.0/4294967296.0,1,-nbitq), 
to_sfixed(538155775.0/4294967296.0,1,-nbitq), 
to_sfixed(-1013129052.0/4294967296.0,1,-nbitq), 
to_sfixed(-199262530.0/4294967296.0,1,-nbitq), 
to_sfixed(86980262.0/4294967296.0,1,-nbitq), 
to_sfixed(213735978.0/4294967296.0,1,-nbitq), 
to_sfixed(277385425.0/4294967296.0,1,-nbitq), 
to_sfixed(-720305390.0/4294967296.0,1,-nbitq), 
to_sfixed(243432717.0/4294967296.0,1,-nbitq), 
to_sfixed(-253016140.0/4294967296.0,1,-nbitq), 
to_sfixed(-70874640.0/4294967296.0,1,-nbitq), 
to_sfixed(95478729.0/4294967296.0,1,-nbitq), 
to_sfixed(422037714.0/4294967296.0,1,-nbitq), 
to_sfixed(-145869381.0/4294967296.0,1,-nbitq), 
to_sfixed(334115441.0/4294967296.0,1,-nbitq), 
to_sfixed(193909746.0/4294967296.0,1,-nbitq), 
to_sfixed(-349741397.0/4294967296.0,1,-nbitq), 
to_sfixed(-1102229100.0/4294967296.0,1,-nbitq), 
to_sfixed(-254739467.0/4294967296.0,1,-nbitq), 
to_sfixed(-415113676.0/4294967296.0,1,-nbitq), 
to_sfixed(-157173234.0/4294967296.0,1,-nbitq), 
to_sfixed(253712754.0/4294967296.0,1,-nbitq), 
to_sfixed(-193079030.0/4294967296.0,1,-nbitq), 
to_sfixed(-756345829.0/4294967296.0,1,-nbitq), 
to_sfixed(919118181.0/4294967296.0,1,-nbitq), 
to_sfixed(627648339.0/4294967296.0,1,-nbitq), 
to_sfixed(-486765251.0/4294967296.0,1,-nbitq), 
to_sfixed(801393897.0/4294967296.0,1,-nbitq), 
to_sfixed(-93299137.0/4294967296.0,1,-nbitq), 
to_sfixed(594445582.0/4294967296.0,1,-nbitq), 
to_sfixed(27270666.0/4294967296.0,1,-nbitq), 
to_sfixed(-354330513.0/4294967296.0,1,-nbitq), 
to_sfixed(-11269638.0/4294967296.0,1,-nbitq), 
to_sfixed(353461642.0/4294967296.0,1,-nbitq), 
to_sfixed(-206425581.0/4294967296.0,1,-nbitq), 
to_sfixed(-33027750.0/4294967296.0,1,-nbitq), 
to_sfixed(-330412946.0/4294967296.0,1,-nbitq), 
to_sfixed(-334356371.0/4294967296.0,1,-nbitq), 
to_sfixed(-828141488.0/4294967296.0,1,-nbitq), 
to_sfixed(10618655.0/4294967296.0,1,-nbitq), 
to_sfixed(-226096554.0/4294967296.0,1,-nbitq), 
to_sfixed(357721649.0/4294967296.0,1,-nbitq), 
to_sfixed(-560685557.0/4294967296.0,1,-nbitq), 
to_sfixed(624674190.0/4294967296.0,1,-nbitq), 
to_sfixed(-92031923.0/4294967296.0,1,-nbitq), 
to_sfixed(-701930792.0/4294967296.0,1,-nbitq), 
to_sfixed(-285402754.0/4294967296.0,1,-nbitq), 
to_sfixed(133245098.0/4294967296.0,1,-nbitq), 
to_sfixed(-781387607.0/4294967296.0,1,-nbitq), 
to_sfixed(157130664.0/4294967296.0,1,-nbitq), 
to_sfixed(1004891276.0/4294967296.0,1,-nbitq), 
to_sfixed(-233801482.0/4294967296.0,1,-nbitq), 
to_sfixed(204451690.0/4294967296.0,1,-nbitq), 
to_sfixed(-225125619.0/4294967296.0,1,-nbitq), 
to_sfixed(-507941016.0/4294967296.0,1,-nbitq), 
to_sfixed(-640258847.0/4294967296.0,1,-nbitq), 
to_sfixed(-170794697.0/4294967296.0,1,-nbitq), 
to_sfixed(-670583145.0/4294967296.0,1,-nbitq), 
to_sfixed(-56599721.0/4294967296.0,1,-nbitq), 
to_sfixed(100321003.0/4294967296.0,1,-nbitq), 
to_sfixed(-251129237.0/4294967296.0,1,-nbitq), 
to_sfixed(-46829182.0/4294967296.0,1,-nbitq), 
to_sfixed(160761293.0/4294967296.0,1,-nbitq), 
to_sfixed(931474301.0/4294967296.0,1,-nbitq), 
to_sfixed(-367587220.0/4294967296.0,1,-nbitq), 
to_sfixed(-50546781.0/4294967296.0,1,-nbitq), 
to_sfixed(23619704.0/4294967296.0,1,-nbitq), 
to_sfixed(157148181.0/4294967296.0,1,-nbitq), 
to_sfixed(-112936565.0/4294967296.0,1,-nbitq), 
to_sfixed(459259424.0/4294967296.0,1,-nbitq), 
to_sfixed(-474436273.0/4294967296.0,1,-nbitq), 
to_sfixed(342609614.0/4294967296.0,1,-nbitq), 
to_sfixed(-158339830.0/4294967296.0,1,-nbitq), 
to_sfixed(87966201.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-498353203.0/4294967296.0,1,-nbitq), 
to_sfixed(1496516119.0/4294967296.0,1,-nbitq), 
to_sfixed(-1088610251.0/4294967296.0,1,-nbitq), 
to_sfixed(-1034675960.0/4294967296.0,1,-nbitq), 
to_sfixed(-534552633.0/4294967296.0,1,-nbitq), 
to_sfixed(-325168964.0/4294967296.0,1,-nbitq), 
to_sfixed(-16921277.0/4294967296.0,1,-nbitq), 
to_sfixed(268523549.0/4294967296.0,1,-nbitq), 
to_sfixed(-669360037.0/4294967296.0,1,-nbitq), 
to_sfixed(-85717965.0/4294967296.0,1,-nbitq), 
to_sfixed(435588511.0/4294967296.0,1,-nbitq), 
to_sfixed(553285634.0/4294967296.0,1,-nbitq), 
to_sfixed(776957225.0/4294967296.0,1,-nbitq), 
to_sfixed(-513164828.0/4294967296.0,1,-nbitq), 
to_sfixed(-21053124.0/4294967296.0,1,-nbitq), 
to_sfixed(-257387965.0/4294967296.0,1,-nbitq), 
to_sfixed(-228344220.0/4294967296.0,1,-nbitq), 
to_sfixed(27745925.0/4294967296.0,1,-nbitq), 
to_sfixed(454444619.0/4294967296.0,1,-nbitq), 
to_sfixed(-312024116.0/4294967296.0,1,-nbitq), 
to_sfixed(375570085.0/4294967296.0,1,-nbitq), 
to_sfixed(-15517935.0/4294967296.0,1,-nbitq), 
to_sfixed(17632053.0/4294967296.0,1,-nbitq), 
to_sfixed(-1097612477.0/4294967296.0,1,-nbitq), 
to_sfixed(140871341.0/4294967296.0,1,-nbitq), 
to_sfixed(470128556.0/4294967296.0,1,-nbitq), 
to_sfixed(18549342.0/4294967296.0,1,-nbitq), 
to_sfixed(42589531.0/4294967296.0,1,-nbitq), 
to_sfixed(-170428437.0/4294967296.0,1,-nbitq), 
to_sfixed(-9046120.0/4294967296.0,1,-nbitq), 
to_sfixed(461320312.0/4294967296.0,1,-nbitq), 
to_sfixed(840020162.0/4294967296.0,1,-nbitq), 
to_sfixed(74261399.0/4294967296.0,1,-nbitq), 
to_sfixed(-2532650.0/4294967296.0,1,-nbitq), 
to_sfixed(-534593801.0/4294967296.0,1,-nbitq), 
to_sfixed(210002502.0/4294967296.0,1,-nbitq), 
to_sfixed(-293147818.0/4294967296.0,1,-nbitq), 
to_sfixed(-204094078.0/4294967296.0,1,-nbitq), 
to_sfixed(436167627.0/4294967296.0,1,-nbitq), 
to_sfixed(-158264914.0/4294967296.0,1,-nbitq), 
to_sfixed(-8537826.0/4294967296.0,1,-nbitq), 
to_sfixed(-103447401.0/4294967296.0,1,-nbitq), 
to_sfixed(-186075583.0/4294967296.0,1,-nbitq), 
to_sfixed(-1087497546.0/4294967296.0,1,-nbitq), 
to_sfixed(-652096480.0/4294967296.0,1,-nbitq), 
to_sfixed(-602759245.0/4294967296.0,1,-nbitq), 
to_sfixed(-360618473.0/4294967296.0,1,-nbitq), 
to_sfixed(354704441.0/4294967296.0,1,-nbitq), 
to_sfixed(-744234850.0/4294967296.0,1,-nbitq), 
to_sfixed(-131203042.0/4294967296.0,1,-nbitq), 
to_sfixed(-168110291.0/4294967296.0,1,-nbitq), 
to_sfixed(-363275692.0/4294967296.0,1,-nbitq), 
to_sfixed(-368659066.0/4294967296.0,1,-nbitq), 
to_sfixed(440854105.0/4294967296.0,1,-nbitq), 
to_sfixed(-655614010.0/4294967296.0,1,-nbitq), 
to_sfixed(129096129.0/4294967296.0,1,-nbitq), 
to_sfixed(708947270.0/4294967296.0,1,-nbitq), 
to_sfixed(-221418865.0/4294967296.0,1,-nbitq), 
to_sfixed(-390529778.0/4294967296.0,1,-nbitq), 
to_sfixed(241197264.0/4294967296.0,1,-nbitq), 
to_sfixed(-369264100.0/4294967296.0,1,-nbitq), 
to_sfixed(-887680217.0/4294967296.0,1,-nbitq), 
to_sfixed(-518807393.0/4294967296.0,1,-nbitq), 
to_sfixed(-606444553.0/4294967296.0,1,-nbitq), 
to_sfixed(364024652.0/4294967296.0,1,-nbitq), 
to_sfixed(257836712.0/4294967296.0,1,-nbitq), 
to_sfixed(-106069981.0/4294967296.0,1,-nbitq), 
to_sfixed(-732153991.0/4294967296.0,1,-nbitq), 
to_sfixed(-265074023.0/4294967296.0,1,-nbitq), 
to_sfixed(281811277.0/4294967296.0,1,-nbitq), 
to_sfixed(-208575559.0/4294967296.0,1,-nbitq), 
to_sfixed(275725099.0/4294967296.0,1,-nbitq), 
to_sfixed(457594690.0/4294967296.0,1,-nbitq), 
to_sfixed(415490387.0/4294967296.0,1,-nbitq), 
to_sfixed(-227643314.0/4294967296.0,1,-nbitq), 
to_sfixed(474250454.0/4294967296.0,1,-nbitq), 
to_sfixed(-818349693.0/4294967296.0,1,-nbitq), 
to_sfixed(1690555.0/4294967296.0,1,-nbitq), 
to_sfixed(-102659976.0/4294967296.0,1,-nbitq), 
to_sfixed(-70746797.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-84418724.0/4294967296.0,1,-nbitq), 
to_sfixed(673022806.0/4294967296.0,1,-nbitq), 
to_sfixed(-857546084.0/4294967296.0,1,-nbitq), 
to_sfixed(-780021761.0/4294967296.0,1,-nbitq), 
to_sfixed(-575801462.0/4294967296.0,1,-nbitq), 
to_sfixed(-398743500.0/4294967296.0,1,-nbitq), 
to_sfixed(-273033946.0/4294967296.0,1,-nbitq), 
to_sfixed(576952747.0/4294967296.0,1,-nbitq), 
to_sfixed(-282071153.0/4294967296.0,1,-nbitq), 
to_sfixed(-61497800.0/4294967296.0,1,-nbitq), 
to_sfixed(677556987.0/4294967296.0,1,-nbitq), 
to_sfixed(42408504.0/4294967296.0,1,-nbitq), 
to_sfixed(623861674.0/4294967296.0,1,-nbitq), 
to_sfixed(-442829998.0/4294967296.0,1,-nbitq), 
to_sfixed(7252657.0/4294967296.0,1,-nbitq), 
to_sfixed(-156031563.0/4294967296.0,1,-nbitq), 
to_sfixed(46700716.0/4294967296.0,1,-nbitq), 
to_sfixed(-150581582.0/4294967296.0,1,-nbitq), 
to_sfixed(475359093.0/4294967296.0,1,-nbitq), 
to_sfixed(-28438135.0/4294967296.0,1,-nbitq), 
to_sfixed(-42457369.0/4294967296.0,1,-nbitq), 
to_sfixed(-202462971.0/4294967296.0,1,-nbitq), 
to_sfixed(-167714982.0/4294967296.0,1,-nbitq), 
to_sfixed(-622114340.0/4294967296.0,1,-nbitq), 
to_sfixed(-203703134.0/4294967296.0,1,-nbitq), 
to_sfixed(553511551.0/4294967296.0,1,-nbitq), 
to_sfixed(-205303472.0/4294967296.0,1,-nbitq), 
to_sfixed(254517086.0/4294967296.0,1,-nbitq), 
to_sfixed(-39485394.0/4294967296.0,1,-nbitq), 
to_sfixed(168490654.0/4294967296.0,1,-nbitq), 
to_sfixed(249602113.0/4294967296.0,1,-nbitq), 
to_sfixed(533618009.0/4294967296.0,1,-nbitq), 
to_sfixed(7752720.0/4294967296.0,1,-nbitq), 
to_sfixed(167589904.0/4294967296.0,1,-nbitq), 
to_sfixed(-209269534.0/4294967296.0,1,-nbitq), 
to_sfixed(-62349642.0/4294967296.0,1,-nbitq), 
to_sfixed(-44207915.0/4294967296.0,1,-nbitq), 
to_sfixed(-313190724.0/4294967296.0,1,-nbitq), 
to_sfixed(331238094.0/4294967296.0,1,-nbitq), 
to_sfixed(-228611842.0/4294967296.0,1,-nbitq), 
to_sfixed(-29236785.0/4294967296.0,1,-nbitq), 
to_sfixed(-529085030.0/4294967296.0,1,-nbitq), 
to_sfixed(-393556349.0/4294967296.0,1,-nbitq), 
to_sfixed(-622452334.0/4294967296.0,1,-nbitq), 
to_sfixed(-619693449.0/4294967296.0,1,-nbitq), 
to_sfixed(-435831788.0/4294967296.0,1,-nbitq), 
to_sfixed(-396362342.0/4294967296.0,1,-nbitq), 
to_sfixed(239201209.0/4294967296.0,1,-nbitq), 
to_sfixed(-282132138.0/4294967296.0,1,-nbitq), 
to_sfixed(274726055.0/4294967296.0,1,-nbitq), 
to_sfixed(-272872920.0/4294967296.0,1,-nbitq), 
to_sfixed(-74401625.0/4294967296.0,1,-nbitq), 
to_sfixed(-93927915.0/4294967296.0,1,-nbitq), 
to_sfixed(204749957.0/4294967296.0,1,-nbitq), 
to_sfixed(-158127428.0/4294967296.0,1,-nbitq), 
to_sfixed(20238601.0/4294967296.0,1,-nbitq), 
to_sfixed(303819636.0/4294967296.0,1,-nbitq), 
to_sfixed(-264217078.0/4294967296.0,1,-nbitq), 
to_sfixed(88928292.0/4294967296.0,1,-nbitq), 
to_sfixed(208520806.0/4294967296.0,1,-nbitq), 
to_sfixed(-434073084.0/4294967296.0,1,-nbitq), 
to_sfixed(-581932323.0/4294967296.0,1,-nbitq), 
to_sfixed(531168579.0/4294967296.0,1,-nbitq), 
to_sfixed(-636314953.0/4294967296.0,1,-nbitq), 
to_sfixed(423720940.0/4294967296.0,1,-nbitq), 
to_sfixed(235079914.0/4294967296.0,1,-nbitq), 
to_sfixed(-331118935.0/4294967296.0,1,-nbitq), 
to_sfixed(-503784447.0/4294967296.0,1,-nbitq), 
to_sfixed(-258003418.0/4294967296.0,1,-nbitq), 
to_sfixed(213128189.0/4294967296.0,1,-nbitq), 
to_sfixed(445532304.0/4294967296.0,1,-nbitq), 
to_sfixed(-170884741.0/4294967296.0,1,-nbitq), 
to_sfixed(-32979545.0/4294967296.0,1,-nbitq), 
to_sfixed(219186707.0/4294967296.0,1,-nbitq), 
to_sfixed(250814459.0/4294967296.0,1,-nbitq), 
to_sfixed(382402012.0/4294967296.0,1,-nbitq), 
to_sfixed(-988722120.0/4294967296.0,1,-nbitq), 
to_sfixed(-520389273.0/4294967296.0,1,-nbitq), 
to_sfixed(-569309971.0/4294967296.0,1,-nbitq), 
to_sfixed(-364434914.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-180962894.0/4294967296.0,1,-nbitq), 
to_sfixed(756354269.0/4294967296.0,1,-nbitq), 
to_sfixed(-94952417.0/4294967296.0,1,-nbitq), 
to_sfixed(-225879764.0/4294967296.0,1,-nbitq), 
to_sfixed(-25410383.0/4294967296.0,1,-nbitq), 
to_sfixed(-504302648.0/4294967296.0,1,-nbitq), 
to_sfixed(41290644.0/4294967296.0,1,-nbitq), 
to_sfixed(262106267.0/4294967296.0,1,-nbitq), 
to_sfixed(-690266753.0/4294967296.0,1,-nbitq), 
to_sfixed(295770314.0/4294967296.0,1,-nbitq), 
to_sfixed(761547865.0/4294967296.0,1,-nbitq), 
to_sfixed(123413648.0/4294967296.0,1,-nbitq), 
to_sfixed(459594138.0/4294967296.0,1,-nbitq), 
to_sfixed(-192854091.0/4294967296.0,1,-nbitq), 
to_sfixed(-22416116.0/4294967296.0,1,-nbitq), 
to_sfixed(-405712893.0/4294967296.0,1,-nbitq), 
to_sfixed(379812546.0/4294967296.0,1,-nbitq), 
to_sfixed(-60401616.0/4294967296.0,1,-nbitq), 
to_sfixed(-146371982.0/4294967296.0,1,-nbitq), 
to_sfixed(400641511.0/4294967296.0,1,-nbitq), 
to_sfixed(-105258833.0/4294967296.0,1,-nbitq), 
to_sfixed(-363752757.0/4294967296.0,1,-nbitq), 
to_sfixed(-275730774.0/4294967296.0,1,-nbitq), 
to_sfixed(39596085.0/4294967296.0,1,-nbitq), 
to_sfixed(216847055.0/4294967296.0,1,-nbitq), 
to_sfixed(-300897163.0/4294967296.0,1,-nbitq), 
to_sfixed(-508962045.0/4294967296.0,1,-nbitq), 
to_sfixed(29332820.0/4294967296.0,1,-nbitq), 
to_sfixed(316006471.0/4294967296.0,1,-nbitq), 
to_sfixed(517602893.0/4294967296.0,1,-nbitq), 
to_sfixed(-192871603.0/4294967296.0,1,-nbitq), 
to_sfixed(-163973705.0/4294967296.0,1,-nbitq), 
to_sfixed(495836836.0/4294967296.0,1,-nbitq), 
to_sfixed(-300163541.0/4294967296.0,1,-nbitq), 
to_sfixed(98419917.0/4294967296.0,1,-nbitq), 
to_sfixed(230034590.0/4294967296.0,1,-nbitq), 
to_sfixed(-491572395.0/4294967296.0,1,-nbitq), 
to_sfixed(-177756336.0/4294967296.0,1,-nbitq), 
to_sfixed(247501444.0/4294967296.0,1,-nbitq), 
to_sfixed(42155706.0/4294967296.0,1,-nbitq), 
to_sfixed(-24249377.0/4294967296.0,1,-nbitq), 
to_sfixed(200509204.0/4294967296.0,1,-nbitq), 
to_sfixed(-198226571.0/4294967296.0,1,-nbitq), 
to_sfixed(-327357525.0/4294967296.0,1,-nbitq), 
to_sfixed(-372650240.0/4294967296.0,1,-nbitq), 
to_sfixed(-625173911.0/4294967296.0,1,-nbitq), 
to_sfixed(271279685.0/4294967296.0,1,-nbitq), 
to_sfixed(9599457.0/4294967296.0,1,-nbitq), 
to_sfixed(-489955014.0/4294967296.0,1,-nbitq), 
to_sfixed(-183294496.0/4294967296.0,1,-nbitq), 
to_sfixed(-56179709.0/4294967296.0,1,-nbitq), 
to_sfixed(127735360.0/4294967296.0,1,-nbitq), 
to_sfixed(-215519327.0/4294967296.0,1,-nbitq), 
to_sfixed(-248640445.0/4294967296.0,1,-nbitq), 
to_sfixed(-111049403.0/4294967296.0,1,-nbitq), 
to_sfixed(-593559587.0/4294967296.0,1,-nbitq), 
to_sfixed(-163013065.0/4294967296.0,1,-nbitq), 
to_sfixed(-73604064.0/4294967296.0,1,-nbitq), 
to_sfixed(-284502531.0/4294967296.0,1,-nbitq), 
to_sfixed(10869992.0/4294967296.0,1,-nbitq), 
to_sfixed(-298488578.0/4294967296.0,1,-nbitq), 
to_sfixed(-410967957.0/4294967296.0,1,-nbitq), 
to_sfixed(315089735.0/4294967296.0,1,-nbitq), 
to_sfixed(-44587800.0/4294967296.0,1,-nbitq), 
to_sfixed(-164984511.0/4294967296.0,1,-nbitq), 
to_sfixed(210084052.0/4294967296.0,1,-nbitq), 
to_sfixed(165218784.0/4294967296.0,1,-nbitq), 
to_sfixed(235572277.0/4294967296.0,1,-nbitq), 
to_sfixed(76314741.0/4294967296.0,1,-nbitq), 
to_sfixed(276549026.0/4294967296.0,1,-nbitq), 
to_sfixed(-102360065.0/4294967296.0,1,-nbitq), 
to_sfixed(-346794819.0/4294967296.0,1,-nbitq), 
to_sfixed(639215664.0/4294967296.0,1,-nbitq), 
to_sfixed(-19632399.0/4294967296.0,1,-nbitq), 
to_sfixed(-101613440.0/4294967296.0,1,-nbitq), 
to_sfixed(255022434.0/4294967296.0,1,-nbitq), 
to_sfixed(-676541371.0/4294967296.0,1,-nbitq), 
to_sfixed(-483476205.0/4294967296.0,1,-nbitq), 
to_sfixed(-490585772.0/4294967296.0,1,-nbitq), 
to_sfixed(-114225891.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-213123270.0/4294967296.0,1,-nbitq), 
to_sfixed(-39327258.0/4294967296.0,1,-nbitq), 
to_sfixed(-269181580.0/4294967296.0,1,-nbitq), 
to_sfixed(-289382630.0/4294967296.0,1,-nbitq), 
to_sfixed(-70685748.0/4294967296.0,1,-nbitq), 
to_sfixed(-122713747.0/4294967296.0,1,-nbitq), 
to_sfixed(-38328978.0/4294967296.0,1,-nbitq), 
to_sfixed(233754571.0/4294967296.0,1,-nbitq), 
to_sfixed(-5753662.0/4294967296.0,1,-nbitq), 
to_sfixed(-13940963.0/4294967296.0,1,-nbitq), 
to_sfixed(-27413231.0/4294967296.0,1,-nbitq), 
to_sfixed(199923958.0/4294967296.0,1,-nbitq), 
to_sfixed(-230492398.0/4294967296.0,1,-nbitq), 
to_sfixed(-273594545.0/4294967296.0,1,-nbitq), 
to_sfixed(-436898640.0/4294967296.0,1,-nbitq), 
to_sfixed(-508188312.0/4294967296.0,1,-nbitq), 
to_sfixed(-187586167.0/4294967296.0,1,-nbitq), 
to_sfixed(-203693803.0/4294967296.0,1,-nbitq), 
to_sfixed(-94115826.0/4294967296.0,1,-nbitq), 
to_sfixed(-189172144.0/4294967296.0,1,-nbitq), 
to_sfixed(-221206132.0/4294967296.0,1,-nbitq), 
to_sfixed(245907084.0/4294967296.0,1,-nbitq), 
to_sfixed(-344105206.0/4294967296.0,1,-nbitq), 
to_sfixed(178825764.0/4294967296.0,1,-nbitq), 
to_sfixed(363273719.0/4294967296.0,1,-nbitq), 
to_sfixed(-217714882.0/4294967296.0,1,-nbitq), 
to_sfixed(-152075718.0/4294967296.0,1,-nbitq), 
to_sfixed(116547732.0/4294967296.0,1,-nbitq), 
to_sfixed(577019553.0/4294967296.0,1,-nbitq), 
to_sfixed(-334887683.0/4294967296.0,1,-nbitq), 
to_sfixed(-509288221.0/4294967296.0,1,-nbitq), 
to_sfixed(319005522.0/4294967296.0,1,-nbitq), 
to_sfixed(155521997.0/4294967296.0,1,-nbitq), 
to_sfixed(-286914683.0/4294967296.0,1,-nbitq), 
to_sfixed(-391530150.0/4294967296.0,1,-nbitq), 
to_sfixed(217857027.0/4294967296.0,1,-nbitq), 
to_sfixed(11791041.0/4294967296.0,1,-nbitq), 
to_sfixed(-440508669.0/4294967296.0,1,-nbitq), 
to_sfixed(267037898.0/4294967296.0,1,-nbitq), 
to_sfixed(3823234.0/4294967296.0,1,-nbitq), 
to_sfixed(446642029.0/4294967296.0,1,-nbitq), 
to_sfixed(288183528.0/4294967296.0,1,-nbitq), 
to_sfixed(-74705745.0/4294967296.0,1,-nbitq), 
to_sfixed(-547643996.0/4294967296.0,1,-nbitq), 
to_sfixed(313417133.0/4294967296.0,1,-nbitq), 
to_sfixed(-467106957.0/4294967296.0,1,-nbitq), 
to_sfixed(-411816566.0/4294967296.0,1,-nbitq), 
to_sfixed(-206259840.0/4294967296.0,1,-nbitq), 
to_sfixed(220221569.0/4294967296.0,1,-nbitq), 
to_sfixed(-457211802.0/4294967296.0,1,-nbitq), 
to_sfixed(51035780.0/4294967296.0,1,-nbitq), 
to_sfixed(-220594155.0/4294967296.0,1,-nbitq), 
to_sfixed(-123126893.0/4294967296.0,1,-nbitq), 
to_sfixed(190258259.0/4294967296.0,1,-nbitq), 
to_sfixed(146388002.0/4294967296.0,1,-nbitq), 
to_sfixed(178027955.0/4294967296.0,1,-nbitq), 
to_sfixed(-93079010.0/4294967296.0,1,-nbitq), 
to_sfixed(310331136.0/4294967296.0,1,-nbitq), 
to_sfixed(355912175.0/4294967296.0,1,-nbitq), 
to_sfixed(93645840.0/4294967296.0,1,-nbitq), 
to_sfixed(278789311.0/4294967296.0,1,-nbitq), 
to_sfixed(-335815222.0/4294967296.0,1,-nbitq), 
to_sfixed(-61461443.0/4294967296.0,1,-nbitq), 
to_sfixed(-163865108.0/4294967296.0,1,-nbitq), 
to_sfixed(318804286.0/4294967296.0,1,-nbitq), 
to_sfixed(-93965875.0/4294967296.0,1,-nbitq), 
to_sfixed(783424994.0/4294967296.0,1,-nbitq), 
to_sfixed(360679903.0/4294967296.0,1,-nbitq), 
to_sfixed(112660578.0/4294967296.0,1,-nbitq), 
to_sfixed(336017084.0/4294967296.0,1,-nbitq), 
to_sfixed(272107737.0/4294967296.0,1,-nbitq), 
to_sfixed(214433426.0/4294967296.0,1,-nbitq), 
to_sfixed(-215855966.0/4294967296.0,1,-nbitq), 
to_sfixed(262204281.0/4294967296.0,1,-nbitq), 
to_sfixed(392863964.0/4294967296.0,1,-nbitq), 
to_sfixed(-119906070.0/4294967296.0,1,-nbitq), 
to_sfixed(-397509752.0/4294967296.0,1,-nbitq), 
to_sfixed(176214038.0/4294967296.0,1,-nbitq), 
to_sfixed(173164912.0/4294967296.0,1,-nbitq), 
to_sfixed(390744309.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(369031006.0/4294967296.0,1,-nbitq), 
to_sfixed(-328108539.0/4294967296.0,1,-nbitq), 
to_sfixed(-357290772.0/4294967296.0,1,-nbitq), 
to_sfixed(-91684655.0/4294967296.0,1,-nbitq), 
to_sfixed(162744411.0/4294967296.0,1,-nbitq), 
to_sfixed(-414178677.0/4294967296.0,1,-nbitq), 
to_sfixed(321911761.0/4294967296.0,1,-nbitq), 
to_sfixed(48887236.0/4294967296.0,1,-nbitq), 
to_sfixed(293558112.0/4294967296.0,1,-nbitq), 
to_sfixed(391667315.0/4294967296.0,1,-nbitq), 
to_sfixed(556777401.0/4294967296.0,1,-nbitq), 
to_sfixed(-47695212.0/4294967296.0,1,-nbitq), 
to_sfixed(286145833.0/4294967296.0,1,-nbitq), 
to_sfixed(138371819.0/4294967296.0,1,-nbitq), 
to_sfixed(-349216966.0/4294967296.0,1,-nbitq), 
to_sfixed(-311748944.0/4294967296.0,1,-nbitq), 
to_sfixed(308159526.0/4294967296.0,1,-nbitq), 
to_sfixed(87547889.0/4294967296.0,1,-nbitq), 
to_sfixed(-294834722.0/4294967296.0,1,-nbitq), 
to_sfixed(-327909862.0/4294967296.0,1,-nbitq), 
to_sfixed(38502865.0/4294967296.0,1,-nbitq), 
to_sfixed(31672866.0/4294967296.0,1,-nbitq), 
to_sfixed(156529387.0/4294967296.0,1,-nbitq), 
to_sfixed(-18397843.0/4294967296.0,1,-nbitq), 
to_sfixed(-166785283.0/4294967296.0,1,-nbitq), 
to_sfixed(461006200.0/4294967296.0,1,-nbitq), 
to_sfixed(-271125643.0/4294967296.0,1,-nbitq), 
to_sfixed(-106740252.0/4294967296.0,1,-nbitq), 
to_sfixed(507262043.0/4294967296.0,1,-nbitq), 
to_sfixed(-36731964.0/4294967296.0,1,-nbitq), 
to_sfixed(8781829.0/4294967296.0,1,-nbitq), 
to_sfixed(-321024905.0/4294967296.0,1,-nbitq), 
to_sfixed(470075887.0/4294967296.0,1,-nbitq), 
to_sfixed(-519722334.0/4294967296.0,1,-nbitq), 
to_sfixed(-92237371.0/4294967296.0,1,-nbitq), 
to_sfixed(-480976372.0/4294967296.0,1,-nbitq), 
to_sfixed(-213595908.0/4294967296.0,1,-nbitq), 
to_sfixed(121329090.0/4294967296.0,1,-nbitq), 
to_sfixed(123055684.0/4294967296.0,1,-nbitq), 
to_sfixed(-54813278.0/4294967296.0,1,-nbitq), 
to_sfixed(222378819.0/4294967296.0,1,-nbitq), 
to_sfixed(-91446686.0/4294967296.0,1,-nbitq), 
to_sfixed(-410278179.0/4294967296.0,1,-nbitq), 
to_sfixed(301706597.0/4294967296.0,1,-nbitq), 
to_sfixed(301684452.0/4294967296.0,1,-nbitq), 
to_sfixed(29912054.0/4294967296.0,1,-nbitq), 
to_sfixed(-109503236.0/4294967296.0,1,-nbitq), 
to_sfixed(120195548.0/4294967296.0,1,-nbitq), 
to_sfixed(-350149888.0/4294967296.0,1,-nbitq), 
to_sfixed(-252565988.0/4294967296.0,1,-nbitq), 
to_sfixed(86392000.0/4294967296.0,1,-nbitq), 
to_sfixed(277416543.0/4294967296.0,1,-nbitq), 
to_sfixed(147374000.0/4294967296.0,1,-nbitq), 
to_sfixed(200709979.0/4294967296.0,1,-nbitq), 
to_sfixed(304659879.0/4294967296.0,1,-nbitq), 
to_sfixed(179517011.0/4294967296.0,1,-nbitq), 
to_sfixed(528905963.0/4294967296.0,1,-nbitq), 
to_sfixed(-243720684.0/4294967296.0,1,-nbitq), 
to_sfixed(-331101824.0/4294967296.0,1,-nbitq), 
to_sfixed(-4741.0/4294967296.0,1,-nbitq), 
to_sfixed(180028163.0/4294967296.0,1,-nbitq), 
to_sfixed(-176157505.0/4294967296.0,1,-nbitq), 
to_sfixed(-295241114.0/4294967296.0,1,-nbitq), 
to_sfixed(-119391226.0/4294967296.0,1,-nbitq), 
to_sfixed(107843291.0/4294967296.0,1,-nbitq), 
to_sfixed(-324434620.0/4294967296.0,1,-nbitq), 
to_sfixed(529673823.0/4294967296.0,1,-nbitq), 
to_sfixed(421714267.0/4294967296.0,1,-nbitq), 
to_sfixed(376286670.0/4294967296.0,1,-nbitq), 
to_sfixed(339842471.0/4294967296.0,1,-nbitq), 
to_sfixed(-427992999.0/4294967296.0,1,-nbitq), 
to_sfixed(351871306.0/4294967296.0,1,-nbitq), 
to_sfixed(357761267.0/4294967296.0,1,-nbitq), 
to_sfixed(108258320.0/4294967296.0,1,-nbitq), 
to_sfixed(433662702.0/4294967296.0,1,-nbitq), 
to_sfixed(-367179233.0/4294967296.0,1,-nbitq), 
to_sfixed(1163892.0/4294967296.0,1,-nbitq), 
to_sfixed(-185606621.0/4294967296.0,1,-nbitq), 
to_sfixed(-85215000.0/4294967296.0,1,-nbitq), 
to_sfixed(328479868.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(380810048.0/4294967296.0,1,-nbitq), 
to_sfixed(-425346505.0/4294967296.0,1,-nbitq), 
to_sfixed(-362094083.0/4294967296.0,1,-nbitq), 
to_sfixed(-120704871.0/4294967296.0,1,-nbitq), 
to_sfixed(79694051.0/4294967296.0,1,-nbitq), 
to_sfixed(216089711.0/4294967296.0,1,-nbitq), 
to_sfixed(-8893137.0/4294967296.0,1,-nbitq), 
to_sfixed(-279651250.0/4294967296.0,1,-nbitq), 
to_sfixed(-73148090.0/4294967296.0,1,-nbitq), 
to_sfixed(-292463699.0/4294967296.0,1,-nbitq), 
to_sfixed(302660184.0/4294967296.0,1,-nbitq), 
to_sfixed(144692062.0/4294967296.0,1,-nbitq), 
to_sfixed(270715540.0/4294967296.0,1,-nbitq), 
to_sfixed(-452426565.0/4294967296.0,1,-nbitq), 
to_sfixed(-427078195.0/4294967296.0,1,-nbitq), 
to_sfixed(10060192.0/4294967296.0,1,-nbitq), 
to_sfixed(390551394.0/4294967296.0,1,-nbitq), 
to_sfixed(297407498.0/4294967296.0,1,-nbitq), 
to_sfixed(381642720.0/4294967296.0,1,-nbitq), 
to_sfixed(-342533973.0/4294967296.0,1,-nbitq), 
to_sfixed(-242881926.0/4294967296.0,1,-nbitq), 
to_sfixed(-201012495.0/4294967296.0,1,-nbitq), 
to_sfixed(-80961425.0/4294967296.0,1,-nbitq), 
to_sfixed(-309636062.0/4294967296.0,1,-nbitq), 
to_sfixed(89078123.0/4294967296.0,1,-nbitq), 
to_sfixed(-92414763.0/4294967296.0,1,-nbitq), 
to_sfixed(385589405.0/4294967296.0,1,-nbitq), 
to_sfixed(-261370107.0/4294967296.0,1,-nbitq), 
to_sfixed(254089991.0/4294967296.0,1,-nbitq), 
to_sfixed(-427956188.0/4294967296.0,1,-nbitq), 
to_sfixed(-420216447.0/4294967296.0,1,-nbitq), 
to_sfixed(-231504132.0/4294967296.0,1,-nbitq), 
to_sfixed(-43366318.0/4294967296.0,1,-nbitq), 
to_sfixed(-12614986.0/4294967296.0,1,-nbitq), 
to_sfixed(190680963.0/4294967296.0,1,-nbitq), 
to_sfixed(-207591725.0/4294967296.0,1,-nbitq), 
to_sfixed(187911417.0/4294967296.0,1,-nbitq), 
to_sfixed(283723019.0/4294967296.0,1,-nbitq), 
to_sfixed(407346488.0/4294967296.0,1,-nbitq), 
to_sfixed(226889554.0/4294967296.0,1,-nbitq), 
to_sfixed(-271028418.0/4294967296.0,1,-nbitq), 
to_sfixed(107719305.0/4294967296.0,1,-nbitq), 
to_sfixed(305321187.0/4294967296.0,1,-nbitq), 
to_sfixed(17564539.0/4294967296.0,1,-nbitq), 
to_sfixed(-39060779.0/4294967296.0,1,-nbitq), 
to_sfixed(403462037.0/4294967296.0,1,-nbitq), 
to_sfixed(131380379.0/4294967296.0,1,-nbitq), 
to_sfixed(-436613394.0/4294967296.0,1,-nbitq), 
to_sfixed(139071148.0/4294967296.0,1,-nbitq), 
to_sfixed(-219028210.0/4294967296.0,1,-nbitq), 
to_sfixed(-264556082.0/4294967296.0,1,-nbitq), 
to_sfixed(62414346.0/4294967296.0,1,-nbitq), 
to_sfixed(-192557532.0/4294967296.0,1,-nbitq), 
to_sfixed(198808376.0/4294967296.0,1,-nbitq), 
to_sfixed(112540335.0/4294967296.0,1,-nbitq), 
to_sfixed(-260839502.0/4294967296.0,1,-nbitq), 
to_sfixed(44125082.0/4294967296.0,1,-nbitq), 
to_sfixed(132756912.0/4294967296.0,1,-nbitq), 
to_sfixed(389533554.0/4294967296.0,1,-nbitq), 
to_sfixed(111745458.0/4294967296.0,1,-nbitq), 
to_sfixed(-219873542.0/4294967296.0,1,-nbitq), 
to_sfixed(423063664.0/4294967296.0,1,-nbitq), 
to_sfixed(-21429616.0/4294967296.0,1,-nbitq), 
to_sfixed(-75607767.0/4294967296.0,1,-nbitq), 
to_sfixed(419096755.0/4294967296.0,1,-nbitq), 
to_sfixed(-158574721.0/4294967296.0,1,-nbitq), 
to_sfixed(402697309.0/4294967296.0,1,-nbitq), 
to_sfixed(300221780.0/4294967296.0,1,-nbitq), 
to_sfixed(-39093912.0/4294967296.0,1,-nbitq), 
to_sfixed(200012886.0/4294967296.0,1,-nbitq), 
to_sfixed(-243525543.0/4294967296.0,1,-nbitq), 
to_sfixed(202114478.0/4294967296.0,1,-nbitq), 
to_sfixed(-382747665.0/4294967296.0,1,-nbitq), 
to_sfixed(-82974749.0/4294967296.0,1,-nbitq), 
to_sfixed(-139982527.0/4294967296.0,1,-nbitq), 
to_sfixed(103551939.0/4294967296.0,1,-nbitq), 
to_sfixed(87718240.0/4294967296.0,1,-nbitq), 
to_sfixed(-62125662.0/4294967296.0,1,-nbitq), 
to_sfixed(-131014162.0/4294967296.0,1,-nbitq), 
to_sfixed(-106167049.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(383177581.0/4294967296.0,1,-nbitq), 
to_sfixed(-69593107.0/4294967296.0,1,-nbitq), 
to_sfixed(140861099.0/4294967296.0,1,-nbitq), 
to_sfixed(-283360036.0/4294967296.0,1,-nbitq), 
to_sfixed(392926057.0/4294967296.0,1,-nbitq), 
to_sfixed(-333576678.0/4294967296.0,1,-nbitq), 
to_sfixed(-296144402.0/4294967296.0,1,-nbitq), 
to_sfixed(194640749.0/4294967296.0,1,-nbitq), 
to_sfixed(42465909.0/4294967296.0,1,-nbitq), 
to_sfixed(195379821.0/4294967296.0,1,-nbitq), 
to_sfixed(-41786315.0/4294967296.0,1,-nbitq), 
to_sfixed(486031414.0/4294967296.0,1,-nbitq), 
to_sfixed(-350853117.0/4294967296.0,1,-nbitq), 
to_sfixed(-249160217.0/4294967296.0,1,-nbitq), 
to_sfixed(-296114679.0/4294967296.0,1,-nbitq), 
to_sfixed(-162498987.0/4294967296.0,1,-nbitq), 
to_sfixed(10359349.0/4294967296.0,1,-nbitq), 
to_sfixed(-398075853.0/4294967296.0,1,-nbitq), 
to_sfixed(-280155782.0/4294967296.0,1,-nbitq), 
to_sfixed(224269194.0/4294967296.0,1,-nbitq), 
to_sfixed(-50030998.0/4294967296.0,1,-nbitq), 
to_sfixed(-157371274.0/4294967296.0,1,-nbitq), 
to_sfixed(485932224.0/4294967296.0,1,-nbitq), 
to_sfixed(416926153.0/4294967296.0,1,-nbitq), 
to_sfixed(-270715520.0/4294967296.0,1,-nbitq), 
to_sfixed(-132883559.0/4294967296.0,1,-nbitq), 
to_sfixed(-300772467.0/4294967296.0,1,-nbitq), 
to_sfixed(-514743730.0/4294967296.0,1,-nbitq), 
to_sfixed(81839557.0/4294967296.0,1,-nbitq), 
to_sfixed(-278825120.0/4294967296.0,1,-nbitq), 
to_sfixed(-1775960.0/4294967296.0,1,-nbitq), 
to_sfixed(54092328.0/4294967296.0,1,-nbitq), 
to_sfixed(191937613.0/4294967296.0,1,-nbitq), 
to_sfixed(-168419933.0/4294967296.0,1,-nbitq), 
to_sfixed(-151158197.0/4294967296.0,1,-nbitq), 
to_sfixed(12777461.0/4294967296.0,1,-nbitq), 
to_sfixed(51725485.0/4294967296.0,1,-nbitq), 
to_sfixed(111482921.0/4294967296.0,1,-nbitq), 
to_sfixed(-18299395.0/4294967296.0,1,-nbitq), 
to_sfixed(-301868159.0/4294967296.0,1,-nbitq), 
to_sfixed(-390107064.0/4294967296.0,1,-nbitq), 
to_sfixed(461628298.0/4294967296.0,1,-nbitq), 
to_sfixed(460995128.0/4294967296.0,1,-nbitq), 
to_sfixed(96327072.0/4294967296.0,1,-nbitq), 
to_sfixed(200205023.0/4294967296.0,1,-nbitq), 
to_sfixed(281069202.0/4294967296.0,1,-nbitq), 
to_sfixed(23127846.0/4294967296.0,1,-nbitq), 
to_sfixed(140044223.0/4294967296.0,1,-nbitq), 
to_sfixed(-102428652.0/4294967296.0,1,-nbitq), 
to_sfixed(75281086.0/4294967296.0,1,-nbitq), 
to_sfixed(13407876.0/4294967296.0,1,-nbitq), 
to_sfixed(409354101.0/4294967296.0,1,-nbitq), 
to_sfixed(191413663.0/4294967296.0,1,-nbitq), 
to_sfixed(98503371.0/4294967296.0,1,-nbitq), 
to_sfixed(120991694.0/4294967296.0,1,-nbitq), 
to_sfixed(-259441584.0/4294967296.0,1,-nbitq), 
to_sfixed(275550930.0/4294967296.0,1,-nbitq), 
to_sfixed(-210219397.0/4294967296.0,1,-nbitq), 
to_sfixed(-196590971.0/4294967296.0,1,-nbitq), 
to_sfixed(221259268.0/4294967296.0,1,-nbitq), 
to_sfixed(75570635.0/4294967296.0,1,-nbitq), 
to_sfixed(20186161.0/4294967296.0,1,-nbitq), 
to_sfixed(147285039.0/4294967296.0,1,-nbitq), 
to_sfixed(257796909.0/4294967296.0,1,-nbitq), 
to_sfixed(396485731.0/4294967296.0,1,-nbitq), 
to_sfixed(-353786821.0/4294967296.0,1,-nbitq), 
to_sfixed(376773659.0/4294967296.0,1,-nbitq), 
to_sfixed(-51035037.0/4294967296.0,1,-nbitq), 
to_sfixed(449026026.0/4294967296.0,1,-nbitq), 
to_sfixed(-205996933.0/4294967296.0,1,-nbitq), 
to_sfixed(-483505115.0/4294967296.0,1,-nbitq), 
to_sfixed(-311936146.0/4294967296.0,1,-nbitq), 
to_sfixed(-461832372.0/4294967296.0,1,-nbitq), 
to_sfixed(269832527.0/4294967296.0,1,-nbitq), 
to_sfixed(425161634.0/4294967296.0,1,-nbitq), 
to_sfixed(-249119382.0/4294967296.0,1,-nbitq), 
to_sfixed(269501525.0/4294967296.0,1,-nbitq), 
to_sfixed(289868502.0/4294967296.0,1,-nbitq), 
to_sfixed(242901077.0/4294967296.0,1,-nbitq), 
to_sfixed(-239092492.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(25865933.0/4294967296.0,1,-nbitq), 
to_sfixed(-162661015.0/4294967296.0,1,-nbitq), 
to_sfixed(512600581.0/4294967296.0,1,-nbitq), 
to_sfixed(-524046323.0/4294967296.0,1,-nbitq), 
to_sfixed(346096686.0/4294967296.0,1,-nbitq), 
to_sfixed(153191369.0/4294967296.0,1,-nbitq), 
to_sfixed(-151764852.0/4294967296.0,1,-nbitq), 
to_sfixed(-138919530.0/4294967296.0,1,-nbitq), 
to_sfixed(129460651.0/4294967296.0,1,-nbitq), 
to_sfixed(313818585.0/4294967296.0,1,-nbitq), 
to_sfixed(179983574.0/4294967296.0,1,-nbitq), 
to_sfixed(-254858991.0/4294967296.0,1,-nbitq), 
to_sfixed(-26838814.0/4294967296.0,1,-nbitq), 
to_sfixed(326955553.0/4294967296.0,1,-nbitq), 
to_sfixed(-68713464.0/4294967296.0,1,-nbitq), 
to_sfixed(122205901.0/4294967296.0,1,-nbitq), 
to_sfixed(116381613.0/4294967296.0,1,-nbitq), 
to_sfixed(-248426353.0/4294967296.0,1,-nbitq), 
to_sfixed(-432504.0/4294967296.0,1,-nbitq), 
to_sfixed(-202648703.0/4294967296.0,1,-nbitq), 
to_sfixed(189917525.0/4294967296.0,1,-nbitq), 
to_sfixed(344198543.0/4294967296.0,1,-nbitq), 
to_sfixed(145301057.0/4294967296.0,1,-nbitq), 
to_sfixed(13924372.0/4294967296.0,1,-nbitq), 
to_sfixed(-30210623.0/4294967296.0,1,-nbitq), 
to_sfixed(581362899.0/4294967296.0,1,-nbitq), 
to_sfixed(123117618.0/4294967296.0,1,-nbitq), 
to_sfixed(-281556886.0/4294967296.0,1,-nbitq), 
to_sfixed(325084790.0/4294967296.0,1,-nbitq), 
to_sfixed(-161795384.0/4294967296.0,1,-nbitq), 
to_sfixed(208995782.0/4294967296.0,1,-nbitq), 
to_sfixed(189247499.0/4294967296.0,1,-nbitq), 
to_sfixed(108908135.0/4294967296.0,1,-nbitq), 
to_sfixed(180600146.0/4294967296.0,1,-nbitq), 
to_sfixed(-195708670.0/4294967296.0,1,-nbitq), 
to_sfixed(312945760.0/4294967296.0,1,-nbitq), 
to_sfixed(28570367.0/4294967296.0,1,-nbitq), 
to_sfixed(192717153.0/4294967296.0,1,-nbitq), 
to_sfixed(327902800.0/4294967296.0,1,-nbitq), 
to_sfixed(-126303167.0/4294967296.0,1,-nbitq), 
to_sfixed(159516744.0/4294967296.0,1,-nbitq), 
to_sfixed(-70149184.0/4294967296.0,1,-nbitq), 
to_sfixed(-200445397.0/4294967296.0,1,-nbitq), 
to_sfixed(362534624.0/4294967296.0,1,-nbitq), 
to_sfixed(207725253.0/4294967296.0,1,-nbitq), 
to_sfixed(-39149224.0/4294967296.0,1,-nbitq), 
to_sfixed(273147374.0/4294967296.0,1,-nbitq), 
to_sfixed(-502362017.0/4294967296.0,1,-nbitq), 
to_sfixed(314399758.0/4294967296.0,1,-nbitq), 
to_sfixed(26839136.0/4294967296.0,1,-nbitq), 
to_sfixed(402441939.0/4294967296.0,1,-nbitq), 
to_sfixed(-272731292.0/4294967296.0,1,-nbitq), 
to_sfixed(-453161836.0/4294967296.0,1,-nbitq), 
to_sfixed(71504475.0/4294967296.0,1,-nbitq), 
to_sfixed(303433181.0/4294967296.0,1,-nbitq), 
to_sfixed(55644725.0/4294967296.0,1,-nbitq), 
to_sfixed(-6563745.0/4294967296.0,1,-nbitq), 
to_sfixed(91936368.0/4294967296.0,1,-nbitq), 
to_sfixed(117481358.0/4294967296.0,1,-nbitq), 
to_sfixed(137438377.0/4294967296.0,1,-nbitq), 
to_sfixed(111829568.0/4294967296.0,1,-nbitq), 
to_sfixed(54941983.0/4294967296.0,1,-nbitq), 
to_sfixed(163371865.0/4294967296.0,1,-nbitq), 
to_sfixed(483612538.0/4294967296.0,1,-nbitq), 
to_sfixed(49497106.0/4294967296.0,1,-nbitq), 
to_sfixed(22313989.0/4294967296.0,1,-nbitq), 
to_sfixed(656660289.0/4294967296.0,1,-nbitq), 
to_sfixed(198479482.0/4294967296.0,1,-nbitq), 
to_sfixed(57222428.0/4294967296.0,1,-nbitq), 
to_sfixed(-222678878.0/4294967296.0,1,-nbitq), 
to_sfixed(-37502683.0/4294967296.0,1,-nbitq), 
to_sfixed(-141489777.0/4294967296.0,1,-nbitq), 
to_sfixed(-430474070.0/4294967296.0,1,-nbitq), 
to_sfixed(-37067234.0/4294967296.0,1,-nbitq), 
to_sfixed(381207860.0/4294967296.0,1,-nbitq), 
to_sfixed(39616224.0/4294967296.0,1,-nbitq), 
to_sfixed(-328853395.0/4294967296.0,1,-nbitq), 
to_sfixed(135547075.0/4294967296.0,1,-nbitq), 
to_sfixed(-102192455.0/4294967296.0,1,-nbitq), 
to_sfixed(-343753519.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-266567153.0/4294967296.0,1,-nbitq), 
to_sfixed(331743030.0/4294967296.0,1,-nbitq), 
to_sfixed(308874968.0/4294967296.0,1,-nbitq), 
to_sfixed(-14205480.0/4294967296.0,1,-nbitq), 
to_sfixed(153823380.0/4294967296.0,1,-nbitq), 
to_sfixed(-24211920.0/4294967296.0,1,-nbitq), 
to_sfixed(185553419.0/4294967296.0,1,-nbitq), 
to_sfixed(257140022.0/4294967296.0,1,-nbitq), 
to_sfixed(-96251135.0/4294967296.0,1,-nbitq), 
to_sfixed(177588093.0/4294967296.0,1,-nbitq), 
to_sfixed(-43754034.0/4294967296.0,1,-nbitq), 
to_sfixed(-461751104.0/4294967296.0,1,-nbitq), 
to_sfixed(743079995.0/4294967296.0,1,-nbitq), 
to_sfixed(279221944.0/4294967296.0,1,-nbitq), 
to_sfixed(-42474691.0/4294967296.0,1,-nbitq), 
to_sfixed(77822647.0/4294967296.0,1,-nbitq), 
to_sfixed(191625364.0/4294967296.0,1,-nbitq), 
to_sfixed(59323084.0/4294967296.0,1,-nbitq), 
to_sfixed(-247853228.0/4294967296.0,1,-nbitq), 
to_sfixed(145813839.0/4294967296.0,1,-nbitq), 
to_sfixed(-276199252.0/4294967296.0,1,-nbitq), 
to_sfixed(112390041.0/4294967296.0,1,-nbitq), 
to_sfixed(-372677002.0/4294967296.0,1,-nbitq), 
to_sfixed(74695072.0/4294967296.0,1,-nbitq), 
to_sfixed(-248568333.0/4294967296.0,1,-nbitq), 
to_sfixed(448855467.0/4294967296.0,1,-nbitq), 
to_sfixed(122238130.0/4294967296.0,1,-nbitq), 
to_sfixed(-151048766.0/4294967296.0,1,-nbitq), 
to_sfixed(-146662695.0/4294967296.0,1,-nbitq), 
to_sfixed(505215177.0/4294967296.0,1,-nbitq), 
to_sfixed(161738323.0/4294967296.0,1,-nbitq), 
to_sfixed(84584320.0/4294967296.0,1,-nbitq), 
to_sfixed(-339516142.0/4294967296.0,1,-nbitq), 
to_sfixed(-82770827.0/4294967296.0,1,-nbitq), 
to_sfixed(123377566.0/4294967296.0,1,-nbitq), 
to_sfixed(286067096.0/4294967296.0,1,-nbitq), 
to_sfixed(-42481549.0/4294967296.0,1,-nbitq), 
to_sfixed(-199979824.0/4294967296.0,1,-nbitq), 
to_sfixed(181276575.0/4294967296.0,1,-nbitq), 
to_sfixed(-28676473.0/4294967296.0,1,-nbitq), 
to_sfixed(-106641646.0/4294967296.0,1,-nbitq), 
to_sfixed(314976641.0/4294967296.0,1,-nbitq), 
to_sfixed(-123483129.0/4294967296.0,1,-nbitq), 
to_sfixed(159111053.0/4294967296.0,1,-nbitq), 
to_sfixed(219974046.0/4294967296.0,1,-nbitq), 
to_sfixed(-352287209.0/4294967296.0,1,-nbitq), 
to_sfixed(220961649.0/4294967296.0,1,-nbitq), 
to_sfixed(-438796724.0/4294967296.0,1,-nbitq), 
to_sfixed(-317177564.0/4294967296.0,1,-nbitq), 
to_sfixed(246988962.0/4294967296.0,1,-nbitq), 
to_sfixed(-185153347.0/4294967296.0,1,-nbitq), 
to_sfixed(127859725.0/4294967296.0,1,-nbitq), 
to_sfixed(130280227.0/4294967296.0,1,-nbitq), 
to_sfixed(375703817.0/4294967296.0,1,-nbitq), 
to_sfixed(-40634652.0/4294967296.0,1,-nbitq), 
to_sfixed(-217546731.0/4294967296.0,1,-nbitq), 
to_sfixed(-22067987.0/4294967296.0,1,-nbitq), 
to_sfixed(-177702012.0/4294967296.0,1,-nbitq), 
to_sfixed(356452658.0/4294967296.0,1,-nbitq), 
to_sfixed(339980292.0/4294967296.0,1,-nbitq), 
to_sfixed(124034520.0/4294967296.0,1,-nbitq), 
to_sfixed(-289223945.0/4294967296.0,1,-nbitq), 
to_sfixed(-228906512.0/4294967296.0,1,-nbitq), 
to_sfixed(402515669.0/4294967296.0,1,-nbitq), 
to_sfixed(-143213411.0/4294967296.0,1,-nbitq), 
to_sfixed(44915663.0/4294967296.0,1,-nbitq), 
to_sfixed(118640575.0/4294967296.0,1,-nbitq), 
to_sfixed(122660023.0/4294967296.0,1,-nbitq), 
to_sfixed(314178647.0/4294967296.0,1,-nbitq), 
to_sfixed(390436198.0/4294967296.0,1,-nbitq), 
to_sfixed(127082213.0/4294967296.0,1,-nbitq), 
to_sfixed(189504992.0/4294967296.0,1,-nbitq), 
to_sfixed(-172756874.0/4294967296.0,1,-nbitq), 
to_sfixed(384893312.0/4294967296.0,1,-nbitq), 
to_sfixed(-48708686.0/4294967296.0,1,-nbitq), 
to_sfixed(-10104050.0/4294967296.0,1,-nbitq), 
to_sfixed(214696324.0/4294967296.0,1,-nbitq), 
to_sfixed(279895897.0/4294967296.0,1,-nbitq), 
to_sfixed(106471255.0/4294967296.0,1,-nbitq), 
to_sfixed(213562184.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-288191564.0/4294967296.0,1,-nbitq), 
to_sfixed(355791929.0/4294967296.0,1,-nbitq), 
to_sfixed(156836606.0/4294967296.0,1,-nbitq), 
to_sfixed(19907661.0/4294967296.0,1,-nbitq), 
to_sfixed(233442895.0/4294967296.0,1,-nbitq), 
to_sfixed(188263299.0/4294967296.0,1,-nbitq), 
to_sfixed(273565468.0/4294967296.0,1,-nbitq), 
to_sfixed(-527298620.0/4294967296.0,1,-nbitq), 
to_sfixed(-605730703.0/4294967296.0,1,-nbitq), 
to_sfixed(160423833.0/4294967296.0,1,-nbitq), 
to_sfixed(-22499948.0/4294967296.0,1,-nbitq), 
to_sfixed(-385173080.0/4294967296.0,1,-nbitq), 
to_sfixed(793583798.0/4294967296.0,1,-nbitq), 
to_sfixed(1102529564.0/4294967296.0,1,-nbitq), 
to_sfixed(313463611.0/4294967296.0,1,-nbitq), 
to_sfixed(-485017294.0/4294967296.0,1,-nbitq), 
to_sfixed(241013035.0/4294967296.0,1,-nbitq), 
to_sfixed(300596306.0/4294967296.0,1,-nbitq), 
to_sfixed(55492169.0/4294967296.0,1,-nbitq), 
to_sfixed(65479207.0/4294967296.0,1,-nbitq), 
to_sfixed(96931126.0/4294967296.0,1,-nbitq), 
to_sfixed(-391669482.0/4294967296.0,1,-nbitq), 
to_sfixed(4150366.0/4294967296.0,1,-nbitq), 
to_sfixed(649864254.0/4294967296.0,1,-nbitq), 
to_sfixed(-225540414.0/4294967296.0,1,-nbitq), 
to_sfixed(893578556.0/4294967296.0,1,-nbitq), 
to_sfixed(123772392.0/4294967296.0,1,-nbitq), 
to_sfixed(-144168417.0/4294967296.0,1,-nbitq), 
to_sfixed(226796427.0/4294967296.0,1,-nbitq), 
to_sfixed(-63511118.0/4294967296.0,1,-nbitq), 
to_sfixed(435961042.0/4294967296.0,1,-nbitq), 
to_sfixed(-146240292.0/4294967296.0,1,-nbitq), 
to_sfixed(-526555589.0/4294967296.0,1,-nbitq), 
to_sfixed(-55731559.0/4294967296.0,1,-nbitq), 
to_sfixed(-327923905.0/4294967296.0,1,-nbitq), 
to_sfixed(293662623.0/4294967296.0,1,-nbitq), 
to_sfixed(103576737.0/4294967296.0,1,-nbitq), 
to_sfixed(-3924549.0/4294967296.0,1,-nbitq), 
to_sfixed(-421965581.0/4294967296.0,1,-nbitq), 
to_sfixed(456049430.0/4294967296.0,1,-nbitq), 
to_sfixed(-394430997.0/4294967296.0,1,-nbitq), 
to_sfixed(-227562176.0/4294967296.0,1,-nbitq), 
to_sfixed(-51698831.0/4294967296.0,1,-nbitq), 
to_sfixed(488368143.0/4294967296.0,1,-nbitq), 
to_sfixed(102047314.0/4294967296.0,1,-nbitq), 
to_sfixed(420417776.0/4294967296.0,1,-nbitq), 
to_sfixed(94637538.0/4294967296.0,1,-nbitq), 
to_sfixed(-543819928.0/4294967296.0,1,-nbitq), 
to_sfixed(118405114.0/4294967296.0,1,-nbitq), 
to_sfixed(-573432472.0/4294967296.0,1,-nbitq), 
to_sfixed(-288871534.0/4294967296.0,1,-nbitq), 
to_sfixed(-603089449.0/4294967296.0,1,-nbitq), 
to_sfixed(-264429247.0/4294967296.0,1,-nbitq), 
to_sfixed(-199159881.0/4294967296.0,1,-nbitq), 
to_sfixed(524413158.0/4294967296.0,1,-nbitq), 
to_sfixed(144420587.0/4294967296.0,1,-nbitq), 
to_sfixed(-109100107.0/4294967296.0,1,-nbitq), 
to_sfixed(-81963222.0/4294967296.0,1,-nbitq), 
to_sfixed(48491549.0/4294967296.0,1,-nbitq), 
to_sfixed(413313887.0/4294967296.0,1,-nbitq), 
to_sfixed(-408646716.0/4294967296.0,1,-nbitq), 
to_sfixed(219309928.0/4294967296.0,1,-nbitq), 
to_sfixed(-202218602.0/4294967296.0,1,-nbitq), 
to_sfixed(581520843.0/4294967296.0,1,-nbitq), 
to_sfixed(205521965.0/4294967296.0,1,-nbitq), 
to_sfixed(-66203205.0/4294967296.0,1,-nbitq), 
to_sfixed(316034035.0/4294967296.0,1,-nbitq), 
to_sfixed(-15045284.0/4294967296.0,1,-nbitq), 
to_sfixed(-53606328.0/4294967296.0,1,-nbitq), 
to_sfixed(319565621.0/4294967296.0,1,-nbitq), 
to_sfixed(162295944.0/4294967296.0,1,-nbitq), 
to_sfixed(371759514.0/4294967296.0,1,-nbitq), 
to_sfixed(-430208585.0/4294967296.0,1,-nbitq), 
to_sfixed(417538747.0/4294967296.0,1,-nbitq), 
to_sfixed(396727564.0/4294967296.0,1,-nbitq), 
to_sfixed(100319991.0/4294967296.0,1,-nbitq), 
to_sfixed(-119401026.0/4294967296.0,1,-nbitq), 
to_sfixed(97902744.0/4294967296.0,1,-nbitq), 
to_sfixed(197890549.0/4294967296.0,1,-nbitq), 
to_sfixed(188348596.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(283099121.0/4294967296.0,1,-nbitq), 
to_sfixed(420518599.0/4294967296.0,1,-nbitq), 
to_sfixed(418023405.0/4294967296.0,1,-nbitq), 
to_sfixed(-325166825.0/4294967296.0,1,-nbitq), 
to_sfixed(152767800.0/4294967296.0,1,-nbitq), 
to_sfixed(-94379153.0/4294967296.0,1,-nbitq), 
to_sfixed(-257438543.0/4294967296.0,1,-nbitq), 
to_sfixed(-291330509.0/4294967296.0,1,-nbitq), 
to_sfixed(-186486502.0/4294967296.0,1,-nbitq), 
to_sfixed(244513392.0/4294967296.0,1,-nbitq), 
to_sfixed(225761114.0/4294967296.0,1,-nbitq), 
to_sfixed(-272604046.0/4294967296.0,1,-nbitq), 
to_sfixed(1274755436.0/4294967296.0,1,-nbitq), 
to_sfixed(1567361456.0/4294967296.0,1,-nbitq), 
to_sfixed(-374513733.0/4294967296.0,1,-nbitq), 
to_sfixed(274137008.0/4294967296.0,1,-nbitq), 
to_sfixed(267127852.0/4294967296.0,1,-nbitq), 
to_sfixed(-60818197.0/4294967296.0,1,-nbitq), 
to_sfixed(-259672829.0/4294967296.0,1,-nbitq), 
to_sfixed(584497769.0/4294967296.0,1,-nbitq), 
to_sfixed(-417206310.0/4294967296.0,1,-nbitq), 
to_sfixed(-79620092.0/4294967296.0,1,-nbitq), 
to_sfixed(-192113690.0/4294967296.0,1,-nbitq), 
to_sfixed(950370178.0/4294967296.0,1,-nbitq), 
to_sfixed(-169583698.0/4294967296.0,1,-nbitq), 
to_sfixed(540027275.0/4294967296.0,1,-nbitq), 
to_sfixed(-408610697.0/4294967296.0,1,-nbitq), 
to_sfixed(353355808.0/4294967296.0,1,-nbitq), 
to_sfixed(218483418.0/4294967296.0,1,-nbitq), 
to_sfixed(11591952.0/4294967296.0,1,-nbitq), 
to_sfixed(-129994491.0/4294967296.0,1,-nbitq), 
to_sfixed(385998920.0/4294967296.0,1,-nbitq), 
to_sfixed(-402682799.0/4294967296.0,1,-nbitq), 
to_sfixed(-691300669.0/4294967296.0,1,-nbitq), 
to_sfixed(50652041.0/4294967296.0,1,-nbitq), 
to_sfixed(-226461680.0/4294967296.0,1,-nbitq), 
to_sfixed(-424260821.0/4294967296.0,1,-nbitq), 
to_sfixed(53932008.0/4294967296.0,1,-nbitq), 
to_sfixed(-321560764.0/4294967296.0,1,-nbitq), 
to_sfixed(-19703544.0/4294967296.0,1,-nbitq), 
to_sfixed(-395538897.0/4294967296.0,1,-nbitq), 
to_sfixed(85984324.0/4294967296.0,1,-nbitq), 
to_sfixed(-196214446.0/4294967296.0,1,-nbitq), 
to_sfixed(220474711.0/4294967296.0,1,-nbitq), 
to_sfixed(244701783.0/4294967296.0,1,-nbitq), 
to_sfixed(264573370.0/4294967296.0,1,-nbitq), 
to_sfixed(-160152125.0/4294967296.0,1,-nbitq), 
to_sfixed(-543178744.0/4294967296.0,1,-nbitq), 
to_sfixed(-272089725.0/4294967296.0,1,-nbitq), 
to_sfixed(-495048281.0/4294967296.0,1,-nbitq), 
to_sfixed(-200641970.0/4294967296.0,1,-nbitq), 
to_sfixed(30279637.0/4294967296.0,1,-nbitq), 
to_sfixed(415612766.0/4294967296.0,1,-nbitq), 
to_sfixed(191302806.0/4294967296.0,1,-nbitq), 
to_sfixed(106350263.0/4294967296.0,1,-nbitq), 
to_sfixed(-196531061.0/4294967296.0,1,-nbitq), 
to_sfixed(173101932.0/4294967296.0,1,-nbitq), 
to_sfixed(90978365.0/4294967296.0,1,-nbitq), 
to_sfixed(-125032707.0/4294967296.0,1,-nbitq), 
to_sfixed(279974893.0/4294967296.0,1,-nbitq), 
to_sfixed(-264065694.0/4294967296.0,1,-nbitq), 
to_sfixed(423908578.0/4294967296.0,1,-nbitq), 
to_sfixed(-266376145.0/4294967296.0,1,-nbitq), 
to_sfixed(581489563.0/4294967296.0,1,-nbitq), 
to_sfixed(-77730387.0/4294967296.0,1,-nbitq), 
to_sfixed(7400680.0/4294967296.0,1,-nbitq), 
to_sfixed(-57914261.0/4294967296.0,1,-nbitq), 
to_sfixed(662008136.0/4294967296.0,1,-nbitq), 
to_sfixed(-199659646.0/4294967296.0,1,-nbitq), 
to_sfixed(92419509.0/4294967296.0,1,-nbitq), 
to_sfixed(1120787690.0/4294967296.0,1,-nbitq), 
to_sfixed(37649164.0/4294967296.0,1,-nbitq), 
to_sfixed(-304546680.0/4294967296.0,1,-nbitq), 
to_sfixed(196227958.0/4294967296.0,1,-nbitq), 
to_sfixed(-290257487.0/4294967296.0,1,-nbitq), 
to_sfixed(261311328.0/4294967296.0,1,-nbitq), 
to_sfixed(160635801.0/4294967296.0,1,-nbitq), 
to_sfixed(195793962.0/4294967296.0,1,-nbitq), 
to_sfixed(-117344607.0/4294967296.0,1,-nbitq), 
to_sfixed(127220374.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-99191834.0/4294967296.0,1,-nbitq), 
to_sfixed(-203158595.0/4294967296.0,1,-nbitq), 
to_sfixed(523721422.0/4294967296.0,1,-nbitq), 
to_sfixed(16621394.0/4294967296.0,1,-nbitq), 
to_sfixed(148505344.0/4294967296.0,1,-nbitq), 
to_sfixed(-235629301.0/4294967296.0,1,-nbitq), 
to_sfixed(-172466006.0/4294967296.0,1,-nbitq), 
to_sfixed(84588616.0/4294967296.0,1,-nbitq), 
to_sfixed(-164957809.0/4294967296.0,1,-nbitq), 
to_sfixed(-200652877.0/4294967296.0,1,-nbitq), 
to_sfixed(317773670.0/4294967296.0,1,-nbitq), 
to_sfixed(274730382.0/4294967296.0,1,-nbitq), 
to_sfixed(1537788719.0/4294967296.0,1,-nbitq), 
to_sfixed(1136581278.0/4294967296.0,1,-nbitq), 
to_sfixed(108895312.0/4294967296.0,1,-nbitq), 
to_sfixed(-499826275.0/4294967296.0,1,-nbitq), 
to_sfixed(163602628.0/4294967296.0,1,-nbitq), 
to_sfixed(36211088.0/4294967296.0,1,-nbitq), 
to_sfixed(-505904375.0/4294967296.0,1,-nbitq), 
to_sfixed(431550989.0/4294967296.0,1,-nbitq), 
to_sfixed(-179038416.0/4294967296.0,1,-nbitq), 
to_sfixed(-362371887.0/4294967296.0,1,-nbitq), 
to_sfixed(106168782.0/4294967296.0,1,-nbitq), 
to_sfixed(656744145.0/4294967296.0,1,-nbitq), 
to_sfixed(87498913.0/4294967296.0,1,-nbitq), 
to_sfixed(922382984.0/4294967296.0,1,-nbitq), 
to_sfixed(77859444.0/4294967296.0,1,-nbitq), 
to_sfixed(276011869.0/4294967296.0,1,-nbitq), 
to_sfixed(229587752.0/4294967296.0,1,-nbitq), 
to_sfixed(2339428.0/4294967296.0,1,-nbitq), 
to_sfixed(-4731639.0/4294967296.0,1,-nbitq), 
to_sfixed(-49855496.0/4294967296.0,1,-nbitq), 
to_sfixed(-216574197.0/4294967296.0,1,-nbitq), 
to_sfixed(-444510194.0/4294967296.0,1,-nbitq), 
to_sfixed(-203672963.0/4294967296.0,1,-nbitq), 
to_sfixed(383626170.0/4294967296.0,1,-nbitq), 
to_sfixed(-212510155.0/4294967296.0,1,-nbitq), 
to_sfixed(-485072846.0/4294967296.0,1,-nbitq), 
to_sfixed(-355081560.0/4294967296.0,1,-nbitq), 
to_sfixed(-14739589.0/4294967296.0,1,-nbitq), 
to_sfixed(156723116.0/4294967296.0,1,-nbitq), 
to_sfixed(-725762678.0/4294967296.0,1,-nbitq), 
to_sfixed(-17918000.0/4294967296.0,1,-nbitq), 
to_sfixed(-189327999.0/4294967296.0,1,-nbitq), 
to_sfixed(446214191.0/4294967296.0,1,-nbitq), 
to_sfixed(341883120.0/4294967296.0,1,-nbitq), 
to_sfixed(-227796558.0/4294967296.0,1,-nbitq), 
to_sfixed(-888443377.0/4294967296.0,1,-nbitq), 
to_sfixed(-231807841.0/4294967296.0,1,-nbitq), 
to_sfixed(109288590.0/4294967296.0,1,-nbitq), 
to_sfixed(-120491374.0/4294967296.0,1,-nbitq), 
to_sfixed(-280216045.0/4294967296.0,1,-nbitq), 
to_sfixed(610964377.0/4294967296.0,1,-nbitq), 
to_sfixed(-263455381.0/4294967296.0,1,-nbitq), 
to_sfixed(479770151.0/4294967296.0,1,-nbitq), 
to_sfixed(534739203.0/4294967296.0,1,-nbitq), 
to_sfixed(118107643.0/4294967296.0,1,-nbitq), 
to_sfixed(101159866.0/4294967296.0,1,-nbitq), 
to_sfixed(-79246661.0/4294967296.0,1,-nbitq), 
to_sfixed(-331233387.0/4294967296.0,1,-nbitq), 
to_sfixed(299915541.0/4294967296.0,1,-nbitq), 
to_sfixed(-266173417.0/4294967296.0,1,-nbitq), 
to_sfixed(-1618585061.0/4294967296.0,1,-nbitq), 
to_sfixed(161839114.0/4294967296.0,1,-nbitq), 
to_sfixed(-134012312.0/4294967296.0,1,-nbitq), 
to_sfixed(-360019691.0/4294967296.0,1,-nbitq), 
to_sfixed(321237212.0/4294967296.0,1,-nbitq), 
to_sfixed(971870948.0/4294967296.0,1,-nbitq), 
to_sfixed(-346420731.0/4294967296.0,1,-nbitq), 
to_sfixed(-243991150.0/4294967296.0,1,-nbitq), 
to_sfixed(82275612.0/4294967296.0,1,-nbitq), 
to_sfixed(-242583957.0/4294967296.0,1,-nbitq), 
to_sfixed(-84053098.0/4294967296.0,1,-nbitq), 
to_sfixed(-257860734.0/4294967296.0,1,-nbitq), 
to_sfixed(417080389.0/4294967296.0,1,-nbitq), 
to_sfixed(620839924.0/4294967296.0,1,-nbitq), 
to_sfixed(740672801.0/4294967296.0,1,-nbitq), 
to_sfixed(-167219924.0/4294967296.0,1,-nbitq), 
to_sfixed(300762120.0/4294967296.0,1,-nbitq), 
to_sfixed(-302921256.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(136119120.0/4294967296.0,1,-nbitq), 
to_sfixed(93854089.0/4294967296.0,1,-nbitq), 
to_sfixed(-733693508.0/4294967296.0,1,-nbitq), 
to_sfixed(-446799263.0/4294967296.0,1,-nbitq), 
to_sfixed(-142524869.0/4294967296.0,1,-nbitq), 
to_sfixed(789483295.0/4294967296.0,1,-nbitq), 
to_sfixed(202357681.0/4294967296.0,1,-nbitq), 
to_sfixed(157805531.0/4294967296.0,1,-nbitq), 
to_sfixed(-592269354.0/4294967296.0,1,-nbitq), 
to_sfixed(134540186.0/4294967296.0,1,-nbitq), 
to_sfixed(-440619085.0/4294967296.0,1,-nbitq), 
to_sfixed(48214809.0/4294967296.0,1,-nbitq), 
to_sfixed(1561310719.0/4294967296.0,1,-nbitq), 
to_sfixed(1232221503.0/4294967296.0,1,-nbitq), 
to_sfixed(143665300.0/4294967296.0,1,-nbitq), 
to_sfixed(-722114969.0/4294967296.0,1,-nbitq), 
to_sfixed(-354508151.0/4294967296.0,1,-nbitq), 
to_sfixed(45378755.0/4294967296.0,1,-nbitq), 
to_sfixed(-281578548.0/4294967296.0,1,-nbitq), 
to_sfixed(438292074.0/4294967296.0,1,-nbitq), 
to_sfixed(323173669.0/4294967296.0,1,-nbitq), 
to_sfixed(-840689639.0/4294967296.0,1,-nbitq), 
to_sfixed(-199594106.0/4294967296.0,1,-nbitq), 
to_sfixed(253744405.0/4294967296.0,1,-nbitq), 
to_sfixed(289569263.0/4294967296.0,1,-nbitq), 
to_sfixed(1315423599.0/4294967296.0,1,-nbitq), 
to_sfixed(-300072744.0/4294967296.0,1,-nbitq), 
to_sfixed(-46698246.0/4294967296.0,1,-nbitq), 
to_sfixed(183786945.0/4294967296.0,1,-nbitq), 
to_sfixed(146003787.0/4294967296.0,1,-nbitq), 
to_sfixed(-115265810.0/4294967296.0,1,-nbitq), 
to_sfixed(201880213.0/4294967296.0,1,-nbitq), 
to_sfixed(-550304907.0/4294967296.0,1,-nbitq), 
to_sfixed(453091219.0/4294967296.0,1,-nbitq), 
to_sfixed(-241788551.0/4294967296.0,1,-nbitq), 
to_sfixed(504030703.0/4294967296.0,1,-nbitq), 
to_sfixed(-445904563.0/4294967296.0,1,-nbitq), 
to_sfixed(-743542377.0/4294967296.0,1,-nbitq), 
to_sfixed(123366933.0/4294967296.0,1,-nbitq), 
to_sfixed(418634405.0/4294967296.0,1,-nbitq), 
to_sfixed(113701730.0/4294967296.0,1,-nbitq), 
to_sfixed(-429583461.0/4294967296.0,1,-nbitq), 
to_sfixed(46792650.0/4294967296.0,1,-nbitq), 
to_sfixed(385325270.0/4294967296.0,1,-nbitq), 
to_sfixed(-500607257.0/4294967296.0,1,-nbitq), 
to_sfixed(469095239.0/4294967296.0,1,-nbitq), 
to_sfixed(276896414.0/4294967296.0,1,-nbitq), 
to_sfixed(-637244255.0/4294967296.0,1,-nbitq), 
to_sfixed(290451464.0/4294967296.0,1,-nbitq), 
to_sfixed(244518549.0/4294967296.0,1,-nbitq), 
to_sfixed(112669532.0/4294967296.0,1,-nbitq), 
to_sfixed(234974593.0/4294967296.0,1,-nbitq), 
to_sfixed(521465164.0/4294967296.0,1,-nbitq), 
to_sfixed(-892870401.0/4294967296.0,1,-nbitq), 
to_sfixed(840262670.0/4294967296.0,1,-nbitq), 
to_sfixed(708252800.0/4294967296.0,1,-nbitq), 
to_sfixed(143760367.0/4294967296.0,1,-nbitq), 
to_sfixed(139760267.0/4294967296.0,1,-nbitq), 
to_sfixed(251398020.0/4294967296.0,1,-nbitq), 
to_sfixed(441619792.0/4294967296.0,1,-nbitq), 
to_sfixed(-279844249.0/4294967296.0,1,-nbitq), 
to_sfixed(-41428468.0/4294967296.0,1,-nbitq), 
to_sfixed(-1520555469.0/4294967296.0,1,-nbitq), 
to_sfixed(-740462179.0/4294967296.0,1,-nbitq), 
to_sfixed(-447417151.0/4294967296.0,1,-nbitq), 
to_sfixed(-457413943.0/4294967296.0,1,-nbitq), 
to_sfixed(326874044.0/4294967296.0,1,-nbitq), 
to_sfixed(1494327708.0/4294967296.0,1,-nbitq), 
to_sfixed(35687753.0/4294967296.0,1,-nbitq), 
to_sfixed(-1408891087.0/4294967296.0,1,-nbitq), 
to_sfixed(394360457.0/4294967296.0,1,-nbitq), 
to_sfixed(-538088827.0/4294967296.0,1,-nbitq), 
to_sfixed(141309953.0/4294967296.0,1,-nbitq), 
to_sfixed(162788010.0/4294967296.0,1,-nbitq), 
to_sfixed(-211376222.0/4294967296.0,1,-nbitq), 
to_sfixed(748414788.0/4294967296.0,1,-nbitq), 
to_sfixed(373211323.0/4294967296.0,1,-nbitq), 
to_sfixed(-251553847.0/4294967296.0,1,-nbitq), 
to_sfixed(1091415272.0/4294967296.0,1,-nbitq), 
to_sfixed(-174000155.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-34840568.0/4294967296.0,1,-nbitq), 
to_sfixed(-177952964.0/4294967296.0,1,-nbitq), 
to_sfixed(-2620433104.0/4294967296.0,1,-nbitq), 
to_sfixed(-508771024.0/4294967296.0,1,-nbitq), 
to_sfixed(358007285.0/4294967296.0,1,-nbitq), 
to_sfixed(1538565221.0/4294967296.0,1,-nbitq), 
to_sfixed(534237594.0/4294967296.0,1,-nbitq), 
to_sfixed(398608379.0/4294967296.0,1,-nbitq), 
to_sfixed(-479832066.0/4294967296.0,1,-nbitq), 
to_sfixed(365701618.0/4294967296.0,1,-nbitq), 
to_sfixed(-1262832451.0/4294967296.0,1,-nbitq), 
to_sfixed(-88990327.0/4294967296.0,1,-nbitq), 
to_sfixed(2045998301.0/4294967296.0,1,-nbitq), 
to_sfixed(986372027.0/4294967296.0,1,-nbitq), 
to_sfixed(-83059209.0/4294967296.0,1,-nbitq), 
to_sfixed(-844640181.0/4294967296.0,1,-nbitq), 
to_sfixed(176930566.0/4294967296.0,1,-nbitq), 
to_sfixed(-210507801.0/4294967296.0,1,-nbitq), 
to_sfixed(509899718.0/4294967296.0,1,-nbitq), 
to_sfixed(672622114.0/4294967296.0,1,-nbitq), 
to_sfixed(118548342.0/4294967296.0,1,-nbitq), 
to_sfixed(-386556031.0/4294967296.0,1,-nbitq), 
to_sfixed(-985885609.0/4294967296.0,1,-nbitq), 
to_sfixed(326250788.0/4294967296.0,1,-nbitq), 
to_sfixed(-221408572.0/4294967296.0,1,-nbitq), 
to_sfixed(671892653.0/4294967296.0,1,-nbitq), 
to_sfixed(-50855036.0/4294967296.0,1,-nbitq), 
to_sfixed(279672497.0/4294967296.0,1,-nbitq), 
to_sfixed(545263491.0/4294967296.0,1,-nbitq), 
to_sfixed(608768056.0/4294967296.0,1,-nbitq), 
to_sfixed(-237432866.0/4294967296.0,1,-nbitq), 
to_sfixed(66971861.0/4294967296.0,1,-nbitq), 
to_sfixed(229635065.0/4294967296.0,1,-nbitq), 
to_sfixed(911066938.0/4294967296.0,1,-nbitq), 
to_sfixed(2213874.0/4294967296.0,1,-nbitq), 
to_sfixed(-637499494.0/4294967296.0,1,-nbitq), 
to_sfixed(120067662.0/4294967296.0,1,-nbitq), 
to_sfixed(68444409.0/4294967296.0,1,-nbitq), 
to_sfixed(-419074892.0/4294967296.0,1,-nbitq), 
to_sfixed(207265749.0/4294967296.0,1,-nbitq), 
to_sfixed(-939820544.0/4294967296.0,1,-nbitq), 
to_sfixed(-579842230.0/4294967296.0,1,-nbitq), 
to_sfixed(249560244.0/4294967296.0,1,-nbitq), 
to_sfixed(809851904.0/4294967296.0,1,-nbitq), 
to_sfixed(-176935567.0/4294967296.0,1,-nbitq), 
to_sfixed(701221811.0/4294967296.0,1,-nbitq), 
to_sfixed(-291644770.0/4294967296.0,1,-nbitq), 
to_sfixed(-848328547.0/4294967296.0,1,-nbitq), 
to_sfixed(-58243072.0/4294967296.0,1,-nbitq), 
to_sfixed(529391331.0/4294967296.0,1,-nbitq), 
to_sfixed(-3000369.0/4294967296.0,1,-nbitq), 
to_sfixed(391866744.0/4294967296.0,1,-nbitq), 
to_sfixed(597178344.0/4294967296.0,1,-nbitq), 
to_sfixed(-554771337.0/4294967296.0,1,-nbitq), 
to_sfixed(615119547.0/4294967296.0,1,-nbitq), 
to_sfixed(637079315.0/4294967296.0,1,-nbitq), 
to_sfixed(393927611.0/4294967296.0,1,-nbitq), 
to_sfixed(746948299.0/4294967296.0,1,-nbitq), 
to_sfixed(-34076380.0/4294967296.0,1,-nbitq), 
to_sfixed(297433814.0/4294967296.0,1,-nbitq), 
to_sfixed(346019157.0/4294967296.0,1,-nbitq), 
to_sfixed(154204804.0/4294967296.0,1,-nbitq), 
to_sfixed(-962050435.0/4294967296.0,1,-nbitq), 
to_sfixed(-904048433.0/4294967296.0,1,-nbitq), 
to_sfixed(-546243945.0/4294967296.0,1,-nbitq), 
to_sfixed(-130724058.0/4294967296.0,1,-nbitq), 
to_sfixed(234658872.0/4294967296.0,1,-nbitq), 
to_sfixed(902888095.0/4294967296.0,1,-nbitq), 
to_sfixed(-195443373.0/4294967296.0,1,-nbitq), 
to_sfixed(-1158443039.0/4294967296.0,1,-nbitq), 
to_sfixed(797799779.0/4294967296.0,1,-nbitq), 
to_sfixed(-159019838.0/4294967296.0,1,-nbitq), 
to_sfixed(-555566544.0/4294967296.0,1,-nbitq), 
to_sfixed(-15551106.0/4294967296.0,1,-nbitq), 
to_sfixed(119299947.0/4294967296.0,1,-nbitq), 
to_sfixed(1133350100.0/4294967296.0,1,-nbitq), 
to_sfixed(-40269593.0/4294967296.0,1,-nbitq), 
to_sfixed(883210.0/4294967296.0,1,-nbitq), 
to_sfixed(843032233.0/4294967296.0,1,-nbitq), 
to_sfixed(408623562.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(189782818.0/4294967296.0,1,-nbitq), 
to_sfixed(-297334839.0/4294967296.0,1,-nbitq), 
to_sfixed(-2068975635.0/4294967296.0,1,-nbitq), 
to_sfixed(-500261792.0/4294967296.0,1,-nbitq), 
to_sfixed(19967395.0/4294967296.0,1,-nbitq), 
to_sfixed(2494638733.0/4294967296.0,1,-nbitq), 
to_sfixed(-238958421.0/4294967296.0,1,-nbitq), 
to_sfixed(1457034635.0/4294967296.0,1,-nbitq), 
to_sfixed(8399924.0/4294967296.0,1,-nbitq), 
to_sfixed(-247162549.0/4294967296.0,1,-nbitq), 
to_sfixed(-1585036328.0/4294967296.0,1,-nbitq), 
to_sfixed(-132618742.0/4294967296.0,1,-nbitq), 
to_sfixed(2140998884.0/4294967296.0,1,-nbitq), 
to_sfixed(928427858.0/4294967296.0,1,-nbitq), 
to_sfixed(-197374751.0/4294967296.0,1,-nbitq), 
to_sfixed(-923419353.0/4294967296.0,1,-nbitq), 
to_sfixed(-140638056.0/4294967296.0,1,-nbitq), 
to_sfixed(387274658.0/4294967296.0,1,-nbitq), 
to_sfixed(125264282.0/4294967296.0,1,-nbitq), 
to_sfixed(476447026.0/4294967296.0,1,-nbitq), 
to_sfixed(-402711273.0/4294967296.0,1,-nbitq), 
to_sfixed(-991786236.0/4294967296.0,1,-nbitq), 
to_sfixed(-1517764359.0/4294967296.0,1,-nbitq), 
to_sfixed(482702919.0/4294967296.0,1,-nbitq), 
to_sfixed(205911220.0/4294967296.0,1,-nbitq), 
to_sfixed(223458455.0/4294967296.0,1,-nbitq), 
to_sfixed(-122365272.0/4294967296.0,1,-nbitq), 
to_sfixed(234575479.0/4294967296.0,1,-nbitq), 
to_sfixed(-248090085.0/4294967296.0,1,-nbitq), 
to_sfixed(365073707.0/4294967296.0,1,-nbitq), 
to_sfixed(222557974.0/4294967296.0,1,-nbitq), 
to_sfixed(-414918727.0/4294967296.0,1,-nbitq), 
to_sfixed(-185599715.0/4294967296.0,1,-nbitq), 
to_sfixed(1141230732.0/4294967296.0,1,-nbitq), 
to_sfixed(-20685134.0/4294967296.0,1,-nbitq), 
to_sfixed(-563324557.0/4294967296.0,1,-nbitq), 
to_sfixed(387729722.0/4294967296.0,1,-nbitq), 
to_sfixed(-560625019.0/4294967296.0,1,-nbitq), 
to_sfixed(-301887439.0/4294967296.0,1,-nbitq), 
to_sfixed(118505854.0/4294967296.0,1,-nbitq), 
to_sfixed(-571533341.0/4294967296.0,1,-nbitq), 
to_sfixed(-768417565.0/4294967296.0,1,-nbitq), 
to_sfixed(405205083.0/4294967296.0,1,-nbitq), 
to_sfixed(-476901743.0/4294967296.0,1,-nbitq), 
to_sfixed(-385559062.0/4294967296.0,1,-nbitq), 
to_sfixed(211741719.0/4294967296.0,1,-nbitq), 
to_sfixed(-209515397.0/4294967296.0,1,-nbitq), 
to_sfixed(-333894484.0/4294967296.0,1,-nbitq), 
to_sfixed(353222083.0/4294967296.0,1,-nbitq), 
to_sfixed(217911276.0/4294967296.0,1,-nbitq), 
to_sfixed(78190362.0/4294967296.0,1,-nbitq), 
to_sfixed(-392701611.0/4294967296.0,1,-nbitq), 
to_sfixed(669007479.0/4294967296.0,1,-nbitq), 
to_sfixed(100988410.0/4294967296.0,1,-nbitq), 
to_sfixed(-93091864.0/4294967296.0,1,-nbitq), 
to_sfixed(48305564.0/4294967296.0,1,-nbitq), 
to_sfixed(203005896.0/4294967296.0,1,-nbitq), 
to_sfixed(372358186.0/4294967296.0,1,-nbitq), 
to_sfixed(-251478908.0/4294967296.0,1,-nbitq), 
to_sfixed(-9155072.0/4294967296.0,1,-nbitq), 
to_sfixed(146800508.0/4294967296.0,1,-nbitq), 
to_sfixed(99550633.0/4294967296.0,1,-nbitq), 
to_sfixed(-1032195018.0/4294967296.0,1,-nbitq), 
to_sfixed(-416466220.0/4294967296.0,1,-nbitq), 
to_sfixed(-406848936.0/4294967296.0,1,-nbitq), 
to_sfixed(64734358.0/4294967296.0,1,-nbitq), 
to_sfixed(-407878834.0/4294967296.0,1,-nbitq), 
to_sfixed(1408615598.0/4294967296.0,1,-nbitq), 
to_sfixed(-248374771.0/4294967296.0,1,-nbitq), 
to_sfixed(-1780369083.0/4294967296.0,1,-nbitq), 
to_sfixed(837951909.0/4294967296.0,1,-nbitq), 
to_sfixed(-712049580.0/4294967296.0,1,-nbitq), 
to_sfixed(138920661.0/4294967296.0,1,-nbitq), 
to_sfixed(-74627665.0/4294967296.0,1,-nbitq), 
to_sfixed(275321507.0/4294967296.0,1,-nbitq), 
to_sfixed(1510399501.0/4294967296.0,1,-nbitq), 
to_sfixed(740070275.0/4294967296.0,1,-nbitq), 
to_sfixed(-386162130.0/4294967296.0,1,-nbitq), 
to_sfixed(1535875496.0/4294967296.0,1,-nbitq), 
to_sfixed(343809243.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(470106189.0/4294967296.0,1,-nbitq), 
to_sfixed(-818409445.0/4294967296.0,1,-nbitq), 
to_sfixed(-1335757975.0/4294967296.0,1,-nbitq), 
to_sfixed(331757970.0/4294967296.0,1,-nbitq), 
to_sfixed(844719798.0/4294967296.0,1,-nbitq), 
to_sfixed(391218210.0/4294967296.0,1,-nbitq), 
to_sfixed(354914093.0/4294967296.0,1,-nbitq), 
to_sfixed(892341531.0/4294967296.0,1,-nbitq), 
to_sfixed(28322956.0/4294967296.0,1,-nbitq), 
to_sfixed(105860279.0/4294967296.0,1,-nbitq), 
to_sfixed(-700253722.0/4294967296.0,1,-nbitq), 
to_sfixed(-633489875.0/4294967296.0,1,-nbitq), 
to_sfixed(1746480822.0/4294967296.0,1,-nbitq), 
to_sfixed(313609223.0/4294967296.0,1,-nbitq), 
to_sfixed(331905233.0/4294967296.0,1,-nbitq), 
to_sfixed(-629494103.0/4294967296.0,1,-nbitq), 
to_sfixed(-26613484.0/4294967296.0,1,-nbitq), 
to_sfixed(-40998825.0/4294967296.0,1,-nbitq), 
to_sfixed(-634146813.0/4294967296.0,1,-nbitq), 
to_sfixed(183858542.0/4294967296.0,1,-nbitq), 
to_sfixed(275833146.0/4294967296.0,1,-nbitq), 
to_sfixed(-1400913307.0/4294967296.0,1,-nbitq), 
to_sfixed(-307662448.0/4294967296.0,1,-nbitq), 
to_sfixed(1142976261.0/4294967296.0,1,-nbitq), 
to_sfixed(4444566.0/4294967296.0,1,-nbitq), 
to_sfixed(384688977.0/4294967296.0,1,-nbitq), 
to_sfixed(-59889508.0/4294967296.0,1,-nbitq), 
to_sfixed(727134251.0/4294967296.0,1,-nbitq), 
to_sfixed(413817590.0/4294967296.0,1,-nbitq), 
to_sfixed(531543082.0/4294967296.0,1,-nbitq), 
to_sfixed(136932836.0/4294967296.0,1,-nbitq), 
to_sfixed(-171340961.0/4294967296.0,1,-nbitq), 
to_sfixed(710654732.0/4294967296.0,1,-nbitq), 
to_sfixed(404772976.0/4294967296.0,1,-nbitq), 
to_sfixed(-495069597.0/4294967296.0,1,-nbitq), 
to_sfixed(-1116753207.0/4294967296.0,1,-nbitq), 
to_sfixed(985075782.0/4294967296.0,1,-nbitq), 
to_sfixed(-795940049.0/4294967296.0,1,-nbitq), 
to_sfixed(-525507848.0/4294967296.0,1,-nbitq), 
to_sfixed(-64724515.0/4294967296.0,1,-nbitq), 
to_sfixed(-448261192.0/4294967296.0,1,-nbitq), 
to_sfixed(-700864736.0/4294967296.0,1,-nbitq), 
to_sfixed(1065300833.0/4294967296.0,1,-nbitq), 
to_sfixed(404541871.0/4294967296.0,1,-nbitq), 
to_sfixed(-554618677.0/4294967296.0,1,-nbitq), 
to_sfixed(773871606.0/4294967296.0,1,-nbitq), 
to_sfixed(130992079.0/4294967296.0,1,-nbitq), 
to_sfixed(-382626178.0/4294967296.0,1,-nbitq), 
to_sfixed(-152883085.0/4294967296.0,1,-nbitq), 
to_sfixed(360156301.0/4294967296.0,1,-nbitq), 
to_sfixed(-867925206.0/4294967296.0,1,-nbitq), 
to_sfixed(-343277636.0/4294967296.0,1,-nbitq), 
to_sfixed(216998217.0/4294967296.0,1,-nbitq), 
to_sfixed(808855861.0/4294967296.0,1,-nbitq), 
to_sfixed(105361551.0/4294967296.0,1,-nbitq), 
to_sfixed(-148649550.0/4294967296.0,1,-nbitq), 
to_sfixed(133136331.0/4294967296.0,1,-nbitq), 
to_sfixed(237325006.0/4294967296.0,1,-nbitq), 
to_sfixed(295923347.0/4294967296.0,1,-nbitq), 
to_sfixed(108871633.0/4294967296.0,1,-nbitq), 
to_sfixed(271220470.0/4294967296.0,1,-nbitq), 
to_sfixed(11175882.0/4294967296.0,1,-nbitq), 
to_sfixed(-892339051.0/4294967296.0,1,-nbitq), 
to_sfixed(522050759.0/4294967296.0,1,-nbitq), 
to_sfixed(409587494.0/4294967296.0,1,-nbitq), 
to_sfixed(-189043361.0/4294967296.0,1,-nbitq), 
to_sfixed(-911158018.0/4294967296.0,1,-nbitq), 
to_sfixed(808501787.0/4294967296.0,1,-nbitq), 
to_sfixed(185970718.0/4294967296.0,1,-nbitq), 
to_sfixed(-1159131589.0/4294967296.0,1,-nbitq), 
to_sfixed(1108286645.0/4294967296.0,1,-nbitq), 
to_sfixed(-554617119.0/4294967296.0,1,-nbitq), 
to_sfixed(773227390.0/4294967296.0,1,-nbitq), 
to_sfixed(-214150671.0/4294967296.0,1,-nbitq), 
to_sfixed(98864214.0/4294967296.0,1,-nbitq), 
to_sfixed(2680273849.0/4294967296.0,1,-nbitq), 
to_sfixed(705899698.0/4294967296.0,1,-nbitq), 
to_sfixed(-467268397.0/4294967296.0,1,-nbitq), 
to_sfixed(1947726027.0/4294967296.0,1,-nbitq), 
to_sfixed(-142337782.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-33973434.0/4294967296.0,1,-nbitq), 
to_sfixed(-768554220.0/4294967296.0,1,-nbitq), 
to_sfixed(-422431632.0/4294967296.0,1,-nbitq), 
to_sfixed(1306183145.0/4294967296.0,1,-nbitq), 
to_sfixed(444756572.0/4294967296.0,1,-nbitq), 
to_sfixed(-63642854.0/4294967296.0,1,-nbitq), 
to_sfixed(-53649558.0/4294967296.0,1,-nbitq), 
to_sfixed(-1460074935.0/4294967296.0,1,-nbitq), 
to_sfixed(-131583466.0/4294967296.0,1,-nbitq), 
to_sfixed(106689154.0/4294967296.0,1,-nbitq), 
to_sfixed(-746862732.0/4294967296.0,1,-nbitq), 
to_sfixed(-508410256.0/4294967296.0,1,-nbitq), 
to_sfixed(1877326623.0/4294967296.0,1,-nbitq), 
to_sfixed(-622763862.0/4294967296.0,1,-nbitq), 
to_sfixed(-292985920.0/4294967296.0,1,-nbitq), 
to_sfixed(-355339714.0/4294967296.0,1,-nbitq), 
to_sfixed(260260111.0/4294967296.0,1,-nbitq), 
to_sfixed(-56450085.0/4294967296.0,1,-nbitq), 
to_sfixed(-883003687.0/4294967296.0,1,-nbitq), 
to_sfixed(-1111847205.0/4294967296.0,1,-nbitq), 
to_sfixed(155905480.0/4294967296.0,1,-nbitq), 
to_sfixed(-663286000.0/4294967296.0,1,-nbitq), 
to_sfixed(195909081.0/4294967296.0,1,-nbitq), 
to_sfixed(1484295693.0/4294967296.0,1,-nbitq), 
to_sfixed(-187722959.0/4294967296.0,1,-nbitq), 
to_sfixed(1170860448.0/4294967296.0,1,-nbitq), 
to_sfixed(-390808391.0/4294967296.0,1,-nbitq), 
to_sfixed(544607938.0/4294967296.0,1,-nbitq), 
to_sfixed(1526875852.0/4294967296.0,1,-nbitq), 
to_sfixed(297867917.0/4294967296.0,1,-nbitq), 
to_sfixed(53018838.0/4294967296.0,1,-nbitq), 
to_sfixed(-362586677.0/4294967296.0,1,-nbitq), 
to_sfixed(330060659.0/4294967296.0,1,-nbitq), 
to_sfixed(-252776119.0/4294967296.0,1,-nbitq), 
to_sfixed(-600079112.0/4294967296.0,1,-nbitq), 
to_sfixed(-1295648437.0/4294967296.0,1,-nbitq), 
to_sfixed(559213391.0/4294967296.0,1,-nbitq), 
to_sfixed(129465218.0/4294967296.0,1,-nbitq), 
to_sfixed(69637602.0/4294967296.0,1,-nbitq), 
to_sfixed(-321325170.0/4294967296.0,1,-nbitq), 
to_sfixed(363845919.0/4294967296.0,1,-nbitq), 
to_sfixed(-287526441.0/4294967296.0,1,-nbitq), 
to_sfixed(559701995.0/4294967296.0,1,-nbitq), 
to_sfixed(395550934.0/4294967296.0,1,-nbitq), 
to_sfixed(-592692981.0/4294967296.0,1,-nbitq), 
to_sfixed(293019407.0/4294967296.0,1,-nbitq), 
to_sfixed(106722958.0/4294967296.0,1,-nbitq), 
to_sfixed(-353865517.0/4294967296.0,1,-nbitq), 
to_sfixed(-96580619.0/4294967296.0,1,-nbitq), 
to_sfixed(289610640.0/4294967296.0,1,-nbitq), 
to_sfixed(-768381619.0/4294967296.0,1,-nbitq), 
to_sfixed(-94787331.0/4294967296.0,1,-nbitq), 
to_sfixed(422430063.0/4294967296.0,1,-nbitq), 
to_sfixed(-59944257.0/4294967296.0,1,-nbitq), 
to_sfixed(-311706917.0/4294967296.0,1,-nbitq), 
to_sfixed(712018093.0/4294967296.0,1,-nbitq), 
to_sfixed(288168034.0/4294967296.0,1,-nbitq), 
to_sfixed(814506881.0/4294967296.0,1,-nbitq), 
to_sfixed(125850698.0/4294967296.0,1,-nbitq), 
to_sfixed(-171322155.0/4294967296.0,1,-nbitq), 
to_sfixed(428084669.0/4294967296.0,1,-nbitq), 
to_sfixed(135890934.0/4294967296.0,1,-nbitq), 
to_sfixed(-435962177.0/4294967296.0,1,-nbitq), 
to_sfixed(1247910203.0/4294967296.0,1,-nbitq), 
to_sfixed(522861378.0/4294967296.0,1,-nbitq), 
to_sfixed(-349014100.0/4294967296.0,1,-nbitq), 
to_sfixed(-209055506.0/4294967296.0,1,-nbitq), 
to_sfixed(854059482.0/4294967296.0,1,-nbitq), 
to_sfixed(-306505054.0/4294967296.0,1,-nbitq), 
to_sfixed(-745181324.0/4294967296.0,1,-nbitq), 
to_sfixed(1396743685.0/4294967296.0,1,-nbitq), 
to_sfixed(-69835326.0/4294967296.0,1,-nbitq), 
to_sfixed(488576513.0/4294967296.0,1,-nbitq), 
to_sfixed(-344282634.0/4294967296.0,1,-nbitq), 
to_sfixed(310594049.0/4294967296.0,1,-nbitq), 
to_sfixed(2262036401.0/4294967296.0,1,-nbitq), 
to_sfixed(503219473.0/4294967296.0,1,-nbitq), 
to_sfixed(-230881082.0/4294967296.0,1,-nbitq), 
to_sfixed(2443836154.0/4294967296.0,1,-nbitq), 
to_sfixed(267117374.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(378917437.0/4294967296.0,1,-nbitq), 
to_sfixed(-246252166.0/4294967296.0,1,-nbitq), 
to_sfixed(493952213.0/4294967296.0,1,-nbitq), 
to_sfixed(521680463.0/4294967296.0,1,-nbitq), 
to_sfixed(171909046.0/4294967296.0,1,-nbitq), 
to_sfixed(10982209.0/4294967296.0,1,-nbitq), 
to_sfixed(-144840345.0/4294967296.0,1,-nbitq), 
to_sfixed(-2240628394.0/4294967296.0,1,-nbitq), 
to_sfixed(863677149.0/4294967296.0,1,-nbitq), 
to_sfixed(168193749.0/4294967296.0,1,-nbitq), 
to_sfixed(672546292.0/4294967296.0,1,-nbitq), 
to_sfixed(-518546669.0/4294967296.0,1,-nbitq), 
to_sfixed(1465505998.0/4294967296.0,1,-nbitq), 
to_sfixed(-1859762878.0/4294967296.0,1,-nbitq), 
to_sfixed(-124441877.0/4294967296.0,1,-nbitq), 
to_sfixed(-934864221.0/4294967296.0,1,-nbitq), 
to_sfixed(-147903033.0/4294967296.0,1,-nbitq), 
to_sfixed(35617614.0/4294967296.0,1,-nbitq), 
to_sfixed(108826434.0/4294967296.0,1,-nbitq), 
to_sfixed(-681807623.0/4294967296.0,1,-nbitq), 
to_sfixed(278816620.0/4294967296.0,1,-nbitq), 
to_sfixed(-16773627.0/4294967296.0,1,-nbitq), 
to_sfixed(-394160255.0/4294967296.0,1,-nbitq), 
to_sfixed(1733206448.0/4294967296.0,1,-nbitq), 
to_sfixed(-70614046.0/4294967296.0,1,-nbitq), 
to_sfixed(1299265150.0/4294967296.0,1,-nbitq), 
to_sfixed(287615728.0/4294967296.0,1,-nbitq), 
to_sfixed(915612017.0/4294967296.0,1,-nbitq), 
to_sfixed(-1257151620.0/4294967296.0,1,-nbitq), 
to_sfixed(-701029072.0/4294967296.0,1,-nbitq), 
to_sfixed(1003165472.0/4294967296.0,1,-nbitq), 
to_sfixed(-623401033.0/4294967296.0,1,-nbitq), 
to_sfixed(204660065.0/4294967296.0,1,-nbitq), 
to_sfixed(-670845441.0/4294967296.0,1,-nbitq), 
to_sfixed(-471432749.0/4294967296.0,1,-nbitq), 
to_sfixed(-33020571.0/4294967296.0,1,-nbitq), 
to_sfixed(800748964.0/4294967296.0,1,-nbitq), 
to_sfixed(273461162.0/4294967296.0,1,-nbitq), 
to_sfixed(579649900.0/4294967296.0,1,-nbitq), 
to_sfixed(227796899.0/4294967296.0,1,-nbitq), 
to_sfixed(1428177829.0/4294967296.0,1,-nbitq), 
to_sfixed(-196162120.0/4294967296.0,1,-nbitq), 
to_sfixed(762205931.0/4294967296.0,1,-nbitq), 
to_sfixed(-185273134.0/4294967296.0,1,-nbitq), 
to_sfixed(-611285738.0/4294967296.0,1,-nbitq), 
to_sfixed(508456000.0/4294967296.0,1,-nbitq), 
to_sfixed(-196497156.0/4294967296.0,1,-nbitq), 
to_sfixed(-1049250970.0/4294967296.0,1,-nbitq), 
to_sfixed(-161786067.0/4294967296.0,1,-nbitq), 
to_sfixed(-272690009.0/4294967296.0,1,-nbitq), 
to_sfixed(-393509339.0/4294967296.0,1,-nbitq), 
to_sfixed(-428091980.0/4294967296.0,1,-nbitq), 
to_sfixed(-178819177.0/4294967296.0,1,-nbitq), 
to_sfixed(-968339563.0/4294967296.0,1,-nbitq), 
to_sfixed(357289015.0/4294967296.0,1,-nbitq), 
to_sfixed(160376984.0/4294967296.0,1,-nbitq), 
to_sfixed(465243137.0/4294967296.0,1,-nbitq), 
to_sfixed(807184153.0/4294967296.0,1,-nbitq), 
to_sfixed(207275427.0/4294967296.0,1,-nbitq), 
to_sfixed(178847368.0/4294967296.0,1,-nbitq), 
to_sfixed(67184328.0/4294967296.0,1,-nbitq), 
to_sfixed(-142439502.0/4294967296.0,1,-nbitq), 
to_sfixed(-26771416.0/4294967296.0,1,-nbitq), 
to_sfixed(858421089.0/4294967296.0,1,-nbitq), 
to_sfixed(298399878.0/4294967296.0,1,-nbitq), 
to_sfixed(138244300.0/4294967296.0,1,-nbitq), 
to_sfixed(321650357.0/4294967296.0,1,-nbitq), 
to_sfixed(1349142120.0/4294967296.0,1,-nbitq), 
to_sfixed(-89770613.0/4294967296.0,1,-nbitq), 
to_sfixed(-498812761.0/4294967296.0,1,-nbitq), 
to_sfixed(1039566701.0/4294967296.0,1,-nbitq), 
to_sfixed(155432056.0/4294967296.0,1,-nbitq), 
to_sfixed(665959012.0/4294967296.0,1,-nbitq), 
to_sfixed(-333018494.0/4294967296.0,1,-nbitq), 
to_sfixed(333162352.0/4294967296.0,1,-nbitq), 
to_sfixed(2144562379.0/4294967296.0,1,-nbitq), 
to_sfixed(1333917616.0/4294967296.0,1,-nbitq), 
to_sfixed(23927858.0/4294967296.0,1,-nbitq), 
to_sfixed(1943411483.0/4294967296.0,1,-nbitq), 
to_sfixed(-292442751.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-37332087.0/4294967296.0,1,-nbitq), 
to_sfixed(-1136031906.0/4294967296.0,1,-nbitq), 
to_sfixed(553417963.0/4294967296.0,1,-nbitq), 
to_sfixed(607364474.0/4294967296.0,1,-nbitq), 
to_sfixed(-27056940.0/4294967296.0,1,-nbitq), 
to_sfixed(-486796800.0/4294967296.0,1,-nbitq), 
to_sfixed(-468702094.0/4294967296.0,1,-nbitq), 
to_sfixed(-923052996.0/4294967296.0,1,-nbitq), 
to_sfixed(-39341889.0/4294967296.0,1,-nbitq), 
to_sfixed(-176106022.0/4294967296.0,1,-nbitq), 
to_sfixed(192953122.0/4294967296.0,1,-nbitq), 
to_sfixed(-778527874.0/4294967296.0,1,-nbitq), 
to_sfixed(950351424.0/4294967296.0,1,-nbitq), 
to_sfixed(92211872.0/4294967296.0,1,-nbitq), 
to_sfixed(-229895165.0/4294967296.0,1,-nbitq), 
to_sfixed(-828939273.0/4294967296.0,1,-nbitq), 
to_sfixed(-115016046.0/4294967296.0,1,-nbitq), 
to_sfixed(-33466561.0/4294967296.0,1,-nbitq), 
to_sfixed(1774190811.0/4294967296.0,1,-nbitq), 
to_sfixed(-141069613.0/4294967296.0,1,-nbitq), 
to_sfixed(-130582562.0/4294967296.0,1,-nbitq), 
to_sfixed(271826389.0/4294967296.0,1,-nbitq), 
to_sfixed(-73873720.0/4294967296.0,1,-nbitq), 
to_sfixed(-108204443.0/4294967296.0,1,-nbitq), 
to_sfixed(-241905676.0/4294967296.0,1,-nbitq), 
to_sfixed(2012031512.0/4294967296.0,1,-nbitq), 
to_sfixed(-12698347.0/4294967296.0,1,-nbitq), 
to_sfixed(83898477.0/4294967296.0,1,-nbitq), 
to_sfixed(-2573807063.0/4294967296.0,1,-nbitq), 
to_sfixed(-1038741257.0/4294967296.0,1,-nbitq), 
to_sfixed(816571459.0/4294967296.0,1,-nbitq), 
to_sfixed(1861222345.0/4294967296.0,1,-nbitq), 
to_sfixed(171745628.0/4294967296.0,1,-nbitq), 
to_sfixed(50167605.0/4294967296.0,1,-nbitq), 
to_sfixed(80799063.0/4294967296.0,1,-nbitq), 
to_sfixed(805407751.0/4294967296.0,1,-nbitq), 
to_sfixed(-16077595.0/4294967296.0,1,-nbitq), 
to_sfixed(1837411484.0/4294967296.0,1,-nbitq), 
to_sfixed(600376920.0/4294967296.0,1,-nbitq), 
to_sfixed(-34328111.0/4294967296.0,1,-nbitq), 
to_sfixed(1794747434.0/4294967296.0,1,-nbitq), 
to_sfixed(170876425.0/4294967296.0,1,-nbitq), 
to_sfixed(1042908574.0/4294967296.0,1,-nbitq), 
to_sfixed(-663557037.0/4294967296.0,1,-nbitq), 
to_sfixed(-870282266.0/4294967296.0,1,-nbitq), 
to_sfixed(-30515462.0/4294967296.0,1,-nbitq), 
to_sfixed(-236217625.0/4294967296.0,1,-nbitq), 
to_sfixed(-327707579.0/4294967296.0,1,-nbitq), 
to_sfixed(254136709.0/4294967296.0,1,-nbitq), 
to_sfixed(-1206888494.0/4294967296.0,1,-nbitq), 
to_sfixed(385106392.0/4294967296.0,1,-nbitq), 
to_sfixed(-633671892.0/4294967296.0,1,-nbitq), 
to_sfixed(-734947327.0/4294967296.0,1,-nbitq), 
to_sfixed(-1047834479.0/4294967296.0,1,-nbitq), 
to_sfixed(-312454277.0/4294967296.0,1,-nbitq), 
to_sfixed(16123399.0/4294967296.0,1,-nbitq), 
to_sfixed(181393989.0/4294967296.0,1,-nbitq), 
to_sfixed(-195330960.0/4294967296.0,1,-nbitq), 
to_sfixed(247015397.0/4294967296.0,1,-nbitq), 
to_sfixed(-2788587.0/4294967296.0,1,-nbitq), 
to_sfixed(51635918.0/4294967296.0,1,-nbitq), 
to_sfixed(-410428740.0/4294967296.0,1,-nbitq), 
to_sfixed(-83079673.0/4294967296.0,1,-nbitq), 
to_sfixed(467082450.0/4294967296.0,1,-nbitq), 
to_sfixed(345311307.0/4294967296.0,1,-nbitq), 
to_sfixed(338357884.0/4294967296.0,1,-nbitq), 
to_sfixed(570433591.0/4294967296.0,1,-nbitq), 
to_sfixed(-444136018.0/4294967296.0,1,-nbitq), 
to_sfixed(-12650214.0/4294967296.0,1,-nbitq), 
to_sfixed(-1654571029.0/4294967296.0,1,-nbitq), 
to_sfixed(-300452235.0/4294967296.0,1,-nbitq), 
to_sfixed(199456671.0/4294967296.0,1,-nbitq), 
to_sfixed(-62582331.0/4294967296.0,1,-nbitq), 
to_sfixed(369238153.0/4294967296.0,1,-nbitq), 
to_sfixed(444579606.0/4294967296.0,1,-nbitq), 
to_sfixed(1541779538.0/4294967296.0,1,-nbitq), 
to_sfixed(860916079.0/4294967296.0,1,-nbitq), 
to_sfixed(-743287418.0/4294967296.0,1,-nbitq), 
to_sfixed(1419837054.0/4294967296.0,1,-nbitq), 
to_sfixed(-319511092.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-386507352.0/4294967296.0,1,-nbitq), 
to_sfixed(-470830563.0/4294967296.0,1,-nbitq), 
to_sfixed(1018362000.0/4294967296.0,1,-nbitq), 
to_sfixed(-155124369.0/4294967296.0,1,-nbitq), 
to_sfixed(-651504546.0/4294967296.0,1,-nbitq), 
to_sfixed(-387961324.0/4294967296.0,1,-nbitq), 
to_sfixed(-576859912.0/4294967296.0,1,-nbitq), 
to_sfixed(1118666545.0/4294967296.0,1,-nbitq), 
to_sfixed(690521743.0/4294967296.0,1,-nbitq), 
to_sfixed(66232377.0/4294967296.0,1,-nbitq), 
to_sfixed(306975453.0/4294967296.0,1,-nbitq), 
to_sfixed(-1020123128.0/4294967296.0,1,-nbitq), 
to_sfixed(1113554613.0/4294967296.0,1,-nbitq), 
to_sfixed(229524239.0/4294967296.0,1,-nbitq), 
to_sfixed(-311170307.0/4294967296.0,1,-nbitq), 
to_sfixed(-1483504756.0/4294967296.0,1,-nbitq), 
to_sfixed(-216737815.0/4294967296.0,1,-nbitq), 
to_sfixed(94867649.0/4294967296.0,1,-nbitq), 
to_sfixed(146027399.0/4294967296.0,1,-nbitq), 
to_sfixed(410918627.0/4294967296.0,1,-nbitq), 
to_sfixed(210688873.0/4294967296.0,1,-nbitq), 
to_sfixed(868693375.0/4294967296.0,1,-nbitq), 
to_sfixed(552882088.0/4294967296.0,1,-nbitq), 
to_sfixed(-2694687203.0/4294967296.0,1,-nbitq), 
to_sfixed(-161680052.0/4294967296.0,1,-nbitq), 
to_sfixed(824229594.0/4294967296.0,1,-nbitq), 
to_sfixed(202336401.0/4294967296.0,1,-nbitq), 
to_sfixed(-1420839138.0/4294967296.0,1,-nbitq), 
to_sfixed(-1506548938.0/4294967296.0,1,-nbitq), 
to_sfixed(-554891206.0/4294967296.0,1,-nbitq), 
to_sfixed(-84045578.0/4294967296.0,1,-nbitq), 
to_sfixed(1211250674.0/4294967296.0,1,-nbitq), 
to_sfixed(-327235169.0/4294967296.0,1,-nbitq), 
to_sfixed(181121848.0/4294967296.0,1,-nbitq), 
to_sfixed(-420954858.0/4294967296.0,1,-nbitq), 
to_sfixed(260293196.0/4294967296.0,1,-nbitq), 
to_sfixed(533170232.0/4294967296.0,1,-nbitq), 
to_sfixed(1259247351.0/4294967296.0,1,-nbitq), 
to_sfixed(-5792029.0/4294967296.0,1,-nbitq), 
to_sfixed(489784223.0/4294967296.0,1,-nbitq), 
to_sfixed(353582896.0/4294967296.0,1,-nbitq), 
to_sfixed(481478567.0/4294967296.0,1,-nbitq), 
to_sfixed(479763736.0/4294967296.0,1,-nbitq), 
to_sfixed(-265207123.0/4294967296.0,1,-nbitq), 
to_sfixed(-1074586994.0/4294967296.0,1,-nbitq), 
to_sfixed(399452261.0/4294967296.0,1,-nbitq), 
to_sfixed(-132151032.0/4294967296.0,1,-nbitq), 
to_sfixed(-179315224.0/4294967296.0,1,-nbitq), 
to_sfixed(144845883.0/4294967296.0,1,-nbitq), 
to_sfixed(-1319288546.0/4294967296.0,1,-nbitq), 
to_sfixed(381422113.0/4294967296.0,1,-nbitq), 
to_sfixed(-1321511823.0/4294967296.0,1,-nbitq), 
to_sfixed(-894218505.0/4294967296.0,1,-nbitq), 
to_sfixed(-1386454593.0/4294967296.0,1,-nbitq), 
to_sfixed(-172615411.0/4294967296.0,1,-nbitq), 
to_sfixed(-469457084.0/4294967296.0,1,-nbitq), 
to_sfixed(398355337.0/4294967296.0,1,-nbitq), 
to_sfixed(298191108.0/4294967296.0,1,-nbitq), 
to_sfixed(373472122.0/4294967296.0,1,-nbitq), 
to_sfixed(135030544.0/4294967296.0,1,-nbitq), 
to_sfixed(397012956.0/4294967296.0,1,-nbitq), 
to_sfixed(758381335.0/4294967296.0,1,-nbitq), 
to_sfixed(-323549844.0/4294967296.0,1,-nbitq), 
to_sfixed(154795040.0/4294967296.0,1,-nbitq), 
to_sfixed(73790606.0/4294967296.0,1,-nbitq), 
to_sfixed(-60302405.0/4294967296.0,1,-nbitq), 
to_sfixed(330165697.0/4294967296.0,1,-nbitq), 
to_sfixed(-31624551.0/4294967296.0,1,-nbitq), 
to_sfixed(-286861202.0/4294967296.0,1,-nbitq), 
to_sfixed(-1167506904.0/4294967296.0,1,-nbitq), 
to_sfixed(-202238764.0/4294967296.0,1,-nbitq), 
to_sfixed(530616744.0/4294967296.0,1,-nbitq), 
to_sfixed(146465419.0/4294967296.0,1,-nbitq), 
to_sfixed(-169737285.0/4294967296.0,1,-nbitq), 
to_sfixed(162822820.0/4294967296.0,1,-nbitq), 
to_sfixed(1128285726.0/4294967296.0,1,-nbitq), 
to_sfixed(1185107750.0/4294967296.0,1,-nbitq), 
to_sfixed(-29454116.0/4294967296.0,1,-nbitq), 
to_sfixed(-107258883.0/4294967296.0,1,-nbitq), 
to_sfixed(-262748304.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(208724346.0/4294967296.0,1,-nbitq), 
to_sfixed(2047939492.0/4294967296.0,1,-nbitq), 
to_sfixed(-107513280.0/4294967296.0,1,-nbitq), 
to_sfixed(-351923582.0/4294967296.0,1,-nbitq), 
to_sfixed(-1133612980.0/4294967296.0,1,-nbitq), 
to_sfixed(-160990843.0/4294967296.0,1,-nbitq), 
to_sfixed(-417067994.0/4294967296.0,1,-nbitq), 
to_sfixed(926452157.0/4294967296.0,1,-nbitq), 
to_sfixed(-76805792.0/4294967296.0,1,-nbitq), 
to_sfixed(363686029.0/4294967296.0,1,-nbitq), 
to_sfixed(-444354896.0/4294967296.0,1,-nbitq), 
to_sfixed(-2066515489.0/4294967296.0,1,-nbitq), 
to_sfixed(397210372.0/4294967296.0,1,-nbitq), 
to_sfixed(544911401.0/4294967296.0,1,-nbitq), 
to_sfixed(44651568.0/4294967296.0,1,-nbitq), 
to_sfixed(-476218586.0/4294967296.0,1,-nbitq), 
to_sfixed(21125337.0/4294967296.0,1,-nbitq), 
to_sfixed(333688470.0/4294967296.0,1,-nbitq), 
to_sfixed(-436120885.0/4294967296.0,1,-nbitq), 
to_sfixed(468063069.0/4294967296.0,1,-nbitq), 
to_sfixed(-135316662.0/4294967296.0,1,-nbitq), 
to_sfixed(303285652.0/4294967296.0,1,-nbitq), 
to_sfixed(684391493.0/4294967296.0,1,-nbitq), 
to_sfixed(-2509017775.0/4294967296.0,1,-nbitq), 
to_sfixed(-331099382.0/4294967296.0,1,-nbitq), 
to_sfixed(-51253153.0/4294967296.0,1,-nbitq), 
to_sfixed(95051661.0/4294967296.0,1,-nbitq), 
to_sfixed(-1317679075.0/4294967296.0,1,-nbitq), 
to_sfixed(-883309848.0/4294967296.0,1,-nbitq), 
to_sfixed(-599223411.0/4294967296.0,1,-nbitq), 
to_sfixed(-1237729987.0/4294967296.0,1,-nbitq), 
to_sfixed(1163208722.0/4294967296.0,1,-nbitq), 
to_sfixed(-211176567.0/4294967296.0,1,-nbitq), 
to_sfixed(420316265.0/4294967296.0,1,-nbitq), 
to_sfixed(684745815.0/4294967296.0,1,-nbitq), 
to_sfixed(189830426.0/4294967296.0,1,-nbitq), 
to_sfixed(-803276132.0/4294967296.0,1,-nbitq), 
to_sfixed(1027524260.0/4294967296.0,1,-nbitq), 
to_sfixed(257870432.0/4294967296.0,1,-nbitq), 
to_sfixed(432210941.0/4294967296.0,1,-nbitq), 
to_sfixed(-263085164.0/4294967296.0,1,-nbitq), 
to_sfixed(665818839.0/4294967296.0,1,-nbitq), 
to_sfixed(-1251050530.0/4294967296.0,1,-nbitq), 
to_sfixed(-777223200.0/4294967296.0,1,-nbitq), 
to_sfixed(-1534278869.0/4294967296.0,1,-nbitq), 
to_sfixed(-584962648.0/4294967296.0,1,-nbitq), 
to_sfixed(-102185578.0/4294967296.0,1,-nbitq), 
to_sfixed(-162891639.0/4294967296.0,1,-nbitq), 
to_sfixed(781766644.0/4294967296.0,1,-nbitq), 
to_sfixed(-178311573.0/4294967296.0,1,-nbitq), 
to_sfixed(-268895368.0/4294967296.0,1,-nbitq), 
to_sfixed(-722731245.0/4294967296.0,1,-nbitq), 
to_sfixed(-122850197.0/4294967296.0,1,-nbitq), 
to_sfixed(-1863774905.0/4294967296.0,1,-nbitq), 
to_sfixed(534302172.0/4294967296.0,1,-nbitq), 
to_sfixed(-957377295.0/4294967296.0,1,-nbitq), 
to_sfixed(650801602.0/4294967296.0,1,-nbitq), 
to_sfixed(1206930236.0/4294967296.0,1,-nbitq), 
to_sfixed(28532277.0/4294967296.0,1,-nbitq), 
to_sfixed(-243907667.0/4294967296.0,1,-nbitq), 
to_sfixed(-290117857.0/4294967296.0,1,-nbitq), 
to_sfixed(637219502.0/4294967296.0,1,-nbitq), 
to_sfixed(-343295045.0/4294967296.0,1,-nbitq), 
to_sfixed(-448963036.0/4294967296.0,1,-nbitq), 
to_sfixed(131087006.0/4294967296.0,1,-nbitq), 
to_sfixed(-274081041.0/4294967296.0,1,-nbitq), 
to_sfixed(1092946335.0/4294967296.0,1,-nbitq), 
to_sfixed(57836916.0/4294967296.0,1,-nbitq), 
to_sfixed(-23214845.0/4294967296.0,1,-nbitq), 
to_sfixed(-309084193.0/4294967296.0,1,-nbitq), 
to_sfixed(-1090816777.0/4294967296.0,1,-nbitq), 
to_sfixed(-294440505.0/4294967296.0,1,-nbitq), 
to_sfixed(516054619.0/4294967296.0,1,-nbitq), 
to_sfixed(275645751.0/4294967296.0,1,-nbitq), 
to_sfixed(24011769.0/4294967296.0,1,-nbitq), 
to_sfixed(234294561.0/4294967296.0,1,-nbitq), 
to_sfixed(662561692.0/4294967296.0,1,-nbitq), 
to_sfixed(107086401.0/4294967296.0,1,-nbitq), 
to_sfixed(-447648182.0/4294967296.0,1,-nbitq), 
to_sfixed(229802048.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(31258720.0/4294967296.0,1,-nbitq), 
to_sfixed(1721775210.0/4294967296.0,1,-nbitq), 
to_sfixed(-65904832.0/4294967296.0,1,-nbitq), 
to_sfixed(-741224097.0/4294967296.0,1,-nbitq), 
to_sfixed(32356417.0/4294967296.0,1,-nbitq), 
to_sfixed(262381397.0/4294967296.0,1,-nbitq), 
to_sfixed(-279010489.0/4294967296.0,1,-nbitq), 
to_sfixed(405507677.0/4294967296.0,1,-nbitq), 
to_sfixed(-805709584.0/4294967296.0,1,-nbitq), 
to_sfixed(416176120.0/4294967296.0,1,-nbitq), 
to_sfixed(-443765269.0/4294967296.0,1,-nbitq), 
to_sfixed(-1988091986.0/4294967296.0,1,-nbitq), 
to_sfixed(842693212.0/4294967296.0,1,-nbitq), 
to_sfixed(215500570.0/4294967296.0,1,-nbitq), 
to_sfixed(157658003.0/4294967296.0,1,-nbitq), 
to_sfixed(-943184919.0/4294967296.0,1,-nbitq), 
to_sfixed(-375875927.0/4294967296.0,1,-nbitq), 
to_sfixed(-255091713.0/4294967296.0,1,-nbitq), 
to_sfixed(714396012.0/4294967296.0,1,-nbitq), 
to_sfixed(530534687.0/4294967296.0,1,-nbitq), 
to_sfixed(-38429024.0/4294967296.0,1,-nbitq), 
to_sfixed(548003482.0/4294967296.0,1,-nbitq), 
to_sfixed(282722675.0/4294967296.0,1,-nbitq), 
to_sfixed(-322146215.0/4294967296.0,1,-nbitq), 
to_sfixed(225912948.0/4294967296.0,1,-nbitq), 
to_sfixed(-720512192.0/4294967296.0,1,-nbitq), 
to_sfixed(-205460974.0/4294967296.0,1,-nbitq), 
to_sfixed(-558879599.0/4294967296.0,1,-nbitq), 
to_sfixed(28429553.0/4294967296.0,1,-nbitq), 
to_sfixed(-529623443.0/4294967296.0,1,-nbitq), 
to_sfixed(-644662792.0/4294967296.0,1,-nbitq), 
to_sfixed(870835167.0/4294967296.0,1,-nbitq), 
to_sfixed(-522087698.0/4294967296.0,1,-nbitq), 
to_sfixed(986423375.0/4294967296.0,1,-nbitq), 
to_sfixed(-161193381.0/4294967296.0,1,-nbitq), 
to_sfixed(476940974.0/4294967296.0,1,-nbitq), 
to_sfixed(-364892976.0/4294967296.0,1,-nbitq), 
to_sfixed(578166986.0/4294967296.0,1,-nbitq), 
to_sfixed(-329508388.0/4294967296.0,1,-nbitq), 
to_sfixed(-42798629.0/4294967296.0,1,-nbitq), 
to_sfixed(-548266181.0/4294967296.0,1,-nbitq), 
to_sfixed(929068220.0/4294967296.0,1,-nbitq), 
to_sfixed(-985811212.0/4294967296.0,1,-nbitq), 
to_sfixed(-257654823.0/4294967296.0,1,-nbitq), 
to_sfixed(-1360289252.0/4294967296.0,1,-nbitq), 
to_sfixed(635074914.0/4294967296.0,1,-nbitq), 
to_sfixed(333350951.0/4294967296.0,1,-nbitq), 
to_sfixed(88904725.0/4294967296.0,1,-nbitq), 
to_sfixed(339243804.0/4294967296.0,1,-nbitq), 
to_sfixed(355425547.0/4294967296.0,1,-nbitq), 
to_sfixed(163471303.0/4294967296.0,1,-nbitq), 
to_sfixed(-710571863.0/4294967296.0,1,-nbitq), 
to_sfixed(467024218.0/4294967296.0,1,-nbitq), 
to_sfixed(-1085724635.0/4294967296.0,1,-nbitq), 
to_sfixed(124432548.0/4294967296.0,1,-nbitq), 
to_sfixed(-1534306391.0/4294967296.0,1,-nbitq), 
to_sfixed(15471196.0/4294967296.0,1,-nbitq), 
to_sfixed(340463141.0/4294967296.0,1,-nbitq), 
to_sfixed(398109277.0/4294967296.0,1,-nbitq), 
to_sfixed(-101897217.0/4294967296.0,1,-nbitq), 
to_sfixed(-35767730.0/4294967296.0,1,-nbitq), 
to_sfixed(263572155.0/4294967296.0,1,-nbitq), 
to_sfixed(-172632853.0/4294967296.0,1,-nbitq), 
to_sfixed(-431233154.0/4294967296.0,1,-nbitq), 
to_sfixed(123330087.0/4294967296.0,1,-nbitq), 
to_sfixed(167533337.0/4294967296.0,1,-nbitq), 
to_sfixed(-631062065.0/4294967296.0,1,-nbitq), 
to_sfixed(112445975.0/4294967296.0,1,-nbitq), 
to_sfixed(149500859.0/4294967296.0,1,-nbitq), 
to_sfixed(-391706372.0/4294967296.0,1,-nbitq), 
to_sfixed(-1094033026.0/4294967296.0,1,-nbitq), 
to_sfixed(-227454526.0/4294967296.0,1,-nbitq), 
to_sfixed(-632175339.0/4294967296.0,1,-nbitq), 
to_sfixed(373943603.0/4294967296.0,1,-nbitq), 
to_sfixed(-79363229.0/4294967296.0,1,-nbitq), 
to_sfixed(-435835603.0/4294967296.0,1,-nbitq), 
to_sfixed(468087213.0/4294967296.0,1,-nbitq), 
to_sfixed(241681586.0/4294967296.0,1,-nbitq), 
to_sfixed(-719639511.0/4294967296.0,1,-nbitq), 
to_sfixed(-311085211.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(321751657.0/4294967296.0,1,-nbitq), 
to_sfixed(706627778.0/4294967296.0,1,-nbitq), 
to_sfixed(-472995753.0/4294967296.0,1,-nbitq), 
to_sfixed(-1126753890.0/4294967296.0,1,-nbitq), 
to_sfixed(125106130.0/4294967296.0,1,-nbitq), 
to_sfixed(69318550.0/4294967296.0,1,-nbitq), 
to_sfixed(222056857.0/4294967296.0,1,-nbitq), 
to_sfixed(-27041166.0/4294967296.0,1,-nbitq), 
to_sfixed(-923167299.0/4294967296.0,1,-nbitq), 
to_sfixed(-268062683.0/4294967296.0,1,-nbitq), 
to_sfixed(-844789001.0/4294967296.0,1,-nbitq), 
to_sfixed(-1374664007.0/4294967296.0,1,-nbitq), 
to_sfixed(1280554319.0/4294967296.0,1,-nbitq), 
to_sfixed(717150953.0/4294967296.0,1,-nbitq), 
to_sfixed(231407767.0/4294967296.0,1,-nbitq), 
to_sfixed(-1609759094.0/4294967296.0,1,-nbitq), 
to_sfixed(244102401.0/4294967296.0,1,-nbitq), 
to_sfixed(-118956233.0/4294967296.0,1,-nbitq), 
to_sfixed(-42151441.0/4294967296.0,1,-nbitq), 
to_sfixed(475785189.0/4294967296.0,1,-nbitq), 
to_sfixed(-344080654.0/4294967296.0,1,-nbitq), 
to_sfixed(-324839837.0/4294967296.0,1,-nbitq), 
to_sfixed(388056056.0/4294967296.0,1,-nbitq), 
to_sfixed(978038.0/4294967296.0,1,-nbitq), 
to_sfixed(227371079.0/4294967296.0,1,-nbitq), 
to_sfixed(-760477397.0/4294967296.0,1,-nbitq), 
to_sfixed(127469698.0/4294967296.0,1,-nbitq), 
to_sfixed(-791811114.0/4294967296.0,1,-nbitq), 
to_sfixed(671431164.0/4294967296.0,1,-nbitq), 
to_sfixed(-580883367.0/4294967296.0,1,-nbitq), 
to_sfixed(-349099026.0/4294967296.0,1,-nbitq), 
to_sfixed(1048417008.0/4294967296.0,1,-nbitq), 
to_sfixed(-482376308.0/4294967296.0,1,-nbitq), 
to_sfixed(467232585.0/4294967296.0,1,-nbitq), 
to_sfixed(-210657412.0/4294967296.0,1,-nbitq), 
to_sfixed(383511962.0/4294967296.0,1,-nbitq), 
to_sfixed(-518411003.0/4294967296.0,1,-nbitq), 
to_sfixed(-363219398.0/4294967296.0,1,-nbitq), 
to_sfixed(-36638383.0/4294967296.0,1,-nbitq), 
to_sfixed(190350907.0/4294967296.0,1,-nbitq), 
to_sfixed(-440040998.0/4294967296.0,1,-nbitq), 
to_sfixed(943996738.0/4294967296.0,1,-nbitq), 
to_sfixed(-1210744734.0/4294967296.0,1,-nbitq), 
to_sfixed(-623122609.0/4294967296.0,1,-nbitq), 
to_sfixed(-621731576.0/4294967296.0,1,-nbitq), 
to_sfixed(58974739.0/4294967296.0,1,-nbitq), 
to_sfixed(179950698.0/4294967296.0,1,-nbitq), 
to_sfixed(27587747.0/4294967296.0,1,-nbitq), 
to_sfixed(177367651.0/4294967296.0,1,-nbitq), 
to_sfixed(-95103230.0/4294967296.0,1,-nbitq), 
to_sfixed(-265064732.0/4294967296.0,1,-nbitq), 
to_sfixed(-588729146.0/4294967296.0,1,-nbitq), 
to_sfixed(-515367219.0/4294967296.0,1,-nbitq), 
to_sfixed(-1208869340.0/4294967296.0,1,-nbitq), 
to_sfixed(145908469.0/4294967296.0,1,-nbitq), 
to_sfixed(-1665060760.0/4294967296.0,1,-nbitq), 
to_sfixed(747797602.0/4294967296.0,1,-nbitq), 
to_sfixed(198211274.0/4294967296.0,1,-nbitq), 
to_sfixed(85694022.0/4294967296.0,1,-nbitq), 
to_sfixed(75425833.0/4294967296.0,1,-nbitq), 
to_sfixed(-146020946.0/4294967296.0,1,-nbitq), 
to_sfixed(91339305.0/4294967296.0,1,-nbitq), 
to_sfixed(387579011.0/4294967296.0,1,-nbitq), 
to_sfixed(-204766891.0/4294967296.0,1,-nbitq), 
to_sfixed(-312658462.0/4294967296.0,1,-nbitq), 
to_sfixed(-272024568.0/4294967296.0,1,-nbitq), 
to_sfixed(-907912155.0/4294967296.0,1,-nbitq), 
to_sfixed(-846543826.0/4294967296.0,1,-nbitq), 
to_sfixed(-59355557.0/4294967296.0,1,-nbitq), 
to_sfixed(-1080334456.0/4294967296.0,1,-nbitq), 
to_sfixed(-43119241.0/4294967296.0,1,-nbitq), 
to_sfixed(304855507.0/4294967296.0,1,-nbitq), 
to_sfixed(-1640358044.0/4294967296.0,1,-nbitq), 
to_sfixed(216139348.0/4294967296.0,1,-nbitq), 
to_sfixed(364761254.0/4294967296.0,1,-nbitq), 
to_sfixed(-304589929.0/4294967296.0,1,-nbitq), 
to_sfixed(9862104.0/4294967296.0,1,-nbitq), 
to_sfixed(125056934.0/4294967296.0,1,-nbitq), 
to_sfixed(-1146417160.0/4294967296.0,1,-nbitq), 
to_sfixed(413570670.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(135969936.0/4294967296.0,1,-nbitq), 
to_sfixed(870801656.0/4294967296.0,1,-nbitq), 
to_sfixed(-210393725.0/4294967296.0,1,-nbitq), 
to_sfixed(-1464767721.0/4294967296.0,1,-nbitq), 
to_sfixed(449901742.0/4294967296.0,1,-nbitq), 
to_sfixed(334127678.0/4294967296.0,1,-nbitq), 
to_sfixed(-92751245.0/4294967296.0,1,-nbitq), 
to_sfixed(-597933528.0/4294967296.0,1,-nbitq), 
to_sfixed(-974418774.0/4294967296.0,1,-nbitq), 
to_sfixed(229552268.0/4294967296.0,1,-nbitq), 
to_sfixed(-768865967.0/4294967296.0,1,-nbitq), 
to_sfixed(-1222858507.0/4294967296.0,1,-nbitq), 
to_sfixed(568792848.0/4294967296.0,1,-nbitq), 
to_sfixed(414287953.0/4294967296.0,1,-nbitq), 
to_sfixed(164576008.0/4294967296.0,1,-nbitq), 
to_sfixed(-747389226.0/4294967296.0,1,-nbitq), 
to_sfixed(-381553737.0/4294967296.0,1,-nbitq), 
to_sfixed(429764197.0/4294967296.0,1,-nbitq), 
to_sfixed(488373845.0/4294967296.0,1,-nbitq), 
to_sfixed(-70855289.0/4294967296.0,1,-nbitq), 
to_sfixed(336402329.0/4294967296.0,1,-nbitq), 
to_sfixed(-110379441.0/4294967296.0,1,-nbitq), 
to_sfixed(-36315283.0/4294967296.0,1,-nbitq), 
to_sfixed(85760816.0/4294967296.0,1,-nbitq), 
to_sfixed(-332368751.0/4294967296.0,1,-nbitq), 
to_sfixed(683913230.0/4294967296.0,1,-nbitq), 
to_sfixed(-462884695.0/4294967296.0,1,-nbitq), 
to_sfixed(127997045.0/4294967296.0,1,-nbitq), 
to_sfixed(501422086.0/4294967296.0,1,-nbitq), 
to_sfixed(-739583428.0/4294967296.0,1,-nbitq), 
to_sfixed(-235488744.0/4294967296.0,1,-nbitq), 
to_sfixed(736445193.0/4294967296.0,1,-nbitq), 
to_sfixed(-453389017.0/4294967296.0,1,-nbitq), 
to_sfixed(677601854.0/4294967296.0,1,-nbitq), 
to_sfixed(-146755948.0/4294967296.0,1,-nbitq), 
to_sfixed(391485624.0/4294967296.0,1,-nbitq), 
to_sfixed(-737098981.0/4294967296.0,1,-nbitq), 
to_sfixed(-221002155.0/4294967296.0,1,-nbitq), 
to_sfixed(295919327.0/4294967296.0,1,-nbitq), 
to_sfixed(-146665209.0/4294967296.0,1,-nbitq), 
to_sfixed(-724707229.0/4294967296.0,1,-nbitq), 
to_sfixed(762121601.0/4294967296.0,1,-nbitq), 
to_sfixed(-364477890.0/4294967296.0,1,-nbitq), 
to_sfixed(382300417.0/4294967296.0,1,-nbitq), 
to_sfixed(-800644284.0/4294967296.0,1,-nbitq), 
to_sfixed(1690809946.0/4294967296.0,1,-nbitq), 
to_sfixed(411704729.0/4294967296.0,1,-nbitq), 
to_sfixed(507860027.0/4294967296.0,1,-nbitq), 
to_sfixed(551807109.0/4294967296.0,1,-nbitq), 
to_sfixed(-521342845.0/4294967296.0,1,-nbitq), 
to_sfixed(-163788969.0/4294967296.0,1,-nbitq), 
to_sfixed(-1051080725.0/4294967296.0,1,-nbitq), 
to_sfixed(-77175392.0/4294967296.0,1,-nbitq), 
to_sfixed(421204812.0/4294967296.0,1,-nbitq), 
to_sfixed(-600652232.0/4294967296.0,1,-nbitq), 
to_sfixed(-1051489111.0/4294967296.0,1,-nbitq), 
to_sfixed(-64279843.0/4294967296.0,1,-nbitq), 
to_sfixed(206205894.0/4294967296.0,1,-nbitq), 
to_sfixed(211350125.0/4294967296.0,1,-nbitq), 
to_sfixed(-176945611.0/4294967296.0,1,-nbitq), 
to_sfixed(189323774.0/4294967296.0,1,-nbitq), 
to_sfixed(673249725.0/4294967296.0,1,-nbitq), 
to_sfixed(351080921.0/4294967296.0,1,-nbitq), 
to_sfixed(-1178750814.0/4294967296.0,1,-nbitq), 
to_sfixed(-131081694.0/4294967296.0,1,-nbitq), 
to_sfixed(112409807.0/4294967296.0,1,-nbitq), 
to_sfixed(-1662529481.0/4294967296.0,1,-nbitq), 
to_sfixed(-1107076586.0/4294967296.0,1,-nbitq), 
to_sfixed(-194972678.0/4294967296.0,1,-nbitq), 
to_sfixed(-1383693776.0/4294967296.0,1,-nbitq), 
to_sfixed(-16621586.0/4294967296.0,1,-nbitq), 
to_sfixed(-408068894.0/4294967296.0,1,-nbitq), 
to_sfixed(-1381570474.0/4294967296.0,1,-nbitq), 
to_sfixed(310803926.0/4294967296.0,1,-nbitq), 
to_sfixed(78369623.0/4294967296.0,1,-nbitq), 
to_sfixed(285039035.0/4294967296.0,1,-nbitq), 
to_sfixed(198453112.0/4294967296.0,1,-nbitq), 
to_sfixed(-56543889.0/4294967296.0,1,-nbitq), 
to_sfixed(-567836449.0/4294967296.0,1,-nbitq), 
to_sfixed(347231128.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-97735132.0/4294967296.0,1,-nbitq), 
to_sfixed(1009574603.0/4294967296.0,1,-nbitq), 
to_sfixed(-1316683917.0/4294967296.0,1,-nbitq), 
to_sfixed(-1648242928.0/4294967296.0,1,-nbitq), 
to_sfixed(426448920.0/4294967296.0,1,-nbitq), 
to_sfixed(-228481192.0/4294967296.0,1,-nbitq), 
to_sfixed(-22230430.0/4294967296.0,1,-nbitq), 
to_sfixed(-236984961.0/4294967296.0,1,-nbitq), 
to_sfixed(-454599299.0/4294967296.0,1,-nbitq), 
to_sfixed(-60754831.0/4294967296.0,1,-nbitq), 
to_sfixed(-703366915.0/4294967296.0,1,-nbitq), 
to_sfixed(-531092553.0/4294967296.0,1,-nbitq), 
to_sfixed(1247366168.0/4294967296.0,1,-nbitq), 
to_sfixed(-297866154.0/4294967296.0,1,-nbitq), 
to_sfixed(-150512553.0/4294967296.0,1,-nbitq), 
to_sfixed(-782151999.0/4294967296.0,1,-nbitq), 
to_sfixed(146398327.0/4294967296.0,1,-nbitq), 
to_sfixed(-364483431.0/4294967296.0,1,-nbitq), 
to_sfixed(41439792.0/4294967296.0,1,-nbitq), 
to_sfixed(479316035.0/4294967296.0,1,-nbitq), 
to_sfixed(356239136.0/4294967296.0,1,-nbitq), 
to_sfixed(-251632030.0/4294967296.0,1,-nbitq), 
to_sfixed(274243101.0/4294967296.0,1,-nbitq), 
to_sfixed(263441019.0/4294967296.0,1,-nbitq), 
to_sfixed(-81901464.0/4294967296.0,1,-nbitq), 
to_sfixed(1209639188.0/4294967296.0,1,-nbitq), 
to_sfixed(-830533084.0/4294967296.0,1,-nbitq), 
to_sfixed(211859324.0/4294967296.0,1,-nbitq), 
to_sfixed(139711801.0/4294967296.0,1,-nbitq), 
to_sfixed(-474534169.0/4294967296.0,1,-nbitq), 
to_sfixed(-441110492.0/4294967296.0,1,-nbitq), 
to_sfixed(607014103.0/4294967296.0,1,-nbitq), 
to_sfixed(238450503.0/4294967296.0,1,-nbitq), 
to_sfixed(612823061.0/4294967296.0,1,-nbitq), 
to_sfixed(-292085926.0/4294967296.0,1,-nbitq), 
to_sfixed(390855576.0/4294967296.0,1,-nbitq), 
to_sfixed(-108185628.0/4294967296.0,1,-nbitq), 
to_sfixed(138630687.0/4294967296.0,1,-nbitq), 
to_sfixed(374718408.0/4294967296.0,1,-nbitq), 
to_sfixed(-209735385.0/4294967296.0,1,-nbitq), 
to_sfixed(49133432.0/4294967296.0,1,-nbitq), 
to_sfixed(603791018.0/4294967296.0,1,-nbitq), 
to_sfixed(-790175840.0/4294967296.0,1,-nbitq), 
to_sfixed(-555069191.0/4294967296.0,1,-nbitq), 
to_sfixed(-586110966.0/4294967296.0,1,-nbitq), 
to_sfixed(228934419.0/4294967296.0,1,-nbitq), 
to_sfixed(-366484801.0/4294967296.0,1,-nbitq), 
to_sfixed(1997705.0/4294967296.0,1,-nbitq), 
to_sfixed(-444318520.0/4294967296.0,1,-nbitq), 
to_sfixed(513925917.0/4294967296.0,1,-nbitq), 
to_sfixed(98484564.0/4294967296.0,1,-nbitq), 
to_sfixed(-810000225.0/4294967296.0,1,-nbitq), 
to_sfixed(177217259.0/4294967296.0,1,-nbitq), 
to_sfixed(634187966.0/4294967296.0,1,-nbitq), 
to_sfixed(-59435313.0/4294967296.0,1,-nbitq), 
to_sfixed(-238945110.0/4294967296.0,1,-nbitq), 
to_sfixed(314671399.0/4294967296.0,1,-nbitq), 
to_sfixed(166777657.0/4294967296.0,1,-nbitq), 
to_sfixed(120417518.0/4294967296.0,1,-nbitq), 
to_sfixed(356315800.0/4294967296.0,1,-nbitq), 
to_sfixed(384557563.0/4294967296.0,1,-nbitq), 
to_sfixed(-227620651.0/4294967296.0,1,-nbitq), 
to_sfixed(-22403272.0/4294967296.0,1,-nbitq), 
to_sfixed(-913301816.0/4294967296.0,1,-nbitq), 
to_sfixed(-97127894.0/4294967296.0,1,-nbitq), 
to_sfixed(-397143683.0/4294967296.0,1,-nbitq), 
to_sfixed(-620859875.0/4294967296.0,1,-nbitq), 
to_sfixed(-1022515605.0/4294967296.0,1,-nbitq), 
to_sfixed(-246032074.0/4294967296.0,1,-nbitq), 
to_sfixed(-616465724.0/4294967296.0,1,-nbitq), 
to_sfixed(227438202.0/4294967296.0,1,-nbitq), 
to_sfixed(-400486399.0/4294967296.0,1,-nbitq), 
to_sfixed(-1046683764.0/4294967296.0,1,-nbitq), 
to_sfixed(-153350559.0/4294967296.0,1,-nbitq), 
to_sfixed(338080504.0/4294967296.0,1,-nbitq), 
to_sfixed(467050275.0/4294967296.0,1,-nbitq), 
to_sfixed(-451290365.0/4294967296.0,1,-nbitq), 
to_sfixed(125969609.0/4294967296.0,1,-nbitq), 
to_sfixed(-204244803.0/4294967296.0,1,-nbitq), 
to_sfixed(156092481.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-205971380.0/4294967296.0,1,-nbitq), 
to_sfixed(1157792990.0/4294967296.0,1,-nbitq), 
to_sfixed(-1424370977.0/4294967296.0,1,-nbitq), 
to_sfixed(-1777244846.0/4294967296.0,1,-nbitq), 
to_sfixed(193306616.0/4294967296.0,1,-nbitq), 
to_sfixed(-63508008.0/4294967296.0,1,-nbitq), 
to_sfixed(-279848789.0/4294967296.0,1,-nbitq), 
to_sfixed(307305414.0/4294967296.0,1,-nbitq), 
to_sfixed(-144905339.0/4294967296.0,1,-nbitq), 
to_sfixed(199751220.0/4294967296.0,1,-nbitq), 
to_sfixed(150348962.0/4294967296.0,1,-nbitq), 
to_sfixed(-160674137.0/4294967296.0,1,-nbitq), 
to_sfixed(1023878864.0/4294967296.0,1,-nbitq), 
to_sfixed(-821668795.0/4294967296.0,1,-nbitq), 
to_sfixed(-26601612.0/4294967296.0,1,-nbitq), 
to_sfixed(-486183851.0/4294967296.0,1,-nbitq), 
to_sfixed(-146347763.0/4294967296.0,1,-nbitq), 
to_sfixed(368164902.0/4294967296.0,1,-nbitq), 
to_sfixed(401086587.0/4294967296.0,1,-nbitq), 
to_sfixed(305924216.0/4294967296.0,1,-nbitq), 
to_sfixed(372055646.0/4294967296.0,1,-nbitq), 
to_sfixed(-53679817.0/4294967296.0,1,-nbitq), 
to_sfixed(-818466872.0/4294967296.0,1,-nbitq), 
to_sfixed(-176886203.0/4294967296.0,1,-nbitq), 
to_sfixed(-106368698.0/4294967296.0,1,-nbitq), 
to_sfixed(715265846.0/4294967296.0,1,-nbitq), 
to_sfixed(-117414205.0/4294967296.0,1,-nbitq), 
to_sfixed(173737207.0/4294967296.0,1,-nbitq), 
to_sfixed(262364816.0/4294967296.0,1,-nbitq), 
to_sfixed(-945050000.0/4294967296.0,1,-nbitq), 
to_sfixed(947875631.0/4294967296.0,1,-nbitq), 
to_sfixed(822372406.0/4294967296.0,1,-nbitq), 
to_sfixed(-396358282.0/4294967296.0,1,-nbitq), 
to_sfixed(260841069.0/4294967296.0,1,-nbitq), 
to_sfixed(-1668211.0/4294967296.0,1,-nbitq), 
to_sfixed(556169634.0/4294967296.0,1,-nbitq), 
to_sfixed(451142451.0/4294967296.0,1,-nbitq), 
to_sfixed(-523387645.0/4294967296.0,1,-nbitq), 
to_sfixed(362820992.0/4294967296.0,1,-nbitq), 
to_sfixed(92594218.0/4294967296.0,1,-nbitq), 
to_sfixed(35870402.0/4294967296.0,1,-nbitq), 
to_sfixed(182593923.0/4294967296.0,1,-nbitq), 
to_sfixed(-728762725.0/4294967296.0,1,-nbitq), 
to_sfixed(-114845965.0/4294967296.0,1,-nbitq), 
to_sfixed(-143278207.0/4294967296.0,1,-nbitq), 
to_sfixed(868734163.0/4294967296.0,1,-nbitq), 
to_sfixed(-210500482.0/4294967296.0,1,-nbitq), 
to_sfixed(128907334.0/4294967296.0,1,-nbitq), 
to_sfixed(-346091554.0/4294967296.0,1,-nbitq), 
to_sfixed(413341452.0/4294967296.0,1,-nbitq), 
to_sfixed(-129005603.0/4294967296.0,1,-nbitq), 
to_sfixed(-1024851781.0/4294967296.0,1,-nbitq), 
to_sfixed(326824955.0/4294967296.0,1,-nbitq), 
to_sfixed(396565327.0/4294967296.0,1,-nbitq), 
to_sfixed(-804070645.0/4294967296.0,1,-nbitq), 
to_sfixed(127037091.0/4294967296.0,1,-nbitq), 
to_sfixed(548977607.0/4294967296.0,1,-nbitq), 
to_sfixed(-24103812.0/4294967296.0,1,-nbitq), 
to_sfixed(202221093.0/4294967296.0,1,-nbitq), 
to_sfixed(-44055092.0/4294967296.0,1,-nbitq), 
to_sfixed(-289194541.0/4294967296.0,1,-nbitq), 
to_sfixed(-930982215.0/4294967296.0,1,-nbitq), 
to_sfixed(92104588.0/4294967296.0,1,-nbitq), 
to_sfixed(-803515598.0/4294967296.0,1,-nbitq), 
to_sfixed(-131279671.0/4294967296.0,1,-nbitq), 
to_sfixed(-32213997.0/4294967296.0,1,-nbitq), 
to_sfixed(-474395733.0/4294967296.0,1,-nbitq), 
to_sfixed(-56069246.0/4294967296.0,1,-nbitq), 
to_sfixed(50384085.0/4294967296.0,1,-nbitq), 
to_sfixed(-235192502.0/4294967296.0,1,-nbitq), 
to_sfixed(461189716.0/4294967296.0,1,-nbitq), 
to_sfixed(236242063.0/4294967296.0,1,-nbitq), 
to_sfixed(-177363896.0/4294967296.0,1,-nbitq), 
to_sfixed(170960148.0/4294967296.0,1,-nbitq), 
to_sfixed(-183224176.0/4294967296.0,1,-nbitq), 
to_sfixed(544741157.0/4294967296.0,1,-nbitq), 
to_sfixed(-703613705.0/4294967296.0,1,-nbitq), 
to_sfixed(164737961.0/4294967296.0,1,-nbitq), 
to_sfixed(-363275061.0/4294967296.0,1,-nbitq), 
to_sfixed(-166248762.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(122547960.0/4294967296.0,1,-nbitq), 
to_sfixed(1304761811.0/4294967296.0,1,-nbitq), 
to_sfixed(-1287693883.0/4294967296.0,1,-nbitq), 
to_sfixed(-760707226.0/4294967296.0,1,-nbitq), 
to_sfixed(118400430.0/4294967296.0,1,-nbitq), 
to_sfixed(-429076358.0/4294967296.0,1,-nbitq), 
to_sfixed(197558192.0/4294967296.0,1,-nbitq), 
to_sfixed(408304405.0/4294967296.0,1,-nbitq), 
to_sfixed(-65936060.0/4294967296.0,1,-nbitq), 
to_sfixed(283657890.0/4294967296.0,1,-nbitq), 
to_sfixed(47728559.0/4294967296.0,1,-nbitq), 
to_sfixed(333459437.0/4294967296.0,1,-nbitq), 
to_sfixed(535777646.0/4294967296.0,1,-nbitq), 
to_sfixed(-94436046.0/4294967296.0,1,-nbitq), 
to_sfixed(-70000329.0/4294967296.0,1,-nbitq), 
to_sfixed(-630830671.0/4294967296.0,1,-nbitq), 
to_sfixed(69639238.0/4294967296.0,1,-nbitq), 
to_sfixed(8468119.0/4294967296.0,1,-nbitq), 
to_sfixed(726682218.0/4294967296.0,1,-nbitq), 
to_sfixed(3342294.0/4294967296.0,1,-nbitq), 
to_sfixed(-390381807.0/4294967296.0,1,-nbitq), 
to_sfixed(512077958.0/4294967296.0,1,-nbitq), 
to_sfixed(-481723471.0/4294967296.0,1,-nbitq), 
to_sfixed(-731825308.0/4294967296.0,1,-nbitq), 
to_sfixed(-38792467.0/4294967296.0,1,-nbitq), 
to_sfixed(185744128.0/4294967296.0,1,-nbitq), 
to_sfixed(-169052838.0/4294967296.0,1,-nbitq), 
to_sfixed(335606117.0/4294967296.0,1,-nbitq), 
to_sfixed(263129055.0/4294967296.0,1,-nbitq), 
to_sfixed(-1085438709.0/4294967296.0,1,-nbitq), 
to_sfixed(545705505.0/4294967296.0,1,-nbitq), 
to_sfixed(607306897.0/4294967296.0,1,-nbitq), 
to_sfixed(57437417.0/4294967296.0,1,-nbitq), 
to_sfixed(133881808.0/4294967296.0,1,-nbitq), 
to_sfixed(550277726.0/4294967296.0,1,-nbitq), 
to_sfixed(511561681.0/4294967296.0,1,-nbitq), 
to_sfixed(-331983375.0/4294967296.0,1,-nbitq), 
to_sfixed(-804354017.0/4294967296.0,1,-nbitq), 
to_sfixed(469876239.0/4294967296.0,1,-nbitq), 
to_sfixed(62458117.0/4294967296.0,1,-nbitq), 
to_sfixed(83201110.0/4294967296.0,1,-nbitq), 
to_sfixed(112887535.0/4294967296.0,1,-nbitq), 
to_sfixed(-306337395.0/4294967296.0,1,-nbitq), 
to_sfixed(-827502746.0/4294967296.0,1,-nbitq), 
to_sfixed(-843380757.0/4294967296.0,1,-nbitq), 
to_sfixed(336463413.0/4294967296.0,1,-nbitq), 
to_sfixed(-117409376.0/4294967296.0,1,-nbitq), 
to_sfixed(-655419001.0/4294967296.0,1,-nbitq), 
to_sfixed(23670618.0/4294967296.0,1,-nbitq), 
to_sfixed(216247344.0/4294967296.0,1,-nbitq), 
to_sfixed(48295312.0/4294967296.0,1,-nbitq), 
to_sfixed(-372340990.0/4294967296.0,1,-nbitq), 
to_sfixed(-293828749.0/4294967296.0,1,-nbitq), 
to_sfixed(742453381.0/4294967296.0,1,-nbitq), 
to_sfixed(-827961309.0/4294967296.0,1,-nbitq), 
to_sfixed(93741020.0/4294967296.0,1,-nbitq), 
to_sfixed(111016264.0/4294967296.0,1,-nbitq), 
to_sfixed(288142136.0/4294967296.0,1,-nbitq), 
to_sfixed(-330397760.0/4294967296.0,1,-nbitq), 
to_sfixed(376192292.0/4294967296.0,1,-nbitq), 
to_sfixed(70356194.0/4294967296.0,1,-nbitq), 
to_sfixed(-947295666.0/4294967296.0,1,-nbitq), 
to_sfixed(-86573964.0/4294967296.0,1,-nbitq), 
to_sfixed(-733883692.0/4294967296.0,1,-nbitq), 
to_sfixed(-36892936.0/4294967296.0,1,-nbitq), 
to_sfixed(392700359.0/4294967296.0,1,-nbitq), 
to_sfixed(-281539702.0/4294967296.0,1,-nbitq), 
to_sfixed(77351491.0/4294967296.0,1,-nbitq), 
to_sfixed(110326525.0/4294967296.0,1,-nbitq), 
to_sfixed(439534857.0/4294967296.0,1,-nbitq), 
to_sfixed(82398065.0/4294967296.0,1,-nbitq), 
to_sfixed(249552081.0/4294967296.0,1,-nbitq), 
to_sfixed(273131525.0/4294967296.0,1,-nbitq), 
to_sfixed(-284706260.0/4294967296.0,1,-nbitq), 
to_sfixed(499671208.0/4294967296.0,1,-nbitq), 
to_sfixed(171807439.0/4294967296.0,1,-nbitq), 
to_sfixed(-939829652.0/4294967296.0,1,-nbitq), 
to_sfixed(-382422679.0/4294967296.0,1,-nbitq), 
to_sfixed(105303513.0/4294967296.0,1,-nbitq), 
to_sfixed(166736862.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-1612125.0/4294967296.0,1,-nbitq), 
to_sfixed(741531094.0/4294967296.0,1,-nbitq), 
to_sfixed(-806506403.0/4294967296.0,1,-nbitq), 
to_sfixed(-678014367.0/4294967296.0,1,-nbitq), 
to_sfixed(-524748022.0/4294967296.0,1,-nbitq), 
to_sfixed(-430120647.0/4294967296.0,1,-nbitq), 
to_sfixed(156284848.0/4294967296.0,1,-nbitq), 
to_sfixed(96745016.0/4294967296.0,1,-nbitq), 
to_sfixed(-271006036.0/4294967296.0,1,-nbitq), 
to_sfixed(-281354140.0/4294967296.0,1,-nbitq), 
to_sfixed(717715348.0/4294967296.0,1,-nbitq), 
to_sfixed(669718584.0/4294967296.0,1,-nbitq), 
to_sfixed(151812445.0/4294967296.0,1,-nbitq), 
to_sfixed(-200506545.0/4294967296.0,1,-nbitq), 
to_sfixed(306388426.0/4294967296.0,1,-nbitq), 
to_sfixed(-656350452.0/4294967296.0,1,-nbitq), 
to_sfixed(77465533.0/4294967296.0,1,-nbitq), 
to_sfixed(-297760771.0/4294967296.0,1,-nbitq), 
to_sfixed(192748397.0/4294967296.0,1,-nbitq), 
to_sfixed(480417539.0/4294967296.0,1,-nbitq), 
to_sfixed(286974136.0/4294967296.0,1,-nbitq), 
to_sfixed(-366455905.0/4294967296.0,1,-nbitq), 
to_sfixed(-531624800.0/4294967296.0,1,-nbitq), 
to_sfixed(-620015939.0/4294967296.0,1,-nbitq), 
to_sfixed(292490020.0/4294967296.0,1,-nbitq), 
to_sfixed(495941189.0/4294967296.0,1,-nbitq), 
to_sfixed(-460351708.0/4294967296.0,1,-nbitq), 
to_sfixed(200318910.0/4294967296.0,1,-nbitq), 
to_sfixed(-268498696.0/4294967296.0,1,-nbitq), 
to_sfixed(-350637472.0/4294967296.0,1,-nbitq), 
to_sfixed(203877196.0/4294967296.0,1,-nbitq), 
to_sfixed(923889179.0/4294967296.0,1,-nbitq), 
to_sfixed(229751101.0/4294967296.0,1,-nbitq), 
to_sfixed(167107296.0/4294967296.0,1,-nbitq), 
to_sfixed(-258294768.0/4294967296.0,1,-nbitq), 
to_sfixed(379342864.0/4294967296.0,1,-nbitq), 
to_sfixed(-767421550.0/4294967296.0,1,-nbitq), 
to_sfixed(-255956970.0/4294967296.0,1,-nbitq), 
to_sfixed(57900815.0/4294967296.0,1,-nbitq), 
to_sfixed(-268321594.0/4294967296.0,1,-nbitq), 
to_sfixed(-110054571.0/4294967296.0,1,-nbitq), 
to_sfixed(-605305381.0/4294967296.0,1,-nbitq), 
to_sfixed(100656114.0/4294967296.0,1,-nbitq), 
to_sfixed(-1108824363.0/4294967296.0,1,-nbitq), 
to_sfixed(-93171771.0/4294967296.0,1,-nbitq), 
to_sfixed(-567613725.0/4294967296.0,1,-nbitq), 
to_sfixed(307629159.0/4294967296.0,1,-nbitq), 
to_sfixed(138776361.0/4294967296.0,1,-nbitq), 
to_sfixed(-515132652.0/4294967296.0,1,-nbitq), 
to_sfixed(65003177.0/4294967296.0,1,-nbitq), 
to_sfixed(-108594153.0/4294967296.0,1,-nbitq), 
to_sfixed(-359393987.0/4294967296.0,1,-nbitq), 
to_sfixed(-227998693.0/4294967296.0,1,-nbitq), 
to_sfixed(411746307.0/4294967296.0,1,-nbitq), 
to_sfixed(-233250631.0/4294967296.0,1,-nbitq), 
to_sfixed(55107608.0/4294967296.0,1,-nbitq), 
to_sfixed(539651213.0/4294967296.0,1,-nbitq), 
to_sfixed(-566325215.0/4294967296.0,1,-nbitq), 
to_sfixed(-287977203.0/4294967296.0,1,-nbitq), 
to_sfixed(-224981918.0/4294967296.0,1,-nbitq), 
to_sfixed(-241807866.0/4294967296.0,1,-nbitq), 
to_sfixed(-643256463.0/4294967296.0,1,-nbitq), 
to_sfixed(386539592.0/4294967296.0,1,-nbitq), 
to_sfixed(-466993827.0/4294967296.0,1,-nbitq), 
to_sfixed(-336709842.0/4294967296.0,1,-nbitq), 
to_sfixed(-217679081.0/4294967296.0,1,-nbitq), 
to_sfixed(-451869393.0/4294967296.0,1,-nbitq), 
to_sfixed(-784403018.0/4294967296.0,1,-nbitq), 
to_sfixed(-50393741.0/4294967296.0,1,-nbitq), 
to_sfixed(205603623.0/4294967296.0,1,-nbitq), 
to_sfixed(295019116.0/4294967296.0,1,-nbitq), 
to_sfixed(216998710.0/4294967296.0,1,-nbitq), 
to_sfixed(-212311134.0/4294967296.0,1,-nbitq), 
to_sfixed(6366725.0/4294967296.0,1,-nbitq), 
to_sfixed(130078600.0/4294967296.0,1,-nbitq), 
to_sfixed(426240.0/4294967296.0,1,-nbitq), 
to_sfixed(-523993974.0/4294967296.0,1,-nbitq), 
to_sfixed(-396257003.0/4294967296.0,1,-nbitq), 
to_sfixed(-466270629.0/4294967296.0,1,-nbitq), 
to_sfixed(-197666263.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(224329911.0/4294967296.0,1,-nbitq), 
to_sfixed(775810243.0/4294967296.0,1,-nbitq), 
to_sfixed(-864731774.0/4294967296.0,1,-nbitq), 
to_sfixed(93749000.0/4294967296.0,1,-nbitq), 
to_sfixed(-256637671.0/4294967296.0,1,-nbitq), 
to_sfixed(-30715714.0/4294967296.0,1,-nbitq), 
to_sfixed(138488663.0/4294967296.0,1,-nbitq), 
to_sfixed(382190799.0/4294967296.0,1,-nbitq), 
to_sfixed(-269119692.0/4294967296.0,1,-nbitq), 
to_sfixed(-233367392.0/4294967296.0,1,-nbitq), 
to_sfixed(893641765.0/4294967296.0,1,-nbitq), 
to_sfixed(18864935.0/4294967296.0,1,-nbitq), 
to_sfixed(497349000.0/4294967296.0,1,-nbitq), 
to_sfixed(-914037819.0/4294967296.0,1,-nbitq), 
to_sfixed(74286149.0/4294967296.0,1,-nbitq), 
to_sfixed(-94617957.0/4294967296.0,1,-nbitq), 
to_sfixed(367406114.0/4294967296.0,1,-nbitq), 
to_sfixed(225146462.0/4294967296.0,1,-nbitq), 
to_sfixed(373561667.0/4294967296.0,1,-nbitq), 
to_sfixed(51681274.0/4294967296.0,1,-nbitq), 
to_sfixed(9824620.0/4294967296.0,1,-nbitq), 
to_sfixed(519854870.0/4294967296.0,1,-nbitq), 
to_sfixed(-268043888.0/4294967296.0,1,-nbitq), 
to_sfixed(-666824158.0/4294967296.0,1,-nbitq), 
to_sfixed(306084620.0/4294967296.0,1,-nbitq), 
to_sfixed(528079365.0/4294967296.0,1,-nbitq), 
to_sfixed(-808958257.0/4294967296.0,1,-nbitq), 
to_sfixed(574371049.0/4294967296.0,1,-nbitq), 
to_sfixed(13135085.0/4294967296.0,1,-nbitq), 
to_sfixed(-244051219.0/4294967296.0,1,-nbitq), 
to_sfixed(871762991.0/4294967296.0,1,-nbitq), 
to_sfixed(789835215.0/4294967296.0,1,-nbitq), 
to_sfixed(211529827.0/4294967296.0,1,-nbitq), 
to_sfixed(-110866145.0/4294967296.0,1,-nbitq), 
to_sfixed(163687556.0/4294967296.0,1,-nbitq), 
to_sfixed(57290421.0/4294967296.0,1,-nbitq), 
to_sfixed(-325306254.0/4294967296.0,1,-nbitq), 
to_sfixed(-197357092.0/4294967296.0,1,-nbitq), 
to_sfixed(157579085.0/4294967296.0,1,-nbitq), 
to_sfixed(89013069.0/4294967296.0,1,-nbitq), 
to_sfixed(518909133.0/4294967296.0,1,-nbitq), 
to_sfixed(-215505602.0/4294967296.0,1,-nbitq), 
to_sfixed(-692123006.0/4294967296.0,1,-nbitq), 
to_sfixed(-353591936.0/4294967296.0,1,-nbitq), 
to_sfixed(100544200.0/4294967296.0,1,-nbitq), 
to_sfixed(-492789449.0/4294967296.0,1,-nbitq), 
to_sfixed(177821916.0/4294967296.0,1,-nbitq), 
to_sfixed(-126408993.0/4294967296.0,1,-nbitq), 
to_sfixed(-329995824.0/4294967296.0,1,-nbitq), 
to_sfixed(-9568649.0/4294967296.0,1,-nbitq), 
to_sfixed(-146221208.0/4294967296.0,1,-nbitq), 
to_sfixed(-7315429.0/4294967296.0,1,-nbitq), 
to_sfixed(-231547536.0/4294967296.0,1,-nbitq), 
to_sfixed(405756450.0/4294967296.0,1,-nbitq), 
to_sfixed(-29471808.0/4294967296.0,1,-nbitq), 
to_sfixed(-422614209.0/4294967296.0,1,-nbitq), 
to_sfixed(-104863476.0/4294967296.0,1,-nbitq), 
to_sfixed(-266281540.0/4294967296.0,1,-nbitq), 
to_sfixed(-6828222.0/4294967296.0,1,-nbitq), 
to_sfixed(238049659.0/4294967296.0,1,-nbitq), 
to_sfixed(-457491703.0/4294967296.0,1,-nbitq), 
to_sfixed(-694478629.0/4294967296.0,1,-nbitq), 
to_sfixed(-162877313.0/4294967296.0,1,-nbitq), 
to_sfixed(97475106.0/4294967296.0,1,-nbitq), 
to_sfixed(-280076397.0/4294967296.0,1,-nbitq), 
to_sfixed(196277720.0/4294967296.0,1,-nbitq), 
to_sfixed(-673561573.0/4294967296.0,1,-nbitq), 
to_sfixed(-193683392.0/4294967296.0,1,-nbitq), 
to_sfixed(-319463926.0/4294967296.0,1,-nbitq), 
to_sfixed(-136962112.0/4294967296.0,1,-nbitq), 
to_sfixed(372438751.0/4294967296.0,1,-nbitq), 
to_sfixed(180459219.0/4294967296.0,1,-nbitq), 
to_sfixed(34717672.0/4294967296.0,1,-nbitq), 
to_sfixed(-191728710.0/4294967296.0,1,-nbitq), 
to_sfixed(-198560076.0/4294967296.0,1,-nbitq), 
to_sfixed(173704376.0/4294967296.0,1,-nbitq), 
to_sfixed(-447807997.0/4294967296.0,1,-nbitq), 
to_sfixed(-229868929.0/4294967296.0,1,-nbitq), 
to_sfixed(-42519760.0/4294967296.0,1,-nbitq), 
to_sfixed(-296480755.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-155101972.0/4294967296.0,1,-nbitq), 
to_sfixed(298754496.0/4294967296.0,1,-nbitq), 
to_sfixed(-423706469.0/4294967296.0,1,-nbitq), 
to_sfixed(271908722.0/4294967296.0,1,-nbitq), 
to_sfixed(193869808.0/4294967296.0,1,-nbitq), 
to_sfixed(179194551.0/4294967296.0,1,-nbitq), 
to_sfixed(50650858.0/4294967296.0,1,-nbitq), 
to_sfixed(49072357.0/4294967296.0,1,-nbitq), 
to_sfixed(-587076974.0/4294967296.0,1,-nbitq), 
to_sfixed(212567255.0/4294967296.0,1,-nbitq), 
to_sfixed(755476058.0/4294967296.0,1,-nbitq), 
to_sfixed(30260481.0/4294967296.0,1,-nbitq), 
to_sfixed(438230094.0/4294967296.0,1,-nbitq), 
to_sfixed(-1126868143.0/4294967296.0,1,-nbitq), 
to_sfixed(349516689.0/4294967296.0,1,-nbitq), 
to_sfixed(-487009121.0/4294967296.0,1,-nbitq), 
to_sfixed(-33105618.0/4294967296.0,1,-nbitq), 
to_sfixed(154330165.0/4294967296.0,1,-nbitq), 
to_sfixed(550929244.0/4294967296.0,1,-nbitq), 
to_sfixed(112423032.0/4294967296.0,1,-nbitq), 
to_sfixed(-38237197.0/4294967296.0,1,-nbitq), 
to_sfixed(281560816.0/4294967296.0,1,-nbitq), 
to_sfixed(-490206324.0/4294967296.0,1,-nbitq), 
to_sfixed(147095930.0/4294967296.0,1,-nbitq), 
to_sfixed(-67601754.0/4294967296.0,1,-nbitq), 
to_sfixed(305209513.0/4294967296.0,1,-nbitq), 
to_sfixed(-564714395.0/4294967296.0,1,-nbitq), 
to_sfixed(473177965.0/4294967296.0,1,-nbitq), 
to_sfixed(137195687.0/4294967296.0,1,-nbitq), 
to_sfixed(238640793.0/4294967296.0,1,-nbitq), 
to_sfixed(-295078633.0/4294967296.0,1,-nbitq), 
to_sfixed(92159587.0/4294967296.0,1,-nbitq), 
to_sfixed(129606119.0/4294967296.0,1,-nbitq), 
to_sfixed(-382781404.0/4294967296.0,1,-nbitq), 
to_sfixed(99136703.0/4294967296.0,1,-nbitq), 
to_sfixed(-289729396.0/4294967296.0,1,-nbitq), 
to_sfixed(-518060031.0/4294967296.0,1,-nbitq), 
to_sfixed(72379293.0/4294967296.0,1,-nbitq), 
to_sfixed(386896255.0/4294967296.0,1,-nbitq), 
to_sfixed(63227149.0/4294967296.0,1,-nbitq), 
to_sfixed(224613768.0/4294967296.0,1,-nbitq), 
to_sfixed(-248817368.0/4294967296.0,1,-nbitq), 
to_sfixed(34134100.0/4294967296.0,1,-nbitq), 
to_sfixed(-210603810.0/4294967296.0,1,-nbitq), 
to_sfixed(24851307.0/4294967296.0,1,-nbitq), 
to_sfixed(-312833007.0/4294967296.0,1,-nbitq), 
to_sfixed(80044960.0/4294967296.0,1,-nbitq), 
to_sfixed(-155431625.0/4294967296.0,1,-nbitq), 
to_sfixed(44185709.0/4294967296.0,1,-nbitq), 
to_sfixed(-365542134.0/4294967296.0,1,-nbitq), 
to_sfixed(13895629.0/4294967296.0,1,-nbitq), 
to_sfixed(-175396192.0/4294967296.0,1,-nbitq), 
to_sfixed(51667824.0/4294967296.0,1,-nbitq), 
to_sfixed(11205805.0/4294967296.0,1,-nbitq), 
to_sfixed(118768126.0/4294967296.0,1,-nbitq), 
to_sfixed(-227459094.0/4294967296.0,1,-nbitq), 
to_sfixed(181193221.0/4294967296.0,1,-nbitq), 
to_sfixed(109635314.0/4294967296.0,1,-nbitq), 
to_sfixed(383327075.0/4294967296.0,1,-nbitq), 
to_sfixed(140771177.0/4294967296.0,1,-nbitq), 
to_sfixed(331744796.0/4294967296.0,1,-nbitq), 
to_sfixed(-440960935.0/4294967296.0,1,-nbitq), 
to_sfixed(174948920.0/4294967296.0,1,-nbitq), 
to_sfixed(-579665819.0/4294967296.0,1,-nbitq), 
to_sfixed(293010842.0/4294967296.0,1,-nbitq), 
to_sfixed(132545259.0/4294967296.0,1,-nbitq), 
to_sfixed(348375740.0/4294967296.0,1,-nbitq), 
to_sfixed(3758276.0/4294967296.0,1,-nbitq), 
to_sfixed(412586109.0/4294967296.0,1,-nbitq), 
to_sfixed(70723139.0/4294967296.0,1,-nbitq), 
to_sfixed(323900510.0/4294967296.0,1,-nbitq), 
to_sfixed(223101358.0/4294967296.0,1,-nbitq), 
to_sfixed(-116186194.0/4294967296.0,1,-nbitq), 
to_sfixed(-167008835.0/4294967296.0,1,-nbitq), 
to_sfixed(153799233.0/4294967296.0,1,-nbitq), 
to_sfixed(156326028.0/4294967296.0,1,-nbitq), 
to_sfixed(-439792293.0/4294967296.0,1,-nbitq), 
to_sfixed(54003945.0/4294967296.0,1,-nbitq), 
to_sfixed(-766486253.0/4294967296.0,1,-nbitq), 
to_sfixed(-219179595.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(204980528.0/4294967296.0,1,-nbitq), 
to_sfixed(411080587.0/4294967296.0,1,-nbitq), 
to_sfixed(-389174865.0/4294967296.0,1,-nbitq), 
to_sfixed(-448859944.0/4294967296.0,1,-nbitq), 
to_sfixed(-189873451.0/4294967296.0,1,-nbitq), 
to_sfixed(393821194.0/4294967296.0,1,-nbitq), 
to_sfixed(-317807829.0/4294967296.0,1,-nbitq), 
to_sfixed(109074175.0/4294967296.0,1,-nbitq), 
to_sfixed(-35434293.0/4294967296.0,1,-nbitq), 
to_sfixed(-211932709.0/4294967296.0,1,-nbitq), 
to_sfixed(37084559.0/4294967296.0,1,-nbitq), 
to_sfixed(-381263715.0/4294967296.0,1,-nbitq), 
to_sfixed(-31400830.0/4294967296.0,1,-nbitq), 
to_sfixed(154178163.0/4294967296.0,1,-nbitq), 
to_sfixed(-134322643.0/4294967296.0,1,-nbitq), 
to_sfixed(170738560.0/4294967296.0,1,-nbitq), 
to_sfixed(-302779827.0/4294967296.0,1,-nbitq), 
to_sfixed(-43850528.0/4294967296.0,1,-nbitq), 
to_sfixed(454717466.0/4294967296.0,1,-nbitq), 
to_sfixed(-144546515.0/4294967296.0,1,-nbitq), 
to_sfixed(30643172.0/4294967296.0,1,-nbitq), 
to_sfixed(294061408.0/4294967296.0,1,-nbitq), 
to_sfixed(256851083.0/4294967296.0,1,-nbitq), 
to_sfixed(132801806.0/4294967296.0,1,-nbitq), 
to_sfixed(326036573.0/4294967296.0,1,-nbitq), 
to_sfixed(206137191.0/4294967296.0,1,-nbitq), 
to_sfixed(-212885367.0/4294967296.0,1,-nbitq), 
to_sfixed(-65708433.0/4294967296.0,1,-nbitq), 
to_sfixed(617423847.0/4294967296.0,1,-nbitq), 
to_sfixed(-373646736.0/4294967296.0,1,-nbitq), 
to_sfixed(135845661.0/4294967296.0,1,-nbitq), 
to_sfixed(-75280250.0/4294967296.0,1,-nbitq), 
to_sfixed(-185874595.0/4294967296.0,1,-nbitq), 
to_sfixed(13361365.0/4294967296.0,1,-nbitq), 
to_sfixed(-135983154.0/4294967296.0,1,-nbitq), 
to_sfixed(-22573426.0/4294967296.0,1,-nbitq), 
to_sfixed(56069093.0/4294967296.0,1,-nbitq), 
to_sfixed(-91980965.0/4294967296.0,1,-nbitq), 
to_sfixed(-46770310.0/4294967296.0,1,-nbitq), 
to_sfixed(84467713.0/4294967296.0,1,-nbitq), 
to_sfixed(-97010187.0/4294967296.0,1,-nbitq), 
to_sfixed(405586051.0/4294967296.0,1,-nbitq), 
to_sfixed(-327813435.0/4294967296.0,1,-nbitq), 
to_sfixed(177474585.0/4294967296.0,1,-nbitq), 
to_sfixed(-30632406.0/4294967296.0,1,-nbitq), 
to_sfixed(-316720958.0/4294967296.0,1,-nbitq), 
to_sfixed(69659243.0/4294967296.0,1,-nbitq), 
to_sfixed(-187502271.0/4294967296.0,1,-nbitq), 
to_sfixed(-158936234.0/4294967296.0,1,-nbitq), 
to_sfixed(123090849.0/4294967296.0,1,-nbitq), 
to_sfixed(-297407291.0/4294967296.0,1,-nbitq), 
to_sfixed(325888014.0/4294967296.0,1,-nbitq), 
to_sfixed(-42842126.0/4294967296.0,1,-nbitq), 
to_sfixed(159075933.0/4294967296.0,1,-nbitq), 
to_sfixed(217385325.0/4294967296.0,1,-nbitq), 
to_sfixed(-177062639.0/4294967296.0,1,-nbitq), 
to_sfixed(600151308.0/4294967296.0,1,-nbitq), 
to_sfixed(-154838822.0/4294967296.0,1,-nbitq), 
to_sfixed(280728707.0/4294967296.0,1,-nbitq), 
to_sfixed(-27452376.0/4294967296.0,1,-nbitq), 
to_sfixed(17180441.0/4294967296.0,1,-nbitq), 
to_sfixed(-389020513.0/4294967296.0,1,-nbitq), 
to_sfixed(310219220.0/4294967296.0,1,-nbitq), 
to_sfixed(-81126680.0/4294967296.0,1,-nbitq), 
to_sfixed(236707923.0/4294967296.0,1,-nbitq), 
to_sfixed(-38131398.0/4294967296.0,1,-nbitq), 
to_sfixed(456821081.0/4294967296.0,1,-nbitq), 
to_sfixed(276638065.0/4294967296.0,1,-nbitq), 
to_sfixed(386344131.0/4294967296.0,1,-nbitq), 
to_sfixed(488207095.0/4294967296.0,1,-nbitq), 
to_sfixed(162750536.0/4294967296.0,1,-nbitq), 
to_sfixed(205603420.0/4294967296.0,1,-nbitq), 
to_sfixed(332200730.0/4294967296.0,1,-nbitq), 
to_sfixed(284917216.0/4294967296.0,1,-nbitq), 
to_sfixed(127128568.0/4294967296.0,1,-nbitq), 
to_sfixed(-75458493.0/4294967296.0,1,-nbitq), 
to_sfixed(200790951.0/4294967296.0,1,-nbitq), 
to_sfixed(-285332732.0/4294967296.0,1,-nbitq), 
to_sfixed(39404810.0/4294967296.0,1,-nbitq), 
to_sfixed(181661157.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(312807883.0/4294967296.0,1,-nbitq), 
to_sfixed(-486508003.0/4294967296.0,1,-nbitq), 
to_sfixed(49710877.0/4294967296.0,1,-nbitq), 
to_sfixed(216383464.0/4294967296.0,1,-nbitq), 
to_sfixed(372979838.0/4294967296.0,1,-nbitq), 
to_sfixed(-132359832.0/4294967296.0,1,-nbitq), 
to_sfixed(-123219491.0/4294967296.0,1,-nbitq), 
to_sfixed(-366468600.0/4294967296.0,1,-nbitq), 
to_sfixed(-37313440.0/4294967296.0,1,-nbitq), 
to_sfixed(-151666631.0/4294967296.0,1,-nbitq), 
to_sfixed(344368864.0/4294967296.0,1,-nbitq), 
to_sfixed(416146474.0/4294967296.0,1,-nbitq), 
to_sfixed(309271266.0/4294967296.0,1,-nbitq), 
to_sfixed(-470406695.0/4294967296.0,1,-nbitq), 
to_sfixed(-93931472.0/4294967296.0,1,-nbitq), 
to_sfixed(-230964906.0/4294967296.0,1,-nbitq), 
to_sfixed(149445375.0/4294967296.0,1,-nbitq), 
to_sfixed(121919957.0/4294967296.0,1,-nbitq), 
to_sfixed(325973273.0/4294967296.0,1,-nbitq), 
to_sfixed(331182241.0/4294967296.0,1,-nbitq), 
to_sfixed(-220635255.0/4294967296.0,1,-nbitq), 
to_sfixed(-202274195.0/4294967296.0,1,-nbitq), 
to_sfixed(534453883.0/4294967296.0,1,-nbitq), 
to_sfixed(279767353.0/4294967296.0,1,-nbitq), 
to_sfixed(229407293.0/4294967296.0,1,-nbitq), 
to_sfixed(172328305.0/4294967296.0,1,-nbitq), 
to_sfixed(334452941.0/4294967296.0,1,-nbitq), 
to_sfixed(-230883321.0/4294967296.0,1,-nbitq), 
to_sfixed(543728595.0/4294967296.0,1,-nbitq), 
to_sfixed(165736721.0/4294967296.0,1,-nbitq), 
to_sfixed(-374468711.0/4294967296.0,1,-nbitq), 
to_sfixed(-312487006.0/4294967296.0,1,-nbitq), 
to_sfixed(166551127.0/4294967296.0,1,-nbitq), 
to_sfixed(-132737614.0/4294967296.0,1,-nbitq), 
to_sfixed(130143133.0/4294967296.0,1,-nbitq), 
to_sfixed(-58717242.0/4294967296.0,1,-nbitq), 
to_sfixed(49758436.0/4294967296.0,1,-nbitq), 
to_sfixed(205366784.0/4294967296.0,1,-nbitq), 
to_sfixed(347753966.0/4294967296.0,1,-nbitq), 
to_sfixed(-25322717.0/4294967296.0,1,-nbitq), 
to_sfixed(504132526.0/4294967296.0,1,-nbitq), 
to_sfixed(409556886.0/4294967296.0,1,-nbitq), 
to_sfixed(-316564873.0/4294967296.0,1,-nbitq), 
to_sfixed(-80796289.0/4294967296.0,1,-nbitq), 
to_sfixed(-191549054.0/4294967296.0,1,-nbitq), 
to_sfixed(308795765.0/4294967296.0,1,-nbitq), 
to_sfixed(-266021984.0/4294967296.0,1,-nbitq), 
to_sfixed(-41223735.0/4294967296.0,1,-nbitq), 
to_sfixed(-66522943.0/4294967296.0,1,-nbitq), 
to_sfixed(119705461.0/4294967296.0,1,-nbitq), 
to_sfixed(-163634045.0/4294967296.0,1,-nbitq), 
to_sfixed(-180676080.0/4294967296.0,1,-nbitq), 
to_sfixed(204234119.0/4294967296.0,1,-nbitq), 
to_sfixed(383096168.0/4294967296.0,1,-nbitq), 
to_sfixed(310442283.0/4294967296.0,1,-nbitq), 
to_sfixed(-77495414.0/4294967296.0,1,-nbitq), 
to_sfixed(149518889.0/4294967296.0,1,-nbitq), 
to_sfixed(8615009.0/4294967296.0,1,-nbitq), 
to_sfixed(271318256.0/4294967296.0,1,-nbitq), 
to_sfixed(-218772158.0/4294967296.0,1,-nbitq), 
to_sfixed(219455615.0/4294967296.0,1,-nbitq), 
to_sfixed(-149507736.0/4294967296.0,1,-nbitq), 
to_sfixed(279934104.0/4294967296.0,1,-nbitq), 
to_sfixed(-126252096.0/4294967296.0,1,-nbitq), 
to_sfixed(-245119090.0/4294967296.0,1,-nbitq), 
to_sfixed(-227613378.0/4294967296.0,1,-nbitq), 
to_sfixed(219687713.0/4294967296.0,1,-nbitq), 
to_sfixed(243600470.0/4294967296.0,1,-nbitq), 
to_sfixed(399958117.0/4294967296.0,1,-nbitq), 
to_sfixed(191261185.0/4294967296.0,1,-nbitq), 
to_sfixed(-478095567.0/4294967296.0,1,-nbitq), 
to_sfixed(-219553716.0/4294967296.0,1,-nbitq), 
to_sfixed(41267814.0/4294967296.0,1,-nbitq), 
to_sfixed(402035633.0/4294967296.0,1,-nbitq), 
to_sfixed(206205660.0/4294967296.0,1,-nbitq), 
to_sfixed(111142418.0/4294967296.0,1,-nbitq), 
to_sfixed(-417071188.0/4294967296.0,1,-nbitq), 
to_sfixed(289155904.0/4294967296.0,1,-nbitq), 
to_sfixed(4198170.0/4294967296.0,1,-nbitq), 
to_sfixed(148073942.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-130772313.0/4294967296.0,1,-nbitq), 
to_sfixed(237094044.0/4294967296.0,1,-nbitq), 
to_sfixed(186836204.0/4294967296.0,1,-nbitq), 
to_sfixed(34817186.0/4294967296.0,1,-nbitq), 
to_sfixed(160532184.0/4294967296.0,1,-nbitq), 
to_sfixed(-155767684.0/4294967296.0,1,-nbitq), 
to_sfixed(41302684.0/4294967296.0,1,-nbitq), 
to_sfixed(-403035478.0/4294967296.0,1,-nbitq), 
to_sfixed(-375476428.0/4294967296.0,1,-nbitq), 
to_sfixed(328974454.0/4294967296.0,1,-nbitq), 
to_sfixed(122432494.0/4294967296.0,1,-nbitq), 
to_sfixed(-118409055.0/4294967296.0,1,-nbitq), 
to_sfixed(61393654.0/4294967296.0,1,-nbitq), 
to_sfixed(-459501149.0/4294967296.0,1,-nbitq), 
to_sfixed(353446578.0/4294967296.0,1,-nbitq), 
to_sfixed(-48524085.0/4294967296.0,1,-nbitq), 
to_sfixed(26874573.0/4294967296.0,1,-nbitq), 
to_sfixed(-220373430.0/4294967296.0,1,-nbitq), 
to_sfixed(251327491.0/4294967296.0,1,-nbitq), 
to_sfixed(-437870071.0/4294967296.0,1,-nbitq), 
to_sfixed(376190417.0/4294967296.0,1,-nbitq), 
to_sfixed(243715825.0/4294967296.0,1,-nbitq), 
to_sfixed(13649927.0/4294967296.0,1,-nbitq), 
to_sfixed(78339456.0/4294967296.0,1,-nbitq), 
to_sfixed(106043038.0/4294967296.0,1,-nbitq), 
to_sfixed(-152150692.0/4294967296.0,1,-nbitq), 
to_sfixed(-282671664.0/4294967296.0,1,-nbitq), 
to_sfixed(99219345.0/4294967296.0,1,-nbitq), 
to_sfixed(81147379.0/4294967296.0,1,-nbitq), 
to_sfixed(244005965.0/4294967296.0,1,-nbitq), 
to_sfixed(-71108661.0/4294967296.0,1,-nbitq), 
to_sfixed(-227743627.0/4294967296.0,1,-nbitq), 
to_sfixed(290612194.0/4294967296.0,1,-nbitq), 
to_sfixed(-304782605.0/4294967296.0,1,-nbitq), 
to_sfixed(87972574.0/4294967296.0,1,-nbitq), 
to_sfixed(154128449.0/4294967296.0,1,-nbitq), 
to_sfixed(-54126860.0/4294967296.0,1,-nbitq), 
to_sfixed(314653379.0/4294967296.0,1,-nbitq), 
to_sfixed(-152905970.0/4294967296.0,1,-nbitq), 
to_sfixed(-10442517.0/4294967296.0,1,-nbitq), 
to_sfixed(387573345.0/4294967296.0,1,-nbitq), 
to_sfixed(541595161.0/4294967296.0,1,-nbitq), 
to_sfixed(34203106.0/4294967296.0,1,-nbitq), 
to_sfixed(-379490861.0/4294967296.0,1,-nbitq), 
to_sfixed(322057283.0/4294967296.0,1,-nbitq), 
to_sfixed(301858233.0/4294967296.0,1,-nbitq), 
to_sfixed(167136891.0/4294967296.0,1,-nbitq), 
to_sfixed(-139705100.0/4294967296.0,1,-nbitq), 
to_sfixed(208675247.0/4294967296.0,1,-nbitq), 
to_sfixed(176978670.0/4294967296.0,1,-nbitq), 
to_sfixed(-223797117.0/4294967296.0,1,-nbitq), 
to_sfixed(-242372461.0/4294967296.0,1,-nbitq), 
to_sfixed(-531582216.0/4294967296.0,1,-nbitq), 
to_sfixed(53916753.0/4294967296.0,1,-nbitq), 
to_sfixed(314251791.0/4294967296.0,1,-nbitq), 
to_sfixed(-130243053.0/4294967296.0,1,-nbitq), 
to_sfixed(445533833.0/4294967296.0,1,-nbitq), 
to_sfixed(23524967.0/4294967296.0,1,-nbitq), 
to_sfixed(222960058.0/4294967296.0,1,-nbitq), 
to_sfixed(247945345.0/4294967296.0,1,-nbitq), 
to_sfixed(-141158910.0/4294967296.0,1,-nbitq), 
to_sfixed(-349706028.0/4294967296.0,1,-nbitq), 
to_sfixed(-358713277.0/4294967296.0,1,-nbitq), 
to_sfixed(-300922300.0/4294967296.0,1,-nbitq), 
to_sfixed(-210076783.0/4294967296.0,1,-nbitq), 
to_sfixed(-3124104.0/4294967296.0,1,-nbitq), 
to_sfixed(224152898.0/4294967296.0,1,-nbitq), 
to_sfixed(-49596654.0/4294967296.0,1,-nbitq), 
to_sfixed(85674971.0/4294967296.0,1,-nbitq), 
to_sfixed(365000271.0/4294967296.0,1,-nbitq), 
to_sfixed(286849158.0/4294967296.0,1,-nbitq), 
to_sfixed(-121555451.0/4294967296.0,1,-nbitq), 
to_sfixed(-409036375.0/4294967296.0,1,-nbitq), 
to_sfixed(294054191.0/4294967296.0,1,-nbitq), 
to_sfixed(-192791985.0/4294967296.0,1,-nbitq), 
to_sfixed(-516420937.0/4294967296.0,1,-nbitq), 
to_sfixed(-164961230.0/4294967296.0,1,-nbitq), 
to_sfixed(-203681975.0/4294967296.0,1,-nbitq), 
to_sfixed(-78113117.0/4294967296.0,1,-nbitq), 
to_sfixed(-15935284.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-259989539.0/4294967296.0,1,-nbitq), 
to_sfixed(58285488.0/4294967296.0,1,-nbitq), 
to_sfixed(-76351673.0/4294967296.0,1,-nbitq), 
to_sfixed(-472109555.0/4294967296.0,1,-nbitq), 
to_sfixed(-300981753.0/4294967296.0,1,-nbitq), 
to_sfixed(112047341.0/4294967296.0,1,-nbitq), 
to_sfixed(260301575.0/4294967296.0,1,-nbitq), 
to_sfixed(-298786939.0/4294967296.0,1,-nbitq), 
to_sfixed(97066789.0/4294967296.0,1,-nbitq), 
to_sfixed(-221102260.0/4294967296.0,1,-nbitq), 
to_sfixed(179352586.0/4294967296.0,1,-nbitq), 
to_sfixed(456150059.0/4294967296.0,1,-nbitq), 
to_sfixed(-126644503.0/4294967296.0,1,-nbitq), 
to_sfixed(58326904.0/4294967296.0,1,-nbitq), 
to_sfixed(123522240.0/4294967296.0,1,-nbitq), 
to_sfixed(-142144123.0/4294967296.0,1,-nbitq), 
to_sfixed(-74838367.0/4294967296.0,1,-nbitq), 
to_sfixed(-302123692.0/4294967296.0,1,-nbitq), 
to_sfixed(-235848960.0/4294967296.0,1,-nbitq), 
to_sfixed(-451379935.0/4294967296.0,1,-nbitq), 
to_sfixed(-158482511.0/4294967296.0,1,-nbitq), 
to_sfixed(-240411194.0/4294967296.0,1,-nbitq), 
to_sfixed(-78293451.0/4294967296.0,1,-nbitq), 
to_sfixed(314158207.0/4294967296.0,1,-nbitq), 
to_sfixed(217760558.0/4294967296.0,1,-nbitq), 
to_sfixed(-94811481.0/4294967296.0,1,-nbitq), 
to_sfixed(-110454426.0/4294967296.0,1,-nbitq), 
to_sfixed(-192238628.0/4294967296.0,1,-nbitq), 
to_sfixed(87478347.0/4294967296.0,1,-nbitq), 
to_sfixed(218578423.0/4294967296.0,1,-nbitq), 
to_sfixed(-365424224.0/4294967296.0,1,-nbitq), 
to_sfixed(-49233863.0/4294967296.0,1,-nbitq), 
to_sfixed(-152396902.0/4294967296.0,1,-nbitq), 
to_sfixed(-436302633.0/4294967296.0,1,-nbitq), 
to_sfixed(-9219592.0/4294967296.0,1,-nbitq), 
to_sfixed(-70706803.0/4294967296.0,1,-nbitq), 
to_sfixed(319938408.0/4294967296.0,1,-nbitq), 
to_sfixed(328839178.0/4294967296.0,1,-nbitq), 
to_sfixed(380238650.0/4294967296.0,1,-nbitq), 
to_sfixed(467914473.0/4294967296.0,1,-nbitq), 
to_sfixed(-308633593.0/4294967296.0,1,-nbitq), 
to_sfixed(457220661.0/4294967296.0,1,-nbitq), 
to_sfixed(42589236.0/4294967296.0,1,-nbitq), 
to_sfixed(67781654.0/4294967296.0,1,-nbitq), 
to_sfixed(-155749449.0/4294967296.0,1,-nbitq), 
to_sfixed(379206272.0/4294967296.0,1,-nbitq), 
to_sfixed(-85885528.0/4294967296.0,1,-nbitq), 
to_sfixed(147032352.0/4294967296.0,1,-nbitq), 
to_sfixed(-404382484.0/4294967296.0,1,-nbitq), 
to_sfixed(24655368.0/4294967296.0,1,-nbitq), 
to_sfixed(268545566.0/4294967296.0,1,-nbitq), 
to_sfixed(-35205781.0/4294967296.0,1,-nbitq), 
to_sfixed(-410462326.0/4294967296.0,1,-nbitq), 
to_sfixed(-74210028.0/4294967296.0,1,-nbitq), 
to_sfixed(291207050.0/4294967296.0,1,-nbitq), 
to_sfixed(-396879618.0/4294967296.0,1,-nbitq), 
to_sfixed(440317204.0/4294967296.0,1,-nbitq), 
to_sfixed(-6022048.0/4294967296.0,1,-nbitq), 
to_sfixed(244942094.0/4294967296.0,1,-nbitq), 
to_sfixed(-106149307.0/4294967296.0,1,-nbitq), 
to_sfixed(130847646.0/4294967296.0,1,-nbitq), 
to_sfixed(142596893.0/4294967296.0,1,-nbitq), 
to_sfixed(175538570.0/4294967296.0,1,-nbitq), 
to_sfixed(117437079.0/4294967296.0,1,-nbitq), 
to_sfixed(362925095.0/4294967296.0,1,-nbitq), 
to_sfixed(-80063263.0/4294967296.0,1,-nbitq), 
to_sfixed(345716488.0/4294967296.0,1,-nbitq), 
to_sfixed(-317965016.0/4294967296.0,1,-nbitq), 
to_sfixed(290698047.0/4294967296.0,1,-nbitq), 
to_sfixed(-130640641.0/4294967296.0,1,-nbitq), 
to_sfixed(227711907.0/4294967296.0,1,-nbitq), 
to_sfixed(-28979185.0/4294967296.0,1,-nbitq), 
to_sfixed(-2547188.0/4294967296.0,1,-nbitq), 
to_sfixed(-236731244.0/4294967296.0,1,-nbitq), 
to_sfixed(452039288.0/4294967296.0,1,-nbitq), 
to_sfixed(47878151.0/4294967296.0,1,-nbitq), 
to_sfixed(-70202059.0/4294967296.0,1,-nbitq), 
to_sfixed(-146059530.0/4294967296.0,1,-nbitq), 
to_sfixed(23897367.0/4294967296.0,1,-nbitq), 
to_sfixed(321213199.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(289463922.0/4294967296.0,1,-nbitq), 
to_sfixed(82252796.0/4294967296.0,1,-nbitq), 
to_sfixed(138291817.0/4294967296.0,1,-nbitq), 
to_sfixed(-142071124.0/4294967296.0,1,-nbitq), 
to_sfixed(302753734.0/4294967296.0,1,-nbitq), 
to_sfixed(95809490.0/4294967296.0,1,-nbitq), 
to_sfixed(-249476290.0/4294967296.0,1,-nbitq), 
to_sfixed(123609249.0/4294967296.0,1,-nbitq), 
to_sfixed(-61448401.0/4294967296.0,1,-nbitq), 
to_sfixed(3160258.0/4294967296.0,1,-nbitq), 
to_sfixed(-7281287.0/4294967296.0,1,-nbitq), 
to_sfixed(-180564586.0/4294967296.0,1,-nbitq), 
to_sfixed(350115533.0/4294967296.0,1,-nbitq), 
to_sfixed(35685356.0/4294967296.0,1,-nbitq), 
to_sfixed(187774899.0/4294967296.0,1,-nbitq), 
to_sfixed(-439606963.0/4294967296.0,1,-nbitq), 
to_sfixed(333208087.0/4294967296.0,1,-nbitq), 
to_sfixed(392594161.0/4294967296.0,1,-nbitq), 
to_sfixed(224342332.0/4294967296.0,1,-nbitq), 
to_sfixed(-456370975.0/4294967296.0,1,-nbitq), 
to_sfixed(-5635753.0/4294967296.0,1,-nbitq), 
to_sfixed(342392262.0/4294967296.0,1,-nbitq), 
to_sfixed(-210816377.0/4294967296.0,1,-nbitq), 
to_sfixed(-214185730.0/4294967296.0,1,-nbitq), 
to_sfixed(119832928.0/4294967296.0,1,-nbitq), 
to_sfixed(21310000.0/4294967296.0,1,-nbitq), 
to_sfixed(-273399179.0/4294967296.0,1,-nbitq), 
to_sfixed(183443218.0/4294967296.0,1,-nbitq), 
to_sfixed(219880061.0/4294967296.0,1,-nbitq), 
to_sfixed(362726619.0/4294967296.0,1,-nbitq), 
to_sfixed(-308620183.0/4294967296.0,1,-nbitq), 
to_sfixed(-8247967.0/4294967296.0,1,-nbitq), 
to_sfixed(366352045.0/4294967296.0,1,-nbitq), 
to_sfixed(88894991.0/4294967296.0,1,-nbitq), 
to_sfixed(-153983294.0/4294967296.0,1,-nbitq), 
to_sfixed(66219593.0/4294967296.0,1,-nbitq), 
to_sfixed(193693040.0/4294967296.0,1,-nbitq), 
to_sfixed(-3564999.0/4294967296.0,1,-nbitq), 
to_sfixed(-254768324.0/4294967296.0,1,-nbitq), 
to_sfixed(-60608235.0/4294967296.0,1,-nbitq), 
to_sfixed(30106413.0/4294967296.0,1,-nbitq), 
to_sfixed(115515548.0/4294967296.0,1,-nbitq), 
to_sfixed(8112522.0/4294967296.0,1,-nbitq), 
to_sfixed(335207228.0/4294967296.0,1,-nbitq), 
to_sfixed(-143624185.0/4294967296.0,1,-nbitq), 
to_sfixed(364568029.0/4294967296.0,1,-nbitq), 
to_sfixed(301592925.0/4294967296.0,1,-nbitq), 
to_sfixed(-528098118.0/4294967296.0,1,-nbitq), 
to_sfixed(361775412.0/4294967296.0,1,-nbitq), 
to_sfixed(-31341032.0/4294967296.0,1,-nbitq), 
to_sfixed(389551823.0/4294967296.0,1,-nbitq), 
to_sfixed(93197741.0/4294967296.0,1,-nbitq), 
to_sfixed(113498697.0/4294967296.0,1,-nbitq), 
to_sfixed(-406629639.0/4294967296.0,1,-nbitq), 
to_sfixed(406123715.0/4294967296.0,1,-nbitq), 
to_sfixed(244777034.0/4294967296.0,1,-nbitq), 
to_sfixed(-161813532.0/4294967296.0,1,-nbitq), 
to_sfixed(215825509.0/4294967296.0,1,-nbitq), 
to_sfixed(28909364.0/4294967296.0,1,-nbitq), 
to_sfixed(-26850841.0/4294967296.0,1,-nbitq), 
to_sfixed(225849222.0/4294967296.0,1,-nbitq), 
to_sfixed(118075390.0/4294967296.0,1,-nbitq), 
to_sfixed(-48990838.0/4294967296.0,1,-nbitq), 
to_sfixed(29989380.0/4294967296.0,1,-nbitq), 
to_sfixed(397128388.0/4294967296.0,1,-nbitq), 
to_sfixed(-334998202.0/4294967296.0,1,-nbitq), 
to_sfixed(265614747.0/4294967296.0,1,-nbitq), 
to_sfixed(72343781.0/4294967296.0,1,-nbitq), 
to_sfixed(282359397.0/4294967296.0,1,-nbitq), 
to_sfixed(-120797631.0/4294967296.0,1,-nbitq), 
to_sfixed(345216671.0/4294967296.0,1,-nbitq), 
to_sfixed(-52044798.0/4294967296.0,1,-nbitq), 
to_sfixed(153494230.0/4294967296.0,1,-nbitq), 
to_sfixed(178438048.0/4294967296.0,1,-nbitq), 
to_sfixed(125585233.0/4294967296.0,1,-nbitq), 
to_sfixed(113787629.0/4294967296.0,1,-nbitq), 
to_sfixed(-309710055.0/4294967296.0,1,-nbitq), 
to_sfixed(74720910.0/4294967296.0,1,-nbitq), 
to_sfixed(-385202349.0/4294967296.0,1,-nbitq), 
to_sfixed(248405986.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-19082961.0/4294967296.0,1,-nbitq), 
to_sfixed(299865253.0/4294967296.0,1,-nbitq), 
to_sfixed(248261500.0/4294967296.0,1,-nbitq), 
to_sfixed(-523456260.0/4294967296.0,1,-nbitq), 
to_sfixed(279981020.0/4294967296.0,1,-nbitq), 
to_sfixed(128079876.0/4294967296.0,1,-nbitq), 
to_sfixed(84828443.0/4294967296.0,1,-nbitq), 
to_sfixed(-104260257.0/4294967296.0,1,-nbitq), 
to_sfixed(-241164714.0/4294967296.0,1,-nbitq), 
to_sfixed(-84551043.0/4294967296.0,1,-nbitq), 
to_sfixed(188481968.0/4294967296.0,1,-nbitq), 
to_sfixed(72260603.0/4294967296.0,1,-nbitq), 
to_sfixed(-93698349.0/4294967296.0,1,-nbitq), 
to_sfixed(681385030.0/4294967296.0,1,-nbitq), 
to_sfixed(-421017830.0/4294967296.0,1,-nbitq), 
to_sfixed(-400418154.0/4294967296.0,1,-nbitq), 
to_sfixed(-273337119.0/4294967296.0,1,-nbitq), 
to_sfixed(-183535399.0/4294967296.0,1,-nbitq), 
to_sfixed(189296789.0/4294967296.0,1,-nbitq), 
to_sfixed(-131116633.0/4294967296.0,1,-nbitq), 
to_sfixed(222182271.0/4294967296.0,1,-nbitq), 
to_sfixed(399806245.0/4294967296.0,1,-nbitq), 
to_sfixed(-134945130.0/4294967296.0,1,-nbitq), 
to_sfixed(531377456.0/4294967296.0,1,-nbitq), 
to_sfixed(-182563734.0/4294967296.0,1,-nbitq), 
to_sfixed(-4583969.0/4294967296.0,1,-nbitq), 
to_sfixed(-185996844.0/4294967296.0,1,-nbitq), 
to_sfixed(-432229585.0/4294967296.0,1,-nbitq), 
to_sfixed(348527731.0/4294967296.0,1,-nbitq), 
to_sfixed(83802560.0/4294967296.0,1,-nbitq), 
to_sfixed(-86773790.0/4294967296.0,1,-nbitq), 
to_sfixed(-295498930.0/4294967296.0,1,-nbitq), 
to_sfixed(312556383.0/4294967296.0,1,-nbitq), 
to_sfixed(-388971859.0/4294967296.0,1,-nbitq), 
to_sfixed(-15932381.0/4294967296.0,1,-nbitq), 
to_sfixed(-306696609.0/4294967296.0,1,-nbitq), 
to_sfixed(271068254.0/4294967296.0,1,-nbitq), 
to_sfixed(-193344485.0/4294967296.0,1,-nbitq), 
to_sfixed(249863231.0/4294967296.0,1,-nbitq), 
to_sfixed(469753017.0/4294967296.0,1,-nbitq), 
to_sfixed(-175739414.0/4294967296.0,1,-nbitq), 
to_sfixed(-300807014.0/4294967296.0,1,-nbitq), 
to_sfixed(-234104440.0/4294967296.0,1,-nbitq), 
to_sfixed(462088418.0/4294967296.0,1,-nbitq), 
to_sfixed(395118486.0/4294967296.0,1,-nbitq), 
to_sfixed(-49918266.0/4294967296.0,1,-nbitq), 
to_sfixed(126833207.0/4294967296.0,1,-nbitq), 
to_sfixed(-748925056.0/4294967296.0,1,-nbitq), 
to_sfixed(-204227620.0/4294967296.0,1,-nbitq), 
to_sfixed(84634691.0/4294967296.0,1,-nbitq), 
to_sfixed(45390216.0/4294967296.0,1,-nbitq), 
to_sfixed(-443364076.0/4294967296.0,1,-nbitq), 
to_sfixed(-296255567.0/4294967296.0,1,-nbitq), 
to_sfixed(127192675.0/4294967296.0,1,-nbitq), 
to_sfixed(199223278.0/4294967296.0,1,-nbitq), 
to_sfixed(-423438350.0/4294967296.0,1,-nbitq), 
to_sfixed(446242746.0/4294967296.0,1,-nbitq), 
to_sfixed(-372143138.0/4294967296.0,1,-nbitq), 
to_sfixed(-179797904.0/4294967296.0,1,-nbitq), 
to_sfixed(390075584.0/4294967296.0,1,-nbitq), 
to_sfixed(310575256.0/4294967296.0,1,-nbitq), 
to_sfixed(-149589679.0/4294967296.0,1,-nbitq), 
to_sfixed(-23306995.0/4294967296.0,1,-nbitq), 
to_sfixed(199325578.0/4294967296.0,1,-nbitq), 
to_sfixed(-171381956.0/4294967296.0,1,-nbitq), 
to_sfixed(123136134.0/4294967296.0,1,-nbitq), 
to_sfixed(293202340.0/4294967296.0,1,-nbitq), 
to_sfixed(-165644846.0/4294967296.0,1,-nbitq), 
to_sfixed(290101506.0/4294967296.0,1,-nbitq), 
to_sfixed(405825655.0/4294967296.0,1,-nbitq), 
to_sfixed(72238752.0/4294967296.0,1,-nbitq), 
to_sfixed(-75264799.0/4294967296.0,1,-nbitq), 
to_sfixed(-44413177.0/4294967296.0,1,-nbitq), 
to_sfixed(238923310.0/4294967296.0,1,-nbitq), 
to_sfixed(-59313985.0/4294967296.0,1,-nbitq), 
to_sfixed(136832626.0/4294967296.0,1,-nbitq), 
to_sfixed(-11166357.0/4294967296.0,1,-nbitq), 
to_sfixed(-456371776.0/4294967296.0,1,-nbitq), 
to_sfixed(13915031.0/4294967296.0,1,-nbitq), 
to_sfixed(77860495.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-38064675.0/4294967296.0,1,-nbitq), 
to_sfixed(244211744.0/4294967296.0,1,-nbitq), 
to_sfixed(-359018283.0/4294967296.0,1,-nbitq), 
to_sfixed(183977240.0/4294967296.0,1,-nbitq), 
to_sfixed(548803759.0/4294967296.0,1,-nbitq), 
to_sfixed(268428638.0/4294967296.0,1,-nbitq), 
to_sfixed(284958357.0/4294967296.0,1,-nbitq), 
to_sfixed(-113761343.0/4294967296.0,1,-nbitq), 
to_sfixed(-49464294.0/4294967296.0,1,-nbitq), 
to_sfixed(-30211480.0/4294967296.0,1,-nbitq), 
to_sfixed(280021417.0/4294967296.0,1,-nbitq), 
to_sfixed(-78145964.0/4294967296.0,1,-nbitq), 
to_sfixed(766674601.0/4294967296.0,1,-nbitq), 
to_sfixed(715253550.0/4294967296.0,1,-nbitq), 
to_sfixed(-13829217.0/4294967296.0,1,-nbitq), 
to_sfixed(-407112349.0/4294967296.0,1,-nbitq), 
to_sfixed(-280692061.0/4294967296.0,1,-nbitq), 
to_sfixed(29459304.0/4294967296.0,1,-nbitq), 
to_sfixed(98894797.0/4294967296.0,1,-nbitq), 
to_sfixed(172198182.0/4294967296.0,1,-nbitq), 
to_sfixed(-150599932.0/4294967296.0,1,-nbitq), 
to_sfixed(191888819.0/4294967296.0,1,-nbitq), 
to_sfixed(-468982531.0/4294967296.0,1,-nbitq), 
to_sfixed(223862181.0/4294967296.0,1,-nbitq), 
to_sfixed(111967647.0/4294967296.0,1,-nbitq), 
to_sfixed(530719881.0/4294967296.0,1,-nbitq), 
to_sfixed(103430251.0/4294967296.0,1,-nbitq), 
to_sfixed(-221055416.0/4294967296.0,1,-nbitq), 
to_sfixed(-211719359.0/4294967296.0,1,-nbitq), 
to_sfixed(206582409.0/4294967296.0,1,-nbitq), 
to_sfixed(240337676.0/4294967296.0,1,-nbitq), 
to_sfixed(-339732977.0/4294967296.0,1,-nbitq), 
to_sfixed(216881998.0/4294967296.0,1,-nbitq), 
to_sfixed(173784625.0/4294967296.0,1,-nbitq), 
to_sfixed(340165543.0/4294967296.0,1,-nbitq), 
to_sfixed(-243175925.0/4294967296.0,1,-nbitq), 
to_sfixed(-352358951.0/4294967296.0,1,-nbitq), 
to_sfixed(311492928.0/4294967296.0,1,-nbitq), 
to_sfixed(-16690961.0/4294967296.0,1,-nbitq), 
to_sfixed(422979338.0/4294967296.0,1,-nbitq), 
to_sfixed(74161810.0/4294967296.0,1,-nbitq), 
to_sfixed(-339704129.0/4294967296.0,1,-nbitq), 
to_sfixed(280469036.0/4294967296.0,1,-nbitq), 
to_sfixed(439183569.0/4294967296.0,1,-nbitq), 
to_sfixed(37894603.0/4294967296.0,1,-nbitq), 
to_sfixed(28410094.0/4294967296.0,1,-nbitq), 
to_sfixed(-2411015.0/4294967296.0,1,-nbitq), 
to_sfixed(-557557659.0/4294967296.0,1,-nbitq), 
to_sfixed(469515864.0/4294967296.0,1,-nbitq), 
to_sfixed(21082719.0/4294967296.0,1,-nbitq), 
to_sfixed(7637512.0/4294967296.0,1,-nbitq), 
to_sfixed(76046122.0/4294967296.0,1,-nbitq), 
to_sfixed(45292242.0/4294967296.0,1,-nbitq), 
to_sfixed(83934404.0/4294967296.0,1,-nbitq), 
to_sfixed(675067491.0/4294967296.0,1,-nbitq), 
to_sfixed(220703662.0/4294967296.0,1,-nbitq), 
to_sfixed(84746248.0/4294967296.0,1,-nbitq), 
to_sfixed(92287172.0/4294967296.0,1,-nbitq), 
to_sfixed(263078271.0/4294967296.0,1,-nbitq), 
to_sfixed(-71962459.0/4294967296.0,1,-nbitq), 
to_sfixed(-292453105.0/4294967296.0,1,-nbitq), 
to_sfixed(49468865.0/4294967296.0,1,-nbitq), 
to_sfixed(89882146.0/4294967296.0,1,-nbitq), 
to_sfixed(197425939.0/4294967296.0,1,-nbitq), 
to_sfixed(-20018409.0/4294967296.0,1,-nbitq), 
to_sfixed(16476950.0/4294967296.0,1,-nbitq), 
to_sfixed(42863237.0/4294967296.0,1,-nbitq), 
to_sfixed(292646753.0/4294967296.0,1,-nbitq), 
to_sfixed(265140458.0/4294967296.0,1,-nbitq), 
to_sfixed(554048228.0/4294967296.0,1,-nbitq), 
to_sfixed(279829481.0/4294967296.0,1,-nbitq), 
to_sfixed(136493880.0/4294967296.0,1,-nbitq), 
to_sfixed(-406282693.0/4294967296.0,1,-nbitq), 
to_sfixed(96428104.0/4294967296.0,1,-nbitq), 
to_sfixed(-105564746.0/4294967296.0,1,-nbitq), 
to_sfixed(-450524084.0/4294967296.0,1,-nbitq), 
to_sfixed(-40918072.0/4294967296.0,1,-nbitq), 
to_sfixed(-96091743.0/4294967296.0,1,-nbitq), 
to_sfixed(92342105.0/4294967296.0,1,-nbitq), 
to_sfixed(321151916.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(349913611.0/4294967296.0,1,-nbitq), 
to_sfixed(547784215.0/4294967296.0,1,-nbitq), 
to_sfixed(265099803.0/4294967296.0,1,-nbitq), 
to_sfixed(172366564.0/4294967296.0,1,-nbitq), 
to_sfixed(405928877.0/4294967296.0,1,-nbitq), 
to_sfixed(-116395987.0/4294967296.0,1,-nbitq), 
to_sfixed(261022777.0/4294967296.0,1,-nbitq), 
to_sfixed(197973867.0/4294967296.0,1,-nbitq), 
to_sfixed(-415895184.0/4294967296.0,1,-nbitq), 
to_sfixed(99910070.0/4294967296.0,1,-nbitq), 
to_sfixed(-61844724.0/4294967296.0,1,-nbitq), 
to_sfixed(-451880634.0/4294967296.0,1,-nbitq), 
to_sfixed(783970569.0/4294967296.0,1,-nbitq), 
to_sfixed(1174460703.0/4294967296.0,1,-nbitq), 
to_sfixed(430052675.0/4294967296.0,1,-nbitq), 
to_sfixed(-854352787.0/4294967296.0,1,-nbitq), 
to_sfixed(-269001423.0/4294967296.0,1,-nbitq), 
to_sfixed(13180958.0/4294967296.0,1,-nbitq), 
to_sfixed(-275444065.0/4294967296.0,1,-nbitq), 
to_sfixed(428226941.0/4294967296.0,1,-nbitq), 
to_sfixed(70766470.0/4294967296.0,1,-nbitq), 
to_sfixed(-502632892.0/4294967296.0,1,-nbitq), 
to_sfixed(80527082.0/4294967296.0,1,-nbitq), 
to_sfixed(276539767.0/4294967296.0,1,-nbitq), 
to_sfixed(232744601.0/4294967296.0,1,-nbitq), 
to_sfixed(571875442.0/4294967296.0,1,-nbitq), 
to_sfixed(156388740.0/4294967296.0,1,-nbitq), 
to_sfixed(245475257.0/4294967296.0,1,-nbitq), 
to_sfixed(554551780.0/4294967296.0,1,-nbitq), 
to_sfixed(-432997776.0/4294967296.0,1,-nbitq), 
to_sfixed(-160026246.0/4294967296.0,1,-nbitq), 
to_sfixed(48330004.0/4294967296.0,1,-nbitq), 
to_sfixed(-463677225.0/4294967296.0,1,-nbitq), 
to_sfixed(-268997406.0/4294967296.0,1,-nbitq), 
to_sfixed(51696132.0/4294967296.0,1,-nbitq), 
to_sfixed(324086110.0/4294967296.0,1,-nbitq), 
to_sfixed(521993437.0/4294967296.0,1,-nbitq), 
to_sfixed(-188998816.0/4294967296.0,1,-nbitq), 
to_sfixed(-337633516.0/4294967296.0,1,-nbitq), 
to_sfixed(391438096.0/4294967296.0,1,-nbitq), 
to_sfixed(339562321.0/4294967296.0,1,-nbitq), 
to_sfixed(-586745374.0/4294967296.0,1,-nbitq), 
to_sfixed(-1992590.0/4294967296.0,1,-nbitq), 
to_sfixed(-636605916.0/4294967296.0,1,-nbitq), 
to_sfixed(830976769.0/4294967296.0,1,-nbitq), 
to_sfixed(347772589.0/4294967296.0,1,-nbitq), 
to_sfixed(-249268867.0/4294967296.0,1,-nbitq), 
to_sfixed(-828659711.0/4294967296.0,1,-nbitq), 
to_sfixed(528975673.0/4294967296.0,1,-nbitq), 
to_sfixed(45893534.0/4294967296.0,1,-nbitq), 
to_sfixed(-400116967.0/4294967296.0,1,-nbitq), 
to_sfixed(368355418.0/4294967296.0,1,-nbitq), 
to_sfixed(326539910.0/4294967296.0,1,-nbitq), 
to_sfixed(-283207718.0/4294967296.0,1,-nbitq), 
to_sfixed(1246547351.0/4294967296.0,1,-nbitq), 
to_sfixed(459611268.0/4294967296.0,1,-nbitq), 
to_sfixed(-247812729.0/4294967296.0,1,-nbitq), 
to_sfixed(-294180818.0/4294967296.0,1,-nbitq), 
to_sfixed(341643524.0/4294967296.0,1,-nbitq), 
to_sfixed(342408617.0/4294967296.0,1,-nbitq), 
to_sfixed(243841902.0/4294967296.0,1,-nbitq), 
to_sfixed(-50902222.0/4294967296.0,1,-nbitq), 
to_sfixed(-762364599.0/4294967296.0,1,-nbitq), 
to_sfixed(-233750197.0/4294967296.0,1,-nbitq), 
to_sfixed(-426603781.0/4294967296.0,1,-nbitq), 
to_sfixed(-32715352.0/4294967296.0,1,-nbitq), 
to_sfixed(8392738.0/4294967296.0,1,-nbitq), 
to_sfixed(349003037.0/4294967296.0,1,-nbitq), 
to_sfixed(255470533.0/4294967296.0,1,-nbitq), 
to_sfixed(167486751.0/4294967296.0,1,-nbitq), 
to_sfixed(158408507.0/4294967296.0,1,-nbitq), 
to_sfixed(295637207.0/4294967296.0,1,-nbitq), 
to_sfixed(-456039877.0/4294967296.0,1,-nbitq), 
to_sfixed(-27386358.0/4294967296.0,1,-nbitq), 
to_sfixed(393290178.0/4294967296.0,1,-nbitq), 
to_sfixed(-87818237.0/4294967296.0,1,-nbitq), 
to_sfixed(457247336.0/4294967296.0,1,-nbitq), 
to_sfixed(75165218.0/4294967296.0,1,-nbitq), 
to_sfixed(-300040373.0/4294967296.0,1,-nbitq), 
to_sfixed(329820093.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(261089165.0/4294967296.0,1,-nbitq), 
to_sfixed(1106531446.0/4294967296.0,1,-nbitq), 
to_sfixed(252744220.0/4294967296.0,1,-nbitq), 
to_sfixed(437861655.0/4294967296.0,1,-nbitq), 
to_sfixed(-249838677.0/4294967296.0,1,-nbitq), 
to_sfixed(35636334.0/4294967296.0,1,-nbitq), 
to_sfixed(419857442.0/4294967296.0,1,-nbitq), 
to_sfixed(-555950444.0/4294967296.0,1,-nbitq), 
to_sfixed(-285926413.0/4294967296.0,1,-nbitq), 
to_sfixed(391445642.0/4294967296.0,1,-nbitq), 
to_sfixed(513187356.0/4294967296.0,1,-nbitq), 
to_sfixed(284074752.0/4294967296.0,1,-nbitq), 
to_sfixed(1160311149.0/4294967296.0,1,-nbitq), 
to_sfixed(1324665685.0/4294967296.0,1,-nbitq), 
to_sfixed(-11427340.0/4294967296.0,1,-nbitq), 
to_sfixed(-741520295.0/4294967296.0,1,-nbitq), 
to_sfixed(336593180.0/4294967296.0,1,-nbitq), 
to_sfixed(297256292.0/4294967296.0,1,-nbitq), 
to_sfixed(-247597275.0/4294967296.0,1,-nbitq), 
to_sfixed(457109481.0/4294967296.0,1,-nbitq), 
to_sfixed(-96748136.0/4294967296.0,1,-nbitq), 
to_sfixed(-5731716.0/4294967296.0,1,-nbitq), 
to_sfixed(558843335.0/4294967296.0,1,-nbitq), 
to_sfixed(771453926.0/4294967296.0,1,-nbitq), 
to_sfixed(58505024.0/4294967296.0,1,-nbitq), 
to_sfixed(1443630871.0/4294967296.0,1,-nbitq), 
to_sfixed(-438930012.0/4294967296.0,1,-nbitq), 
to_sfixed(-359474468.0/4294967296.0,1,-nbitq), 
to_sfixed(783169460.0/4294967296.0,1,-nbitq), 
to_sfixed(-58977632.0/4294967296.0,1,-nbitq), 
to_sfixed(-58767056.0/4294967296.0,1,-nbitq), 
to_sfixed(52555065.0/4294967296.0,1,-nbitq), 
to_sfixed(-505354199.0/4294967296.0,1,-nbitq), 
to_sfixed(-51949627.0/4294967296.0,1,-nbitq), 
to_sfixed(-334971102.0/4294967296.0,1,-nbitq), 
to_sfixed(647983574.0/4294967296.0,1,-nbitq), 
to_sfixed(-222362040.0/4294967296.0,1,-nbitq), 
to_sfixed(-136107606.0/4294967296.0,1,-nbitq), 
to_sfixed(-499949199.0/4294967296.0,1,-nbitq), 
to_sfixed(73338341.0/4294967296.0,1,-nbitq), 
to_sfixed(257592902.0/4294967296.0,1,-nbitq), 
to_sfixed(-41317471.0/4294967296.0,1,-nbitq), 
to_sfixed(394663671.0/4294967296.0,1,-nbitq), 
to_sfixed(-252574658.0/4294967296.0,1,-nbitq), 
to_sfixed(273049179.0/4294967296.0,1,-nbitq), 
to_sfixed(1172995719.0/4294967296.0,1,-nbitq), 
to_sfixed(65723472.0/4294967296.0,1,-nbitq), 
to_sfixed(-785008574.0/4294967296.0,1,-nbitq), 
to_sfixed(392782687.0/4294967296.0,1,-nbitq), 
to_sfixed(-435311942.0/4294967296.0,1,-nbitq), 
to_sfixed(344871071.0/4294967296.0,1,-nbitq), 
to_sfixed(128927178.0/4294967296.0,1,-nbitq), 
to_sfixed(838239655.0/4294967296.0,1,-nbitq), 
to_sfixed(-738017016.0/4294967296.0,1,-nbitq), 
to_sfixed(663730430.0/4294967296.0,1,-nbitq), 
to_sfixed(757029383.0/4294967296.0,1,-nbitq), 
to_sfixed(367160582.0/4294967296.0,1,-nbitq), 
to_sfixed(611444975.0/4294967296.0,1,-nbitq), 
to_sfixed(151550230.0/4294967296.0,1,-nbitq), 
to_sfixed(179495981.0/4294967296.0,1,-nbitq), 
to_sfixed(375123201.0/4294967296.0,1,-nbitq), 
to_sfixed(-94982702.0/4294967296.0,1,-nbitq), 
to_sfixed(-900166053.0/4294967296.0,1,-nbitq), 
to_sfixed(-279807562.0/4294967296.0,1,-nbitq), 
to_sfixed(-684490528.0/4294967296.0,1,-nbitq), 
to_sfixed(-14762950.0/4294967296.0,1,-nbitq), 
to_sfixed(-527200332.0/4294967296.0,1,-nbitq), 
to_sfixed(54177462.0/4294967296.0,1,-nbitq), 
to_sfixed(-350700813.0/4294967296.0,1,-nbitq), 
to_sfixed(-506202047.0/4294967296.0,1,-nbitq), 
to_sfixed(661827354.0/4294967296.0,1,-nbitq), 
to_sfixed(178543243.0/4294967296.0,1,-nbitq), 
to_sfixed(-94475918.0/4294967296.0,1,-nbitq), 
to_sfixed(-253111303.0/4294967296.0,1,-nbitq), 
to_sfixed(226814909.0/4294967296.0,1,-nbitq), 
to_sfixed(179152616.0/4294967296.0,1,-nbitq), 
to_sfixed(635539142.0/4294967296.0,1,-nbitq), 
to_sfixed(-219155331.0/4294967296.0,1,-nbitq), 
to_sfixed(-402670391.0/4294967296.0,1,-nbitq), 
to_sfixed(31449027.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-23663694.0/4294967296.0,1,-nbitq), 
to_sfixed(426435576.0/4294967296.0,1,-nbitq), 
to_sfixed(-721355675.0/4294967296.0,1,-nbitq), 
to_sfixed(-78907898.0/4294967296.0,1,-nbitq), 
to_sfixed(114795144.0/4294967296.0,1,-nbitq), 
to_sfixed(263252537.0/4294967296.0,1,-nbitq), 
to_sfixed(-153361187.0/4294967296.0,1,-nbitq), 
to_sfixed(-275745240.0/4294967296.0,1,-nbitq), 
to_sfixed(843087719.0/4294967296.0,1,-nbitq), 
to_sfixed(47159472.0/4294967296.0,1,-nbitq), 
to_sfixed(-9779432.0/4294967296.0,1,-nbitq), 
to_sfixed(77286536.0/4294967296.0,1,-nbitq), 
to_sfixed(1401064555.0/4294967296.0,1,-nbitq), 
to_sfixed(1080058997.0/4294967296.0,1,-nbitq), 
to_sfixed(-335194518.0/4294967296.0,1,-nbitq), 
to_sfixed(-153935705.0/4294967296.0,1,-nbitq), 
to_sfixed(-6301437.0/4294967296.0,1,-nbitq), 
to_sfixed(-190956106.0/4294967296.0,1,-nbitq), 
to_sfixed(-197461447.0/4294967296.0,1,-nbitq), 
to_sfixed(486517916.0/4294967296.0,1,-nbitq), 
to_sfixed(-52480571.0/4294967296.0,1,-nbitq), 
to_sfixed(-396994890.0/4294967296.0,1,-nbitq), 
to_sfixed(60978596.0/4294967296.0,1,-nbitq), 
to_sfixed(247291089.0/4294967296.0,1,-nbitq), 
to_sfixed(-328853444.0/4294967296.0,1,-nbitq), 
to_sfixed(1144316038.0/4294967296.0,1,-nbitq), 
to_sfixed(143979598.0/4294967296.0,1,-nbitq), 
to_sfixed(390249646.0/4294967296.0,1,-nbitq), 
to_sfixed(99876524.0/4294967296.0,1,-nbitq), 
to_sfixed(-246098911.0/4294967296.0,1,-nbitq), 
to_sfixed(-107708666.0/4294967296.0,1,-nbitq), 
to_sfixed(-398882883.0/4294967296.0,1,-nbitq), 
to_sfixed(-447327101.0/4294967296.0,1,-nbitq), 
to_sfixed(-165192527.0/4294967296.0,1,-nbitq), 
to_sfixed(-424785582.0/4294967296.0,1,-nbitq), 
to_sfixed(586567881.0/4294967296.0,1,-nbitq), 
to_sfixed(-39585881.0/4294967296.0,1,-nbitq), 
to_sfixed(-236377492.0/4294967296.0,1,-nbitq), 
to_sfixed(207247704.0/4294967296.0,1,-nbitq), 
to_sfixed(444368062.0/4294967296.0,1,-nbitq), 
to_sfixed(-629053391.0/4294967296.0,1,-nbitq), 
to_sfixed(-478334222.0/4294967296.0,1,-nbitq), 
to_sfixed(-329629944.0/4294967296.0,1,-nbitq), 
to_sfixed(308953921.0/4294967296.0,1,-nbitq), 
to_sfixed(-295362404.0/4294967296.0,1,-nbitq), 
to_sfixed(1343455255.0/4294967296.0,1,-nbitq), 
to_sfixed(-71680250.0/4294967296.0,1,-nbitq), 
to_sfixed(-1192741814.0/4294967296.0,1,-nbitq), 
to_sfixed(137575890.0/4294967296.0,1,-nbitq), 
to_sfixed(-841291406.0/4294967296.0,1,-nbitq), 
to_sfixed(488160829.0/4294967296.0,1,-nbitq), 
to_sfixed(57718334.0/4294967296.0,1,-nbitq), 
to_sfixed(350797988.0/4294967296.0,1,-nbitq), 
to_sfixed(-141326278.0/4294967296.0,1,-nbitq), 
to_sfixed(745496159.0/4294967296.0,1,-nbitq), 
to_sfixed(405704524.0/4294967296.0,1,-nbitq), 
to_sfixed(421270780.0/4294967296.0,1,-nbitq), 
to_sfixed(376853579.0/4294967296.0,1,-nbitq), 
to_sfixed(320389674.0/4294967296.0,1,-nbitq), 
to_sfixed(5344321.0/4294967296.0,1,-nbitq), 
to_sfixed(-168957152.0/4294967296.0,1,-nbitq), 
to_sfixed(-25503350.0/4294967296.0,1,-nbitq), 
to_sfixed(-1006809007.0/4294967296.0,1,-nbitq), 
to_sfixed(-483348256.0/4294967296.0,1,-nbitq), 
to_sfixed(-563242525.0/4294967296.0,1,-nbitq), 
to_sfixed(-137580603.0/4294967296.0,1,-nbitq), 
to_sfixed(-456384856.0/4294967296.0,1,-nbitq), 
to_sfixed(560003832.0/4294967296.0,1,-nbitq), 
to_sfixed(153521071.0/4294967296.0,1,-nbitq), 
to_sfixed(-1604342136.0/4294967296.0,1,-nbitq), 
to_sfixed(-256677767.0/4294967296.0,1,-nbitq), 
to_sfixed(271630785.0/4294967296.0,1,-nbitq), 
to_sfixed(124295213.0/4294967296.0,1,-nbitq), 
to_sfixed(-69114210.0/4294967296.0,1,-nbitq), 
to_sfixed(57390524.0/4294967296.0,1,-nbitq), 
to_sfixed(-174044502.0/4294967296.0,1,-nbitq), 
to_sfixed(386828777.0/4294967296.0,1,-nbitq), 
to_sfixed(14113010.0/4294967296.0,1,-nbitq), 
to_sfixed(-231144725.0/4294967296.0,1,-nbitq), 
to_sfixed(-285876270.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-68266186.0/4294967296.0,1,-nbitq), 
to_sfixed(217283875.0/4294967296.0,1,-nbitq), 
to_sfixed(-1434602754.0/4294967296.0,1,-nbitq), 
to_sfixed(419491274.0/4294967296.0,1,-nbitq), 
to_sfixed(806411644.0/4294967296.0,1,-nbitq), 
to_sfixed(1182631826.0/4294967296.0,1,-nbitq), 
to_sfixed(260950845.0/4294967296.0,1,-nbitq), 
to_sfixed(419343754.0/4294967296.0,1,-nbitq), 
to_sfixed(10301202.0/4294967296.0,1,-nbitq), 
to_sfixed(-158200059.0/4294967296.0,1,-nbitq), 
to_sfixed(-820857702.0/4294967296.0,1,-nbitq), 
to_sfixed(-320170128.0/4294967296.0,1,-nbitq), 
to_sfixed(1404291913.0/4294967296.0,1,-nbitq), 
to_sfixed(509133088.0/4294967296.0,1,-nbitq), 
to_sfixed(-33319373.0/4294967296.0,1,-nbitq), 
to_sfixed(-567012420.0/4294967296.0,1,-nbitq), 
to_sfixed(211417201.0/4294967296.0,1,-nbitq), 
to_sfixed(11826369.0/4294967296.0,1,-nbitq), 
to_sfixed(607710557.0/4294967296.0,1,-nbitq), 
to_sfixed(233187472.0/4294967296.0,1,-nbitq), 
to_sfixed(210252858.0/4294967296.0,1,-nbitq), 
to_sfixed(-673882638.0/4294967296.0,1,-nbitq), 
to_sfixed(-70214869.0/4294967296.0,1,-nbitq), 
to_sfixed(652439712.0/4294967296.0,1,-nbitq), 
to_sfixed(8287633.0/4294967296.0,1,-nbitq), 
to_sfixed(1954279655.0/4294967296.0,1,-nbitq), 
to_sfixed(302946963.0/4294967296.0,1,-nbitq), 
to_sfixed(298082431.0/4294967296.0,1,-nbitq), 
to_sfixed(1023220795.0/4294967296.0,1,-nbitq), 
to_sfixed(-29141373.0/4294967296.0,1,-nbitq), 
to_sfixed(42538673.0/4294967296.0,1,-nbitq), 
to_sfixed(-479886384.0/4294967296.0,1,-nbitq), 
to_sfixed(-237819302.0/4294967296.0,1,-nbitq), 
to_sfixed(559772777.0/4294967296.0,1,-nbitq), 
to_sfixed(-437853714.0/4294967296.0,1,-nbitq), 
to_sfixed(330938843.0/4294967296.0,1,-nbitq), 
to_sfixed(268934644.0/4294967296.0,1,-nbitq), 
to_sfixed(88559287.0/4294967296.0,1,-nbitq), 
to_sfixed(-364144878.0/4294967296.0,1,-nbitq), 
to_sfixed(32538329.0/4294967296.0,1,-nbitq), 
to_sfixed(-446909227.0/4294967296.0,1,-nbitq), 
to_sfixed(-615295902.0/4294967296.0,1,-nbitq), 
to_sfixed(-131792429.0/4294967296.0,1,-nbitq), 
to_sfixed(393368771.0/4294967296.0,1,-nbitq), 
to_sfixed(-119344191.0/4294967296.0,1,-nbitq), 
to_sfixed(695086677.0/4294967296.0,1,-nbitq), 
to_sfixed(149992355.0/4294967296.0,1,-nbitq), 
to_sfixed(-1027072234.0/4294967296.0,1,-nbitq), 
to_sfixed(-119765910.0/4294967296.0,1,-nbitq), 
to_sfixed(-1137689604.0/4294967296.0,1,-nbitq), 
to_sfixed(547205657.0/4294967296.0,1,-nbitq), 
to_sfixed(-135143616.0/4294967296.0,1,-nbitq), 
to_sfixed(145566938.0/4294967296.0,1,-nbitq), 
to_sfixed(-251680524.0/4294967296.0,1,-nbitq), 
to_sfixed(-36972018.0/4294967296.0,1,-nbitq), 
to_sfixed(312987954.0/4294967296.0,1,-nbitq), 
to_sfixed(7179018.0/4294967296.0,1,-nbitq), 
to_sfixed(193423894.0/4294967296.0,1,-nbitq), 
to_sfixed(135151855.0/4294967296.0,1,-nbitq), 
to_sfixed(-117149578.0/4294967296.0,1,-nbitq), 
to_sfixed(-65654049.0/4294967296.0,1,-nbitq), 
to_sfixed(283152480.0/4294967296.0,1,-nbitq), 
to_sfixed(-767994310.0/4294967296.0,1,-nbitq), 
to_sfixed(340328367.0/4294967296.0,1,-nbitq), 
to_sfixed(51840743.0/4294967296.0,1,-nbitq), 
to_sfixed(-397317153.0/4294967296.0,1,-nbitq), 
to_sfixed(-756685615.0/4294967296.0,1,-nbitq), 
to_sfixed(190560976.0/4294967296.0,1,-nbitq), 
to_sfixed(-64032971.0/4294967296.0,1,-nbitq), 
to_sfixed(-1915729130.0/4294967296.0,1,-nbitq), 
to_sfixed(226427649.0/4294967296.0,1,-nbitq), 
to_sfixed(-79744374.0/4294967296.0,1,-nbitq), 
to_sfixed(-16375128.0/4294967296.0,1,-nbitq), 
to_sfixed(8930073.0/4294967296.0,1,-nbitq), 
to_sfixed(137055793.0/4294967296.0,1,-nbitq), 
to_sfixed(-343821300.0/4294967296.0,1,-nbitq), 
to_sfixed(920496193.0/4294967296.0,1,-nbitq), 
to_sfixed(56790644.0/4294967296.0,1,-nbitq), 
to_sfixed(-196934191.0/4294967296.0,1,-nbitq), 
to_sfixed(-320829591.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(159562866.0/4294967296.0,1,-nbitq), 
to_sfixed(54182391.0/4294967296.0,1,-nbitq), 
to_sfixed(-834570247.0/4294967296.0,1,-nbitq), 
to_sfixed(920184417.0/4294967296.0,1,-nbitq), 
to_sfixed(712237853.0/4294967296.0,1,-nbitq), 
to_sfixed(1997018117.0/4294967296.0,1,-nbitq), 
to_sfixed(-71919666.0/4294967296.0,1,-nbitq), 
to_sfixed(963659598.0/4294967296.0,1,-nbitq), 
to_sfixed(-364033722.0/4294967296.0,1,-nbitq), 
to_sfixed(-283347157.0/4294967296.0,1,-nbitq), 
to_sfixed(-1519820059.0/4294967296.0,1,-nbitq), 
to_sfixed(-138888334.0/4294967296.0,1,-nbitq), 
to_sfixed(1697230267.0/4294967296.0,1,-nbitq), 
to_sfixed(729028784.0/4294967296.0,1,-nbitq), 
to_sfixed(243233558.0/4294967296.0,1,-nbitq), 
to_sfixed(-1533212706.0/4294967296.0,1,-nbitq), 
to_sfixed(-4961400.0/4294967296.0,1,-nbitq), 
to_sfixed(125795892.0/4294967296.0,1,-nbitq), 
to_sfixed(-378708427.0/4294967296.0,1,-nbitq), 
to_sfixed(579542616.0/4294967296.0,1,-nbitq), 
to_sfixed(297074706.0/4294967296.0,1,-nbitq), 
to_sfixed(-714215394.0/4294967296.0,1,-nbitq), 
to_sfixed(-144534559.0/4294967296.0,1,-nbitq), 
to_sfixed(1364686633.0/4294967296.0,1,-nbitq), 
to_sfixed(-275055830.0/4294967296.0,1,-nbitq), 
to_sfixed(1676020548.0/4294967296.0,1,-nbitq), 
to_sfixed(-137179515.0/4294967296.0,1,-nbitq), 
to_sfixed(344900.0/4294967296.0,1,-nbitq), 
to_sfixed(42190805.0/4294967296.0,1,-nbitq), 
to_sfixed(236512232.0/4294967296.0,1,-nbitq), 
to_sfixed(271802211.0/4294967296.0,1,-nbitq), 
to_sfixed(-481651547.0/4294967296.0,1,-nbitq), 
to_sfixed(-291478530.0/4294967296.0,1,-nbitq), 
to_sfixed(-41077148.0/4294967296.0,1,-nbitq), 
to_sfixed(97013070.0/4294967296.0,1,-nbitq), 
to_sfixed(70303321.0/4294967296.0,1,-nbitq), 
to_sfixed(510640485.0/4294967296.0,1,-nbitq), 
to_sfixed(-1242746373.0/4294967296.0,1,-nbitq), 
to_sfixed(-606031797.0/4294967296.0,1,-nbitq), 
to_sfixed(-281604272.0/4294967296.0,1,-nbitq), 
to_sfixed(-189798908.0/4294967296.0,1,-nbitq), 
to_sfixed(-935505604.0/4294967296.0,1,-nbitq), 
to_sfixed(37061650.0/4294967296.0,1,-nbitq), 
to_sfixed(100513268.0/4294967296.0,1,-nbitq), 
to_sfixed(-90862289.0/4294967296.0,1,-nbitq), 
to_sfixed(432561049.0/4294967296.0,1,-nbitq), 
to_sfixed(-114846369.0/4294967296.0,1,-nbitq), 
to_sfixed(-948503700.0/4294967296.0,1,-nbitq), 
to_sfixed(-106472071.0/4294967296.0,1,-nbitq), 
to_sfixed(-1239073434.0/4294967296.0,1,-nbitq), 
to_sfixed(452120442.0/4294967296.0,1,-nbitq), 
to_sfixed(2336559.0/4294967296.0,1,-nbitq), 
to_sfixed(-589052821.0/4294967296.0,1,-nbitq), 
to_sfixed(347841350.0/4294967296.0,1,-nbitq), 
to_sfixed(-166279568.0/4294967296.0,1,-nbitq), 
to_sfixed(396311641.0/4294967296.0,1,-nbitq), 
to_sfixed(572689135.0/4294967296.0,1,-nbitq), 
to_sfixed(-517840091.0/4294967296.0,1,-nbitq), 
to_sfixed(27618320.0/4294967296.0,1,-nbitq), 
to_sfixed(-214425650.0/4294967296.0,1,-nbitq), 
to_sfixed(76430223.0/4294967296.0,1,-nbitq), 
to_sfixed(-240754712.0/4294967296.0,1,-nbitq), 
to_sfixed(-718131021.0/4294967296.0,1,-nbitq), 
to_sfixed(493692565.0/4294967296.0,1,-nbitq), 
to_sfixed(77078577.0/4294967296.0,1,-nbitq), 
to_sfixed(-400899483.0/4294967296.0,1,-nbitq), 
to_sfixed(-316148157.0/4294967296.0,1,-nbitq), 
to_sfixed(86269041.0/4294967296.0,1,-nbitq), 
to_sfixed(224854744.0/4294967296.0,1,-nbitq), 
to_sfixed(-1952065866.0/4294967296.0,1,-nbitq), 
to_sfixed(175885357.0/4294967296.0,1,-nbitq), 
to_sfixed(207872606.0/4294967296.0,1,-nbitq), 
to_sfixed(241521992.0/4294967296.0,1,-nbitq), 
to_sfixed(396867113.0/4294967296.0,1,-nbitq), 
to_sfixed(424685614.0/4294967296.0,1,-nbitq), 
to_sfixed(307983494.0/4294967296.0,1,-nbitq), 
to_sfixed(1311827366.0/4294967296.0,1,-nbitq), 
to_sfixed(436401424.0/4294967296.0,1,-nbitq), 
to_sfixed(36611932.0/4294967296.0,1,-nbitq), 
to_sfixed(207590784.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-208324544.0/4294967296.0,1,-nbitq), 
to_sfixed(-379332575.0/4294967296.0,1,-nbitq), 
to_sfixed(-582619054.0/4294967296.0,1,-nbitq), 
to_sfixed(938282396.0/4294967296.0,1,-nbitq), 
to_sfixed(211237786.0/4294967296.0,1,-nbitq), 
to_sfixed(600812826.0/4294967296.0,1,-nbitq), 
to_sfixed(-221767179.0/4294967296.0,1,-nbitq), 
to_sfixed(659683430.0/4294967296.0,1,-nbitq), 
to_sfixed(-120153385.0/4294967296.0,1,-nbitq), 
to_sfixed(225333774.0/4294967296.0,1,-nbitq), 
to_sfixed(-1816778737.0/4294967296.0,1,-nbitq), 
to_sfixed(-107198686.0/4294967296.0,1,-nbitq), 
to_sfixed(1758732083.0/4294967296.0,1,-nbitq), 
to_sfixed(-509410309.0/4294967296.0,1,-nbitq), 
to_sfixed(420097946.0/4294967296.0,1,-nbitq), 
to_sfixed(-1345461395.0/4294967296.0,1,-nbitq), 
to_sfixed(-337632160.0/4294967296.0,1,-nbitq), 
to_sfixed(115923771.0/4294967296.0,1,-nbitq), 
to_sfixed(-568982140.0/4294967296.0,1,-nbitq), 
to_sfixed(183668487.0/4294967296.0,1,-nbitq), 
to_sfixed(111527314.0/4294967296.0,1,-nbitq), 
to_sfixed(-560377199.0/4294967296.0,1,-nbitq), 
to_sfixed(396277843.0/4294967296.0,1,-nbitq), 
to_sfixed(1970930207.0/4294967296.0,1,-nbitq), 
to_sfixed(29126625.0/4294967296.0,1,-nbitq), 
to_sfixed(1075080246.0/4294967296.0,1,-nbitq), 
to_sfixed(530260793.0/4294967296.0,1,-nbitq), 
to_sfixed(332985969.0/4294967296.0,1,-nbitq), 
to_sfixed(372240703.0/4294967296.0,1,-nbitq), 
to_sfixed(-573112935.0/4294967296.0,1,-nbitq), 
to_sfixed(-54960900.0/4294967296.0,1,-nbitq), 
to_sfixed(-563039634.0/4294967296.0,1,-nbitq), 
to_sfixed(224983305.0/4294967296.0,1,-nbitq), 
to_sfixed(265438417.0/4294967296.0,1,-nbitq), 
to_sfixed(-46837140.0/4294967296.0,1,-nbitq), 
to_sfixed(-253959077.0/4294967296.0,1,-nbitq), 
to_sfixed(1347535664.0/4294967296.0,1,-nbitq), 
to_sfixed(-1295417145.0/4294967296.0,1,-nbitq), 
to_sfixed(-24502922.0/4294967296.0,1,-nbitq), 
to_sfixed(-297088260.0/4294967296.0,1,-nbitq), 
to_sfixed(-56745065.0/4294967296.0,1,-nbitq), 
to_sfixed(-510246648.0/4294967296.0,1,-nbitq), 
to_sfixed(362837070.0/4294967296.0,1,-nbitq), 
to_sfixed(37989630.0/4294967296.0,1,-nbitq), 
to_sfixed(-166846111.0/4294967296.0,1,-nbitq), 
to_sfixed(512260454.0/4294967296.0,1,-nbitq), 
to_sfixed(-208341899.0/4294967296.0,1,-nbitq), 
to_sfixed(-913321164.0/4294967296.0,1,-nbitq), 
to_sfixed(-37285292.0/4294967296.0,1,-nbitq), 
to_sfixed(-1304739740.0/4294967296.0,1,-nbitq), 
to_sfixed(-321397950.0/4294967296.0,1,-nbitq), 
to_sfixed(327327202.0/4294967296.0,1,-nbitq), 
to_sfixed(-452983371.0/4294967296.0,1,-nbitq), 
to_sfixed(449457193.0/4294967296.0,1,-nbitq), 
to_sfixed(469461383.0/4294967296.0,1,-nbitq), 
to_sfixed(513570979.0/4294967296.0,1,-nbitq), 
to_sfixed(221109149.0/4294967296.0,1,-nbitq), 
to_sfixed(341353059.0/4294967296.0,1,-nbitq), 
to_sfixed(-25206977.0/4294967296.0,1,-nbitq), 
to_sfixed(-169007478.0/4294967296.0,1,-nbitq), 
to_sfixed(383453562.0/4294967296.0,1,-nbitq), 
to_sfixed(105195733.0/4294967296.0,1,-nbitq), 
to_sfixed(-696220080.0/4294967296.0,1,-nbitq), 
to_sfixed(915128822.0/4294967296.0,1,-nbitq), 
to_sfixed(-18149286.0/4294967296.0,1,-nbitq), 
to_sfixed(45932220.0/4294967296.0,1,-nbitq), 
to_sfixed(-600752616.0/4294967296.0,1,-nbitq), 
to_sfixed(849271288.0/4294967296.0,1,-nbitq), 
to_sfixed(-327286319.0/4294967296.0,1,-nbitq), 
to_sfixed(-839482474.0/4294967296.0,1,-nbitq), 
to_sfixed(-186501755.0/4294967296.0,1,-nbitq), 
to_sfixed(-534692416.0/4294967296.0,1,-nbitq), 
to_sfixed(963865541.0/4294967296.0,1,-nbitq), 
to_sfixed(878664.0/4294967296.0,1,-nbitq), 
to_sfixed(112139127.0/4294967296.0,1,-nbitq), 
to_sfixed(374570969.0/4294967296.0,1,-nbitq), 
to_sfixed(1541649809.0/4294967296.0,1,-nbitq), 
to_sfixed(230662561.0/4294967296.0,1,-nbitq), 
to_sfixed(926513992.0/4294967296.0,1,-nbitq), 
to_sfixed(185363323.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(270331433.0/4294967296.0,1,-nbitq), 
to_sfixed(-197678424.0/4294967296.0,1,-nbitq), 
to_sfixed(-69766761.0/4294967296.0,1,-nbitq), 
to_sfixed(351639074.0/4294967296.0,1,-nbitq), 
to_sfixed(-26998972.0/4294967296.0,1,-nbitq), 
to_sfixed(-881692021.0/4294967296.0,1,-nbitq), 
to_sfixed(377544885.0/4294967296.0,1,-nbitq), 
to_sfixed(-1461602648.0/4294967296.0,1,-nbitq), 
to_sfixed(719321644.0/4294967296.0,1,-nbitq), 
to_sfixed(-64957812.0/4294967296.0,1,-nbitq), 
to_sfixed(-1559498838.0/4294967296.0,1,-nbitq), 
to_sfixed(-604872521.0/4294967296.0,1,-nbitq), 
to_sfixed(1312729027.0/4294967296.0,1,-nbitq), 
to_sfixed(-981967773.0/4294967296.0,1,-nbitq), 
to_sfixed(327209706.0/4294967296.0,1,-nbitq), 
to_sfixed(-825621379.0/4294967296.0,1,-nbitq), 
to_sfixed(229817813.0/4294967296.0,1,-nbitq), 
to_sfixed(353019142.0/4294967296.0,1,-nbitq), 
to_sfixed(362421690.0/4294967296.0,1,-nbitq), 
to_sfixed(-817788556.0/4294967296.0,1,-nbitq), 
to_sfixed(41959842.0/4294967296.0,1,-nbitq), 
to_sfixed(-56369676.0/4294967296.0,1,-nbitq), 
to_sfixed(-135223745.0/4294967296.0,1,-nbitq), 
to_sfixed(1691192082.0/4294967296.0,1,-nbitq), 
to_sfixed(-247213408.0/4294967296.0,1,-nbitq), 
to_sfixed(295411478.0/4294967296.0,1,-nbitq), 
to_sfixed(146079603.0/4294967296.0,1,-nbitq), 
to_sfixed(951022821.0/4294967296.0,1,-nbitq), 
to_sfixed(1372298867.0/4294967296.0,1,-nbitq), 
to_sfixed(-613689993.0/4294967296.0,1,-nbitq), 
to_sfixed(361824708.0/4294967296.0,1,-nbitq), 
to_sfixed(-782081053.0/4294967296.0,1,-nbitq), 
to_sfixed(-85871540.0/4294967296.0,1,-nbitq), 
to_sfixed(646404062.0/4294967296.0,1,-nbitq), 
to_sfixed(-21577900.0/4294967296.0,1,-nbitq), 
to_sfixed(-784864463.0/4294967296.0,1,-nbitq), 
to_sfixed(651235076.0/4294967296.0,1,-nbitq), 
to_sfixed(-385390856.0/4294967296.0,1,-nbitq), 
to_sfixed(132123481.0/4294967296.0,1,-nbitq), 
to_sfixed(-220482037.0/4294967296.0,1,-nbitq), 
to_sfixed(658445440.0/4294967296.0,1,-nbitq), 
to_sfixed(-549019035.0/4294967296.0,1,-nbitq), 
to_sfixed(-5495734.0/4294967296.0,1,-nbitq), 
to_sfixed(-485909833.0/4294967296.0,1,-nbitq), 
to_sfixed(-161317864.0/4294967296.0,1,-nbitq), 
to_sfixed(-174983614.0/4294967296.0,1,-nbitq), 
to_sfixed(-422116248.0/4294967296.0,1,-nbitq), 
to_sfixed(-1208654836.0/4294967296.0,1,-nbitq), 
to_sfixed(-166958290.0/4294967296.0,1,-nbitq), 
to_sfixed(-1176808852.0/4294967296.0,1,-nbitq), 
to_sfixed(-249438944.0/4294967296.0,1,-nbitq), 
to_sfixed(368346364.0/4294967296.0,1,-nbitq), 
to_sfixed(19707951.0/4294967296.0,1,-nbitq), 
to_sfixed(793101562.0/4294967296.0,1,-nbitq), 
to_sfixed(156896353.0/4294967296.0,1,-nbitq), 
to_sfixed(906117992.0/4294967296.0,1,-nbitq), 
to_sfixed(324866000.0/4294967296.0,1,-nbitq), 
to_sfixed(1215770273.0/4294967296.0,1,-nbitq), 
to_sfixed(-80391366.0/4294967296.0,1,-nbitq), 
to_sfixed(-276496585.0/4294967296.0,1,-nbitq), 
to_sfixed(556872060.0/4294967296.0,1,-nbitq), 
to_sfixed(435378823.0/4294967296.0,1,-nbitq), 
to_sfixed(536931597.0/4294967296.0,1,-nbitq), 
to_sfixed(910563418.0/4294967296.0,1,-nbitq), 
to_sfixed(190826358.0/4294967296.0,1,-nbitq), 
to_sfixed(210776754.0/4294967296.0,1,-nbitq), 
to_sfixed(-624391014.0/4294967296.0,1,-nbitq), 
to_sfixed(654071090.0/4294967296.0,1,-nbitq), 
to_sfixed(-231074517.0/4294967296.0,1,-nbitq), 
to_sfixed(-738942320.0/4294967296.0,1,-nbitq), 
to_sfixed(-3411121.0/4294967296.0,1,-nbitq), 
to_sfixed(-12296554.0/4294967296.0,1,-nbitq), 
to_sfixed(639614207.0/4294967296.0,1,-nbitq), 
to_sfixed(-107959401.0/4294967296.0,1,-nbitq), 
to_sfixed(36443196.0/4294967296.0,1,-nbitq), 
to_sfixed(503941132.0/4294967296.0,1,-nbitq), 
to_sfixed(1086908362.0/4294967296.0,1,-nbitq), 
to_sfixed(139056817.0/4294967296.0,1,-nbitq), 
to_sfixed(1570603153.0/4294967296.0,1,-nbitq), 
to_sfixed(-229452232.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(81097897.0/4294967296.0,1,-nbitq), 
to_sfixed(-652619097.0/4294967296.0,1,-nbitq), 
to_sfixed(-130355288.0/4294967296.0,1,-nbitq), 
to_sfixed(716361865.0/4294967296.0,1,-nbitq), 
to_sfixed(725423759.0/4294967296.0,1,-nbitq), 
to_sfixed(-836391034.0/4294967296.0,1,-nbitq), 
to_sfixed(123408690.0/4294967296.0,1,-nbitq), 
to_sfixed(-2086487820.0/4294967296.0,1,-nbitq), 
to_sfixed(885428393.0/4294967296.0,1,-nbitq), 
to_sfixed(-345550110.0/4294967296.0,1,-nbitq), 
to_sfixed(-1033646056.0/4294967296.0,1,-nbitq), 
to_sfixed(-13763122.0/4294967296.0,1,-nbitq), 
to_sfixed(1967872995.0/4294967296.0,1,-nbitq), 
to_sfixed(-1510647791.0/4294967296.0,1,-nbitq), 
to_sfixed(202300374.0/4294967296.0,1,-nbitq), 
to_sfixed(-1464250985.0/4294967296.0,1,-nbitq), 
to_sfixed(64134681.0/4294967296.0,1,-nbitq), 
to_sfixed(86877420.0/4294967296.0,1,-nbitq), 
to_sfixed(820044234.0/4294967296.0,1,-nbitq), 
to_sfixed(-857412642.0/4294967296.0,1,-nbitq), 
to_sfixed(110173968.0/4294967296.0,1,-nbitq), 
to_sfixed(381198892.0/4294967296.0,1,-nbitq), 
to_sfixed(-423883619.0/4294967296.0,1,-nbitq), 
to_sfixed(807087585.0/4294967296.0,1,-nbitq), 
to_sfixed(-44457065.0/4294967296.0,1,-nbitq), 
to_sfixed(555050059.0/4294967296.0,1,-nbitq), 
to_sfixed(-803916626.0/4294967296.0,1,-nbitq), 
to_sfixed(1292239482.0/4294967296.0,1,-nbitq), 
to_sfixed(-74304509.0/4294967296.0,1,-nbitq), 
to_sfixed(-514488353.0/4294967296.0,1,-nbitq), 
to_sfixed(906168932.0/4294967296.0,1,-nbitq), 
to_sfixed(-274424823.0/4294967296.0,1,-nbitq), 
to_sfixed(163127199.0/4294967296.0,1,-nbitq), 
to_sfixed(245460318.0/4294967296.0,1,-nbitq), 
to_sfixed(-195881290.0/4294967296.0,1,-nbitq), 
to_sfixed(-75253213.0/4294967296.0,1,-nbitq), 
to_sfixed(739566198.0/4294967296.0,1,-nbitq), 
to_sfixed(627773468.0/4294967296.0,1,-nbitq), 
to_sfixed(-16903401.0/4294967296.0,1,-nbitq), 
to_sfixed(157513083.0/4294967296.0,1,-nbitq), 
to_sfixed(920471092.0/4294967296.0,1,-nbitq), 
to_sfixed(-342095432.0/4294967296.0,1,-nbitq), 
to_sfixed(670116236.0/4294967296.0,1,-nbitq), 
to_sfixed(-279281869.0/4294967296.0,1,-nbitq), 
to_sfixed(-815272620.0/4294967296.0,1,-nbitq), 
to_sfixed(-212770377.0/4294967296.0,1,-nbitq), 
to_sfixed(-348781653.0/4294967296.0,1,-nbitq), 
to_sfixed(-1248157366.0/4294967296.0,1,-nbitq), 
to_sfixed(-540956400.0/4294967296.0,1,-nbitq), 
to_sfixed(-1491585009.0/4294967296.0,1,-nbitq), 
to_sfixed(-48131254.0/4294967296.0,1,-nbitq), 
to_sfixed(285842119.0/4294967296.0,1,-nbitq), 
to_sfixed(-429657132.0/4294967296.0,1,-nbitq), 
to_sfixed(43796278.0/4294967296.0,1,-nbitq), 
to_sfixed(141058420.0/4294967296.0,1,-nbitq), 
to_sfixed(632279923.0/4294967296.0,1,-nbitq), 
to_sfixed(594700458.0/4294967296.0,1,-nbitq), 
to_sfixed(949520026.0/4294967296.0,1,-nbitq), 
to_sfixed(-204732848.0/4294967296.0,1,-nbitq), 
to_sfixed(-231126872.0/4294967296.0,1,-nbitq), 
to_sfixed(-40027539.0/4294967296.0,1,-nbitq), 
to_sfixed(-157440402.0/4294967296.0,1,-nbitq), 
to_sfixed(690317591.0/4294967296.0,1,-nbitq), 
to_sfixed(718126378.0/4294967296.0,1,-nbitq), 
to_sfixed(-299604376.0/4294967296.0,1,-nbitq), 
to_sfixed(-99808469.0/4294967296.0,1,-nbitq), 
to_sfixed(-374954632.0/4294967296.0,1,-nbitq), 
to_sfixed(-80482952.0/4294967296.0,1,-nbitq), 
to_sfixed(171267153.0/4294967296.0,1,-nbitq), 
to_sfixed(-711735503.0/4294967296.0,1,-nbitq), 
to_sfixed(364709246.0/4294967296.0,1,-nbitq), 
to_sfixed(-15132044.0/4294967296.0,1,-nbitq), 
to_sfixed(260715686.0/4294967296.0,1,-nbitq), 
to_sfixed(329286330.0/4294967296.0,1,-nbitq), 
to_sfixed(337919099.0/4294967296.0,1,-nbitq), 
to_sfixed(1461315050.0/4294967296.0,1,-nbitq), 
to_sfixed(893584323.0/4294967296.0,1,-nbitq), 
to_sfixed(668196535.0/4294967296.0,1,-nbitq), 
to_sfixed(1806324814.0/4294967296.0,1,-nbitq), 
to_sfixed(142693441.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-406405702.0/4294967296.0,1,-nbitq), 
to_sfixed(-1142049303.0/4294967296.0,1,-nbitq), 
to_sfixed(464836968.0/4294967296.0,1,-nbitq), 
to_sfixed(628843241.0/4294967296.0,1,-nbitq), 
to_sfixed(534894830.0/4294967296.0,1,-nbitq), 
to_sfixed(-68073443.0/4294967296.0,1,-nbitq), 
to_sfixed(-235750379.0/4294967296.0,1,-nbitq), 
to_sfixed(-313740993.0/4294967296.0,1,-nbitq), 
to_sfixed(1028622737.0/4294967296.0,1,-nbitq), 
to_sfixed(93040421.0/4294967296.0,1,-nbitq), 
to_sfixed(348613610.0/4294967296.0,1,-nbitq), 
to_sfixed(-480821312.0/4294967296.0,1,-nbitq), 
to_sfixed(1228704929.0/4294967296.0,1,-nbitq), 
to_sfixed(-785886664.0/4294967296.0,1,-nbitq), 
to_sfixed(329500999.0/4294967296.0,1,-nbitq), 
to_sfixed(-1899952512.0/4294967296.0,1,-nbitq), 
to_sfixed(-150459022.0/4294967296.0,1,-nbitq), 
to_sfixed(220179525.0/4294967296.0,1,-nbitq), 
to_sfixed(1084577037.0/4294967296.0,1,-nbitq), 
to_sfixed(254458687.0/4294967296.0,1,-nbitq), 
to_sfixed(115727065.0/4294967296.0,1,-nbitq), 
to_sfixed(320558326.0/4294967296.0,1,-nbitq), 
to_sfixed(-554883446.0/4294967296.0,1,-nbitq), 
to_sfixed(-502376407.0/4294967296.0,1,-nbitq), 
to_sfixed(441329275.0/4294967296.0,1,-nbitq), 
to_sfixed(813037496.0/4294967296.0,1,-nbitq), 
to_sfixed(-96279543.0/4294967296.0,1,-nbitq), 
to_sfixed(731685040.0/4294967296.0,1,-nbitq), 
to_sfixed(-1613022372.0/4294967296.0,1,-nbitq), 
to_sfixed(-331387392.0/4294967296.0,1,-nbitq), 
to_sfixed(1184010674.0/4294967296.0,1,-nbitq), 
to_sfixed(1069770464.0/4294967296.0,1,-nbitq), 
to_sfixed(-626571322.0/4294967296.0,1,-nbitq), 
to_sfixed(374907819.0/4294967296.0,1,-nbitq), 
to_sfixed(630620569.0/4294967296.0,1,-nbitq), 
to_sfixed(885369440.0/4294967296.0,1,-nbitq), 
to_sfixed(428115479.0/4294967296.0,1,-nbitq), 
to_sfixed(1114285070.0/4294967296.0,1,-nbitq), 
to_sfixed(392845445.0/4294967296.0,1,-nbitq), 
to_sfixed(-123597819.0/4294967296.0,1,-nbitq), 
to_sfixed(1731381059.0/4294967296.0,1,-nbitq), 
to_sfixed(-207439104.0/4294967296.0,1,-nbitq), 
to_sfixed(933550114.0/4294967296.0,1,-nbitq), 
to_sfixed(-1105900614.0/4294967296.0,1,-nbitq), 
to_sfixed(-948632270.0/4294967296.0,1,-nbitq), 
to_sfixed(-641563980.0/4294967296.0,1,-nbitq), 
to_sfixed(-193187991.0/4294967296.0,1,-nbitq), 
to_sfixed(-1161132976.0/4294967296.0,1,-nbitq), 
to_sfixed(-606551188.0/4294967296.0,1,-nbitq), 
to_sfixed(-1483967845.0/4294967296.0,1,-nbitq), 
to_sfixed(-433205037.0/4294967296.0,1,-nbitq), 
to_sfixed(124110744.0/4294967296.0,1,-nbitq), 
to_sfixed(-533855196.0/4294967296.0,1,-nbitq), 
to_sfixed(-592771874.0/4294967296.0,1,-nbitq), 
to_sfixed(-388451270.0/4294967296.0,1,-nbitq), 
to_sfixed(818595719.0/4294967296.0,1,-nbitq), 
to_sfixed(457354589.0/4294967296.0,1,-nbitq), 
to_sfixed(-235186934.0/4294967296.0,1,-nbitq), 
to_sfixed(102956820.0/4294967296.0,1,-nbitq), 
to_sfixed(256736387.0/4294967296.0,1,-nbitq), 
to_sfixed(-157377620.0/4294967296.0,1,-nbitq), 
to_sfixed(305746534.0/4294967296.0,1,-nbitq), 
to_sfixed(96076285.0/4294967296.0,1,-nbitq), 
to_sfixed(319823092.0/4294967296.0,1,-nbitq), 
to_sfixed(-78047694.0/4294967296.0,1,-nbitq), 
to_sfixed(394318287.0/4294967296.0,1,-nbitq), 
to_sfixed(417220192.0/4294967296.0,1,-nbitq), 
to_sfixed(-1431357024.0/4294967296.0,1,-nbitq), 
to_sfixed(-5709043.0/4294967296.0,1,-nbitq), 
to_sfixed(-910595206.0/4294967296.0,1,-nbitq), 
to_sfixed(-618651694.0/4294967296.0,1,-nbitq), 
to_sfixed(-380737492.0/4294967296.0,1,-nbitq), 
to_sfixed(466329539.0/4294967296.0,1,-nbitq), 
to_sfixed(336614152.0/4294967296.0,1,-nbitq), 
to_sfixed(368336789.0/4294967296.0,1,-nbitq), 
to_sfixed(941509003.0/4294967296.0,1,-nbitq), 
to_sfixed(778685523.0/4294967296.0,1,-nbitq), 
to_sfixed(-196310760.0/4294967296.0,1,-nbitq), 
to_sfixed(904065815.0/4294967296.0,1,-nbitq), 
to_sfixed(324895564.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(155806803.0/4294967296.0,1,-nbitq), 
to_sfixed(-702805631.0/4294967296.0,1,-nbitq), 
to_sfixed(1581243002.0/4294967296.0,1,-nbitq), 
to_sfixed(165905042.0/4294967296.0,1,-nbitq), 
to_sfixed(78188166.0/4294967296.0,1,-nbitq), 
to_sfixed(-343633241.0/4294967296.0,1,-nbitq), 
to_sfixed(24608192.0/4294967296.0,1,-nbitq), 
to_sfixed(79984964.0/4294967296.0,1,-nbitq), 
to_sfixed(944000454.0/4294967296.0,1,-nbitq), 
to_sfixed(157118474.0/4294967296.0,1,-nbitq), 
to_sfixed(153640124.0/4294967296.0,1,-nbitq), 
to_sfixed(-329903375.0/4294967296.0,1,-nbitq), 
to_sfixed(882871136.0/4294967296.0,1,-nbitq), 
to_sfixed(529298838.0/4294967296.0,1,-nbitq), 
to_sfixed(-147365534.0/4294967296.0,1,-nbitq), 
to_sfixed(-1416770144.0/4294967296.0,1,-nbitq), 
to_sfixed(-290761706.0/4294967296.0,1,-nbitq), 
to_sfixed(-6235167.0/4294967296.0,1,-nbitq), 
to_sfixed(462348015.0/4294967296.0,1,-nbitq), 
to_sfixed(395852296.0/4294967296.0,1,-nbitq), 
to_sfixed(-263184110.0/4294967296.0,1,-nbitq), 
to_sfixed(997297026.0/4294967296.0,1,-nbitq), 
to_sfixed(169257254.0/4294967296.0,1,-nbitq), 
to_sfixed(-2079852398.0/4294967296.0,1,-nbitq), 
to_sfixed(-179279479.0/4294967296.0,1,-nbitq), 
to_sfixed(992134394.0/4294967296.0,1,-nbitq), 
to_sfixed(-361538295.0/4294967296.0,1,-nbitq), 
to_sfixed(15372764.0/4294967296.0,1,-nbitq), 
to_sfixed(-1716437519.0/4294967296.0,1,-nbitq), 
to_sfixed(-263253276.0/4294967296.0,1,-nbitq), 
to_sfixed(959598502.0/4294967296.0,1,-nbitq), 
to_sfixed(726631455.0/4294967296.0,1,-nbitq), 
to_sfixed(-587633130.0/4294967296.0,1,-nbitq), 
to_sfixed(-124122885.0/4294967296.0,1,-nbitq), 
to_sfixed(809789979.0/4294967296.0,1,-nbitq), 
to_sfixed(573809271.0/4294967296.0,1,-nbitq), 
to_sfixed(64532816.0/4294967296.0,1,-nbitq), 
to_sfixed(1187414651.0/4294967296.0,1,-nbitq), 
to_sfixed(410416163.0/4294967296.0,1,-nbitq), 
to_sfixed(129801779.0/4294967296.0,1,-nbitq), 
to_sfixed(31952280.0/4294967296.0,1,-nbitq), 
to_sfixed(-220600552.0/4294967296.0,1,-nbitq), 
to_sfixed(509568246.0/4294967296.0,1,-nbitq), 
to_sfixed(-261441837.0/4294967296.0,1,-nbitq), 
to_sfixed(-1380683683.0/4294967296.0,1,-nbitq), 
to_sfixed(-638977734.0/4294967296.0,1,-nbitq), 
to_sfixed(-214134526.0/4294967296.0,1,-nbitq), 
to_sfixed(-1356023223.0/4294967296.0,1,-nbitq), 
to_sfixed(175086072.0/4294967296.0,1,-nbitq), 
to_sfixed(-1020229056.0/4294967296.0,1,-nbitq), 
to_sfixed(155220544.0/4294967296.0,1,-nbitq), 
to_sfixed(-789881066.0/4294967296.0,1,-nbitq), 
to_sfixed(-220382195.0/4294967296.0,1,-nbitq), 
to_sfixed(-429458740.0/4294967296.0,1,-nbitq), 
to_sfixed(-785999225.0/4294967296.0,1,-nbitq), 
to_sfixed(788854596.0/4294967296.0,1,-nbitq), 
to_sfixed(440535093.0/4294967296.0,1,-nbitq), 
to_sfixed(217316350.0/4294967296.0,1,-nbitq), 
to_sfixed(347896707.0/4294967296.0,1,-nbitq), 
to_sfixed(-68617961.0/4294967296.0,1,-nbitq), 
to_sfixed(-63368749.0/4294967296.0,1,-nbitq), 
to_sfixed(345691114.0/4294967296.0,1,-nbitq), 
to_sfixed(-177285914.0/4294967296.0,1,-nbitq), 
to_sfixed(-429218003.0/4294967296.0,1,-nbitq), 
to_sfixed(-87577521.0/4294967296.0,1,-nbitq), 
to_sfixed(143420137.0/4294967296.0,1,-nbitq), 
to_sfixed(638543981.0/4294967296.0,1,-nbitq), 
to_sfixed(-905796442.0/4294967296.0,1,-nbitq), 
to_sfixed(101606185.0/4294967296.0,1,-nbitq), 
to_sfixed(-1055203853.0/4294967296.0,1,-nbitq), 
to_sfixed(-939047213.0/4294967296.0,1,-nbitq), 
to_sfixed(-198313434.0/4294967296.0,1,-nbitq), 
to_sfixed(1229604042.0/4294967296.0,1,-nbitq), 
to_sfixed(-6038597.0/4294967296.0,1,-nbitq), 
to_sfixed(185826558.0/4294967296.0,1,-nbitq), 
to_sfixed(865345152.0/4294967296.0,1,-nbitq), 
to_sfixed(640962369.0/4294967296.0,1,-nbitq), 
to_sfixed(-223160465.0/4294967296.0,1,-nbitq), 
to_sfixed(1264466547.0/4294967296.0,1,-nbitq), 
to_sfixed(-41543565.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-181914165.0/4294967296.0,1,-nbitq), 
to_sfixed(1357792003.0/4294967296.0,1,-nbitq), 
to_sfixed(921929734.0/4294967296.0,1,-nbitq), 
to_sfixed(130876411.0/4294967296.0,1,-nbitq), 
to_sfixed(12923892.0/4294967296.0,1,-nbitq), 
to_sfixed(116603973.0/4294967296.0,1,-nbitq), 
to_sfixed(21242295.0/4294967296.0,1,-nbitq), 
to_sfixed(689790034.0/4294967296.0,1,-nbitq), 
to_sfixed(229805972.0/4294967296.0,1,-nbitq), 
to_sfixed(376052023.0/4294967296.0,1,-nbitq), 
to_sfixed(-84797210.0/4294967296.0,1,-nbitq), 
to_sfixed(-965462677.0/4294967296.0,1,-nbitq), 
to_sfixed(1673190943.0/4294967296.0,1,-nbitq), 
to_sfixed(64845005.0/4294967296.0,1,-nbitq), 
to_sfixed(64494656.0/4294967296.0,1,-nbitq), 
to_sfixed(-1278208464.0/4294967296.0,1,-nbitq), 
to_sfixed(-319162246.0/4294967296.0,1,-nbitq), 
to_sfixed(287669519.0/4294967296.0,1,-nbitq), 
to_sfixed(391089465.0/4294967296.0,1,-nbitq), 
to_sfixed(222232654.0/4294967296.0,1,-nbitq), 
to_sfixed(375972047.0/4294967296.0,1,-nbitq), 
to_sfixed(1093260323.0/4294967296.0,1,-nbitq), 
to_sfixed(479941984.0/4294967296.0,1,-nbitq), 
to_sfixed(-2528499312.0/4294967296.0,1,-nbitq), 
to_sfixed(-40125051.0/4294967296.0,1,-nbitq), 
to_sfixed(850405719.0/4294967296.0,1,-nbitq), 
to_sfixed(-181121864.0/4294967296.0,1,-nbitq), 
to_sfixed(-815831561.0/4294967296.0,1,-nbitq), 
to_sfixed(-1648257651.0/4294967296.0,1,-nbitq), 
to_sfixed(-618530281.0/4294967296.0,1,-nbitq), 
to_sfixed(905727385.0/4294967296.0,1,-nbitq), 
to_sfixed(992596291.0/4294967296.0,1,-nbitq), 
to_sfixed(-555552995.0/4294967296.0,1,-nbitq), 
to_sfixed(156731890.0/4294967296.0,1,-nbitq), 
to_sfixed(1080230763.0/4294967296.0,1,-nbitq), 
to_sfixed(501427411.0/4294967296.0,1,-nbitq), 
to_sfixed(-705703220.0/4294967296.0,1,-nbitq), 
to_sfixed(541896473.0/4294967296.0,1,-nbitq), 
to_sfixed(374704365.0/4294967296.0,1,-nbitq), 
to_sfixed(508342972.0/4294967296.0,1,-nbitq), 
to_sfixed(-1003435593.0/4294967296.0,1,-nbitq), 
to_sfixed(940856838.0/4294967296.0,1,-nbitq), 
to_sfixed(-677469772.0/4294967296.0,1,-nbitq), 
to_sfixed(257238184.0/4294967296.0,1,-nbitq), 
to_sfixed(-865739639.0/4294967296.0,1,-nbitq), 
to_sfixed(771016839.0/4294967296.0,1,-nbitq), 
to_sfixed(-371223624.0/4294967296.0,1,-nbitq), 
to_sfixed(-1119953808.0/4294967296.0,1,-nbitq), 
to_sfixed(-156763383.0/4294967296.0,1,-nbitq), 
to_sfixed(-1350006988.0/4294967296.0,1,-nbitq), 
to_sfixed(-67142363.0/4294967296.0,1,-nbitq), 
to_sfixed(2321538.0/4294967296.0,1,-nbitq), 
to_sfixed(-111018495.0/4294967296.0,1,-nbitq), 
to_sfixed(440287731.0/4294967296.0,1,-nbitq), 
to_sfixed(638515314.0/4294967296.0,1,-nbitq), 
to_sfixed(781662674.0/4294967296.0,1,-nbitq), 
to_sfixed(305629531.0/4294967296.0,1,-nbitq), 
to_sfixed(367366804.0/4294967296.0,1,-nbitq), 
to_sfixed(361062757.0/4294967296.0,1,-nbitq), 
to_sfixed(291207102.0/4294967296.0,1,-nbitq), 
to_sfixed(-212859842.0/4294967296.0,1,-nbitq), 
to_sfixed(223279777.0/4294967296.0,1,-nbitq), 
to_sfixed(-591241474.0/4294967296.0,1,-nbitq), 
to_sfixed(-1908753.0/4294967296.0,1,-nbitq), 
to_sfixed(-485198807.0/4294967296.0,1,-nbitq), 
to_sfixed(382828563.0/4294967296.0,1,-nbitq), 
to_sfixed(692193935.0/4294967296.0,1,-nbitq), 
to_sfixed(44793793.0/4294967296.0,1,-nbitq), 
to_sfixed(-258071059.0/4294967296.0,1,-nbitq), 
to_sfixed(-1184421576.0/4294967296.0,1,-nbitq), 
to_sfixed(-856384024.0/4294967296.0,1,-nbitq), 
to_sfixed(99846310.0/4294967296.0,1,-nbitq), 
to_sfixed(1035311093.0/4294967296.0,1,-nbitq), 
to_sfixed(-183597126.0/4294967296.0,1,-nbitq), 
to_sfixed(538899915.0/4294967296.0,1,-nbitq), 
to_sfixed(928543662.0/4294967296.0,1,-nbitq), 
to_sfixed(924837226.0/4294967296.0,1,-nbitq), 
to_sfixed(-61205341.0/4294967296.0,1,-nbitq), 
to_sfixed(307003597.0/4294967296.0,1,-nbitq), 
to_sfixed(-210791010.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-457285744.0/4294967296.0,1,-nbitq), 
to_sfixed(1455185636.0/4294967296.0,1,-nbitq), 
to_sfixed(827924449.0/4294967296.0,1,-nbitq), 
to_sfixed(-691706267.0/4294967296.0,1,-nbitq), 
to_sfixed(45984271.0/4294967296.0,1,-nbitq), 
to_sfixed(-523544256.0/4294967296.0,1,-nbitq), 
to_sfixed(-341940659.0/4294967296.0,1,-nbitq), 
to_sfixed(782874492.0/4294967296.0,1,-nbitq), 
to_sfixed(258128785.0/4294967296.0,1,-nbitq), 
to_sfixed(400084547.0/4294967296.0,1,-nbitq), 
to_sfixed(682581118.0/4294967296.0,1,-nbitq), 
to_sfixed(-1034991671.0/4294967296.0,1,-nbitq), 
to_sfixed(838810347.0/4294967296.0,1,-nbitq), 
to_sfixed(1049212490.0/4294967296.0,1,-nbitq), 
to_sfixed(-70046512.0/4294967296.0,1,-nbitq), 
to_sfixed(-809778773.0/4294967296.0,1,-nbitq), 
to_sfixed(396471587.0/4294967296.0,1,-nbitq), 
to_sfixed(149073458.0/4294967296.0,1,-nbitq), 
to_sfixed(192800615.0/4294967296.0,1,-nbitq), 
to_sfixed(910521862.0/4294967296.0,1,-nbitq), 
to_sfixed(-63675369.0/4294967296.0,1,-nbitq), 
to_sfixed(252668877.0/4294967296.0,1,-nbitq), 
to_sfixed(792367672.0/4294967296.0,1,-nbitq), 
to_sfixed(-835879554.0/4294967296.0,1,-nbitq), 
to_sfixed(13570741.0/4294967296.0,1,-nbitq), 
to_sfixed(-387984945.0/4294967296.0,1,-nbitq), 
to_sfixed(436305203.0/4294967296.0,1,-nbitq), 
to_sfixed(-737857856.0/4294967296.0,1,-nbitq), 
to_sfixed(-775077042.0/4294967296.0,1,-nbitq), 
to_sfixed(-420955598.0/4294967296.0,1,-nbitq), 
to_sfixed(-640328811.0/4294967296.0,1,-nbitq), 
to_sfixed(819908760.0/4294967296.0,1,-nbitq), 
to_sfixed(-662118607.0/4294967296.0,1,-nbitq), 
to_sfixed(475852414.0/4294967296.0,1,-nbitq), 
to_sfixed(96012041.0/4294967296.0,1,-nbitq), 
to_sfixed(471570727.0/4294967296.0,1,-nbitq), 
to_sfixed(-456909978.0/4294967296.0,1,-nbitq), 
to_sfixed(334792462.0/4294967296.0,1,-nbitq), 
to_sfixed(-449320649.0/4294967296.0,1,-nbitq), 
to_sfixed(296819627.0/4294967296.0,1,-nbitq), 
to_sfixed(-1001961467.0/4294967296.0,1,-nbitq), 
to_sfixed(606849125.0/4294967296.0,1,-nbitq), 
to_sfixed(-511606422.0/4294967296.0,1,-nbitq), 
to_sfixed(-878132638.0/4294967296.0,1,-nbitq), 
to_sfixed(-1071422295.0/4294967296.0,1,-nbitq), 
to_sfixed(138709320.0/4294967296.0,1,-nbitq), 
to_sfixed(-353075202.0/4294967296.0,1,-nbitq), 
to_sfixed(-1363974427.0/4294967296.0,1,-nbitq), 
to_sfixed(35002761.0/4294967296.0,1,-nbitq), 
to_sfixed(-347409914.0/4294967296.0,1,-nbitq), 
to_sfixed(60395208.0/4294967296.0,1,-nbitq), 
to_sfixed(28683748.0/4294967296.0,1,-nbitq), 
to_sfixed(405405880.0/4294967296.0,1,-nbitq), 
to_sfixed(145852169.0/4294967296.0,1,-nbitq), 
to_sfixed(305925641.0/4294967296.0,1,-nbitq), 
to_sfixed(-809106705.0/4294967296.0,1,-nbitq), 
to_sfixed(851848833.0/4294967296.0,1,-nbitq), 
to_sfixed(680317333.0/4294967296.0,1,-nbitq), 
to_sfixed(-202529410.0/4294967296.0,1,-nbitq), 
to_sfixed(12119857.0/4294967296.0,1,-nbitq), 
to_sfixed(171118945.0/4294967296.0,1,-nbitq), 
to_sfixed(-471046812.0/4294967296.0,1,-nbitq), 
to_sfixed(136318667.0/4294967296.0,1,-nbitq), 
to_sfixed(-554826817.0/4294967296.0,1,-nbitq), 
to_sfixed(-250674527.0/4294967296.0,1,-nbitq), 
to_sfixed(-151700101.0/4294967296.0,1,-nbitq), 
to_sfixed(-150689117.0/4294967296.0,1,-nbitq), 
to_sfixed(-711196662.0/4294967296.0,1,-nbitq), 
to_sfixed(-174829030.0/4294967296.0,1,-nbitq), 
to_sfixed(-1246471279.0/4294967296.0,1,-nbitq), 
to_sfixed(-1279278375.0/4294967296.0,1,-nbitq), 
to_sfixed(-616113910.0/4294967296.0,1,-nbitq), 
to_sfixed(508270737.0/4294967296.0,1,-nbitq), 
to_sfixed(292805416.0/4294967296.0,1,-nbitq), 
to_sfixed(52989125.0/4294967296.0,1,-nbitq), 
to_sfixed(939994841.0/4294967296.0,1,-nbitq), 
to_sfixed(697328715.0/4294967296.0,1,-nbitq), 
to_sfixed(547676568.0/4294967296.0,1,-nbitq), 
to_sfixed(-30329609.0/4294967296.0,1,-nbitq), 
to_sfixed(-327663710.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-347791409.0/4294967296.0,1,-nbitq), 
to_sfixed(885788021.0/4294967296.0,1,-nbitq), 
to_sfixed(165658569.0/4294967296.0,1,-nbitq), 
to_sfixed(-745706781.0/4294967296.0,1,-nbitq), 
to_sfixed(896362839.0/4294967296.0,1,-nbitq), 
to_sfixed(-749960531.0/4294967296.0,1,-nbitq), 
to_sfixed(-282532585.0/4294967296.0,1,-nbitq), 
to_sfixed(172466081.0/4294967296.0,1,-nbitq), 
to_sfixed(753644476.0/4294967296.0,1,-nbitq), 
to_sfixed(-410788147.0/4294967296.0,1,-nbitq), 
to_sfixed(469983197.0/4294967296.0,1,-nbitq), 
to_sfixed(-990316178.0/4294967296.0,1,-nbitq), 
to_sfixed(1128770639.0/4294967296.0,1,-nbitq), 
to_sfixed(732306628.0/4294967296.0,1,-nbitq), 
to_sfixed(253299430.0/4294967296.0,1,-nbitq), 
to_sfixed(-225962020.0/4294967296.0,1,-nbitq), 
to_sfixed(352677276.0/4294967296.0,1,-nbitq), 
to_sfixed(-254410119.0/4294967296.0,1,-nbitq), 
to_sfixed(16125951.0/4294967296.0,1,-nbitq), 
to_sfixed(551275168.0/4294967296.0,1,-nbitq), 
to_sfixed(57230858.0/4294967296.0,1,-nbitq), 
to_sfixed(-611999206.0/4294967296.0,1,-nbitq), 
to_sfixed(546002726.0/4294967296.0,1,-nbitq), 
to_sfixed(-27378159.0/4294967296.0,1,-nbitq), 
to_sfixed(363527534.0/4294967296.0,1,-nbitq), 
to_sfixed(-1149816326.0/4294967296.0,1,-nbitq), 
to_sfixed(121212998.0/4294967296.0,1,-nbitq), 
to_sfixed(-693030882.0/4294967296.0,1,-nbitq), 
to_sfixed(564701295.0/4294967296.0,1,-nbitq), 
to_sfixed(-734727340.0/4294967296.0,1,-nbitq), 
to_sfixed(-410405954.0/4294967296.0,1,-nbitq), 
to_sfixed(432269139.0/4294967296.0,1,-nbitq), 
to_sfixed(-987239211.0/4294967296.0,1,-nbitq), 
to_sfixed(261701108.0/4294967296.0,1,-nbitq), 
to_sfixed(-728281350.0/4294967296.0,1,-nbitq), 
to_sfixed(870266331.0/4294967296.0,1,-nbitq), 
to_sfixed(-508441320.0/4294967296.0,1,-nbitq), 
to_sfixed(-210711640.0/4294967296.0,1,-nbitq), 
to_sfixed(-420965473.0/4294967296.0,1,-nbitq), 
to_sfixed(387952373.0/4294967296.0,1,-nbitq), 
to_sfixed(-495383659.0/4294967296.0,1,-nbitq), 
to_sfixed(1508812119.0/4294967296.0,1,-nbitq), 
to_sfixed(-123278852.0/4294967296.0,1,-nbitq), 
to_sfixed(-836490095.0/4294967296.0,1,-nbitq), 
to_sfixed(-1417888884.0/4294967296.0,1,-nbitq), 
to_sfixed(658339155.0/4294967296.0,1,-nbitq), 
to_sfixed(91995723.0/4294967296.0,1,-nbitq), 
to_sfixed(-552822565.0/4294967296.0,1,-nbitq), 
to_sfixed(363124916.0/4294967296.0,1,-nbitq), 
to_sfixed(-23244483.0/4294967296.0,1,-nbitq), 
to_sfixed(-83381524.0/4294967296.0,1,-nbitq), 
to_sfixed(235576160.0/4294967296.0,1,-nbitq), 
to_sfixed(14455025.0/4294967296.0,1,-nbitq), 
to_sfixed(1017120775.0/4294967296.0,1,-nbitq), 
to_sfixed(1045373451.0/4294967296.0,1,-nbitq), 
to_sfixed(-1564213752.0/4294967296.0,1,-nbitq), 
to_sfixed(173887613.0/4294967296.0,1,-nbitq), 
to_sfixed(912113178.0/4294967296.0,1,-nbitq), 
to_sfixed(-14654816.0/4294967296.0,1,-nbitq), 
to_sfixed(-26211792.0/4294967296.0,1,-nbitq), 
to_sfixed(38640191.0/4294967296.0,1,-nbitq), 
to_sfixed(252818971.0/4294967296.0,1,-nbitq), 
to_sfixed(785183476.0/4294967296.0,1,-nbitq), 
to_sfixed(-322470801.0/4294967296.0,1,-nbitq), 
to_sfixed(282564855.0/4294967296.0,1,-nbitq), 
to_sfixed(-503084353.0/4294967296.0,1,-nbitq), 
to_sfixed(-999303509.0/4294967296.0,1,-nbitq), 
to_sfixed(-302530174.0/4294967296.0,1,-nbitq), 
to_sfixed(110668957.0/4294967296.0,1,-nbitq), 
to_sfixed(-1017306501.0/4294967296.0,1,-nbitq), 
to_sfixed(-162158987.0/4294967296.0,1,-nbitq), 
to_sfixed(-170757494.0/4294967296.0,1,-nbitq), 
to_sfixed(-737323135.0/4294967296.0,1,-nbitq), 
to_sfixed(-223019507.0/4294967296.0,1,-nbitq), 
to_sfixed(518956109.0/4294967296.0,1,-nbitq), 
to_sfixed(-521902392.0/4294967296.0,1,-nbitq), 
to_sfixed(379878231.0/4294967296.0,1,-nbitq), 
to_sfixed(423708198.0/4294967296.0,1,-nbitq), 
to_sfixed(-570484816.0/4294967296.0,1,-nbitq), 
to_sfixed(217770394.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(360260804.0/4294967296.0,1,-nbitq), 
to_sfixed(1048205807.0/4294967296.0,1,-nbitq), 
to_sfixed(-748467261.0/4294967296.0,1,-nbitq), 
to_sfixed(-1900988125.0/4294967296.0,1,-nbitq), 
to_sfixed(205600281.0/4294967296.0,1,-nbitq), 
to_sfixed(-415351955.0/4294967296.0,1,-nbitq), 
to_sfixed(-187469726.0/4294967296.0,1,-nbitq), 
to_sfixed(-594031945.0/4294967296.0,1,-nbitq), 
to_sfixed(-528474641.0/4294967296.0,1,-nbitq), 
to_sfixed(155824315.0/4294967296.0,1,-nbitq), 
to_sfixed(-138638749.0/4294967296.0,1,-nbitq), 
to_sfixed(-1374676546.0/4294967296.0,1,-nbitq), 
to_sfixed(261449919.0/4294967296.0,1,-nbitq), 
to_sfixed(370619869.0/4294967296.0,1,-nbitq), 
to_sfixed(461877125.0/4294967296.0,1,-nbitq), 
to_sfixed(-726771279.0/4294967296.0,1,-nbitq), 
to_sfixed(-376777427.0/4294967296.0,1,-nbitq), 
to_sfixed(3846187.0/4294967296.0,1,-nbitq), 
to_sfixed(409061859.0/4294967296.0,1,-nbitq), 
to_sfixed(193873196.0/4294967296.0,1,-nbitq), 
to_sfixed(153410386.0/4294967296.0,1,-nbitq), 
to_sfixed(-26646420.0/4294967296.0,1,-nbitq), 
to_sfixed(437978990.0/4294967296.0,1,-nbitq), 
to_sfixed(-28448988.0/4294967296.0,1,-nbitq), 
to_sfixed(374260125.0/4294967296.0,1,-nbitq), 
to_sfixed(-188610965.0/4294967296.0,1,-nbitq), 
to_sfixed(177740469.0/4294967296.0,1,-nbitq), 
to_sfixed(-300146696.0/4294967296.0,1,-nbitq), 
to_sfixed(1094772607.0/4294967296.0,1,-nbitq), 
to_sfixed(-411043477.0/4294967296.0,1,-nbitq), 
to_sfixed(-156322680.0/4294967296.0,1,-nbitq), 
to_sfixed(784112427.0/4294967296.0,1,-nbitq), 
to_sfixed(-686825207.0/4294967296.0,1,-nbitq), 
to_sfixed(-166204319.0/4294967296.0,1,-nbitq), 
to_sfixed(-568022240.0/4294967296.0,1,-nbitq), 
to_sfixed(-89162225.0/4294967296.0,1,-nbitq), 
to_sfixed(-653131000.0/4294967296.0,1,-nbitq), 
to_sfixed(-293969821.0/4294967296.0,1,-nbitq), 
to_sfixed(-392611967.0/4294967296.0,1,-nbitq), 
to_sfixed(488491344.0/4294967296.0,1,-nbitq), 
to_sfixed(-481181391.0/4294967296.0,1,-nbitq), 
to_sfixed(505961228.0/4294967296.0,1,-nbitq), 
to_sfixed(635103040.0/4294967296.0,1,-nbitq), 
to_sfixed(189117694.0/4294967296.0,1,-nbitq), 
to_sfixed(-1009268668.0/4294967296.0,1,-nbitq), 
to_sfixed(1246322922.0/4294967296.0,1,-nbitq), 
to_sfixed(67437758.0/4294967296.0,1,-nbitq), 
to_sfixed(-559403184.0/4294967296.0,1,-nbitq), 
to_sfixed(-313970575.0/4294967296.0,1,-nbitq), 
to_sfixed(-223340656.0/4294967296.0,1,-nbitq), 
to_sfixed(304751790.0/4294967296.0,1,-nbitq), 
to_sfixed(-201301629.0/4294967296.0,1,-nbitq), 
to_sfixed(-184824602.0/4294967296.0,1,-nbitq), 
to_sfixed(1211439708.0/4294967296.0,1,-nbitq), 
to_sfixed(467754728.0/4294967296.0,1,-nbitq), 
to_sfixed(-1083819263.0/4294967296.0,1,-nbitq), 
to_sfixed(368552401.0/4294967296.0,1,-nbitq), 
to_sfixed(582648020.0/4294967296.0,1,-nbitq), 
to_sfixed(162330240.0/4294967296.0,1,-nbitq), 
to_sfixed(-350483697.0/4294967296.0,1,-nbitq), 
to_sfixed(195307695.0/4294967296.0,1,-nbitq), 
to_sfixed(-97626211.0/4294967296.0,1,-nbitq), 
to_sfixed(949892601.0/4294967296.0,1,-nbitq), 
to_sfixed(130020268.0/4294967296.0,1,-nbitq), 
to_sfixed(-104567205.0/4294967296.0,1,-nbitq), 
to_sfixed(136576309.0/4294967296.0,1,-nbitq), 
to_sfixed(-1443086687.0/4294967296.0,1,-nbitq), 
to_sfixed(-277964688.0/4294967296.0,1,-nbitq), 
to_sfixed(67708726.0/4294967296.0,1,-nbitq), 
to_sfixed(-1272104770.0/4294967296.0,1,-nbitq), 
to_sfixed(166362562.0/4294967296.0,1,-nbitq), 
to_sfixed(71428734.0/4294967296.0,1,-nbitq), 
to_sfixed(-829257870.0/4294967296.0,1,-nbitq), 
to_sfixed(233576203.0/4294967296.0,1,-nbitq), 
to_sfixed(475391940.0/4294967296.0,1,-nbitq), 
to_sfixed(36272218.0/4294967296.0,1,-nbitq), 
to_sfixed(-326468770.0/4294967296.0,1,-nbitq), 
to_sfixed(243395208.0/4294967296.0,1,-nbitq), 
to_sfixed(-617260246.0/4294967296.0,1,-nbitq), 
to_sfixed(50396879.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(232277335.0/4294967296.0,1,-nbitq), 
to_sfixed(780267647.0/4294967296.0,1,-nbitq), 
to_sfixed(-1013847585.0/4294967296.0,1,-nbitq), 
to_sfixed(-1278040931.0/4294967296.0,1,-nbitq), 
to_sfixed(943119119.0/4294967296.0,1,-nbitq), 
to_sfixed(-767192494.0/4294967296.0,1,-nbitq), 
to_sfixed(-170321132.0/4294967296.0,1,-nbitq), 
to_sfixed(-606449182.0/4294967296.0,1,-nbitq), 
to_sfixed(126366995.0/4294967296.0,1,-nbitq), 
to_sfixed(186430875.0/4294967296.0,1,-nbitq), 
to_sfixed(-339506320.0/4294967296.0,1,-nbitq), 
to_sfixed(-1608127952.0/4294967296.0,1,-nbitq), 
to_sfixed(508980604.0/4294967296.0,1,-nbitq), 
to_sfixed(699012530.0/4294967296.0,1,-nbitq), 
to_sfixed(475488646.0/4294967296.0,1,-nbitq), 
to_sfixed(-240729751.0/4294967296.0,1,-nbitq), 
to_sfixed(325014732.0/4294967296.0,1,-nbitq), 
to_sfixed(48670812.0/4294967296.0,1,-nbitq), 
to_sfixed(629615373.0/4294967296.0,1,-nbitq), 
to_sfixed(115037337.0/4294967296.0,1,-nbitq), 
to_sfixed(139723444.0/4294967296.0,1,-nbitq), 
to_sfixed(-226034438.0/4294967296.0,1,-nbitq), 
to_sfixed(119962267.0/4294967296.0,1,-nbitq), 
to_sfixed(527765520.0/4294967296.0,1,-nbitq), 
to_sfixed(-300471443.0/4294967296.0,1,-nbitq), 
to_sfixed(709985133.0/4294967296.0,1,-nbitq), 
to_sfixed(10184128.0/4294967296.0,1,-nbitq), 
to_sfixed(-433065615.0/4294967296.0,1,-nbitq), 
to_sfixed(322431663.0/4294967296.0,1,-nbitq), 
to_sfixed(-637038888.0/4294967296.0,1,-nbitq), 
to_sfixed(-673607182.0/4294967296.0,1,-nbitq), 
to_sfixed(642014772.0/4294967296.0,1,-nbitq), 
to_sfixed(-632325978.0/4294967296.0,1,-nbitq), 
to_sfixed(-71860094.0/4294967296.0,1,-nbitq), 
to_sfixed(21238581.0/4294967296.0,1,-nbitq), 
to_sfixed(434263063.0/4294967296.0,1,-nbitq), 
to_sfixed(91436579.0/4294967296.0,1,-nbitq), 
to_sfixed(-5225378.0/4294967296.0,1,-nbitq), 
to_sfixed(-140623142.0/4294967296.0,1,-nbitq), 
to_sfixed(586362057.0/4294967296.0,1,-nbitq), 
to_sfixed(-144110641.0/4294967296.0,1,-nbitq), 
to_sfixed(639263509.0/4294967296.0,1,-nbitq), 
to_sfixed(148954211.0/4294967296.0,1,-nbitq), 
to_sfixed(-142339915.0/4294967296.0,1,-nbitq), 
to_sfixed(-486630020.0/4294967296.0,1,-nbitq), 
to_sfixed(548830262.0/4294967296.0,1,-nbitq), 
to_sfixed(148309133.0/4294967296.0,1,-nbitq), 
to_sfixed(-553842050.0/4294967296.0,1,-nbitq), 
to_sfixed(-7738422.0/4294967296.0,1,-nbitq), 
to_sfixed(268801072.0/4294967296.0,1,-nbitq), 
to_sfixed(244527068.0/4294967296.0,1,-nbitq), 
to_sfixed(-486164901.0/4294967296.0,1,-nbitq), 
to_sfixed(-485881712.0/4294967296.0,1,-nbitq), 
to_sfixed(618951150.0/4294967296.0,1,-nbitq), 
to_sfixed(-81396712.0/4294967296.0,1,-nbitq), 
to_sfixed(-204411671.0/4294967296.0,1,-nbitq), 
to_sfixed(103543832.0/4294967296.0,1,-nbitq), 
to_sfixed(918020028.0/4294967296.0,1,-nbitq), 
to_sfixed(-47640834.0/4294967296.0,1,-nbitq), 
to_sfixed(340939783.0/4294967296.0,1,-nbitq), 
to_sfixed(236544246.0/4294967296.0,1,-nbitq), 
to_sfixed(-357656490.0/4294967296.0,1,-nbitq), 
to_sfixed(71109588.0/4294967296.0,1,-nbitq), 
to_sfixed(-254692391.0/4294967296.0,1,-nbitq), 
to_sfixed(-395829496.0/4294967296.0,1,-nbitq), 
to_sfixed(-343586115.0/4294967296.0,1,-nbitq), 
to_sfixed(-1113765276.0/4294967296.0,1,-nbitq), 
to_sfixed(-479446679.0/4294967296.0,1,-nbitq), 
to_sfixed(298504347.0/4294967296.0,1,-nbitq), 
to_sfixed(-857967708.0/4294967296.0,1,-nbitq), 
to_sfixed(-280824281.0/4294967296.0,1,-nbitq), 
to_sfixed(405874777.0/4294967296.0,1,-nbitq), 
to_sfixed(-1033304453.0/4294967296.0,1,-nbitq), 
to_sfixed(383200287.0/4294967296.0,1,-nbitq), 
to_sfixed(148826991.0/4294967296.0,1,-nbitq), 
to_sfixed(618565733.0/4294967296.0,1,-nbitq), 
to_sfixed(68743131.0/4294967296.0,1,-nbitq), 
to_sfixed(312453779.0/4294967296.0,1,-nbitq), 
to_sfixed(-439592019.0/4294967296.0,1,-nbitq), 
to_sfixed(279023674.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-198582203.0/4294967296.0,1,-nbitq), 
to_sfixed(643143933.0/4294967296.0,1,-nbitq), 
to_sfixed(-718345204.0/4294967296.0,1,-nbitq), 
to_sfixed(-301799862.0/4294967296.0,1,-nbitq), 
to_sfixed(745953267.0/4294967296.0,1,-nbitq), 
to_sfixed(-274755998.0/4294967296.0,1,-nbitq), 
to_sfixed(-299555389.0/4294967296.0,1,-nbitq), 
to_sfixed(40674696.0/4294967296.0,1,-nbitq), 
to_sfixed(252281187.0/4294967296.0,1,-nbitq), 
to_sfixed(-354244864.0/4294967296.0,1,-nbitq), 
to_sfixed(-415709860.0/4294967296.0,1,-nbitq), 
to_sfixed(-525355621.0/4294967296.0,1,-nbitq), 
to_sfixed(1224220660.0/4294967296.0,1,-nbitq), 
to_sfixed(-430765266.0/4294967296.0,1,-nbitq), 
to_sfixed(387820090.0/4294967296.0,1,-nbitq), 
to_sfixed(-86852975.0/4294967296.0,1,-nbitq), 
to_sfixed(-86637883.0/4294967296.0,1,-nbitq), 
to_sfixed(-296900861.0/4294967296.0,1,-nbitq), 
to_sfixed(180853941.0/4294967296.0,1,-nbitq), 
to_sfixed(-36745753.0/4294967296.0,1,-nbitq), 
to_sfixed(245926256.0/4294967296.0,1,-nbitq), 
to_sfixed(639134208.0/4294967296.0,1,-nbitq), 
to_sfixed(-598123029.0/4294967296.0,1,-nbitq), 
to_sfixed(111851259.0/4294967296.0,1,-nbitq), 
to_sfixed(-269458870.0/4294967296.0,1,-nbitq), 
to_sfixed(910720432.0/4294967296.0,1,-nbitq), 
to_sfixed(-530917807.0/4294967296.0,1,-nbitq), 
to_sfixed(212817846.0/4294967296.0,1,-nbitq), 
to_sfixed(39623028.0/4294967296.0,1,-nbitq), 
to_sfixed(-111658832.0/4294967296.0,1,-nbitq), 
to_sfixed(-374349645.0/4294967296.0,1,-nbitq), 
to_sfixed(721457714.0/4294967296.0,1,-nbitq), 
to_sfixed(-160566633.0/4294967296.0,1,-nbitq), 
to_sfixed(-29422167.0/4294967296.0,1,-nbitq), 
to_sfixed(-99553762.0/4294967296.0,1,-nbitq), 
to_sfixed(636370939.0/4294967296.0,1,-nbitq), 
to_sfixed(224736962.0/4294967296.0,1,-nbitq), 
to_sfixed(-671712048.0/4294967296.0,1,-nbitq), 
to_sfixed(174014314.0/4294967296.0,1,-nbitq), 
to_sfixed(-70893002.0/4294967296.0,1,-nbitq), 
to_sfixed(305755730.0/4294967296.0,1,-nbitq), 
to_sfixed(580446749.0/4294967296.0,1,-nbitq), 
to_sfixed(-306288488.0/4294967296.0,1,-nbitq), 
to_sfixed(-475143538.0/4294967296.0,1,-nbitq), 
to_sfixed(-329609110.0/4294967296.0,1,-nbitq), 
to_sfixed(891315879.0/4294967296.0,1,-nbitq), 
to_sfixed(-245336236.0/4294967296.0,1,-nbitq), 
to_sfixed(-181618898.0/4294967296.0,1,-nbitq), 
to_sfixed(-232782406.0/4294967296.0,1,-nbitq), 
to_sfixed(443023524.0/4294967296.0,1,-nbitq), 
to_sfixed(324796980.0/4294967296.0,1,-nbitq), 
to_sfixed(-1209068637.0/4294967296.0,1,-nbitq), 
to_sfixed(330399877.0/4294967296.0,1,-nbitq), 
to_sfixed(254327357.0/4294967296.0,1,-nbitq), 
to_sfixed(121314488.0/4294967296.0,1,-nbitq), 
to_sfixed(-130573819.0/4294967296.0,1,-nbitq), 
to_sfixed(2396182.0/4294967296.0,1,-nbitq), 
to_sfixed(31435769.0/4294967296.0,1,-nbitq), 
to_sfixed(33825019.0/4294967296.0,1,-nbitq), 
to_sfixed(-197052426.0/4294967296.0,1,-nbitq), 
to_sfixed(-174938330.0/4294967296.0,1,-nbitq), 
to_sfixed(-653418474.0/4294967296.0,1,-nbitq), 
to_sfixed(-423581827.0/4294967296.0,1,-nbitq), 
to_sfixed(180585549.0/4294967296.0,1,-nbitq), 
to_sfixed(252296030.0/4294967296.0,1,-nbitq), 
to_sfixed(56616356.0/4294967296.0,1,-nbitq), 
to_sfixed(-74562927.0/4294967296.0,1,-nbitq), 
to_sfixed(129294170.0/4294967296.0,1,-nbitq), 
to_sfixed(132122718.0/4294967296.0,1,-nbitq), 
to_sfixed(-290433184.0/4294967296.0,1,-nbitq), 
to_sfixed(89509954.0/4294967296.0,1,-nbitq), 
to_sfixed(192137758.0/4294967296.0,1,-nbitq), 
to_sfixed(-246376168.0/4294967296.0,1,-nbitq), 
to_sfixed(278928482.0/4294967296.0,1,-nbitq), 
to_sfixed(511155033.0/4294967296.0,1,-nbitq), 
to_sfixed(386273913.0/4294967296.0,1,-nbitq), 
to_sfixed(410146931.0/4294967296.0,1,-nbitq), 
to_sfixed(30325045.0/4294967296.0,1,-nbitq), 
to_sfixed(-509214316.0/4294967296.0,1,-nbitq), 
to_sfixed(-22245973.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-521161493.0/4294967296.0,1,-nbitq), 
to_sfixed(897464663.0/4294967296.0,1,-nbitq), 
to_sfixed(-509156561.0/4294967296.0,1,-nbitq), 
to_sfixed(-757724745.0/4294967296.0,1,-nbitq), 
to_sfixed(189675556.0/4294967296.0,1,-nbitq), 
to_sfixed(-310475855.0/4294967296.0,1,-nbitq), 
to_sfixed(163237464.0/4294967296.0,1,-nbitq), 
to_sfixed(748741944.0/4294967296.0,1,-nbitq), 
to_sfixed(66598689.0/4294967296.0,1,-nbitq), 
to_sfixed(-35714705.0/4294967296.0,1,-nbitq), 
to_sfixed(341848493.0/4294967296.0,1,-nbitq), 
to_sfixed(-107947506.0/4294967296.0,1,-nbitq), 
to_sfixed(248511120.0/4294967296.0,1,-nbitq), 
to_sfixed(-112755388.0/4294967296.0,1,-nbitq), 
to_sfixed(-342676590.0/4294967296.0,1,-nbitq), 
to_sfixed(-391376724.0/4294967296.0,1,-nbitq), 
to_sfixed(21306638.0/4294967296.0,1,-nbitq), 
to_sfixed(331694001.0/4294967296.0,1,-nbitq), 
to_sfixed(386341540.0/4294967296.0,1,-nbitq), 
to_sfixed(17482258.0/4294967296.0,1,-nbitq), 
to_sfixed(-7513505.0/4294967296.0,1,-nbitq), 
to_sfixed(-78005066.0/4294967296.0,1,-nbitq), 
to_sfixed(-614814259.0/4294967296.0,1,-nbitq), 
to_sfixed(140284941.0/4294967296.0,1,-nbitq), 
to_sfixed(289210018.0/4294967296.0,1,-nbitq), 
to_sfixed(754986921.0/4294967296.0,1,-nbitq), 
to_sfixed(-603251650.0/4294967296.0,1,-nbitq), 
to_sfixed(840521690.0/4294967296.0,1,-nbitq), 
to_sfixed(278850668.0/4294967296.0,1,-nbitq), 
to_sfixed(-555134127.0/4294967296.0,1,-nbitq), 
to_sfixed(-155365430.0/4294967296.0,1,-nbitq), 
to_sfixed(189439054.0/4294967296.0,1,-nbitq), 
to_sfixed(146741683.0/4294967296.0,1,-nbitq), 
to_sfixed(-327920544.0/4294967296.0,1,-nbitq), 
to_sfixed(215268271.0/4294967296.0,1,-nbitq), 
to_sfixed(661742863.0/4294967296.0,1,-nbitq), 
to_sfixed(372969212.0/4294967296.0,1,-nbitq), 
to_sfixed(54393356.0/4294967296.0,1,-nbitq), 
to_sfixed(93647732.0/4294967296.0,1,-nbitq), 
to_sfixed(-3088195.0/4294967296.0,1,-nbitq), 
to_sfixed(397452999.0/4294967296.0,1,-nbitq), 
to_sfixed(6393135.0/4294967296.0,1,-nbitq), 
to_sfixed(-104453156.0/4294967296.0,1,-nbitq), 
to_sfixed(-776217638.0/4294967296.0,1,-nbitq), 
to_sfixed(-341423127.0/4294967296.0,1,-nbitq), 
to_sfixed(-54427223.0/4294967296.0,1,-nbitq), 
to_sfixed(-51314470.0/4294967296.0,1,-nbitq), 
to_sfixed(-359107184.0/4294967296.0,1,-nbitq), 
to_sfixed(-292107064.0/4294967296.0,1,-nbitq), 
to_sfixed(-300148995.0/4294967296.0,1,-nbitq), 
to_sfixed(52336571.0/4294967296.0,1,-nbitq), 
to_sfixed(-155451927.0/4294967296.0,1,-nbitq), 
to_sfixed(-261891568.0/4294967296.0,1,-nbitq), 
to_sfixed(684714716.0/4294967296.0,1,-nbitq), 
to_sfixed(24716215.0/4294967296.0,1,-nbitq), 
to_sfixed(-232884973.0/4294967296.0,1,-nbitq), 
to_sfixed(573945966.0/4294967296.0,1,-nbitq), 
to_sfixed(21391541.0/4294967296.0,1,-nbitq), 
to_sfixed(282157865.0/4294967296.0,1,-nbitq), 
to_sfixed(111238088.0/4294967296.0,1,-nbitq), 
to_sfixed(301212756.0/4294967296.0,1,-nbitq), 
to_sfixed(-494691106.0/4294967296.0,1,-nbitq), 
to_sfixed(472637824.0/4294967296.0,1,-nbitq), 
to_sfixed(22333995.0/4294967296.0,1,-nbitq), 
to_sfixed(-13933223.0/4294967296.0,1,-nbitq), 
to_sfixed(-225422256.0/4294967296.0,1,-nbitq), 
to_sfixed(-548037278.0/4294967296.0,1,-nbitq), 
to_sfixed(-386763084.0/4294967296.0,1,-nbitq), 
to_sfixed(185798500.0/4294967296.0,1,-nbitq), 
to_sfixed(386941092.0/4294967296.0,1,-nbitq), 
to_sfixed(287331132.0/4294967296.0,1,-nbitq), 
to_sfixed(-197260639.0/4294967296.0,1,-nbitq), 
to_sfixed(126117980.0/4294967296.0,1,-nbitq), 
to_sfixed(-234928483.0/4294967296.0,1,-nbitq), 
to_sfixed(212146246.0/4294967296.0,1,-nbitq), 
to_sfixed(339442181.0/4294967296.0,1,-nbitq), 
to_sfixed(-675804857.0/4294967296.0,1,-nbitq), 
to_sfixed(-74476708.0/4294967296.0,1,-nbitq), 
to_sfixed(-757851659.0/4294967296.0,1,-nbitq), 
to_sfixed(340766414.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-20282447.0/4294967296.0,1,-nbitq), 
to_sfixed(942464620.0/4294967296.0,1,-nbitq), 
to_sfixed(-739415275.0/4294967296.0,1,-nbitq), 
to_sfixed(-276755093.0/4294967296.0,1,-nbitq), 
to_sfixed(-105298609.0/4294967296.0,1,-nbitq), 
to_sfixed(-197098728.0/4294967296.0,1,-nbitq), 
to_sfixed(42546754.0/4294967296.0,1,-nbitq), 
to_sfixed(-91641132.0/4294967296.0,1,-nbitq), 
to_sfixed(-478418299.0/4294967296.0,1,-nbitq), 
to_sfixed(399474671.0/4294967296.0,1,-nbitq), 
to_sfixed(808719790.0/4294967296.0,1,-nbitq), 
to_sfixed(758449756.0/4294967296.0,1,-nbitq), 
to_sfixed(81644766.0/4294967296.0,1,-nbitq), 
to_sfixed(-332028058.0/4294967296.0,1,-nbitq), 
to_sfixed(11925962.0/4294967296.0,1,-nbitq), 
to_sfixed(-201405325.0/4294967296.0,1,-nbitq), 
to_sfixed(9781901.0/4294967296.0,1,-nbitq), 
to_sfixed(-110175714.0/4294967296.0,1,-nbitq), 
to_sfixed(768627935.0/4294967296.0,1,-nbitq), 
to_sfixed(406886130.0/4294967296.0,1,-nbitq), 
to_sfixed(-147887433.0/4294967296.0,1,-nbitq), 
to_sfixed(341631241.0/4294967296.0,1,-nbitq), 
to_sfixed(-279986963.0/4294967296.0,1,-nbitq), 
to_sfixed(-42092649.0/4294967296.0,1,-nbitq), 
to_sfixed(182568123.0/4294967296.0,1,-nbitq), 
to_sfixed(716323461.0/4294967296.0,1,-nbitq), 
to_sfixed(-797434975.0/4294967296.0,1,-nbitq), 
to_sfixed(492947047.0/4294967296.0,1,-nbitq), 
to_sfixed(-350699702.0/4294967296.0,1,-nbitq), 
to_sfixed(-100051085.0/4294967296.0,1,-nbitq), 
to_sfixed(256291885.0/4294967296.0,1,-nbitq), 
to_sfixed(761233538.0/4294967296.0,1,-nbitq), 
to_sfixed(194135190.0/4294967296.0,1,-nbitq), 
to_sfixed(-70899571.0/4294967296.0,1,-nbitq), 
to_sfixed(265502408.0/4294967296.0,1,-nbitq), 
to_sfixed(178900482.0/4294967296.0,1,-nbitq), 
to_sfixed(-383636969.0/4294967296.0,1,-nbitq), 
to_sfixed(-747727376.0/4294967296.0,1,-nbitq), 
to_sfixed(422503572.0/4294967296.0,1,-nbitq), 
to_sfixed(-122846166.0/4294967296.0,1,-nbitq), 
to_sfixed(506007305.0/4294967296.0,1,-nbitq), 
to_sfixed(55078640.0/4294967296.0,1,-nbitq), 
to_sfixed(604921309.0/4294967296.0,1,-nbitq), 
to_sfixed(-718606426.0/4294967296.0,1,-nbitq), 
to_sfixed(290165067.0/4294967296.0,1,-nbitq), 
to_sfixed(-549255486.0/4294967296.0,1,-nbitq), 
to_sfixed(257219867.0/4294967296.0,1,-nbitq), 
to_sfixed(-286384406.0/4294967296.0,1,-nbitq), 
to_sfixed(-799035000.0/4294967296.0,1,-nbitq), 
to_sfixed(-275602019.0/4294967296.0,1,-nbitq), 
to_sfixed(-455293281.0/4294967296.0,1,-nbitq), 
to_sfixed(261134047.0/4294967296.0,1,-nbitq), 
to_sfixed(-461256431.0/4294967296.0,1,-nbitq), 
to_sfixed(380317356.0/4294967296.0,1,-nbitq), 
to_sfixed(15071746.0/4294967296.0,1,-nbitq), 
to_sfixed(-825365422.0/4294967296.0,1,-nbitq), 
to_sfixed(131463601.0/4294967296.0,1,-nbitq), 
to_sfixed(-331840770.0/4294967296.0,1,-nbitq), 
to_sfixed(-27191151.0/4294967296.0,1,-nbitq), 
to_sfixed(292842591.0/4294967296.0,1,-nbitq), 
to_sfixed(-390336145.0/4294967296.0,1,-nbitq), 
to_sfixed(-716309112.0/4294967296.0,1,-nbitq), 
to_sfixed(105157596.0/4294967296.0,1,-nbitq), 
to_sfixed(383657569.0/4294967296.0,1,-nbitq), 
to_sfixed(385936414.0/4294967296.0,1,-nbitq), 
to_sfixed(145171534.0/4294967296.0,1,-nbitq), 
to_sfixed(-627042644.0/4294967296.0,1,-nbitq), 
to_sfixed(-724043169.0/4294967296.0,1,-nbitq), 
to_sfixed(148649171.0/4294967296.0,1,-nbitq), 
to_sfixed(-93027568.0/4294967296.0,1,-nbitq), 
to_sfixed(467966564.0/4294967296.0,1,-nbitq), 
to_sfixed(377358296.0/4294967296.0,1,-nbitq), 
to_sfixed(57367684.0/4294967296.0,1,-nbitq), 
to_sfixed(360015742.0/4294967296.0,1,-nbitq), 
to_sfixed(210685373.0/4294967296.0,1,-nbitq), 
to_sfixed(421888510.0/4294967296.0,1,-nbitq), 
to_sfixed(-244714610.0/4294967296.0,1,-nbitq), 
to_sfixed(-77325232.0/4294967296.0,1,-nbitq), 
to_sfixed(-232711497.0/4294967296.0,1,-nbitq), 
to_sfixed(320198363.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(151221443.0/4294967296.0,1,-nbitq), 
to_sfixed(536864465.0/4294967296.0,1,-nbitq), 
to_sfixed(-334948663.0/4294967296.0,1,-nbitq), 
to_sfixed(39730513.0/4294967296.0,1,-nbitq), 
to_sfixed(-127466420.0/4294967296.0,1,-nbitq), 
to_sfixed(-108719013.0/4294967296.0,1,-nbitq), 
to_sfixed(-454865283.0/4294967296.0,1,-nbitq), 
to_sfixed(359626036.0/4294967296.0,1,-nbitq), 
to_sfixed(-826520744.0/4294967296.0,1,-nbitq), 
to_sfixed(-178838497.0/4294967296.0,1,-nbitq), 
to_sfixed(508488189.0/4294967296.0,1,-nbitq), 
to_sfixed(614952803.0/4294967296.0,1,-nbitq), 
to_sfixed(428823835.0/4294967296.0,1,-nbitq), 
to_sfixed(-1014719004.0/4294967296.0,1,-nbitq), 
to_sfixed(207998703.0/4294967296.0,1,-nbitq), 
to_sfixed(-297375906.0/4294967296.0,1,-nbitq), 
to_sfixed(-50339946.0/4294967296.0,1,-nbitq), 
to_sfixed(76131375.0/4294967296.0,1,-nbitq), 
to_sfixed(573775987.0/4294967296.0,1,-nbitq), 
to_sfixed(-73360158.0/4294967296.0,1,-nbitq), 
to_sfixed(208616518.0/4294967296.0,1,-nbitq), 
to_sfixed(145678036.0/4294967296.0,1,-nbitq), 
to_sfixed(-453817511.0/4294967296.0,1,-nbitq), 
to_sfixed(-770025093.0/4294967296.0,1,-nbitq), 
to_sfixed(-74207957.0/4294967296.0,1,-nbitq), 
to_sfixed(943520621.0/4294967296.0,1,-nbitq), 
to_sfixed(-243333637.0/4294967296.0,1,-nbitq), 
to_sfixed(497539851.0/4294967296.0,1,-nbitq), 
to_sfixed(61484366.0/4294967296.0,1,-nbitq), 
to_sfixed(170375445.0/4294967296.0,1,-nbitq), 
to_sfixed(347644612.0/4294967296.0,1,-nbitq), 
to_sfixed(64650045.0/4294967296.0,1,-nbitq), 
to_sfixed(235926932.0/4294967296.0,1,-nbitq), 
to_sfixed(-245123593.0/4294967296.0,1,-nbitq), 
to_sfixed(144185957.0/4294967296.0,1,-nbitq), 
to_sfixed(50482729.0/4294967296.0,1,-nbitq), 
to_sfixed(-515243523.0/4294967296.0,1,-nbitq), 
to_sfixed(-390326641.0/4294967296.0,1,-nbitq), 
to_sfixed(261612879.0/4294967296.0,1,-nbitq), 
to_sfixed(-77347636.0/4294967296.0,1,-nbitq), 
to_sfixed(278444872.0/4294967296.0,1,-nbitq), 
to_sfixed(-19244971.0/4294967296.0,1,-nbitq), 
to_sfixed(74638707.0/4294967296.0,1,-nbitq), 
to_sfixed(-298771352.0/4294967296.0,1,-nbitq), 
to_sfixed(84541791.0/4294967296.0,1,-nbitq), 
to_sfixed(-560204021.0/4294967296.0,1,-nbitq), 
to_sfixed(-209321694.0/4294967296.0,1,-nbitq), 
to_sfixed(109248016.0/4294967296.0,1,-nbitq), 
to_sfixed(-323669753.0/4294967296.0,1,-nbitq), 
to_sfixed(304698567.0/4294967296.0,1,-nbitq), 
to_sfixed(23876327.0/4294967296.0,1,-nbitq), 
to_sfixed(-69449879.0/4294967296.0,1,-nbitq), 
to_sfixed(-343200944.0/4294967296.0,1,-nbitq), 
to_sfixed(595494687.0/4294967296.0,1,-nbitq), 
to_sfixed(81299679.0/4294967296.0,1,-nbitq), 
to_sfixed(-282955456.0/4294967296.0,1,-nbitq), 
to_sfixed(-393219301.0/4294967296.0,1,-nbitq), 
to_sfixed(-65532918.0/4294967296.0,1,-nbitq), 
to_sfixed(-166105541.0/4294967296.0,1,-nbitq), 
to_sfixed(416120496.0/4294967296.0,1,-nbitq), 
to_sfixed(-94692911.0/4294967296.0,1,-nbitq), 
to_sfixed(-688322293.0/4294967296.0,1,-nbitq), 
to_sfixed(131680186.0/4294967296.0,1,-nbitq), 
to_sfixed(-82831269.0/4294967296.0,1,-nbitq), 
to_sfixed(97687843.0/4294967296.0,1,-nbitq), 
to_sfixed(368919422.0/4294967296.0,1,-nbitq), 
to_sfixed(-438224655.0/4294967296.0,1,-nbitq), 
to_sfixed(-489035253.0/4294967296.0,1,-nbitq), 
to_sfixed(379827575.0/4294967296.0,1,-nbitq), 
to_sfixed(243738542.0/4294967296.0,1,-nbitq), 
to_sfixed(427723949.0/4294967296.0,1,-nbitq), 
to_sfixed(-112221095.0/4294967296.0,1,-nbitq), 
to_sfixed(318858800.0/4294967296.0,1,-nbitq), 
to_sfixed(197981685.0/4294967296.0,1,-nbitq), 
to_sfixed(322745422.0/4294967296.0,1,-nbitq), 
to_sfixed(100700048.0/4294967296.0,1,-nbitq), 
to_sfixed(-677302321.0/4294967296.0,1,-nbitq), 
to_sfixed(209379365.0/4294967296.0,1,-nbitq), 
to_sfixed(-629480638.0/4294967296.0,1,-nbitq), 
to_sfixed(-280079394.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-305558744.0/4294967296.0,1,-nbitq), 
to_sfixed(272221561.0/4294967296.0,1,-nbitq), 
to_sfixed(-320867032.0/4294967296.0,1,-nbitq), 
to_sfixed(123544945.0/4294967296.0,1,-nbitq), 
to_sfixed(-178724234.0/4294967296.0,1,-nbitq), 
to_sfixed(-473462552.0/4294967296.0,1,-nbitq), 
to_sfixed(50202920.0/4294967296.0,1,-nbitq), 
to_sfixed(67375518.0/4294967296.0,1,-nbitq), 
to_sfixed(18824800.0/4294967296.0,1,-nbitq), 
to_sfixed(-334532863.0/4294967296.0,1,-nbitq), 
to_sfixed(299821318.0/4294967296.0,1,-nbitq), 
to_sfixed(233097713.0/4294967296.0,1,-nbitq), 
to_sfixed(705558285.0/4294967296.0,1,-nbitq), 
to_sfixed(-209966859.0/4294967296.0,1,-nbitq), 
to_sfixed(313944836.0/4294967296.0,1,-nbitq), 
to_sfixed(-368043764.0/4294967296.0,1,-nbitq), 
to_sfixed(21630021.0/4294967296.0,1,-nbitq), 
to_sfixed(-96751892.0/4294967296.0,1,-nbitq), 
to_sfixed(427005439.0/4294967296.0,1,-nbitq), 
to_sfixed(241147325.0/4294967296.0,1,-nbitq), 
to_sfixed(351790969.0/4294967296.0,1,-nbitq), 
to_sfixed(-321519529.0/4294967296.0,1,-nbitq), 
to_sfixed(-73438099.0/4294967296.0,1,-nbitq), 
to_sfixed(-206407735.0/4294967296.0,1,-nbitq), 
to_sfixed(188389979.0/4294967296.0,1,-nbitq), 
to_sfixed(378242584.0/4294967296.0,1,-nbitq), 
to_sfixed(-471389461.0/4294967296.0,1,-nbitq), 
to_sfixed(-145748020.0/4294967296.0,1,-nbitq), 
to_sfixed(607665695.0/4294967296.0,1,-nbitq), 
to_sfixed(-37343484.0/4294967296.0,1,-nbitq), 
to_sfixed(32121595.0/4294967296.0,1,-nbitq), 
to_sfixed(3564185.0/4294967296.0,1,-nbitq), 
to_sfixed(503068016.0/4294967296.0,1,-nbitq), 
to_sfixed(-249774693.0/4294967296.0,1,-nbitq), 
to_sfixed(-198710720.0/4294967296.0,1,-nbitq), 
to_sfixed(-78350137.0/4294967296.0,1,-nbitq), 
to_sfixed(187880957.0/4294967296.0,1,-nbitq), 
to_sfixed(-750956211.0/4294967296.0,1,-nbitq), 
to_sfixed(-372883261.0/4294967296.0,1,-nbitq), 
to_sfixed(412252637.0/4294967296.0,1,-nbitq), 
to_sfixed(803275714.0/4294967296.0,1,-nbitq), 
to_sfixed(-121083639.0/4294967296.0,1,-nbitq), 
to_sfixed(-589896442.0/4294967296.0,1,-nbitq), 
to_sfixed(202038942.0/4294967296.0,1,-nbitq), 
to_sfixed(-69702225.0/4294967296.0,1,-nbitq), 
to_sfixed(276973896.0/4294967296.0,1,-nbitq), 
to_sfixed(225905517.0/4294967296.0,1,-nbitq), 
to_sfixed(-108096368.0/4294967296.0,1,-nbitq), 
to_sfixed(-13870871.0/4294967296.0,1,-nbitq), 
to_sfixed(-90688222.0/4294967296.0,1,-nbitq), 
to_sfixed(-312453058.0/4294967296.0,1,-nbitq), 
to_sfixed(-389341578.0/4294967296.0,1,-nbitq), 
to_sfixed(-198741397.0/4294967296.0,1,-nbitq), 
to_sfixed(-92698981.0/4294967296.0,1,-nbitq), 
to_sfixed(287234995.0/4294967296.0,1,-nbitq), 
to_sfixed(321404924.0/4294967296.0,1,-nbitq), 
to_sfixed(10012323.0/4294967296.0,1,-nbitq), 
to_sfixed(-318806485.0/4294967296.0,1,-nbitq), 
to_sfixed(212061685.0/4294967296.0,1,-nbitq), 
to_sfixed(-224424240.0/4294967296.0,1,-nbitq), 
to_sfixed(-513696810.0/4294967296.0,1,-nbitq), 
to_sfixed(83771672.0/4294967296.0,1,-nbitq), 
to_sfixed(143062606.0/4294967296.0,1,-nbitq), 
to_sfixed(-544527279.0/4294967296.0,1,-nbitq), 
to_sfixed(-232951354.0/4294967296.0,1,-nbitq), 
to_sfixed(-316913496.0/4294967296.0,1,-nbitq), 
to_sfixed(470909235.0/4294967296.0,1,-nbitq), 
to_sfixed(-496446665.0/4294967296.0,1,-nbitq), 
to_sfixed(111747731.0/4294967296.0,1,-nbitq), 
to_sfixed(303562858.0/4294967296.0,1,-nbitq), 
to_sfixed(-214396252.0/4294967296.0,1,-nbitq), 
to_sfixed(-170227063.0/4294967296.0,1,-nbitq), 
to_sfixed(-78328242.0/4294967296.0,1,-nbitq), 
to_sfixed(78469589.0/4294967296.0,1,-nbitq), 
to_sfixed(348791918.0/4294967296.0,1,-nbitq), 
to_sfixed(-150482007.0/4294967296.0,1,-nbitq), 
to_sfixed(-247010350.0/4294967296.0,1,-nbitq), 
to_sfixed(17054003.0/4294967296.0,1,-nbitq), 
to_sfixed(-36412573.0/4294967296.0,1,-nbitq), 
to_sfixed(-372520535.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-389366180.0/4294967296.0,1,-nbitq), 
to_sfixed(-34629768.0/4294967296.0,1,-nbitq), 
to_sfixed(-61449122.0/4294967296.0,1,-nbitq), 
to_sfixed(107376433.0/4294967296.0,1,-nbitq), 
to_sfixed(384618997.0/4294967296.0,1,-nbitq), 
to_sfixed(175069501.0/4294967296.0,1,-nbitq), 
to_sfixed(322374101.0/4294967296.0,1,-nbitq), 
to_sfixed(-141512840.0/4294967296.0,1,-nbitq), 
to_sfixed(334916409.0/4294967296.0,1,-nbitq), 
to_sfixed(166936081.0/4294967296.0,1,-nbitq), 
to_sfixed(458155425.0/4294967296.0,1,-nbitq), 
to_sfixed(152419111.0/4294967296.0,1,-nbitq), 
to_sfixed(101353744.0/4294967296.0,1,-nbitq), 
to_sfixed(-335573323.0/4294967296.0,1,-nbitq), 
to_sfixed(23292418.0/4294967296.0,1,-nbitq), 
to_sfixed(-362045458.0/4294967296.0,1,-nbitq), 
to_sfixed(-222370185.0/4294967296.0,1,-nbitq), 
to_sfixed(8641085.0/4294967296.0,1,-nbitq), 
to_sfixed(275103978.0/4294967296.0,1,-nbitq), 
to_sfixed(227307306.0/4294967296.0,1,-nbitq), 
to_sfixed(-276933589.0/4294967296.0,1,-nbitq), 
to_sfixed(62595979.0/4294967296.0,1,-nbitq), 
to_sfixed(252003425.0/4294967296.0,1,-nbitq), 
to_sfixed(306702852.0/4294967296.0,1,-nbitq), 
to_sfixed(280352595.0/4294967296.0,1,-nbitq), 
to_sfixed(-185475244.0/4294967296.0,1,-nbitq), 
to_sfixed(260968376.0/4294967296.0,1,-nbitq), 
to_sfixed(-709585700.0/4294967296.0,1,-nbitq), 
to_sfixed(174950328.0/4294967296.0,1,-nbitq), 
to_sfixed(-564634709.0/4294967296.0,1,-nbitq), 
to_sfixed(-111366044.0/4294967296.0,1,-nbitq), 
to_sfixed(-331414205.0/4294967296.0,1,-nbitq), 
to_sfixed(202365388.0/4294967296.0,1,-nbitq), 
to_sfixed(-119696003.0/4294967296.0,1,-nbitq), 
to_sfixed(36103415.0/4294967296.0,1,-nbitq), 
to_sfixed(-449531796.0/4294967296.0,1,-nbitq), 
to_sfixed(-172242371.0/4294967296.0,1,-nbitq), 
to_sfixed(88664153.0/4294967296.0,1,-nbitq), 
to_sfixed(-332856274.0/4294967296.0,1,-nbitq), 
to_sfixed(436538685.0/4294967296.0,1,-nbitq), 
to_sfixed(-135571679.0/4294967296.0,1,-nbitq), 
to_sfixed(143186100.0/4294967296.0,1,-nbitq), 
to_sfixed(-143331051.0/4294967296.0,1,-nbitq), 
to_sfixed(34332639.0/4294967296.0,1,-nbitq), 
to_sfixed(3761108.0/4294967296.0,1,-nbitq), 
to_sfixed(424706631.0/4294967296.0,1,-nbitq), 
to_sfixed(-330799823.0/4294967296.0,1,-nbitq), 
to_sfixed(-335928532.0/4294967296.0,1,-nbitq), 
to_sfixed(-40180236.0/4294967296.0,1,-nbitq), 
to_sfixed(-1952141.0/4294967296.0,1,-nbitq), 
to_sfixed(-178758058.0/4294967296.0,1,-nbitq), 
to_sfixed(379538539.0/4294967296.0,1,-nbitq), 
to_sfixed(-60964474.0/4294967296.0,1,-nbitq), 
to_sfixed(5994747.0/4294967296.0,1,-nbitq), 
to_sfixed(11428515.0/4294967296.0,1,-nbitq), 
to_sfixed(-1657988.0/4294967296.0,1,-nbitq), 
to_sfixed(286419687.0/4294967296.0,1,-nbitq), 
to_sfixed(-253338178.0/4294967296.0,1,-nbitq), 
to_sfixed(242056493.0/4294967296.0,1,-nbitq), 
to_sfixed(162792282.0/4294967296.0,1,-nbitq), 
to_sfixed(-119572586.0/4294967296.0,1,-nbitq), 
to_sfixed(-33521846.0/4294967296.0,1,-nbitq), 
to_sfixed(-83576695.0/4294967296.0,1,-nbitq), 
to_sfixed(-339317128.0/4294967296.0,1,-nbitq), 
to_sfixed(-263465428.0/4294967296.0,1,-nbitq), 
to_sfixed(116513510.0/4294967296.0,1,-nbitq), 
to_sfixed(325939949.0/4294967296.0,1,-nbitq), 
to_sfixed(-74096919.0/4294967296.0,1,-nbitq), 
to_sfixed(-66297766.0/4294967296.0,1,-nbitq), 
to_sfixed(242024361.0/4294967296.0,1,-nbitq), 
to_sfixed(-150330852.0/4294967296.0,1,-nbitq), 
to_sfixed(38451456.0/4294967296.0,1,-nbitq), 
to_sfixed(-422148423.0/4294967296.0,1,-nbitq), 
to_sfixed(81691889.0/4294967296.0,1,-nbitq), 
to_sfixed(-11575589.0/4294967296.0,1,-nbitq), 
to_sfixed(118507773.0/4294967296.0,1,-nbitq), 
to_sfixed(-280873197.0/4294967296.0,1,-nbitq), 
to_sfixed(-232045997.0/4294967296.0,1,-nbitq), 
to_sfixed(-352405952.0/4294967296.0,1,-nbitq), 
to_sfixed(128513462.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-21476653.0/4294967296.0,1,-nbitq), 
to_sfixed(-226762770.0/4294967296.0,1,-nbitq), 
to_sfixed(-404216913.0/4294967296.0,1,-nbitq), 
to_sfixed(231822459.0/4294967296.0,1,-nbitq), 
to_sfixed(-145562080.0/4294967296.0,1,-nbitq), 
to_sfixed(224089476.0/4294967296.0,1,-nbitq), 
to_sfixed(-299829946.0/4294967296.0,1,-nbitq), 
to_sfixed(-245319836.0/4294967296.0,1,-nbitq), 
to_sfixed(-72712168.0/4294967296.0,1,-nbitq), 
to_sfixed(-188274563.0/4294967296.0,1,-nbitq), 
to_sfixed(119497319.0/4294967296.0,1,-nbitq), 
to_sfixed(-82373828.0/4294967296.0,1,-nbitq), 
to_sfixed(63459343.0/4294967296.0,1,-nbitq), 
to_sfixed(-58739511.0/4294967296.0,1,-nbitq), 
to_sfixed(-332249660.0/4294967296.0,1,-nbitq), 
to_sfixed(194601017.0/4294967296.0,1,-nbitq), 
to_sfixed(-283468706.0/4294967296.0,1,-nbitq), 
to_sfixed(132228105.0/4294967296.0,1,-nbitq), 
to_sfixed(-272291727.0/4294967296.0,1,-nbitq), 
to_sfixed(-393848932.0/4294967296.0,1,-nbitq), 
to_sfixed(99891899.0/4294967296.0,1,-nbitq), 
to_sfixed(332578702.0/4294967296.0,1,-nbitq), 
to_sfixed(299206268.0/4294967296.0,1,-nbitq), 
to_sfixed(-324205706.0/4294967296.0,1,-nbitq), 
to_sfixed(342699092.0/4294967296.0,1,-nbitq), 
to_sfixed(80410036.0/4294967296.0,1,-nbitq), 
to_sfixed(104306341.0/4294967296.0,1,-nbitq), 
to_sfixed(-657964691.0/4294967296.0,1,-nbitq), 
to_sfixed(56699556.0/4294967296.0,1,-nbitq), 
to_sfixed(-49444598.0/4294967296.0,1,-nbitq), 
to_sfixed(154309407.0/4294967296.0,1,-nbitq), 
to_sfixed(175586563.0/4294967296.0,1,-nbitq), 
to_sfixed(301136037.0/4294967296.0,1,-nbitq), 
to_sfixed(-144441943.0/4294967296.0,1,-nbitq), 
to_sfixed(159162604.0/4294967296.0,1,-nbitq), 
to_sfixed(-272350524.0/4294967296.0,1,-nbitq), 
to_sfixed(-117114590.0/4294967296.0,1,-nbitq), 
to_sfixed(-247649524.0/4294967296.0,1,-nbitq), 
to_sfixed(358151333.0/4294967296.0,1,-nbitq), 
to_sfixed(317333096.0/4294967296.0,1,-nbitq), 
to_sfixed(362632882.0/4294967296.0,1,-nbitq), 
to_sfixed(345078275.0/4294967296.0,1,-nbitq), 
to_sfixed(-381410927.0/4294967296.0,1,-nbitq), 
to_sfixed(59564985.0/4294967296.0,1,-nbitq), 
to_sfixed(-112633009.0/4294967296.0,1,-nbitq), 
to_sfixed(-147513594.0/4294967296.0,1,-nbitq), 
to_sfixed(-48569797.0/4294967296.0,1,-nbitq), 
to_sfixed(-343192452.0/4294967296.0,1,-nbitq), 
to_sfixed(-367436988.0/4294967296.0,1,-nbitq), 
to_sfixed(-195188483.0/4294967296.0,1,-nbitq), 
to_sfixed(-136992918.0/4294967296.0,1,-nbitq), 
to_sfixed(67484883.0/4294967296.0,1,-nbitq), 
to_sfixed(-28889342.0/4294967296.0,1,-nbitq), 
to_sfixed(34901889.0/4294967296.0,1,-nbitq), 
to_sfixed(219443447.0/4294967296.0,1,-nbitq), 
to_sfixed(-263587245.0/4294967296.0,1,-nbitq), 
to_sfixed(-160743948.0/4294967296.0,1,-nbitq), 
to_sfixed(-68201327.0/4294967296.0,1,-nbitq), 
to_sfixed(-227090813.0/4294967296.0,1,-nbitq), 
to_sfixed(-48431673.0/4294967296.0,1,-nbitq), 
to_sfixed(-84993207.0/4294967296.0,1,-nbitq), 
to_sfixed(-119489736.0/4294967296.0,1,-nbitq), 
to_sfixed(-419787129.0/4294967296.0,1,-nbitq), 
to_sfixed(36310922.0/4294967296.0,1,-nbitq), 
to_sfixed(419082827.0/4294967296.0,1,-nbitq), 
to_sfixed(-96912011.0/4294967296.0,1,-nbitq), 
to_sfixed(752988237.0/4294967296.0,1,-nbitq), 
to_sfixed(-368529179.0/4294967296.0,1,-nbitq), 
to_sfixed(-3797548.0/4294967296.0,1,-nbitq), 
to_sfixed(130806478.0/4294967296.0,1,-nbitq), 
to_sfixed(301414763.0/4294967296.0,1,-nbitq), 
to_sfixed(267819582.0/4294967296.0,1,-nbitq), 
to_sfixed(-289601094.0/4294967296.0,1,-nbitq), 
to_sfixed(5709033.0/4294967296.0,1,-nbitq), 
to_sfixed(-121873900.0/4294967296.0,1,-nbitq), 
to_sfixed(168737980.0/4294967296.0,1,-nbitq), 
to_sfixed(-111422668.0/4294967296.0,1,-nbitq), 
to_sfixed(266593057.0/4294967296.0,1,-nbitq), 
to_sfixed(-357820052.0/4294967296.0,1,-nbitq), 
to_sfixed(145269620.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-113034337.0/4294967296.0,1,-nbitq), 
to_sfixed(144060042.0/4294967296.0,1,-nbitq), 
to_sfixed(17508759.0/4294967296.0,1,-nbitq), 
to_sfixed(-393340941.0/4294967296.0,1,-nbitq), 
to_sfixed(459197941.0/4294967296.0,1,-nbitq), 
to_sfixed(-38921396.0/4294967296.0,1,-nbitq), 
to_sfixed(33162373.0/4294967296.0,1,-nbitq), 
to_sfixed(304112422.0/4294967296.0,1,-nbitq), 
to_sfixed(268884769.0/4294967296.0,1,-nbitq), 
to_sfixed(-202368453.0/4294967296.0,1,-nbitq), 
to_sfixed(337984291.0/4294967296.0,1,-nbitq), 
to_sfixed(113697179.0/4294967296.0,1,-nbitq), 
to_sfixed(398150406.0/4294967296.0,1,-nbitq), 
to_sfixed(454933910.0/4294967296.0,1,-nbitq), 
to_sfixed(-905090.0/4294967296.0,1,-nbitq), 
to_sfixed(-267868873.0/4294967296.0,1,-nbitq), 
to_sfixed(-166224320.0/4294967296.0,1,-nbitq), 
to_sfixed(-274345121.0/4294967296.0,1,-nbitq), 
to_sfixed(-40567062.0/4294967296.0,1,-nbitq), 
to_sfixed(-302788921.0/4294967296.0,1,-nbitq), 
to_sfixed(-109919584.0/4294967296.0,1,-nbitq), 
to_sfixed(435461195.0/4294967296.0,1,-nbitq), 
to_sfixed(541806732.0/4294967296.0,1,-nbitq), 
to_sfixed(-89544543.0/4294967296.0,1,-nbitq), 
to_sfixed(-208312767.0/4294967296.0,1,-nbitq), 
to_sfixed(251592502.0/4294967296.0,1,-nbitq), 
to_sfixed(-213054318.0/4294967296.0,1,-nbitq), 
to_sfixed(-1973743.0/4294967296.0,1,-nbitq), 
to_sfixed(259359441.0/4294967296.0,1,-nbitq), 
to_sfixed(-23912100.0/4294967296.0,1,-nbitq), 
to_sfixed(-208245379.0/4294967296.0,1,-nbitq), 
to_sfixed(-329102230.0/4294967296.0,1,-nbitq), 
to_sfixed(154802012.0/4294967296.0,1,-nbitq), 
to_sfixed(-196769550.0/4294967296.0,1,-nbitq), 
to_sfixed(398446063.0/4294967296.0,1,-nbitq), 
to_sfixed(-362134662.0/4294967296.0,1,-nbitq), 
to_sfixed(268726058.0/4294967296.0,1,-nbitq), 
to_sfixed(-283238257.0/4294967296.0,1,-nbitq), 
to_sfixed(118349980.0/4294967296.0,1,-nbitq), 
to_sfixed(376208831.0/4294967296.0,1,-nbitq), 
to_sfixed(188180073.0/4294967296.0,1,-nbitq), 
to_sfixed(26179295.0/4294967296.0,1,-nbitq), 
to_sfixed(-312509089.0/4294967296.0,1,-nbitq), 
to_sfixed(268419145.0/4294967296.0,1,-nbitq), 
to_sfixed(-334470189.0/4294967296.0,1,-nbitq), 
to_sfixed(25153217.0/4294967296.0,1,-nbitq), 
to_sfixed(-50221509.0/4294967296.0,1,-nbitq), 
to_sfixed(-11709022.0/4294967296.0,1,-nbitq), 
to_sfixed(-48115422.0/4294967296.0,1,-nbitq), 
to_sfixed(527576335.0/4294967296.0,1,-nbitq), 
to_sfixed(143007373.0/4294967296.0,1,-nbitq), 
to_sfixed(-291331034.0/4294967296.0,1,-nbitq), 
to_sfixed(-473546560.0/4294967296.0,1,-nbitq), 
to_sfixed(-139889475.0/4294967296.0,1,-nbitq), 
to_sfixed(149391860.0/4294967296.0,1,-nbitq), 
to_sfixed(116950160.0/4294967296.0,1,-nbitq), 
to_sfixed(405044289.0/4294967296.0,1,-nbitq), 
to_sfixed(100870048.0/4294967296.0,1,-nbitq), 
to_sfixed(-293769384.0/4294967296.0,1,-nbitq), 
to_sfixed(227172039.0/4294967296.0,1,-nbitq), 
to_sfixed(-360161491.0/4294967296.0,1,-nbitq), 
to_sfixed(29136629.0/4294967296.0,1,-nbitq), 
to_sfixed(-242963253.0/4294967296.0,1,-nbitq), 
to_sfixed(418942102.0/4294967296.0,1,-nbitq), 
to_sfixed(438610159.0/4294967296.0,1,-nbitq), 
to_sfixed(-380294003.0/4294967296.0,1,-nbitq), 
to_sfixed(551927518.0/4294967296.0,1,-nbitq), 
to_sfixed(38478651.0/4294967296.0,1,-nbitq), 
to_sfixed(-62992490.0/4294967296.0,1,-nbitq), 
to_sfixed(363341331.0/4294967296.0,1,-nbitq), 
to_sfixed(-41342655.0/4294967296.0,1,-nbitq), 
to_sfixed(-86687700.0/4294967296.0,1,-nbitq), 
to_sfixed(129610430.0/4294967296.0,1,-nbitq), 
to_sfixed(265188108.0/4294967296.0,1,-nbitq), 
to_sfixed(53068916.0/4294967296.0,1,-nbitq), 
to_sfixed(-135138550.0/4294967296.0,1,-nbitq), 
to_sfixed(-142215106.0/4294967296.0,1,-nbitq), 
to_sfixed(-416128205.0/4294967296.0,1,-nbitq), 
to_sfixed(-420500890.0/4294967296.0,1,-nbitq), 
to_sfixed(70020323.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(136394696.0/4294967296.0,1,-nbitq), 
to_sfixed(118992655.0/4294967296.0,1,-nbitq), 
to_sfixed(-352523471.0/4294967296.0,1,-nbitq), 
to_sfixed(-234002478.0/4294967296.0,1,-nbitq), 
to_sfixed(294892202.0/4294967296.0,1,-nbitq), 
to_sfixed(168979366.0/4294967296.0,1,-nbitq), 
to_sfixed(-133741239.0/4294967296.0,1,-nbitq), 
to_sfixed(-24491711.0/4294967296.0,1,-nbitq), 
to_sfixed(-150826406.0/4294967296.0,1,-nbitq), 
to_sfixed(16117759.0/4294967296.0,1,-nbitq), 
to_sfixed(-394938890.0/4294967296.0,1,-nbitq), 
to_sfixed(397303447.0/4294967296.0,1,-nbitq), 
to_sfixed(-183675571.0/4294967296.0,1,-nbitq), 
to_sfixed(159502063.0/4294967296.0,1,-nbitq), 
to_sfixed(-256891139.0/4294967296.0,1,-nbitq), 
to_sfixed(-366144698.0/4294967296.0,1,-nbitq), 
to_sfixed(-410499650.0/4294967296.0,1,-nbitq), 
to_sfixed(-170163042.0/4294967296.0,1,-nbitq), 
to_sfixed(41932392.0/4294967296.0,1,-nbitq), 
to_sfixed(-47288108.0/4294967296.0,1,-nbitq), 
to_sfixed(43840384.0/4294967296.0,1,-nbitq), 
to_sfixed(40244314.0/4294967296.0,1,-nbitq), 
to_sfixed(51701813.0/4294967296.0,1,-nbitq), 
to_sfixed(155787040.0/4294967296.0,1,-nbitq), 
to_sfixed(168327299.0/4294967296.0,1,-nbitq), 
to_sfixed(-190494521.0/4294967296.0,1,-nbitq), 
to_sfixed(-32655759.0/4294967296.0,1,-nbitq), 
to_sfixed(58382626.0/4294967296.0,1,-nbitq), 
to_sfixed(433064305.0/4294967296.0,1,-nbitq), 
to_sfixed(-186671798.0/4294967296.0,1,-nbitq), 
to_sfixed(-155267661.0/4294967296.0,1,-nbitq), 
to_sfixed(-451967882.0/4294967296.0,1,-nbitq), 
to_sfixed(110397549.0/4294967296.0,1,-nbitq), 
to_sfixed(227107224.0/4294967296.0,1,-nbitq), 
to_sfixed(411236881.0/4294967296.0,1,-nbitq), 
to_sfixed(336750383.0/4294967296.0,1,-nbitq), 
to_sfixed(406647265.0/4294967296.0,1,-nbitq), 
to_sfixed(-89944839.0/4294967296.0,1,-nbitq), 
to_sfixed(-284707798.0/4294967296.0,1,-nbitq), 
to_sfixed(233652817.0/4294967296.0,1,-nbitq), 
to_sfixed(-387042400.0/4294967296.0,1,-nbitq), 
to_sfixed(-15676422.0/4294967296.0,1,-nbitq), 
to_sfixed(272550354.0/4294967296.0,1,-nbitq), 
to_sfixed(302019981.0/4294967296.0,1,-nbitq), 
to_sfixed(-324608933.0/4294967296.0,1,-nbitq), 
to_sfixed(298967993.0/4294967296.0,1,-nbitq), 
to_sfixed(267397566.0/4294967296.0,1,-nbitq), 
to_sfixed(72106730.0/4294967296.0,1,-nbitq), 
to_sfixed(95273110.0/4294967296.0,1,-nbitq), 
to_sfixed(228099577.0/4294967296.0,1,-nbitq), 
to_sfixed(137460900.0/4294967296.0,1,-nbitq), 
to_sfixed(277683155.0/4294967296.0,1,-nbitq), 
to_sfixed(95120325.0/4294967296.0,1,-nbitq), 
to_sfixed(-112028936.0/4294967296.0,1,-nbitq), 
to_sfixed(252527330.0/4294967296.0,1,-nbitq), 
to_sfixed(-351791381.0/4294967296.0,1,-nbitq), 
to_sfixed(358612368.0/4294967296.0,1,-nbitq), 
to_sfixed(174086149.0/4294967296.0,1,-nbitq), 
to_sfixed(194307635.0/4294967296.0,1,-nbitq), 
to_sfixed(345899018.0/4294967296.0,1,-nbitq), 
to_sfixed(-189114859.0/4294967296.0,1,-nbitq), 
to_sfixed(511290597.0/4294967296.0,1,-nbitq), 
to_sfixed(-289815315.0/4294967296.0,1,-nbitq), 
to_sfixed(107507874.0/4294967296.0,1,-nbitq), 
to_sfixed(-358243813.0/4294967296.0,1,-nbitq), 
to_sfixed(-308592721.0/4294967296.0,1,-nbitq), 
to_sfixed(249140480.0/4294967296.0,1,-nbitq), 
to_sfixed(72935265.0/4294967296.0,1,-nbitq), 
to_sfixed(-310799242.0/4294967296.0,1,-nbitq), 
to_sfixed(276015459.0/4294967296.0,1,-nbitq), 
to_sfixed(-42298488.0/4294967296.0,1,-nbitq), 
to_sfixed(-48279221.0/4294967296.0,1,-nbitq), 
to_sfixed(-62482215.0/4294967296.0,1,-nbitq), 
to_sfixed(267221882.0/4294967296.0,1,-nbitq), 
to_sfixed(130291514.0/4294967296.0,1,-nbitq), 
to_sfixed(-343945237.0/4294967296.0,1,-nbitq), 
to_sfixed(-447155282.0/4294967296.0,1,-nbitq), 
to_sfixed(272099564.0/4294967296.0,1,-nbitq), 
to_sfixed(-38845046.0/4294967296.0,1,-nbitq), 
to_sfixed(-72965714.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(109872369.0/4294967296.0,1,-nbitq), 
to_sfixed(-126949223.0/4294967296.0,1,-nbitq), 
to_sfixed(114452087.0/4294967296.0,1,-nbitq), 
to_sfixed(-367628809.0/4294967296.0,1,-nbitq), 
to_sfixed(-24669832.0/4294967296.0,1,-nbitq), 
to_sfixed(218829006.0/4294967296.0,1,-nbitq), 
to_sfixed(41257301.0/4294967296.0,1,-nbitq), 
to_sfixed(-310728328.0/4294967296.0,1,-nbitq), 
to_sfixed(-466879615.0/4294967296.0,1,-nbitq), 
to_sfixed(10270914.0/4294967296.0,1,-nbitq), 
to_sfixed(-68557308.0/4294967296.0,1,-nbitq), 
to_sfixed(-150221496.0/4294967296.0,1,-nbitq), 
to_sfixed(423921043.0/4294967296.0,1,-nbitq), 
to_sfixed(720594739.0/4294967296.0,1,-nbitq), 
to_sfixed(-377345907.0/4294967296.0,1,-nbitq), 
to_sfixed(-188349251.0/4294967296.0,1,-nbitq), 
to_sfixed(30675244.0/4294967296.0,1,-nbitq), 
to_sfixed(337539337.0/4294967296.0,1,-nbitq), 
to_sfixed(500846182.0/4294967296.0,1,-nbitq), 
to_sfixed(-181784885.0/4294967296.0,1,-nbitq), 
to_sfixed(46263260.0/4294967296.0,1,-nbitq), 
to_sfixed(26325752.0/4294967296.0,1,-nbitq), 
to_sfixed(-38817153.0/4294967296.0,1,-nbitq), 
to_sfixed(150241821.0/4294967296.0,1,-nbitq), 
to_sfixed(-64816952.0/4294967296.0,1,-nbitq), 
to_sfixed(-70628162.0/4294967296.0,1,-nbitq), 
to_sfixed(521772.0/4294967296.0,1,-nbitq), 
to_sfixed(19040665.0/4294967296.0,1,-nbitq), 
to_sfixed(80392636.0/4294967296.0,1,-nbitq), 
to_sfixed(408483078.0/4294967296.0,1,-nbitq), 
to_sfixed(-138513287.0/4294967296.0,1,-nbitq), 
to_sfixed(-97043760.0/4294967296.0,1,-nbitq), 
to_sfixed(-156861774.0/4294967296.0,1,-nbitq), 
to_sfixed(-627247435.0/4294967296.0,1,-nbitq), 
to_sfixed(292262609.0/4294967296.0,1,-nbitq), 
to_sfixed(212291722.0/4294967296.0,1,-nbitq), 
to_sfixed(-114358374.0/4294967296.0,1,-nbitq), 
to_sfixed(135588672.0/4294967296.0,1,-nbitq), 
to_sfixed(-177987581.0/4294967296.0,1,-nbitq), 
to_sfixed(65865490.0/4294967296.0,1,-nbitq), 
to_sfixed(-439518896.0/4294967296.0,1,-nbitq), 
to_sfixed(-326021077.0/4294967296.0,1,-nbitq), 
to_sfixed(168217705.0/4294967296.0,1,-nbitq), 
to_sfixed(-146090580.0/4294967296.0,1,-nbitq), 
to_sfixed(422982442.0/4294967296.0,1,-nbitq), 
to_sfixed(-918382.0/4294967296.0,1,-nbitq), 
to_sfixed(150113952.0/4294967296.0,1,-nbitq), 
to_sfixed(-327368368.0/4294967296.0,1,-nbitq), 
to_sfixed(424614615.0/4294967296.0,1,-nbitq), 
to_sfixed(-73032323.0/4294967296.0,1,-nbitq), 
to_sfixed(-22782582.0/4294967296.0,1,-nbitq), 
to_sfixed(-66625100.0/4294967296.0,1,-nbitq), 
to_sfixed(-408055534.0/4294967296.0,1,-nbitq), 
to_sfixed(-124702601.0/4294967296.0,1,-nbitq), 
to_sfixed(-1531040.0/4294967296.0,1,-nbitq), 
to_sfixed(-172424904.0/4294967296.0,1,-nbitq), 
to_sfixed(359472166.0/4294967296.0,1,-nbitq), 
to_sfixed(-409734218.0/4294967296.0,1,-nbitq), 
to_sfixed(-188849784.0/4294967296.0,1,-nbitq), 
to_sfixed(-26700189.0/4294967296.0,1,-nbitq), 
to_sfixed(-277895090.0/4294967296.0,1,-nbitq), 
to_sfixed(222270952.0/4294967296.0,1,-nbitq), 
to_sfixed(263556313.0/4294967296.0,1,-nbitq), 
to_sfixed(94129222.0/4294967296.0,1,-nbitq), 
to_sfixed(-85956259.0/4294967296.0,1,-nbitq), 
to_sfixed(-106158415.0/4294967296.0,1,-nbitq), 
to_sfixed(518773601.0/4294967296.0,1,-nbitq), 
to_sfixed(-65340887.0/4294967296.0,1,-nbitq), 
to_sfixed(50260475.0/4294967296.0,1,-nbitq), 
to_sfixed(-294451048.0/4294967296.0,1,-nbitq), 
to_sfixed(-123486724.0/4294967296.0,1,-nbitq), 
to_sfixed(-210090982.0/4294967296.0,1,-nbitq), 
to_sfixed(-117742753.0/4294967296.0,1,-nbitq), 
to_sfixed(-162492969.0/4294967296.0,1,-nbitq), 
to_sfixed(39747065.0/4294967296.0,1,-nbitq), 
to_sfixed(45472219.0/4294967296.0,1,-nbitq), 
to_sfixed(-41522315.0/4294967296.0,1,-nbitq), 
to_sfixed(-168761636.0/4294967296.0,1,-nbitq), 
to_sfixed(253359090.0/4294967296.0,1,-nbitq), 
to_sfixed(-166768922.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-218815038.0/4294967296.0,1,-nbitq), 
to_sfixed(171820610.0/4294967296.0,1,-nbitq), 
to_sfixed(-614936500.0/4294967296.0,1,-nbitq), 
to_sfixed(355151465.0/4294967296.0,1,-nbitq), 
to_sfixed(-122647888.0/4294967296.0,1,-nbitq), 
to_sfixed(26799847.0/4294967296.0,1,-nbitq), 
to_sfixed(-477417339.0/4294967296.0,1,-nbitq), 
to_sfixed(72597221.0/4294967296.0,1,-nbitq), 
to_sfixed(-339851705.0/4294967296.0,1,-nbitq), 
to_sfixed(51751484.0/4294967296.0,1,-nbitq), 
to_sfixed(-214691229.0/4294967296.0,1,-nbitq), 
to_sfixed(-395284291.0/4294967296.0,1,-nbitq), 
to_sfixed(458230558.0/4294967296.0,1,-nbitq), 
to_sfixed(149177388.0/4294967296.0,1,-nbitq), 
to_sfixed(-64072448.0/4294967296.0,1,-nbitq), 
to_sfixed(-24331829.0/4294967296.0,1,-nbitq), 
to_sfixed(283630617.0/4294967296.0,1,-nbitq), 
to_sfixed(96697691.0/4294967296.0,1,-nbitq), 
to_sfixed(609709650.0/4294967296.0,1,-nbitq), 
to_sfixed(347654056.0/4294967296.0,1,-nbitq), 
to_sfixed(-44174143.0/4294967296.0,1,-nbitq), 
to_sfixed(181727323.0/4294967296.0,1,-nbitq), 
to_sfixed(-174881328.0/4294967296.0,1,-nbitq), 
to_sfixed(510406450.0/4294967296.0,1,-nbitq), 
to_sfixed(98389676.0/4294967296.0,1,-nbitq), 
to_sfixed(616470292.0/4294967296.0,1,-nbitq), 
to_sfixed(-238201847.0/4294967296.0,1,-nbitq), 
to_sfixed(-340749370.0/4294967296.0,1,-nbitq), 
to_sfixed(322120025.0/4294967296.0,1,-nbitq), 
to_sfixed(-105009898.0/4294967296.0,1,-nbitq), 
to_sfixed(-330549115.0/4294967296.0,1,-nbitq), 
to_sfixed(-71819667.0/4294967296.0,1,-nbitq), 
to_sfixed(96528154.0/4294967296.0,1,-nbitq), 
to_sfixed(-421103874.0/4294967296.0,1,-nbitq), 
to_sfixed(113073254.0/4294967296.0,1,-nbitq), 
to_sfixed(-83606060.0/4294967296.0,1,-nbitq), 
to_sfixed(-322705866.0/4294967296.0,1,-nbitq), 
to_sfixed(199082743.0/4294967296.0,1,-nbitq), 
to_sfixed(-357569490.0/4294967296.0,1,-nbitq), 
to_sfixed(-83516034.0/4294967296.0,1,-nbitq), 
to_sfixed(-32285056.0/4294967296.0,1,-nbitq), 
to_sfixed(149548054.0/4294967296.0,1,-nbitq), 
to_sfixed(-127974125.0/4294967296.0,1,-nbitq), 
to_sfixed(484368296.0/4294967296.0,1,-nbitq), 
to_sfixed(142597368.0/4294967296.0,1,-nbitq), 
to_sfixed(506592457.0/4294967296.0,1,-nbitq), 
to_sfixed(22435271.0/4294967296.0,1,-nbitq), 
to_sfixed(-824825670.0/4294967296.0,1,-nbitq), 
to_sfixed(-9517851.0/4294967296.0,1,-nbitq), 
to_sfixed(92664507.0/4294967296.0,1,-nbitq), 
to_sfixed(307662944.0/4294967296.0,1,-nbitq), 
to_sfixed(144347548.0/4294967296.0,1,-nbitq), 
to_sfixed(200380925.0/4294967296.0,1,-nbitq), 
to_sfixed(223596115.0/4294967296.0,1,-nbitq), 
to_sfixed(434870386.0/4294967296.0,1,-nbitq), 
to_sfixed(-324241930.0/4294967296.0,1,-nbitq), 
to_sfixed(-24146953.0/4294967296.0,1,-nbitq), 
to_sfixed(-170005264.0/4294967296.0,1,-nbitq), 
to_sfixed(-131932259.0/4294967296.0,1,-nbitq), 
to_sfixed(176719670.0/4294967296.0,1,-nbitq), 
to_sfixed(328898954.0/4294967296.0,1,-nbitq), 
to_sfixed(564720165.0/4294967296.0,1,-nbitq), 
to_sfixed(-287962360.0/4294967296.0,1,-nbitq), 
to_sfixed(-169536726.0/4294967296.0,1,-nbitq), 
to_sfixed(320513024.0/4294967296.0,1,-nbitq), 
to_sfixed(-291392712.0/4294967296.0,1,-nbitq), 
to_sfixed(-191754463.0/4294967296.0,1,-nbitq), 
to_sfixed(361460347.0/4294967296.0,1,-nbitq), 
to_sfixed(264318686.0/4294967296.0,1,-nbitq), 
to_sfixed(-146624693.0/4294967296.0,1,-nbitq), 
to_sfixed(-261570709.0/4294967296.0,1,-nbitq), 
to_sfixed(5489916.0/4294967296.0,1,-nbitq), 
to_sfixed(-282175342.0/4294967296.0,1,-nbitq), 
to_sfixed(135569993.0/4294967296.0,1,-nbitq), 
to_sfixed(457789121.0/4294967296.0,1,-nbitq), 
to_sfixed(89099364.0/4294967296.0,1,-nbitq), 
to_sfixed(-378419159.0/4294967296.0,1,-nbitq), 
to_sfixed(-170985436.0/4294967296.0,1,-nbitq), 
to_sfixed(-396550896.0/4294967296.0,1,-nbitq), 
to_sfixed(-29591872.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(201162805.0/4294967296.0,1,-nbitq), 
to_sfixed(397201607.0/4294967296.0,1,-nbitq), 
to_sfixed(-325819099.0/4294967296.0,1,-nbitq), 
to_sfixed(455039966.0/4294967296.0,1,-nbitq), 
to_sfixed(475757163.0/4294967296.0,1,-nbitq), 
to_sfixed(-211035034.0/4294967296.0,1,-nbitq), 
to_sfixed(-500287981.0/4294967296.0,1,-nbitq), 
to_sfixed(-526166264.0/4294967296.0,1,-nbitq), 
to_sfixed(-946283354.0/4294967296.0,1,-nbitq), 
to_sfixed(-70684969.0/4294967296.0,1,-nbitq), 
to_sfixed(273700504.0/4294967296.0,1,-nbitq), 
to_sfixed(-632282191.0/4294967296.0,1,-nbitq), 
to_sfixed(857840769.0/4294967296.0,1,-nbitq), 
to_sfixed(906067961.0/4294967296.0,1,-nbitq), 
to_sfixed(155315932.0/4294967296.0,1,-nbitq), 
to_sfixed(-903108055.0/4294967296.0,1,-nbitq), 
to_sfixed(229021084.0/4294967296.0,1,-nbitq), 
to_sfixed(-165545927.0/4294967296.0,1,-nbitq), 
to_sfixed(166382239.0/4294967296.0,1,-nbitq), 
to_sfixed(408544910.0/4294967296.0,1,-nbitq), 
to_sfixed(64870894.0/4294967296.0,1,-nbitq), 
to_sfixed(-385701907.0/4294967296.0,1,-nbitq), 
to_sfixed(-461125722.0/4294967296.0,1,-nbitq), 
to_sfixed(328241754.0/4294967296.0,1,-nbitq), 
to_sfixed(-55674933.0/4294967296.0,1,-nbitq), 
to_sfixed(157855658.0/4294967296.0,1,-nbitq), 
to_sfixed(129499020.0/4294967296.0,1,-nbitq), 
to_sfixed(473936965.0/4294967296.0,1,-nbitq), 
to_sfixed(788403542.0/4294967296.0,1,-nbitq), 
to_sfixed(-59022532.0/4294967296.0,1,-nbitq), 
to_sfixed(50712694.0/4294967296.0,1,-nbitq), 
to_sfixed(5726761.0/4294967296.0,1,-nbitq), 
to_sfixed(-54925375.0/4294967296.0,1,-nbitq), 
to_sfixed(113258139.0/4294967296.0,1,-nbitq), 
to_sfixed(262420936.0/4294967296.0,1,-nbitq), 
to_sfixed(360096436.0/4294967296.0,1,-nbitq), 
to_sfixed(405648594.0/4294967296.0,1,-nbitq), 
to_sfixed(156399402.0/4294967296.0,1,-nbitq), 
to_sfixed(130576479.0/4294967296.0,1,-nbitq), 
to_sfixed(114101625.0/4294967296.0,1,-nbitq), 
to_sfixed(302027559.0/4294967296.0,1,-nbitq), 
to_sfixed(-376178656.0/4294967296.0,1,-nbitq), 
to_sfixed(13798512.0/4294967296.0,1,-nbitq), 
to_sfixed(398477142.0/4294967296.0,1,-nbitq), 
to_sfixed(403752516.0/4294967296.0,1,-nbitq), 
to_sfixed(-80133715.0/4294967296.0,1,-nbitq), 
to_sfixed(-101054576.0/4294967296.0,1,-nbitq), 
to_sfixed(-111939164.0/4294967296.0,1,-nbitq), 
to_sfixed(-211457995.0/4294967296.0,1,-nbitq), 
to_sfixed(-448178979.0/4294967296.0,1,-nbitq), 
to_sfixed(-95445096.0/4294967296.0,1,-nbitq), 
to_sfixed(-41801804.0/4294967296.0,1,-nbitq), 
to_sfixed(847496322.0/4294967296.0,1,-nbitq), 
to_sfixed(-47270540.0/4294967296.0,1,-nbitq), 
to_sfixed(916423980.0/4294967296.0,1,-nbitq), 
to_sfixed(-45653481.0/4294967296.0,1,-nbitq), 
to_sfixed(-54093436.0/4294967296.0,1,-nbitq), 
to_sfixed(-156429418.0/4294967296.0,1,-nbitq), 
to_sfixed(92361915.0/4294967296.0,1,-nbitq), 
to_sfixed(-247789978.0/4294967296.0,1,-nbitq), 
to_sfixed(42607756.0/4294967296.0,1,-nbitq), 
to_sfixed(68450008.0/4294967296.0,1,-nbitq), 
to_sfixed(-317949744.0/4294967296.0,1,-nbitq), 
to_sfixed(522509485.0/4294967296.0,1,-nbitq), 
to_sfixed(-220178472.0/4294967296.0,1,-nbitq), 
to_sfixed(-165790502.0/4294967296.0,1,-nbitq), 
to_sfixed(-67286211.0/4294967296.0,1,-nbitq), 
to_sfixed(596933719.0/4294967296.0,1,-nbitq), 
to_sfixed(-93656274.0/4294967296.0,1,-nbitq), 
to_sfixed(-547104172.0/4294967296.0,1,-nbitq), 
to_sfixed(792228536.0/4294967296.0,1,-nbitq), 
to_sfixed(-10237943.0/4294967296.0,1,-nbitq), 
to_sfixed(-392986556.0/4294967296.0,1,-nbitq), 
to_sfixed(60922313.0/4294967296.0,1,-nbitq), 
to_sfixed(287535380.0/4294967296.0,1,-nbitq), 
to_sfixed(-498567020.0/4294967296.0,1,-nbitq), 
to_sfixed(55003911.0/4294967296.0,1,-nbitq), 
to_sfixed(268962801.0/4294967296.0,1,-nbitq), 
to_sfixed(30240346.0/4294967296.0,1,-nbitq), 
to_sfixed(113031708.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(33169398.0/4294967296.0,1,-nbitq), 
to_sfixed(959573928.0/4294967296.0,1,-nbitq), 
to_sfixed(73458364.0/4294967296.0,1,-nbitq), 
to_sfixed(633691145.0/4294967296.0,1,-nbitq), 
to_sfixed(508431699.0/4294967296.0,1,-nbitq), 
to_sfixed(-195044610.0/4294967296.0,1,-nbitq), 
to_sfixed(377182797.0/4294967296.0,1,-nbitq), 
to_sfixed(-540240795.0/4294967296.0,1,-nbitq), 
to_sfixed(-462949247.0/4294967296.0,1,-nbitq), 
to_sfixed(-268817048.0/4294967296.0,1,-nbitq), 
to_sfixed(314738981.0/4294967296.0,1,-nbitq), 
to_sfixed(-350219526.0/4294967296.0,1,-nbitq), 
to_sfixed(1039389433.0/4294967296.0,1,-nbitq), 
to_sfixed(824877171.0/4294967296.0,1,-nbitq), 
to_sfixed(399130751.0/4294967296.0,1,-nbitq), 
to_sfixed(-888486671.0/4294967296.0,1,-nbitq), 
to_sfixed(148609259.0/4294967296.0,1,-nbitq), 
to_sfixed(-278510301.0/4294967296.0,1,-nbitq), 
to_sfixed(-133712228.0/4294967296.0,1,-nbitq), 
to_sfixed(343309831.0/4294967296.0,1,-nbitq), 
to_sfixed(-15693940.0/4294967296.0,1,-nbitq), 
to_sfixed(123685187.0/4294967296.0,1,-nbitq), 
to_sfixed(-198224278.0/4294967296.0,1,-nbitq), 
to_sfixed(730745364.0/4294967296.0,1,-nbitq), 
to_sfixed(284419878.0/4294967296.0,1,-nbitq), 
to_sfixed(600648993.0/4294967296.0,1,-nbitq), 
to_sfixed(210643093.0/4294967296.0,1,-nbitq), 
to_sfixed(-175256063.0/4294967296.0,1,-nbitq), 
to_sfixed(675136246.0/4294967296.0,1,-nbitq), 
to_sfixed(-15235168.0/4294967296.0,1,-nbitq), 
to_sfixed(-258850880.0/4294967296.0,1,-nbitq), 
to_sfixed(251117290.0/4294967296.0,1,-nbitq), 
to_sfixed(26816871.0/4294967296.0,1,-nbitq), 
to_sfixed(188591697.0/4294967296.0,1,-nbitq), 
to_sfixed(-27204173.0/4294967296.0,1,-nbitq), 
to_sfixed(-5707777.0/4294967296.0,1,-nbitq), 
to_sfixed(306651856.0/4294967296.0,1,-nbitq), 
to_sfixed(936868424.0/4294967296.0,1,-nbitq), 
to_sfixed(-513244282.0/4294967296.0,1,-nbitq), 
to_sfixed(545929598.0/4294967296.0,1,-nbitq), 
to_sfixed(-78334185.0/4294967296.0,1,-nbitq), 
to_sfixed(31034286.0/4294967296.0,1,-nbitq), 
to_sfixed(208840807.0/4294967296.0,1,-nbitq), 
to_sfixed(-59584358.0/4294967296.0,1,-nbitq), 
to_sfixed(580797272.0/4294967296.0,1,-nbitq), 
to_sfixed(493591913.0/4294967296.0,1,-nbitq), 
to_sfixed(-424637809.0/4294967296.0,1,-nbitq), 
to_sfixed(-482381181.0/4294967296.0,1,-nbitq), 
to_sfixed(-11640206.0/4294967296.0,1,-nbitq), 
to_sfixed(-441568331.0/4294967296.0,1,-nbitq), 
to_sfixed(-211814177.0/4294967296.0,1,-nbitq), 
to_sfixed(-147680542.0/4294967296.0,1,-nbitq), 
to_sfixed(464493052.0/4294967296.0,1,-nbitq), 
to_sfixed(-654896685.0/4294967296.0,1,-nbitq), 
to_sfixed(381191167.0/4294967296.0,1,-nbitq), 
to_sfixed(501272558.0/4294967296.0,1,-nbitq), 
to_sfixed(334011158.0/4294967296.0,1,-nbitq), 
to_sfixed(138263585.0/4294967296.0,1,-nbitq), 
to_sfixed(-205137130.0/4294967296.0,1,-nbitq), 
to_sfixed(-312491103.0/4294967296.0,1,-nbitq), 
to_sfixed(351805735.0/4294967296.0,1,-nbitq), 
to_sfixed(-354548767.0/4294967296.0,1,-nbitq), 
to_sfixed(-1462993131.0/4294967296.0,1,-nbitq), 
to_sfixed(282962299.0/4294967296.0,1,-nbitq), 
to_sfixed(-709390728.0/4294967296.0,1,-nbitq), 
to_sfixed(-484972257.0/4294967296.0,1,-nbitq), 
to_sfixed(-40121230.0/4294967296.0,1,-nbitq), 
to_sfixed(110975635.0/4294967296.0,1,-nbitq), 
to_sfixed(5044149.0/4294967296.0,1,-nbitq), 
to_sfixed(-181943913.0/4294967296.0,1,-nbitq), 
to_sfixed(428763939.0/4294967296.0,1,-nbitq), 
to_sfixed(-207365341.0/4294967296.0,1,-nbitq), 
to_sfixed(-347776987.0/4294967296.0,1,-nbitq), 
to_sfixed(259996791.0/4294967296.0,1,-nbitq), 
to_sfixed(419841440.0/4294967296.0,1,-nbitq), 
to_sfixed(69705012.0/4294967296.0,1,-nbitq), 
to_sfixed(331682868.0/4294967296.0,1,-nbitq), 
to_sfixed(410755867.0/4294967296.0,1,-nbitq), 
to_sfixed(196010652.0/4294967296.0,1,-nbitq), 
to_sfixed(310493693.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(316590775.0/4294967296.0,1,-nbitq), 
to_sfixed(420865710.0/4294967296.0,1,-nbitq), 
to_sfixed(-259813659.0/4294967296.0,1,-nbitq), 
to_sfixed(273630603.0/4294967296.0,1,-nbitq), 
to_sfixed(999028505.0/4294967296.0,1,-nbitq), 
to_sfixed(322014180.0/4294967296.0,1,-nbitq), 
to_sfixed(-91057853.0/4294967296.0,1,-nbitq), 
to_sfixed(-439659397.0/4294967296.0,1,-nbitq), 
to_sfixed(262133694.0/4294967296.0,1,-nbitq), 
to_sfixed(236300672.0/4294967296.0,1,-nbitq), 
to_sfixed(-111279202.0/4294967296.0,1,-nbitq), 
to_sfixed(-719885037.0/4294967296.0,1,-nbitq), 
to_sfixed(1383820055.0/4294967296.0,1,-nbitq), 
to_sfixed(695810230.0/4294967296.0,1,-nbitq), 
to_sfixed(109621803.0/4294967296.0,1,-nbitq), 
to_sfixed(-866197842.0/4294967296.0,1,-nbitq), 
to_sfixed(416154925.0/4294967296.0,1,-nbitq), 
to_sfixed(-48179194.0/4294967296.0,1,-nbitq), 
to_sfixed(375145654.0/4294967296.0,1,-nbitq), 
to_sfixed(685507358.0/4294967296.0,1,-nbitq), 
to_sfixed(-325930525.0/4294967296.0,1,-nbitq), 
to_sfixed(-87326757.0/4294967296.0,1,-nbitq), 
to_sfixed(-529608641.0/4294967296.0,1,-nbitq), 
to_sfixed(545357034.0/4294967296.0,1,-nbitq), 
to_sfixed(-75545928.0/4294967296.0,1,-nbitq), 
to_sfixed(873062462.0/4294967296.0,1,-nbitq), 
to_sfixed(-654610160.0/4294967296.0,1,-nbitq), 
to_sfixed(-49429808.0/4294967296.0,1,-nbitq), 
to_sfixed(367981896.0/4294967296.0,1,-nbitq), 
to_sfixed(-570122462.0/4294967296.0,1,-nbitq), 
to_sfixed(-503855968.0/4294967296.0,1,-nbitq), 
to_sfixed(-391285873.0/4294967296.0,1,-nbitq), 
to_sfixed(-46049802.0/4294967296.0,1,-nbitq), 
to_sfixed(-34035605.0/4294967296.0,1,-nbitq), 
to_sfixed(-262420325.0/4294967296.0,1,-nbitq), 
to_sfixed(280409292.0/4294967296.0,1,-nbitq), 
to_sfixed(287099706.0/4294967296.0,1,-nbitq), 
to_sfixed(535917925.0/4294967296.0,1,-nbitq), 
to_sfixed(-609490812.0/4294967296.0,1,-nbitq), 
to_sfixed(367196148.0/4294967296.0,1,-nbitq), 
to_sfixed(-521459508.0/4294967296.0,1,-nbitq), 
to_sfixed(33270549.0/4294967296.0,1,-nbitq), 
to_sfixed(71450968.0/4294967296.0,1,-nbitq), 
to_sfixed(-24088190.0/4294967296.0,1,-nbitq), 
to_sfixed(-453044397.0/4294967296.0,1,-nbitq), 
to_sfixed(999190025.0/4294967296.0,1,-nbitq), 
to_sfixed(-195890181.0/4294967296.0,1,-nbitq), 
to_sfixed(-1515971229.0/4294967296.0,1,-nbitq), 
to_sfixed(92757426.0/4294967296.0,1,-nbitq), 
to_sfixed(-667387104.0/4294967296.0,1,-nbitq), 
to_sfixed(-58650697.0/4294967296.0,1,-nbitq), 
to_sfixed(-210116286.0/4294967296.0,1,-nbitq), 
to_sfixed(782211371.0/4294967296.0,1,-nbitq), 
to_sfixed(-47835411.0/4294967296.0,1,-nbitq), 
to_sfixed(393297601.0/4294967296.0,1,-nbitq), 
to_sfixed(844761973.0/4294967296.0,1,-nbitq), 
to_sfixed(30372198.0/4294967296.0,1,-nbitq), 
to_sfixed(510528708.0/4294967296.0,1,-nbitq), 
to_sfixed(235460084.0/4294967296.0,1,-nbitq), 
to_sfixed(381799734.0/4294967296.0,1,-nbitq), 
to_sfixed(-170754892.0/4294967296.0,1,-nbitq), 
to_sfixed(2356238.0/4294967296.0,1,-nbitq), 
to_sfixed(-1192306946.0/4294967296.0,1,-nbitq), 
to_sfixed(770378292.0/4294967296.0,1,-nbitq), 
to_sfixed(-26567693.0/4294967296.0,1,-nbitq), 
to_sfixed(189599512.0/4294967296.0,1,-nbitq), 
to_sfixed(-886771001.0/4294967296.0,1,-nbitq), 
to_sfixed(376236029.0/4294967296.0,1,-nbitq), 
to_sfixed(136795472.0/4294967296.0,1,-nbitq), 
to_sfixed(-1324995989.0/4294967296.0,1,-nbitq), 
to_sfixed(106595270.0/4294967296.0,1,-nbitq), 
to_sfixed(591198074.0/4294967296.0,1,-nbitq), 
to_sfixed(322521361.0/4294967296.0,1,-nbitq), 
to_sfixed(127551496.0/4294967296.0,1,-nbitq), 
to_sfixed(-115028668.0/4294967296.0,1,-nbitq), 
to_sfixed(-337942545.0/4294967296.0,1,-nbitq), 
to_sfixed(802620876.0/4294967296.0,1,-nbitq), 
to_sfixed(259244245.0/4294967296.0,1,-nbitq), 
to_sfixed(-173109995.0/4294967296.0,1,-nbitq), 
to_sfixed(440488597.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-258301037.0/4294967296.0,1,-nbitq), 
to_sfixed(45931177.0/4294967296.0,1,-nbitq), 
to_sfixed(-940966040.0/4294967296.0,1,-nbitq), 
to_sfixed(-308719171.0/4294967296.0,1,-nbitq), 
to_sfixed(1059292054.0/4294967296.0,1,-nbitq), 
to_sfixed(1966395158.0/4294967296.0,1,-nbitq), 
to_sfixed(324774003.0/4294967296.0,1,-nbitq), 
to_sfixed(516667597.0/4294967296.0,1,-nbitq), 
to_sfixed(332508539.0/4294967296.0,1,-nbitq), 
to_sfixed(-312480415.0/4294967296.0,1,-nbitq), 
to_sfixed(-244560355.0/4294967296.0,1,-nbitq), 
to_sfixed(-288206439.0/4294967296.0,1,-nbitq), 
to_sfixed(1769238056.0/4294967296.0,1,-nbitq), 
to_sfixed(-79227594.0/4294967296.0,1,-nbitq), 
to_sfixed(-106303879.0/4294967296.0,1,-nbitq), 
to_sfixed(-1164221635.0/4294967296.0,1,-nbitq), 
to_sfixed(-236121239.0/4294967296.0,1,-nbitq), 
to_sfixed(-1388234.0/4294967296.0,1,-nbitq), 
to_sfixed(-3907252.0/4294967296.0,1,-nbitq), 
to_sfixed(462610276.0/4294967296.0,1,-nbitq), 
to_sfixed(-193912919.0/4294967296.0,1,-nbitq), 
to_sfixed(-227676351.0/4294967296.0,1,-nbitq), 
to_sfixed(-400805725.0/4294967296.0,1,-nbitq), 
to_sfixed(788989116.0/4294967296.0,1,-nbitq), 
to_sfixed(389020182.0/4294967296.0,1,-nbitq), 
to_sfixed(1005908325.0/4294967296.0,1,-nbitq), 
to_sfixed(-58118639.0/4294967296.0,1,-nbitq), 
to_sfixed(89988448.0/4294967296.0,1,-nbitq), 
to_sfixed(238475065.0/4294967296.0,1,-nbitq), 
to_sfixed(50818754.0/4294967296.0,1,-nbitq), 
to_sfixed(-476187126.0/4294967296.0,1,-nbitq), 
to_sfixed(-424764760.0/4294967296.0,1,-nbitq), 
to_sfixed(283830871.0/4294967296.0,1,-nbitq), 
to_sfixed(-406259826.0/4294967296.0,1,-nbitq), 
to_sfixed(-314160760.0/4294967296.0,1,-nbitq), 
to_sfixed(983961644.0/4294967296.0,1,-nbitq), 
to_sfixed(502363526.0/4294967296.0,1,-nbitq), 
to_sfixed(-251800520.0/4294967296.0,1,-nbitq), 
to_sfixed(-579101777.0/4294967296.0,1,-nbitq), 
to_sfixed(92749877.0/4294967296.0,1,-nbitq), 
to_sfixed(-463283581.0/4294967296.0,1,-nbitq), 
to_sfixed(-592091911.0/4294967296.0,1,-nbitq), 
to_sfixed(108442443.0/4294967296.0,1,-nbitq), 
to_sfixed(234117739.0/4294967296.0,1,-nbitq), 
to_sfixed(-38854407.0/4294967296.0,1,-nbitq), 
to_sfixed(151989052.0/4294967296.0,1,-nbitq), 
to_sfixed(-154164102.0/4294967296.0,1,-nbitq), 
to_sfixed(-503413559.0/4294967296.0,1,-nbitq), 
to_sfixed(-156692423.0/4294967296.0,1,-nbitq), 
to_sfixed(-898664805.0/4294967296.0,1,-nbitq), 
to_sfixed(450457251.0/4294967296.0,1,-nbitq), 
to_sfixed(-272270699.0/4294967296.0,1,-nbitq), 
to_sfixed(262130301.0/4294967296.0,1,-nbitq), 
to_sfixed(-189369421.0/4294967296.0,1,-nbitq), 
to_sfixed(763963238.0/4294967296.0,1,-nbitq), 
to_sfixed(934952836.0/4294967296.0,1,-nbitq), 
to_sfixed(98806019.0/4294967296.0,1,-nbitq), 
to_sfixed(-209879539.0/4294967296.0,1,-nbitq), 
to_sfixed(57426761.0/4294967296.0,1,-nbitq), 
to_sfixed(148516323.0/4294967296.0,1,-nbitq), 
to_sfixed(-69311456.0/4294967296.0,1,-nbitq), 
to_sfixed(21301653.0/4294967296.0,1,-nbitq), 
to_sfixed(-631234688.0/4294967296.0,1,-nbitq), 
to_sfixed(533638607.0/4294967296.0,1,-nbitq), 
to_sfixed(-109078850.0/4294967296.0,1,-nbitq), 
to_sfixed(-85432455.0/4294967296.0,1,-nbitq), 
to_sfixed(-609518070.0/4294967296.0,1,-nbitq), 
to_sfixed(377784417.0/4294967296.0,1,-nbitq), 
to_sfixed(322994096.0/4294967296.0,1,-nbitq), 
to_sfixed(-1589567358.0/4294967296.0,1,-nbitq), 
to_sfixed(-168701273.0/4294967296.0,1,-nbitq), 
to_sfixed(529207220.0/4294967296.0,1,-nbitq), 
to_sfixed(353958936.0/4294967296.0,1,-nbitq), 
to_sfixed(9549730.0/4294967296.0,1,-nbitq), 
to_sfixed(-146660078.0/4294967296.0,1,-nbitq), 
to_sfixed(-462601720.0/4294967296.0,1,-nbitq), 
to_sfixed(1008052025.0/4294967296.0,1,-nbitq), 
to_sfixed(457605479.0/4294967296.0,1,-nbitq), 
to_sfixed(-746521672.0/4294967296.0,1,-nbitq), 
to_sfixed(24760018.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-71989535.0/4294967296.0,1,-nbitq), 
to_sfixed(-127402394.0/4294967296.0,1,-nbitq), 
to_sfixed(-659283719.0/4294967296.0,1,-nbitq), 
to_sfixed(128697790.0/4294967296.0,1,-nbitq), 
to_sfixed(278059152.0/4294967296.0,1,-nbitq), 
to_sfixed(2226077627.0/4294967296.0,1,-nbitq), 
to_sfixed(-187200419.0/4294967296.0,1,-nbitq), 
to_sfixed(577691177.0/4294967296.0,1,-nbitq), 
to_sfixed(228815147.0/4294967296.0,1,-nbitq), 
to_sfixed(-32616158.0/4294967296.0,1,-nbitq), 
to_sfixed(-622996601.0/4294967296.0,1,-nbitq), 
to_sfixed(209306061.0/4294967296.0,1,-nbitq), 
to_sfixed(943628469.0/4294967296.0,1,-nbitq), 
to_sfixed(74327988.0/4294967296.0,1,-nbitq), 
to_sfixed(61970628.0/4294967296.0,1,-nbitq), 
to_sfixed(-1184919382.0/4294967296.0,1,-nbitq), 
to_sfixed(-319350676.0/4294967296.0,1,-nbitq), 
to_sfixed(139195505.0/4294967296.0,1,-nbitq), 
to_sfixed(-29249028.0/4294967296.0,1,-nbitq), 
to_sfixed(517928573.0/4294967296.0,1,-nbitq), 
to_sfixed(72325654.0/4294967296.0,1,-nbitq), 
to_sfixed(-250521957.0/4294967296.0,1,-nbitq), 
to_sfixed(-360374699.0/4294967296.0,1,-nbitq), 
to_sfixed(1147478254.0/4294967296.0,1,-nbitq), 
to_sfixed(-107837884.0/4294967296.0,1,-nbitq), 
to_sfixed(1197476654.0/4294967296.0,1,-nbitq), 
to_sfixed(-269547279.0/4294967296.0,1,-nbitq), 
to_sfixed(91034330.0/4294967296.0,1,-nbitq), 
to_sfixed(359904493.0/4294967296.0,1,-nbitq), 
to_sfixed(21943792.0/4294967296.0,1,-nbitq), 
to_sfixed(-336962655.0/4294967296.0,1,-nbitq), 
to_sfixed(-604454384.0/4294967296.0,1,-nbitq), 
to_sfixed(324281228.0/4294967296.0,1,-nbitq), 
to_sfixed(8006526.0/4294967296.0,1,-nbitq), 
to_sfixed(-783306797.0/4294967296.0,1,-nbitq), 
to_sfixed(-138373808.0/4294967296.0,1,-nbitq), 
to_sfixed(506087019.0/4294967296.0,1,-nbitq), 
to_sfixed(-1107913834.0/4294967296.0,1,-nbitq), 
to_sfixed(-453358135.0/4294967296.0,1,-nbitq), 
to_sfixed(-325367609.0/4294967296.0,1,-nbitq), 
to_sfixed(-694399353.0/4294967296.0,1,-nbitq), 
to_sfixed(-731970152.0/4294967296.0,1,-nbitq), 
to_sfixed(-402099534.0/4294967296.0,1,-nbitq), 
to_sfixed(-281900817.0/4294967296.0,1,-nbitq), 
to_sfixed(270065547.0/4294967296.0,1,-nbitq), 
to_sfixed(-23939729.0/4294967296.0,1,-nbitq), 
to_sfixed(-238685191.0/4294967296.0,1,-nbitq), 
to_sfixed(-837518232.0/4294967296.0,1,-nbitq), 
to_sfixed(-44181188.0/4294967296.0,1,-nbitq), 
to_sfixed(-1256260895.0/4294967296.0,1,-nbitq), 
to_sfixed(-50308326.0/4294967296.0,1,-nbitq), 
to_sfixed(173032009.0/4294967296.0,1,-nbitq), 
to_sfixed(-21920014.0/4294967296.0,1,-nbitq), 
to_sfixed(324673944.0/4294967296.0,1,-nbitq), 
to_sfixed(-167748403.0/4294967296.0,1,-nbitq), 
to_sfixed(1018699747.0/4294967296.0,1,-nbitq), 
to_sfixed(317816055.0/4294967296.0,1,-nbitq), 
to_sfixed(-14649681.0/4294967296.0,1,-nbitq), 
to_sfixed(-393940058.0/4294967296.0,1,-nbitq), 
to_sfixed(-219652098.0/4294967296.0,1,-nbitq), 
to_sfixed(386606449.0/4294967296.0,1,-nbitq), 
to_sfixed(-106676405.0/4294967296.0,1,-nbitq), 
to_sfixed(-430358841.0/4294967296.0,1,-nbitq), 
to_sfixed(945020105.0/4294967296.0,1,-nbitq), 
to_sfixed(166080703.0/4294967296.0,1,-nbitq), 
to_sfixed(62380238.0/4294967296.0,1,-nbitq), 
to_sfixed(-1310053574.0/4294967296.0,1,-nbitq), 
to_sfixed(-418711068.0/4294967296.0,1,-nbitq), 
to_sfixed(-101273870.0/4294967296.0,1,-nbitq), 
to_sfixed(-1438026263.0/4294967296.0,1,-nbitq), 
to_sfixed(-604697012.0/4294967296.0,1,-nbitq), 
to_sfixed(331277491.0/4294967296.0,1,-nbitq), 
to_sfixed(304973721.0/4294967296.0,1,-nbitq), 
to_sfixed(-138954604.0/4294967296.0,1,-nbitq), 
to_sfixed(-146524587.0/4294967296.0,1,-nbitq), 
to_sfixed(-366191299.0/4294967296.0,1,-nbitq), 
to_sfixed(855884692.0/4294967296.0,1,-nbitq), 
to_sfixed(271115585.0/4294967296.0,1,-nbitq), 
to_sfixed(-1239946624.0/4294967296.0,1,-nbitq), 
to_sfixed(233924277.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-1662220.0/4294967296.0,1,-nbitq), 
to_sfixed(-11605530.0/4294967296.0,1,-nbitq), 
to_sfixed(-843321773.0/4294967296.0,1,-nbitq), 
to_sfixed(136031722.0/4294967296.0,1,-nbitq), 
to_sfixed(216506306.0/4294967296.0,1,-nbitq), 
to_sfixed(1204160449.0/4294967296.0,1,-nbitq), 
to_sfixed(119063347.0/4294967296.0,1,-nbitq), 
to_sfixed(301900989.0/4294967296.0,1,-nbitq), 
to_sfixed(325076953.0/4294967296.0,1,-nbitq), 
to_sfixed(61675199.0/4294967296.0,1,-nbitq), 
to_sfixed(-726541929.0/4294967296.0,1,-nbitq), 
to_sfixed(-244832652.0/4294967296.0,1,-nbitq), 
to_sfixed(1250354078.0/4294967296.0,1,-nbitq), 
to_sfixed(-1053840598.0/4294967296.0,1,-nbitq), 
to_sfixed(62432690.0/4294967296.0,1,-nbitq), 
to_sfixed(-964443124.0/4294967296.0,1,-nbitq), 
to_sfixed(-346734854.0/4294967296.0,1,-nbitq), 
to_sfixed(63952005.0/4294967296.0,1,-nbitq), 
to_sfixed(474506921.0/4294967296.0,1,-nbitq), 
to_sfixed(31497784.0/4294967296.0,1,-nbitq), 
to_sfixed(-188069381.0/4294967296.0,1,-nbitq), 
to_sfixed(-143259942.0/4294967296.0,1,-nbitq), 
to_sfixed(-672054468.0/4294967296.0,1,-nbitq), 
to_sfixed(1333030026.0/4294967296.0,1,-nbitq), 
to_sfixed(285587520.0/4294967296.0,1,-nbitq), 
to_sfixed(259933638.0/4294967296.0,1,-nbitq), 
to_sfixed(71513428.0/4294967296.0,1,-nbitq), 
to_sfixed(522888182.0/4294967296.0,1,-nbitq), 
to_sfixed(744960492.0/4294967296.0,1,-nbitq), 
to_sfixed(-413919531.0/4294967296.0,1,-nbitq), 
to_sfixed(13801418.0/4294967296.0,1,-nbitq), 
to_sfixed(-1539682224.0/4294967296.0,1,-nbitq), 
to_sfixed(627945299.0/4294967296.0,1,-nbitq), 
to_sfixed(342962715.0/4294967296.0,1,-nbitq), 
to_sfixed(-511592648.0/4294967296.0,1,-nbitq), 
to_sfixed(-299906550.0/4294967296.0,1,-nbitq), 
to_sfixed(866493650.0/4294967296.0,1,-nbitq), 
to_sfixed(-1234496226.0/4294967296.0,1,-nbitq), 
to_sfixed(318818164.0/4294967296.0,1,-nbitq), 
to_sfixed(396471815.0/4294967296.0,1,-nbitq), 
to_sfixed(36528668.0/4294967296.0,1,-nbitq), 
to_sfixed(-348396201.0/4294967296.0,1,-nbitq), 
to_sfixed(-133562947.0/4294967296.0,1,-nbitq), 
to_sfixed(-743223712.0/4294967296.0,1,-nbitq), 
to_sfixed(-26332110.0/4294967296.0,1,-nbitq), 
to_sfixed(-45758414.0/4294967296.0,1,-nbitq), 
to_sfixed(141948456.0/4294967296.0,1,-nbitq), 
to_sfixed(81880985.0/4294967296.0,1,-nbitq), 
to_sfixed(-78222686.0/4294967296.0,1,-nbitq), 
to_sfixed(-1187895796.0/4294967296.0,1,-nbitq), 
to_sfixed(-103303801.0/4294967296.0,1,-nbitq), 
to_sfixed(692041169.0/4294967296.0,1,-nbitq), 
to_sfixed(-320114014.0/4294967296.0,1,-nbitq), 
to_sfixed(458842012.0/4294967296.0,1,-nbitq), 
to_sfixed(-801961723.0/4294967296.0,1,-nbitq), 
to_sfixed(472761791.0/4294967296.0,1,-nbitq), 
to_sfixed(418954164.0/4294967296.0,1,-nbitq), 
to_sfixed(520053408.0/4294967296.0,1,-nbitq), 
to_sfixed(361289702.0/4294967296.0,1,-nbitq), 
to_sfixed(-363523890.0/4294967296.0,1,-nbitq), 
to_sfixed(-3974903.0/4294967296.0,1,-nbitq), 
to_sfixed(-191715466.0/4294967296.0,1,-nbitq), 
to_sfixed(-556653096.0/4294967296.0,1,-nbitq), 
to_sfixed(1232447265.0/4294967296.0,1,-nbitq), 
to_sfixed(-286156717.0/4294967296.0,1,-nbitq), 
to_sfixed(-88581096.0/4294967296.0,1,-nbitq), 
to_sfixed(-1444474241.0/4294967296.0,1,-nbitq), 
to_sfixed(153946721.0/4294967296.0,1,-nbitq), 
to_sfixed(44799512.0/4294967296.0,1,-nbitq), 
to_sfixed(-85639269.0/4294967296.0,1,-nbitq), 
to_sfixed(-892861078.0/4294967296.0,1,-nbitq), 
to_sfixed(349233407.0/4294967296.0,1,-nbitq), 
to_sfixed(273771395.0/4294967296.0,1,-nbitq), 
to_sfixed(-286912385.0/4294967296.0,1,-nbitq), 
to_sfixed(-301301225.0/4294967296.0,1,-nbitq), 
to_sfixed(-200298669.0/4294967296.0,1,-nbitq), 
to_sfixed(1229889556.0/4294967296.0,1,-nbitq), 
to_sfixed(103538725.0/4294967296.0,1,-nbitq), 
to_sfixed(-689674492.0/4294967296.0,1,-nbitq), 
to_sfixed(243060370.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-282074006.0/4294967296.0,1,-nbitq), 
to_sfixed(-181800153.0/4294967296.0,1,-nbitq), 
to_sfixed(-658468996.0/4294967296.0,1,-nbitq), 
to_sfixed(-368347177.0/4294967296.0,1,-nbitq), 
to_sfixed(202350554.0/4294967296.0,1,-nbitq), 
to_sfixed(-863678867.0/4294967296.0,1,-nbitq), 
to_sfixed(-221835929.0/4294967296.0,1,-nbitq), 
to_sfixed(-765035761.0/4294967296.0,1,-nbitq), 
to_sfixed(1279866020.0/4294967296.0,1,-nbitq), 
to_sfixed(-260920015.0/4294967296.0,1,-nbitq), 
to_sfixed(-1867153612.0/4294967296.0,1,-nbitq), 
to_sfixed(-472241922.0/4294967296.0,1,-nbitq), 
to_sfixed(753396284.0/4294967296.0,1,-nbitq), 
to_sfixed(-517232697.0/4294967296.0,1,-nbitq), 
to_sfixed(-119913104.0/4294967296.0,1,-nbitq), 
to_sfixed(-434446602.0/4294967296.0,1,-nbitq), 
to_sfixed(-182134856.0/4294967296.0,1,-nbitq), 
to_sfixed(-194967178.0/4294967296.0,1,-nbitq), 
to_sfixed(1020237611.0/4294967296.0,1,-nbitq), 
to_sfixed(-360288775.0/4294967296.0,1,-nbitq), 
to_sfixed(108187277.0/4294967296.0,1,-nbitq), 
to_sfixed(265998711.0/4294967296.0,1,-nbitq), 
to_sfixed(-920180099.0/4294967296.0,1,-nbitq), 
to_sfixed(-300269551.0/4294967296.0,1,-nbitq), 
to_sfixed(-341588524.0/4294967296.0,1,-nbitq), 
to_sfixed(122464167.0/4294967296.0,1,-nbitq), 
to_sfixed(123701438.0/4294967296.0,1,-nbitq), 
to_sfixed(1076986546.0/4294967296.0,1,-nbitq), 
to_sfixed(1704062780.0/4294967296.0,1,-nbitq), 
to_sfixed(-1239447569.0/4294967296.0,1,-nbitq), 
to_sfixed(103599001.0/4294967296.0,1,-nbitq), 
to_sfixed(-1311186602.0/4294967296.0,1,-nbitq), 
to_sfixed(129821484.0/4294967296.0,1,-nbitq), 
to_sfixed(144917969.0/4294967296.0,1,-nbitq), 
to_sfixed(-489096726.0/4294967296.0,1,-nbitq), 
to_sfixed(-818586332.0/4294967296.0,1,-nbitq), 
to_sfixed(635267855.0/4294967296.0,1,-nbitq), 
to_sfixed(-429354111.0/4294967296.0,1,-nbitq), 
to_sfixed(549239980.0/4294967296.0,1,-nbitq), 
to_sfixed(363109130.0/4294967296.0,1,-nbitq), 
to_sfixed(-143790749.0/4294967296.0,1,-nbitq), 
to_sfixed(-458755196.0/4294967296.0,1,-nbitq), 
to_sfixed(-70995402.0/4294967296.0,1,-nbitq), 
to_sfixed(53280064.0/4294967296.0,1,-nbitq), 
to_sfixed(364689563.0/4294967296.0,1,-nbitq), 
to_sfixed(-726435374.0/4294967296.0,1,-nbitq), 
to_sfixed(45171449.0/4294967296.0,1,-nbitq), 
to_sfixed(-283742075.0/4294967296.0,1,-nbitq), 
to_sfixed(-307908365.0/4294967296.0,1,-nbitq), 
to_sfixed(-1122777059.0/4294967296.0,1,-nbitq), 
to_sfixed(-791008577.0/4294967296.0,1,-nbitq), 
to_sfixed(290139317.0/4294967296.0,1,-nbitq), 
to_sfixed(-298317776.0/4294967296.0,1,-nbitq), 
to_sfixed(882943771.0/4294967296.0,1,-nbitq), 
to_sfixed(-708347384.0/4294967296.0,1,-nbitq), 
to_sfixed(988121432.0/4294967296.0,1,-nbitq), 
to_sfixed(151255976.0/4294967296.0,1,-nbitq), 
to_sfixed(1342517189.0/4294967296.0,1,-nbitq), 
to_sfixed(417022343.0/4294967296.0,1,-nbitq), 
to_sfixed(-176314062.0/4294967296.0,1,-nbitq), 
to_sfixed(495677731.0/4294967296.0,1,-nbitq), 
to_sfixed(855406531.0/4294967296.0,1,-nbitq), 
to_sfixed(523696642.0/4294967296.0,1,-nbitq), 
to_sfixed(268173917.0/4294967296.0,1,-nbitq), 
to_sfixed(293141475.0/4294967296.0,1,-nbitq), 
to_sfixed(286637923.0/4294967296.0,1,-nbitq), 
to_sfixed(-554624053.0/4294967296.0,1,-nbitq), 
to_sfixed(-69325433.0/4294967296.0,1,-nbitq), 
to_sfixed(-330482102.0/4294967296.0,1,-nbitq), 
to_sfixed(-111956277.0/4294967296.0,1,-nbitq), 
to_sfixed(-474624554.0/4294967296.0,1,-nbitq), 
to_sfixed(-120872016.0/4294967296.0,1,-nbitq), 
to_sfixed(358968056.0/4294967296.0,1,-nbitq), 
to_sfixed(81528304.0/4294967296.0,1,-nbitq), 
to_sfixed(-217281129.0/4294967296.0,1,-nbitq), 
to_sfixed(874140002.0/4294967296.0,1,-nbitq), 
to_sfixed(1718227562.0/4294967296.0,1,-nbitq), 
to_sfixed(557165702.0/4294967296.0,1,-nbitq), 
to_sfixed(-496214127.0/4294967296.0,1,-nbitq), 
to_sfixed(-196882303.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-404765133.0/4294967296.0,1,-nbitq), 
to_sfixed(-545823988.0/4294967296.0,1,-nbitq), 
to_sfixed(-661803036.0/4294967296.0,1,-nbitq), 
to_sfixed(-102252330.0/4294967296.0,1,-nbitq), 
to_sfixed(696837489.0/4294967296.0,1,-nbitq), 
to_sfixed(-598545017.0/4294967296.0,1,-nbitq), 
to_sfixed(-685285641.0/4294967296.0,1,-nbitq), 
to_sfixed(-1487120554.0/4294967296.0,1,-nbitq), 
to_sfixed(846314076.0/4294967296.0,1,-nbitq), 
to_sfixed(78954447.0/4294967296.0,1,-nbitq), 
to_sfixed(-1158941399.0/4294967296.0,1,-nbitq), 
to_sfixed(-209759031.0/4294967296.0,1,-nbitq), 
to_sfixed(552343350.0/4294967296.0,1,-nbitq), 
to_sfixed(-1291223864.0/4294967296.0,1,-nbitq), 
to_sfixed(211040820.0/4294967296.0,1,-nbitq), 
to_sfixed(-1559219930.0/4294967296.0,1,-nbitq), 
to_sfixed(-287571245.0/4294967296.0,1,-nbitq), 
to_sfixed(389353943.0/4294967296.0,1,-nbitq), 
to_sfixed(1210581409.0/4294967296.0,1,-nbitq), 
to_sfixed(-12445031.0/4294967296.0,1,-nbitq), 
to_sfixed(92339503.0/4294967296.0,1,-nbitq), 
to_sfixed(372905185.0/4294967296.0,1,-nbitq), 
to_sfixed(-290524184.0/4294967296.0,1,-nbitq), 
to_sfixed(-131633881.0/4294967296.0,1,-nbitq), 
to_sfixed(-340242583.0/4294967296.0,1,-nbitq), 
to_sfixed(144060261.0/4294967296.0,1,-nbitq), 
to_sfixed(-188451277.0/4294967296.0,1,-nbitq), 
to_sfixed(1218067483.0/4294967296.0,1,-nbitq), 
to_sfixed(420212030.0/4294967296.0,1,-nbitq), 
to_sfixed(-801800080.0/4294967296.0,1,-nbitq), 
to_sfixed(1062724547.0/4294967296.0,1,-nbitq), 
to_sfixed(-199143371.0/4294967296.0,1,-nbitq), 
to_sfixed(30813591.0/4294967296.0,1,-nbitq), 
to_sfixed(188578841.0/4294967296.0,1,-nbitq), 
to_sfixed(-187132986.0/4294967296.0,1,-nbitq), 
to_sfixed(-592131975.0/4294967296.0,1,-nbitq), 
to_sfixed(-283994637.0/4294967296.0,1,-nbitq), 
to_sfixed(-267658004.0/4294967296.0,1,-nbitq), 
to_sfixed(363388471.0/4294967296.0,1,-nbitq), 
to_sfixed(230476141.0/4294967296.0,1,-nbitq), 
to_sfixed(566365492.0/4294967296.0,1,-nbitq), 
to_sfixed(132278101.0/4294967296.0,1,-nbitq), 
to_sfixed(613844966.0/4294967296.0,1,-nbitq), 
to_sfixed(-1049837283.0/4294967296.0,1,-nbitq), 
to_sfixed(114163949.0/4294967296.0,1,-nbitq), 
to_sfixed(-501273678.0/4294967296.0,1,-nbitq), 
to_sfixed(95208614.0/4294967296.0,1,-nbitq), 
to_sfixed(-972269388.0/4294967296.0,1,-nbitq), 
to_sfixed(-362297999.0/4294967296.0,1,-nbitq), 
to_sfixed(-938078907.0/4294967296.0,1,-nbitq), 
to_sfixed(-196095198.0/4294967296.0,1,-nbitq), 
to_sfixed(727153086.0/4294967296.0,1,-nbitq), 
to_sfixed(-229781599.0/4294967296.0,1,-nbitq), 
to_sfixed(816736522.0/4294967296.0,1,-nbitq), 
to_sfixed(-1246316030.0/4294967296.0,1,-nbitq), 
to_sfixed(570207672.0/4294967296.0,1,-nbitq), 
to_sfixed(36671652.0/4294967296.0,1,-nbitq), 
to_sfixed(1054053263.0/4294967296.0,1,-nbitq), 
to_sfixed(-100815945.0/4294967296.0,1,-nbitq), 
to_sfixed(350213082.0/4294967296.0,1,-nbitq), 
to_sfixed(-130878305.0/4294967296.0,1,-nbitq), 
to_sfixed(301624810.0/4294967296.0,1,-nbitq), 
to_sfixed(90986425.0/4294967296.0,1,-nbitq), 
to_sfixed(871469788.0/4294967296.0,1,-nbitq), 
to_sfixed(277944971.0/4294967296.0,1,-nbitq), 
to_sfixed(464878496.0/4294967296.0,1,-nbitq), 
to_sfixed(151282751.0/4294967296.0,1,-nbitq), 
to_sfixed(-690396055.0/4294967296.0,1,-nbitq), 
to_sfixed(-84818811.0/4294967296.0,1,-nbitq), 
to_sfixed(-322511271.0/4294967296.0,1,-nbitq), 
to_sfixed(-862360162.0/4294967296.0,1,-nbitq), 
to_sfixed(-504768384.0/4294967296.0,1,-nbitq), 
to_sfixed(-101533961.0/4294967296.0,1,-nbitq), 
to_sfixed(17727437.0/4294967296.0,1,-nbitq), 
to_sfixed(-430696827.0/4294967296.0,1,-nbitq), 
to_sfixed(771051690.0/4294967296.0,1,-nbitq), 
to_sfixed(503752651.0/4294967296.0,1,-nbitq), 
to_sfixed(900049885.0/4294967296.0,1,-nbitq), 
to_sfixed(-106525257.0/4294967296.0,1,-nbitq), 
to_sfixed(231595831.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-939616781.0/4294967296.0,1,-nbitq), 
to_sfixed(-1251041731.0/4294967296.0,1,-nbitq), 
to_sfixed(-315696039.0/4294967296.0,1,-nbitq), 
to_sfixed(374830862.0/4294967296.0,1,-nbitq), 
to_sfixed(417666930.0/4294967296.0,1,-nbitq), 
to_sfixed(-378551396.0/4294967296.0,1,-nbitq), 
to_sfixed(-258184585.0/4294967296.0,1,-nbitq), 
to_sfixed(-346176627.0/4294967296.0,1,-nbitq), 
to_sfixed(1615986618.0/4294967296.0,1,-nbitq), 
to_sfixed(31232098.0/4294967296.0,1,-nbitq), 
to_sfixed(97486547.0/4294967296.0,1,-nbitq), 
to_sfixed(-570746665.0/4294967296.0,1,-nbitq), 
to_sfixed(795025056.0/4294967296.0,1,-nbitq), 
to_sfixed(-1067113827.0/4294967296.0,1,-nbitq), 
to_sfixed(-173793206.0/4294967296.0,1,-nbitq), 
to_sfixed(-1280760509.0/4294967296.0,1,-nbitq), 
to_sfixed(-294252688.0/4294967296.0,1,-nbitq), 
to_sfixed(196838125.0/4294967296.0,1,-nbitq), 
to_sfixed(632828731.0/4294967296.0,1,-nbitq), 
to_sfixed(-72564764.0/4294967296.0,1,-nbitq), 
to_sfixed(-369394719.0/4294967296.0,1,-nbitq), 
to_sfixed(-74073138.0/4294967296.0,1,-nbitq), 
to_sfixed(-125751937.0/4294967296.0,1,-nbitq), 
to_sfixed(-648339351.0/4294967296.0,1,-nbitq), 
to_sfixed(392557407.0/4294967296.0,1,-nbitq), 
to_sfixed(562141977.0/4294967296.0,1,-nbitq), 
to_sfixed(-635203098.0/4294967296.0,1,-nbitq), 
to_sfixed(517086368.0/4294967296.0,1,-nbitq), 
to_sfixed(-764749289.0/4294967296.0,1,-nbitq), 
to_sfixed(-345628675.0/4294967296.0,1,-nbitq), 
to_sfixed(1057687288.0/4294967296.0,1,-nbitq), 
to_sfixed(617682613.0/4294967296.0,1,-nbitq), 
to_sfixed(-215240971.0/4294967296.0,1,-nbitq), 
to_sfixed(351013081.0/4294967296.0,1,-nbitq), 
to_sfixed(81276559.0/4294967296.0,1,-nbitq), 
to_sfixed(1062116567.0/4294967296.0,1,-nbitq), 
to_sfixed(-47742857.0/4294967296.0,1,-nbitq), 
to_sfixed(-416358324.0/4294967296.0,1,-nbitq), 
to_sfixed(425054239.0/4294967296.0,1,-nbitq), 
to_sfixed(87156053.0/4294967296.0,1,-nbitq), 
to_sfixed(743474176.0/4294967296.0,1,-nbitq), 
to_sfixed(41128568.0/4294967296.0,1,-nbitq), 
to_sfixed(1108393874.0/4294967296.0,1,-nbitq), 
to_sfixed(-4104244.0/4294967296.0,1,-nbitq), 
to_sfixed(-837520191.0/4294967296.0,1,-nbitq), 
to_sfixed(-1330457409.0/4294967296.0,1,-nbitq), 
to_sfixed(128118055.0/4294967296.0,1,-nbitq), 
to_sfixed(-1086866523.0/4294967296.0,1,-nbitq), 
to_sfixed(-606754680.0/4294967296.0,1,-nbitq), 
to_sfixed(-984234909.0/4294967296.0,1,-nbitq), 
to_sfixed(-317060983.0/4294967296.0,1,-nbitq), 
to_sfixed(143019362.0/4294967296.0,1,-nbitq), 
to_sfixed(-682930463.0/4294967296.0,1,-nbitq), 
to_sfixed(1430479858.0/4294967296.0,1,-nbitq), 
to_sfixed(-552778338.0/4294967296.0,1,-nbitq), 
to_sfixed(365698064.0/4294967296.0,1,-nbitq), 
to_sfixed(623031633.0/4294967296.0,1,-nbitq), 
to_sfixed(357916296.0/4294967296.0,1,-nbitq), 
to_sfixed(-177148456.0/4294967296.0,1,-nbitq), 
to_sfixed(-356373786.0/4294967296.0,1,-nbitq), 
to_sfixed(295832500.0/4294967296.0,1,-nbitq), 
to_sfixed(791156514.0/4294967296.0,1,-nbitq), 
to_sfixed(-196068166.0/4294967296.0,1,-nbitq), 
to_sfixed(715814454.0/4294967296.0,1,-nbitq), 
to_sfixed(-144311881.0/4294967296.0,1,-nbitq), 
to_sfixed(55853601.0/4294967296.0,1,-nbitq), 
to_sfixed(774285369.0/4294967296.0,1,-nbitq), 
to_sfixed(-935384430.0/4294967296.0,1,-nbitq), 
to_sfixed(167784749.0/4294967296.0,1,-nbitq), 
to_sfixed(50999383.0/4294967296.0,1,-nbitq), 
to_sfixed(-1146119438.0/4294967296.0,1,-nbitq), 
to_sfixed(-622734052.0/4294967296.0,1,-nbitq), 
to_sfixed(144899107.0/4294967296.0,1,-nbitq), 
to_sfixed(-341782297.0/4294967296.0,1,-nbitq), 
to_sfixed(-440015627.0/4294967296.0,1,-nbitq), 
to_sfixed(870990420.0/4294967296.0,1,-nbitq), 
to_sfixed(971694012.0/4294967296.0,1,-nbitq), 
to_sfixed(167471113.0/4294967296.0,1,-nbitq), 
to_sfixed(26249403.0/4294967296.0,1,-nbitq), 
to_sfixed(-274305855.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-208800674.0/4294967296.0,1,-nbitq), 
to_sfixed(-348800146.0/4294967296.0,1,-nbitq), 
to_sfixed(679541339.0/4294967296.0,1,-nbitq), 
to_sfixed(-162668261.0/4294967296.0,1,-nbitq), 
to_sfixed(95178997.0/4294967296.0,1,-nbitq), 
to_sfixed(-636528897.0/4294967296.0,1,-nbitq), 
to_sfixed(149648816.0/4294967296.0,1,-nbitq), 
to_sfixed(-194300216.0/4294967296.0,1,-nbitq), 
to_sfixed(1398947676.0/4294967296.0,1,-nbitq), 
to_sfixed(-102195452.0/4294967296.0,1,-nbitq), 
to_sfixed(-82876032.0/4294967296.0,1,-nbitq), 
to_sfixed(-1344146521.0/4294967296.0,1,-nbitq), 
to_sfixed(-399399125.0/4294967296.0,1,-nbitq), 
to_sfixed(494699406.0/4294967296.0,1,-nbitq), 
to_sfixed(476853814.0/4294967296.0,1,-nbitq), 
to_sfixed(-797264617.0/4294967296.0,1,-nbitq), 
to_sfixed(-323196752.0/4294967296.0,1,-nbitq), 
to_sfixed(102011558.0/4294967296.0,1,-nbitq), 
to_sfixed(1225489100.0/4294967296.0,1,-nbitq), 
to_sfixed(445187894.0/4294967296.0,1,-nbitq), 
to_sfixed(-295783218.0/4294967296.0,1,-nbitq), 
to_sfixed(864110579.0/4294967296.0,1,-nbitq), 
to_sfixed(106050496.0/4294967296.0,1,-nbitq), 
to_sfixed(-1581033008.0/4294967296.0,1,-nbitq), 
to_sfixed(-286343667.0/4294967296.0,1,-nbitq), 
to_sfixed(289422129.0/4294967296.0,1,-nbitq), 
to_sfixed(-287536405.0/4294967296.0,1,-nbitq), 
to_sfixed(-77135957.0/4294967296.0,1,-nbitq), 
to_sfixed(-1407663048.0/4294967296.0,1,-nbitq), 
to_sfixed(-663104496.0/4294967296.0,1,-nbitq), 
to_sfixed(441142499.0/4294967296.0,1,-nbitq), 
to_sfixed(808242643.0/4294967296.0,1,-nbitq), 
to_sfixed(-477131658.0/4294967296.0,1,-nbitq), 
to_sfixed(120231431.0/4294967296.0,1,-nbitq), 
to_sfixed(264946181.0/4294967296.0,1,-nbitq), 
to_sfixed(708802837.0/4294967296.0,1,-nbitq), 
to_sfixed(-1090156149.0/4294967296.0,1,-nbitq), 
to_sfixed(216389004.0/4294967296.0,1,-nbitq), 
to_sfixed(158323786.0/4294967296.0,1,-nbitq), 
to_sfixed(-73606207.0/4294967296.0,1,-nbitq), 
to_sfixed(26849497.0/4294967296.0,1,-nbitq), 
to_sfixed(290094085.0/4294967296.0,1,-nbitq), 
to_sfixed(1234533627.0/4294967296.0,1,-nbitq), 
to_sfixed(519883131.0/4294967296.0,1,-nbitq), 
to_sfixed(-984985504.0/4294967296.0,1,-nbitq), 
to_sfixed(-1078268218.0/4294967296.0,1,-nbitq), 
to_sfixed(68864540.0/4294967296.0,1,-nbitq), 
to_sfixed(-1420915718.0/4294967296.0,1,-nbitq), 
to_sfixed(-116146828.0/4294967296.0,1,-nbitq), 
to_sfixed(-33707736.0/4294967296.0,1,-nbitq), 
to_sfixed(248724339.0/4294967296.0,1,-nbitq), 
to_sfixed(-419129241.0/4294967296.0,1,-nbitq), 
to_sfixed(-608909973.0/4294967296.0,1,-nbitq), 
to_sfixed(1715152643.0/4294967296.0,1,-nbitq), 
to_sfixed(-202073680.0/4294967296.0,1,-nbitq), 
to_sfixed(717915490.0/4294967296.0,1,-nbitq), 
to_sfixed(462011258.0/4294967296.0,1,-nbitq), 
to_sfixed(-151525746.0/4294967296.0,1,-nbitq), 
to_sfixed(165940672.0/4294967296.0,1,-nbitq), 
to_sfixed(-154371621.0/4294967296.0,1,-nbitq), 
to_sfixed(-315129858.0/4294967296.0,1,-nbitq), 
to_sfixed(201627071.0/4294967296.0,1,-nbitq), 
to_sfixed(295560585.0/4294967296.0,1,-nbitq), 
to_sfixed(900537882.0/4294967296.0,1,-nbitq), 
to_sfixed(220518449.0/4294967296.0,1,-nbitq), 
to_sfixed(-76790357.0/4294967296.0,1,-nbitq), 
to_sfixed(175669507.0/4294967296.0,1,-nbitq), 
to_sfixed(-662143935.0/4294967296.0,1,-nbitq), 
to_sfixed(435041063.0/4294967296.0,1,-nbitq), 
to_sfixed(-1472428656.0/4294967296.0,1,-nbitq), 
to_sfixed(-1161033723.0/4294967296.0,1,-nbitq), 
to_sfixed(-441883062.0/4294967296.0,1,-nbitq), 
to_sfixed(503615737.0/4294967296.0,1,-nbitq), 
to_sfixed(-23266522.0/4294967296.0,1,-nbitq), 
to_sfixed(-7802409.0/4294967296.0,1,-nbitq), 
to_sfixed(419136920.0/4294967296.0,1,-nbitq), 
to_sfixed(994256998.0/4294967296.0,1,-nbitq), 
to_sfixed(-114773860.0/4294967296.0,1,-nbitq), 
to_sfixed(846073463.0/4294967296.0,1,-nbitq), 
to_sfixed(-222755381.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(66543697.0/4294967296.0,1,-nbitq), 
to_sfixed(1077648856.0/4294967296.0,1,-nbitq), 
to_sfixed(457406520.0/4294967296.0,1,-nbitq), 
to_sfixed(-190871414.0/4294967296.0,1,-nbitq), 
to_sfixed(627141319.0/4294967296.0,1,-nbitq), 
to_sfixed(-688007667.0/4294967296.0,1,-nbitq), 
to_sfixed(-443253111.0/4294967296.0,1,-nbitq), 
to_sfixed(442556867.0/4294967296.0,1,-nbitq), 
to_sfixed(1050801011.0/4294967296.0,1,-nbitq), 
to_sfixed(-402337552.0/4294967296.0,1,-nbitq), 
to_sfixed(496950428.0/4294967296.0,1,-nbitq), 
to_sfixed(-329744898.0/4294967296.0,1,-nbitq), 
to_sfixed(839002651.0/4294967296.0,1,-nbitq), 
to_sfixed(888710870.0/4294967296.0,1,-nbitq), 
to_sfixed(339827279.0/4294967296.0,1,-nbitq), 
to_sfixed(-566178727.0/4294967296.0,1,-nbitq), 
to_sfixed(-274652844.0/4294967296.0,1,-nbitq), 
to_sfixed(-295308180.0/4294967296.0,1,-nbitq), 
to_sfixed(204100319.0/4294967296.0,1,-nbitq), 
to_sfixed(283511777.0/4294967296.0,1,-nbitq), 
to_sfixed(-316162440.0/4294967296.0,1,-nbitq), 
to_sfixed(1541206353.0/4294967296.0,1,-nbitq), 
to_sfixed(938190604.0/4294967296.0,1,-nbitq), 
to_sfixed(-2065504992.0/4294967296.0,1,-nbitq), 
to_sfixed(83568328.0/4294967296.0,1,-nbitq), 
to_sfixed(183096798.0/4294967296.0,1,-nbitq), 
to_sfixed(685457264.0/4294967296.0,1,-nbitq), 
to_sfixed(-233012453.0/4294967296.0,1,-nbitq), 
to_sfixed(-1921851782.0/4294967296.0,1,-nbitq), 
to_sfixed(-461799265.0/4294967296.0,1,-nbitq), 
to_sfixed(182607191.0/4294967296.0,1,-nbitq), 
to_sfixed(814825638.0/4294967296.0,1,-nbitq), 
to_sfixed(-3728823.0/4294967296.0,1,-nbitq), 
to_sfixed(-120571845.0/4294967296.0,1,-nbitq), 
to_sfixed(746557862.0/4294967296.0,1,-nbitq), 
to_sfixed(1257058439.0/4294967296.0,1,-nbitq), 
to_sfixed(-407409195.0/4294967296.0,1,-nbitq), 
to_sfixed(-44680397.0/4294967296.0,1,-nbitq), 
to_sfixed(118292166.0/4294967296.0,1,-nbitq), 
to_sfixed(-235140904.0/4294967296.0,1,-nbitq), 
to_sfixed(-455755923.0/4294967296.0,1,-nbitq), 
to_sfixed(333675604.0/4294967296.0,1,-nbitq), 
to_sfixed(97483048.0/4294967296.0,1,-nbitq), 
to_sfixed(283985248.0/4294967296.0,1,-nbitq), 
to_sfixed(-1222951536.0/4294967296.0,1,-nbitq), 
to_sfixed(-289888020.0/4294967296.0,1,-nbitq), 
to_sfixed(-289931393.0/4294967296.0,1,-nbitq), 
to_sfixed(-1105078745.0/4294967296.0,1,-nbitq), 
to_sfixed(-287965539.0/4294967296.0,1,-nbitq), 
to_sfixed(-643083147.0/4294967296.0,1,-nbitq), 
to_sfixed(-229091473.0/4294967296.0,1,-nbitq), 
to_sfixed(-671492461.0/4294967296.0,1,-nbitq), 
to_sfixed(-356169075.0/4294967296.0,1,-nbitq), 
to_sfixed(1642257064.0/4294967296.0,1,-nbitq), 
to_sfixed(166961122.0/4294967296.0,1,-nbitq), 
to_sfixed(581857589.0/4294967296.0,1,-nbitq), 
to_sfixed(295163809.0/4294967296.0,1,-nbitq), 
to_sfixed(40310081.0/4294967296.0,1,-nbitq), 
to_sfixed(105860305.0/4294967296.0,1,-nbitq), 
to_sfixed(-215293928.0/4294967296.0,1,-nbitq), 
to_sfixed(165774418.0/4294967296.0,1,-nbitq), 
to_sfixed(-421634627.0/4294967296.0,1,-nbitq), 
to_sfixed(65301775.0/4294967296.0,1,-nbitq), 
to_sfixed(364891415.0/4294967296.0,1,-nbitq), 
to_sfixed(288458188.0/4294967296.0,1,-nbitq), 
to_sfixed(226200951.0/4294967296.0,1,-nbitq), 
to_sfixed(387754574.0/4294967296.0,1,-nbitq), 
to_sfixed(-79880468.0/4294967296.0,1,-nbitq), 
to_sfixed(-108033007.0/4294967296.0,1,-nbitq), 
to_sfixed(-1041718991.0/4294967296.0,1,-nbitq), 
to_sfixed(-378825924.0/4294967296.0,1,-nbitq), 
to_sfixed(-424468679.0/4294967296.0,1,-nbitq), 
to_sfixed(775385196.0/4294967296.0,1,-nbitq), 
to_sfixed(-225148743.0/4294967296.0,1,-nbitq), 
to_sfixed(80782579.0/4294967296.0,1,-nbitq), 
to_sfixed(743517425.0/4294967296.0,1,-nbitq), 
to_sfixed(1192562266.0/4294967296.0,1,-nbitq), 
to_sfixed(436411796.0/4294967296.0,1,-nbitq), 
to_sfixed(500833365.0/4294967296.0,1,-nbitq), 
to_sfixed(-159269564.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-260212428.0/4294967296.0,1,-nbitq), 
to_sfixed(644912699.0/4294967296.0,1,-nbitq), 
to_sfixed(320232420.0/4294967296.0,1,-nbitq), 
to_sfixed(-438908833.0/4294967296.0,1,-nbitq), 
to_sfixed(81235835.0/4294967296.0,1,-nbitq), 
to_sfixed(-819917282.0/4294967296.0,1,-nbitq), 
to_sfixed(-167957481.0/4294967296.0,1,-nbitq), 
to_sfixed(82543171.0/4294967296.0,1,-nbitq), 
to_sfixed(783817250.0/4294967296.0,1,-nbitq), 
to_sfixed(-346186691.0/4294967296.0,1,-nbitq), 
to_sfixed(1142727046.0/4294967296.0,1,-nbitq), 
to_sfixed(-311575563.0/4294967296.0,1,-nbitq), 
to_sfixed(711510968.0/4294967296.0,1,-nbitq), 
to_sfixed(960063076.0/4294967296.0,1,-nbitq), 
to_sfixed(-52702264.0/4294967296.0,1,-nbitq), 
to_sfixed(-533282265.0/4294967296.0,1,-nbitq), 
to_sfixed(-8106051.0/4294967296.0,1,-nbitq), 
to_sfixed(331696140.0/4294967296.0,1,-nbitq), 
to_sfixed(609496734.0/4294967296.0,1,-nbitq), 
to_sfixed(11048127.0/4294967296.0,1,-nbitq), 
to_sfixed(6404844.0/4294967296.0,1,-nbitq), 
to_sfixed(-76333173.0/4294967296.0,1,-nbitq), 
to_sfixed(240039447.0/4294967296.0,1,-nbitq), 
to_sfixed(-869176851.0/4294967296.0,1,-nbitq), 
to_sfixed(406423840.0/4294967296.0,1,-nbitq), 
to_sfixed(96122917.0/4294967296.0,1,-nbitq), 
to_sfixed(398459189.0/4294967296.0,1,-nbitq), 
to_sfixed(-929732701.0/4294967296.0,1,-nbitq), 
to_sfixed(-1158275888.0/4294967296.0,1,-nbitq), 
to_sfixed(-217919252.0/4294967296.0,1,-nbitq), 
to_sfixed(447613527.0/4294967296.0,1,-nbitq), 
to_sfixed(835267489.0/4294967296.0,1,-nbitq), 
to_sfixed(-660915825.0/4294967296.0,1,-nbitq), 
to_sfixed(-63430116.0/4294967296.0,1,-nbitq), 
to_sfixed(274421188.0/4294967296.0,1,-nbitq), 
to_sfixed(20346246.0/4294967296.0,1,-nbitq), 
to_sfixed(-806037798.0/4294967296.0,1,-nbitq), 
to_sfixed(49380081.0/4294967296.0,1,-nbitq), 
to_sfixed(-227847223.0/4294967296.0,1,-nbitq), 
to_sfixed(20933492.0/4294967296.0,1,-nbitq), 
to_sfixed(62027973.0/4294967296.0,1,-nbitq), 
to_sfixed(1086278574.0/4294967296.0,1,-nbitq), 
to_sfixed(36703507.0/4294967296.0,1,-nbitq), 
to_sfixed(-158015331.0/4294967296.0,1,-nbitq), 
to_sfixed(-681999950.0/4294967296.0,1,-nbitq), 
to_sfixed(-146763780.0/4294967296.0,1,-nbitq), 
to_sfixed(-325074248.0/4294967296.0,1,-nbitq), 
to_sfixed(-408688288.0/4294967296.0,1,-nbitq), 
to_sfixed(279137595.0/4294967296.0,1,-nbitq), 
to_sfixed(-111277594.0/4294967296.0,1,-nbitq), 
to_sfixed(502709610.0/4294967296.0,1,-nbitq), 
to_sfixed(456823244.0/4294967296.0,1,-nbitq), 
to_sfixed(140333453.0/4294967296.0,1,-nbitq), 
to_sfixed(1163515352.0/4294967296.0,1,-nbitq), 
to_sfixed(239935461.0/4294967296.0,1,-nbitq), 
to_sfixed(-670486422.0/4294967296.0,1,-nbitq), 
to_sfixed(-21657135.0/4294967296.0,1,-nbitq), 
to_sfixed(620830150.0/4294967296.0,1,-nbitq), 
to_sfixed(-323724196.0/4294967296.0,1,-nbitq), 
to_sfixed(-47926035.0/4294967296.0,1,-nbitq), 
to_sfixed(-249167354.0/4294967296.0,1,-nbitq), 
to_sfixed(-772035365.0/4294967296.0,1,-nbitq), 
to_sfixed(387411255.0/4294967296.0,1,-nbitq), 
to_sfixed(488925739.0/4294967296.0,1,-nbitq), 
to_sfixed(406210983.0/4294967296.0,1,-nbitq), 
to_sfixed(166080514.0/4294967296.0,1,-nbitq), 
to_sfixed(-630481807.0/4294967296.0,1,-nbitq), 
to_sfixed(-760666351.0/4294967296.0,1,-nbitq), 
to_sfixed(-122754661.0/4294967296.0,1,-nbitq), 
to_sfixed(-1334186142.0/4294967296.0,1,-nbitq), 
to_sfixed(-878710770.0/4294967296.0,1,-nbitq), 
to_sfixed(-364631342.0/4294967296.0,1,-nbitq), 
to_sfixed(290601316.0/4294967296.0,1,-nbitq), 
to_sfixed(355305461.0/4294967296.0,1,-nbitq), 
to_sfixed(-38762606.0/4294967296.0,1,-nbitq), 
to_sfixed(711604828.0/4294967296.0,1,-nbitq), 
to_sfixed(1604282457.0/4294967296.0,1,-nbitq), 
to_sfixed(349058752.0/4294967296.0,1,-nbitq), 
to_sfixed(490916935.0/4294967296.0,1,-nbitq), 
to_sfixed(-219285391.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-294637585.0/4294967296.0,1,-nbitq), 
to_sfixed(542841805.0/4294967296.0,1,-nbitq), 
to_sfixed(-779105349.0/4294967296.0,1,-nbitq), 
to_sfixed(-366940992.0/4294967296.0,1,-nbitq), 
to_sfixed(503779227.0/4294967296.0,1,-nbitq), 
to_sfixed(-1218300526.0/4294967296.0,1,-nbitq), 
to_sfixed(-368332253.0/4294967296.0,1,-nbitq), 
to_sfixed(-171152736.0/4294967296.0,1,-nbitq), 
to_sfixed(849452274.0/4294967296.0,1,-nbitq), 
to_sfixed(-15174293.0/4294967296.0,1,-nbitq), 
to_sfixed(869078434.0/4294967296.0,1,-nbitq), 
to_sfixed(-411370574.0/4294967296.0,1,-nbitq), 
to_sfixed(434400394.0/4294967296.0,1,-nbitq), 
to_sfixed(1238926569.0/4294967296.0,1,-nbitq), 
to_sfixed(-277879294.0/4294967296.0,1,-nbitq), 
to_sfixed(-504738289.0/4294967296.0,1,-nbitq), 
to_sfixed(68484820.0/4294967296.0,1,-nbitq), 
to_sfixed(269060693.0/4294967296.0,1,-nbitq), 
to_sfixed(32952912.0/4294967296.0,1,-nbitq), 
to_sfixed(699738123.0/4294967296.0,1,-nbitq), 
to_sfixed(280511306.0/4294967296.0,1,-nbitq), 
to_sfixed(-163347605.0/4294967296.0,1,-nbitq), 
to_sfixed(667834218.0/4294967296.0,1,-nbitq), 
to_sfixed(-497558565.0/4294967296.0,1,-nbitq), 
to_sfixed(281507274.0/4294967296.0,1,-nbitq), 
to_sfixed(-307184898.0/4294967296.0,1,-nbitq), 
to_sfixed(-195960505.0/4294967296.0,1,-nbitq), 
to_sfixed(-952563682.0/4294967296.0,1,-nbitq), 
to_sfixed(13881684.0/4294967296.0,1,-nbitq), 
to_sfixed(-1071559399.0/4294967296.0,1,-nbitq), 
to_sfixed(-740750579.0/4294967296.0,1,-nbitq), 
to_sfixed(879667906.0/4294967296.0,1,-nbitq), 
to_sfixed(-784241037.0/4294967296.0,1,-nbitq), 
to_sfixed(66914525.0/4294967296.0,1,-nbitq), 
to_sfixed(-113845136.0/4294967296.0,1,-nbitq), 
to_sfixed(466938842.0/4294967296.0,1,-nbitq), 
to_sfixed(75560150.0/4294967296.0,1,-nbitq), 
to_sfixed(80466249.0/4294967296.0,1,-nbitq), 
to_sfixed(252719891.0/4294967296.0,1,-nbitq), 
to_sfixed(-271170165.0/4294967296.0,1,-nbitq), 
to_sfixed(-434266397.0/4294967296.0,1,-nbitq), 
to_sfixed(1320721370.0/4294967296.0,1,-nbitq), 
to_sfixed(317413770.0/4294967296.0,1,-nbitq), 
to_sfixed(42640596.0/4294967296.0,1,-nbitq), 
to_sfixed(-683224543.0/4294967296.0,1,-nbitq), 
to_sfixed(-458198634.0/4294967296.0,1,-nbitq), 
to_sfixed(122622518.0/4294967296.0,1,-nbitq), 
to_sfixed(-724274327.0/4294967296.0,1,-nbitq), 
to_sfixed(-213910498.0/4294967296.0,1,-nbitq), 
to_sfixed(453173681.0/4294967296.0,1,-nbitq), 
to_sfixed(-262047805.0/4294967296.0,1,-nbitq), 
to_sfixed(414697556.0/4294967296.0,1,-nbitq), 
to_sfixed(-420547680.0/4294967296.0,1,-nbitq), 
to_sfixed(1636730887.0/4294967296.0,1,-nbitq), 
to_sfixed(840008565.0/4294967296.0,1,-nbitq), 
to_sfixed(-980076121.0/4294967296.0,1,-nbitq), 
to_sfixed(111113243.0/4294967296.0,1,-nbitq), 
to_sfixed(762629759.0/4294967296.0,1,-nbitq), 
to_sfixed(314641984.0/4294967296.0,1,-nbitq), 
to_sfixed(-358255598.0/4294967296.0,1,-nbitq), 
to_sfixed(-73237526.0/4294967296.0,1,-nbitq), 
to_sfixed(-435137794.0/4294967296.0,1,-nbitq), 
to_sfixed(780530391.0/4294967296.0,1,-nbitq), 
to_sfixed(656073014.0/4294967296.0,1,-nbitq), 
to_sfixed(563494827.0/4294967296.0,1,-nbitq), 
to_sfixed(206834799.0/4294967296.0,1,-nbitq), 
to_sfixed(-869794121.0/4294967296.0,1,-nbitq), 
to_sfixed(-347131861.0/4294967296.0,1,-nbitq), 
to_sfixed(239455263.0/4294967296.0,1,-nbitq), 
to_sfixed(-1335704792.0/4294967296.0,1,-nbitq), 
to_sfixed(116379879.0/4294967296.0,1,-nbitq), 
to_sfixed(21859232.0/4294967296.0,1,-nbitq), 
to_sfixed(-142536776.0/4294967296.0,1,-nbitq), 
to_sfixed(108912466.0/4294967296.0,1,-nbitq), 
to_sfixed(406020351.0/4294967296.0,1,-nbitq), 
to_sfixed(-508692589.0/4294967296.0,1,-nbitq), 
to_sfixed(1497312691.0/4294967296.0,1,-nbitq), 
to_sfixed(-39470189.0/4294967296.0,1,-nbitq), 
to_sfixed(732725006.0/4294967296.0,1,-nbitq), 
to_sfixed(220052334.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-453924839.0/4294967296.0,1,-nbitq), 
to_sfixed(751896160.0/4294967296.0,1,-nbitq), 
to_sfixed(-550844544.0/4294967296.0,1,-nbitq), 
to_sfixed(-870270694.0/4294967296.0,1,-nbitq), 
to_sfixed(-434497700.0/4294967296.0,1,-nbitq), 
to_sfixed(-690448384.0/4294967296.0,1,-nbitq), 
to_sfixed(-2297945.0/4294967296.0,1,-nbitq), 
to_sfixed(-505185218.0/4294967296.0,1,-nbitq), 
to_sfixed(-23178569.0/4294967296.0,1,-nbitq), 
to_sfixed(177214520.0/4294967296.0,1,-nbitq), 
to_sfixed(213321156.0/4294967296.0,1,-nbitq), 
to_sfixed(-803345423.0/4294967296.0,1,-nbitq), 
to_sfixed(867829454.0/4294967296.0,1,-nbitq), 
to_sfixed(590905911.0/4294967296.0,1,-nbitq), 
to_sfixed(-153614472.0/4294967296.0,1,-nbitq), 
to_sfixed(-280684524.0/4294967296.0,1,-nbitq), 
to_sfixed(55480902.0/4294967296.0,1,-nbitq), 
to_sfixed(218741987.0/4294967296.0,1,-nbitq), 
to_sfixed(324281468.0/4294967296.0,1,-nbitq), 
to_sfixed(751800826.0/4294967296.0,1,-nbitq), 
to_sfixed(-62398211.0/4294967296.0,1,-nbitq), 
to_sfixed(-94735810.0/4294967296.0,1,-nbitq), 
to_sfixed(773149934.0/4294967296.0,1,-nbitq), 
to_sfixed(-358988020.0/4294967296.0,1,-nbitq), 
to_sfixed(205659344.0/4294967296.0,1,-nbitq), 
to_sfixed(-84105682.0/4294967296.0,1,-nbitq), 
to_sfixed(195586663.0/4294967296.0,1,-nbitq), 
to_sfixed(-111738935.0/4294967296.0,1,-nbitq), 
to_sfixed(437671709.0/4294967296.0,1,-nbitq), 
to_sfixed(-843575012.0/4294967296.0,1,-nbitq), 
to_sfixed(-279148157.0/4294967296.0,1,-nbitq), 
to_sfixed(480460327.0/4294967296.0,1,-nbitq), 
to_sfixed(-335468586.0/4294967296.0,1,-nbitq), 
to_sfixed(224595642.0/4294967296.0,1,-nbitq), 
to_sfixed(-100557938.0/4294967296.0,1,-nbitq), 
to_sfixed(934983058.0/4294967296.0,1,-nbitq), 
to_sfixed(187323999.0/4294967296.0,1,-nbitq), 
to_sfixed(-335369362.0/4294967296.0,1,-nbitq), 
to_sfixed(-5217410.0/4294967296.0,1,-nbitq), 
to_sfixed(216402075.0/4294967296.0,1,-nbitq), 
to_sfixed(331049896.0/4294967296.0,1,-nbitq), 
to_sfixed(872775337.0/4294967296.0,1,-nbitq), 
to_sfixed(20073242.0/4294967296.0,1,-nbitq), 
to_sfixed(235245464.0/4294967296.0,1,-nbitq), 
to_sfixed(-71245935.0/4294967296.0,1,-nbitq), 
to_sfixed(-488095011.0/4294967296.0,1,-nbitq), 
to_sfixed(-15485248.0/4294967296.0,1,-nbitq), 
to_sfixed(-684531042.0/4294967296.0,1,-nbitq), 
to_sfixed(212962521.0/4294967296.0,1,-nbitq), 
to_sfixed(312618512.0/4294967296.0,1,-nbitq), 
to_sfixed(-152461171.0/4294967296.0,1,-nbitq), 
to_sfixed(-166111350.0/4294967296.0,1,-nbitq), 
to_sfixed(-268493113.0/4294967296.0,1,-nbitq), 
to_sfixed(1250154702.0/4294967296.0,1,-nbitq), 
to_sfixed(797217351.0/4294967296.0,1,-nbitq), 
to_sfixed(-1120287937.0/4294967296.0,1,-nbitq), 
to_sfixed(-246842960.0/4294967296.0,1,-nbitq), 
to_sfixed(464653197.0/4294967296.0,1,-nbitq), 
to_sfixed(275499051.0/4294967296.0,1,-nbitq), 
to_sfixed(-89272396.0/4294967296.0,1,-nbitq), 
to_sfixed(-287378890.0/4294967296.0,1,-nbitq), 
to_sfixed(-840433167.0/4294967296.0,1,-nbitq), 
to_sfixed(443850855.0/4294967296.0,1,-nbitq), 
to_sfixed(1258521335.0/4294967296.0,1,-nbitq), 
to_sfixed(-309063927.0/4294967296.0,1,-nbitq), 
to_sfixed(-146454688.0/4294967296.0,1,-nbitq), 
to_sfixed(-967498114.0/4294967296.0,1,-nbitq), 
to_sfixed(-483356673.0/4294967296.0,1,-nbitq), 
to_sfixed(-375062419.0/4294967296.0,1,-nbitq), 
to_sfixed(-426200933.0/4294967296.0,1,-nbitq), 
to_sfixed(480500978.0/4294967296.0,1,-nbitq), 
to_sfixed(-119699542.0/4294967296.0,1,-nbitq), 
to_sfixed(-529933109.0/4294967296.0,1,-nbitq), 
to_sfixed(-11369803.0/4294967296.0,1,-nbitq), 
to_sfixed(27767866.0/4294967296.0,1,-nbitq), 
to_sfixed(-366777561.0/4294967296.0,1,-nbitq), 
to_sfixed(1114774156.0/4294967296.0,1,-nbitq), 
to_sfixed(592170500.0/4294967296.0,1,-nbitq), 
to_sfixed(-577658066.0/4294967296.0,1,-nbitq), 
to_sfixed(189842636.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(62115459.0/4294967296.0,1,-nbitq), 
to_sfixed(733413852.0/4294967296.0,1,-nbitq), 
to_sfixed(-344686213.0/4294967296.0,1,-nbitq), 
to_sfixed(-330293431.0/4294967296.0,1,-nbitq), 
to_sfixed(481772610.0/4294967296.0,1,-nbitq), 
to_sfixed(-383152102.0/4294967296.0,1,-nbitq), 
to_sfixed(-380746088.0/4294967296.0,1,-nbitq), 
to_sfixed(-209520258.0/4294967296.0,1,-nbitq), 
to_sfixed(243774235.0/4294967296.0,1,-nbitq), 
to_sfixed(-118097080.0/4294967296.0,1,-nbitq), 
to_sfixed(364323923.0/4294967296.0,1,-nbitq), 
to_sfixed(-774041805.0/4294967296.0,1,-nbitq), 
to_sfixed(358396985.0/4294967296.0,1,-nbitq), 
to_sfixed(713473952.0/4294967296.0,1,-nbitq), 
to_sfixed(-88672451.0/4294967296.0,1,-nbitq), 
to_sfixed(-35799777.0/4294967296.0,1,-nbitq), 
to_sfixed(-102269579.0/4294967296.0,1,-nbitq), 
to_sfixed(138472476.0/4294967296.0,1,-nbitq), 
to_sfixed(1080713237.0/4294967296.0,1,-nbitq), 
to_sfixed(451450964.0/4294967296.0,1,-nbitq), 
to_sfixed(-240098940.0/4294967296.0,1,-nbitq), 
to_sfixed(-146745297.0/4294967296.0,1,-nbitq), 
to_sfixed(555706482.0/4294967296.0,1,-nbitq), 
to_sfixed(-567808263.0/4294967296.0,1,-nbitq), 
to_sfixed(184676799.0/4294967296.0,1,-nbitq), 
to_sfixed(653895049.0/4294967296.0,1,-nbitq), 
to_sfixed(-180410940.0/4294967296.0,1,-nbitq), 
to_sfixed(-143753028.0/4294967296.0,1,-nbitq), 
to_sfixed(109194068.0/4294967296.0,1,-nbitq), 
to_sfixed(-69733785.0/4294967296.0,1,-nbitq), 
to_sfixed(159227233.0/4294967296.0,1,-nbitq), 
to_sfixed(60131267.0/4294967296.0,1,-nbitq), 
to_sfixed(-461894457.0/4294967296.0,1,-nbitq), 
to_sfixed(-142067663.0/4294967296.0,1,-nbitq), 
to_sfixed(241074159.0/4294967296.0,1,-nbitq), 
to_sfixed(523494082.0/4294967296.0,1,-nbitq), 
to_sfixed(35989380.0/4294967296.0,1,-nbitq), 
to_sfixed(350751399.0/4294967296.0,1,-nbitq), 
to_sfixed(-14208336.0/4294967296.0,1,-nbitq), 
to_sfixed(58063391.0/4294967296.0,1,-nbitq), 
to_sfixed(304630488.0/4294967296.0,1,-nbitq), 
to_sfixed(551561865.0/4294967296.0,1,-nbitq), 
to_sfixed(303005556.0/4294967296.0,1,-nbitq), 
to_sfixed(397327420.0/4294967296.0,1,-nbitq), 
to_sfixed(-670067149.0/4294967296.0,1,-nbitq), 
to_sfixed(-463467795.0/4294967296.0,1,-nbitq), 
to_sfixed(-383314615.0/4294967296.0,1,-nbitq), 
to_sfixed(-1170978303.0/4294967296.0,1,-nbitq), 
to_sfixed(220988776.0/4294967296.0,1,-nbitq), 
to_sfixed(697231683.0/4294967296.0,1,-nbitq), 
to_sfixed(24240387.0/4294967296.0,1,-nbitq), 
to_sfixed(122990988.0/4294967296.0,1,-nbitq), 
to_sfixed(347295818.0/4294967296.0,1,-nbitq), 
to_sfixed(905093446.0/4294967296.0,1,-nbitq), 
to_sfixed(700260683.0/4294967296.0,1,-nbitq), 
to_sfixed(-593266618.0/4294967296.0,1,-nbitq), 
to_sfixed(104205658.0/4294967296.0,1,-nbitq), 
to_sfixed(412205831.0/4294967296.0,1,-nbitq), 
to_sfixed(-248765139.0/4294967296.0,1,-nbitq), 
to_sfixed(386108185.0/4294967296.0,1,-nbitq), 
to_sfixed(382153802.0/4294967296.0,1,-nbitq), 
to_sfixed(-757606926.0/4294967296.0,1,-nbitq), 
to_sfixed(-193512871.0/4294967296.0,1,-nbitq), 
to_sfixed(243920450.0/4294967296.0,1,-nbitq), 
to_sfixed(233780766.0/4294967296.0,1,-nbitq), 
to_sfixed(-19878345.0/4294967296.0,1,-nbitq), 
to_sfixed(-880464602.0/4294967296.0,1,-nbitq), 
to_sfixed(-416407266.0/4294967296.0,1,-nbitq), 
to_sfixed(345973664.0/4294967296.0,1,-nbitq), 
to_sfixed(-698405507.0/4294967296.0,1,-nbitq), 
to_sfixed(1199370.0/4294967296.0,1,-nbitq), 
to_sfixed(401601724.0/4294967296.0,1,-nbitq), 
to_sfixed(-443661213.0/4294967296.0,1,-nbitq), 
to_sfixed(-12185629.0/4294967296.0,1,-nbitq), 
to_sfixed(100000675.0/4294967296.0,1,-nbitq), 
to_sfixed(191275360.0/4294967296.0,1,-nbitq), 
to_sfixed(-124807700.0/4294967296.0,1,-nbitq), 
to_sfixed(632450016.0/4294967296.0,1,-nbitq), 
to_sfixed(-816491734.0/4294967296.0,1,-nbitq), 
to_sfixed(384862210.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(55624265.0/4294967296.0,1,-nbitq), 
to_sfixed(503486137.0/4294967296.0,1,-nbitq), 
to_sfixed(-931077632.0/4294967296.0,1,-nbitq), 
to_sfixed(-106651558.0/4294967296.0,1,-nbitq), 
to_sfixed(1253087277.0/4294967296.0,1,-nbitq), 
to_sfixed(1125167088.0/4294967296.0,1,-nbitq), 
to_sfixed(-189839004.0/4294967296.0,1,-nbitq), 
to_sfixed(-215063083.0/4294967296.0,1,-nbitq), 
to_sfixed(288792811.0/4294967296.0,1,-nbitq), 
to_sfixed(73655940.0/4294967296.0,1,-nbitq), 
to_sfixed(-438216467.0/4294967296.0,1,-nbitq), 
to_sfixed(-555559157.0/4294967296.0,1,-nbitq), 
to_sfixed(503899824.0/4294967296.0,1,-nbitq), 
to_sfixed(-35136556.0/4294967296.0,1,-nbitq), 
to_sfixed(266791640.0/4294967296.0,1,-nbitq), 
to_sfixed(-759611775.0/4294967296.0,1,-nbitq), 
to_sfixed(59628329.0/4294967296.0,1,-nbitq), 
to_sfixed(66030551.0/4294967296.0,1,-nbitq), 
to_sfixed(-109978013.0/4294967296.0,1,-nbitq), 
to_sfixed(450495688.0/4294967296.0,1,-nbitq), 
to_sfixed(219675596.0/4294967296.0,1,-nbitq), 
to_sfixed(235305585.0/4294967296.0,1,-nbitq), 
to_sfixed(181537890.0/4294967296.0,1,-nbitq), 
to_sfixed(-314204678.0/4294967296.0,1,-nbitq), 
to_sfixed(30715366.0/4294967296.0,1,-nbitq), 
to_sfixed(1253908610.0/4294967296.0,1,-nbitq), 
to_sfixed(-87045322.0/4294967296.0,1,-nbitq), 
to_sfixed(334548247.0/4294967296.0,1,-nbitq), 
to_sfixed(-425759388.0/4294967296.0,1,-nbitq), 
to_sfixed(-1073827.0/4294967296.0,1,-nbitq), 
to_sfixed(-317380486.0/4294967296.0,1,-nbitq), 
to_sfixed(-18519397.0/4294967296.0,1,-nbitq), 
to_sfixed(-106510546.0/4294967296.0,1,-nbitq), 
to_sfixed(-832827188.0/4294967296.0,1,-nbitq), 
to_sfixed(485139982.0/4294967296.0,1,-nbitq), 
to_sfixed(775066244.0/4294967296.0,1,-nbitq), 
to_sfixed(-64336454.0/4294967296.0,1,-nbitq), 
to_sfixed(82486888.0/4294967296.0,1,-nbitq), 
to_sfixed(399150055.0/4294967296.0,1,-nbitq), 
to_sfixed(-60302440.0/4294967296.0,1,-nbitq), 
to_sfixed(582962432.0/4294967296.0,1,-nbitq), 
to_sfixed(226286473.0/4294967296.0,1,-nbitq), 
to_sfixed(90770361.0/4294967296.0,1,-nbitq), 
to_sfixed(-107045969.0/4294967296.0,1,-nbitq), 
to_sfixed(23183680.0/4294967296.0,1,-nbitq), 
to_sfixed(-432220398.0/4294967296.0,1,-nbitq), 
to_sfixed(360983177.0/4294967296.0,1,-nbitq), 
to_sfixed(-657738328.0/4294967296.0,1,-nbitq), 
to_sfixed(-152367167.0/4294967296.0,1,-nbitq), 
to_sfixed(-207944841.0/4294967296.0,1,-nbitq), 
to_sfixed(147935450.0/4294967296.0,1,-nbitq), 
to_sfixed(-363209188.0/4294967296.0,1,-nbitq), 
to_sfixed(289026533.0/4294967296.0,1,-nbitq), 
to_sfixed(681065205.0/4294967296.0,1,-nbitq), 
to_sfixed(231085785.0/4294967296.0,1,-nbitq), 
to_sfixed(-195960643.0/4294967296.0,1,-nbitq), 
to_sfixed(-313390585.0/4294967296.0,1,-nbitq), 
to_sfixed(354862853.0/4294967296.0,1,-nbitq), 
to_sfixed(-74877758.0/4294967296.0,1,-nbitq), 
to_sfixed(136869725.0/4294967296.0,1,-nbitq), 
to_sfixed(37416248.0/4294967296.0,1,-nbitq), 
to_sfixed(-1394346306.0/4294967296.0,1,-nbitq), 
to_sfixed(34527888.0/4294967296.0,1,-nbitq), 
to_sfixed(522214225.0/4294967296.0,1,-nbitq), 
to_sfixed(226206004.0/4294967296.0,1,-nbitq), 
to_sfixed(-9233034.0/4294967296.0,1,-nbitq), 
to_sfixed(-681551539.0/4294967296.0,1,-nbitq), 
to_sfixed(-492252070.0/4294967296.0,1,-nbitq), 
to_sfixed(106581983.0/4294967296.0,1,-nbitq), 
to_sfixed(-389169049.0/4294967296.0,1,-nbitq), 
to_sfixed(394808752.0/4294967296.0,1,-nbitq), 
to_sfixed(217199980.0/4294967296.0,1,-nbitq), 
to_sfixed(-639736445.0/4294967296.0,1,-nbitq), 
to_sfixed(261612033.0/4294967296.0,1,-nbitq), 
to_sfixed(-72393431.0/4294967296.0,1,-nbitq), 
to_sfixed(329003144.0/4294967296.0,1,-nbitq), 
to_sfixed(-262181607.0/4294967296.0,1,-nbitq), 
to_sfixed(-9524916.0/4294967296.0,1,-nbitq), 
to_sfixed(-366671404.0/4294967296.0,1,-nbitq), 
to_sfixed(-199170901.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(198882965.0/4294967296.0,1,-nbitq), 
to_sfixed(877358905.0/4294967296.0,1,-nbitq), 
to_sfixed(-285348404.0/4294967296.0,1,-nbitq), 
to_sfixed(-794521248.0/4294967296.0,1,-nbitq), 
to_sfixed(880617734.0/4294967296.0,1,-nbitq), 
to_sfixed(312874799.0/4294967296.0,1,-nbitq), 
to_sfixed(39505134.0/4294967296.0,1,-nbitq), 
to_sfixed(-137948318.0/4294967296.0,1,-nbitq), 
to_sfixed(-22475753.0/4294967296.0,1,-nbitq), 
to_sfixed(-73219179.0/4294967296.0,1,-nbitq), 
to_sfixed(82146041.0/4294967296.0,1,-nbitq), 
to_sfixed(-192815823.0/4294967296.0,1,-nbitq), 
to_sfixed(-65844264.0/4294967296.0,1,-nbitq), 
to_sfixed(-447037998.0/4294967296.0,1,-nbitq), 
to_sfixed(155809454.0/4294967296.0,1,-nbitq), 
to_sfixed(-865142428.0/4294967296.0,1,-nbitq), 
to_sfixed(-98439203.0/4294967296.0,1,-nbitq), 
to_sfixed(340610629.0/4294967296.0,1,-nbitq), 
to_sfixed(-32695382.0/4294967296.0,1,-nbitq), 
to_sfixed(-46387423.0/4294967296.0,1,-nbitq), 
to_sfixed(226729278.0/4294967296.0,1,-nbitq), 
to_sfixed(-345310439.0/4294967296.0,1,-nbitq), 
to_sfixed(-17605691.0/4294967296.0,1,-nbitq), 
to_sfixed(-529689059.0/4294967296.0,1,-nbitq), 
to_sfixed(282082441.0/4294967296.0,1,-nbitq), 
to_sfixed(481495465.0/4294967296.0,1,-nbitq), 
to_sfixed(-204863570.0/4294967296.0,1,-nbitq), 
to_sfixed(575986135.0/4294967296.0,1,-nbitq), 
to_sfixed(-451108492.0/4294967296.0,1,-nbitq), 
to_sfixed(-454651295.0/4294967296.0,1,-nbitq), 
to_sfixed(-37280319.0/4294967296.0,1,-nbitq), 
to_sfixed(218674969.0/4294967296.0,1,-nbitq), 
to_sfixed(-192464568.0/4294967296.0,1,-nbitq), 
to_sfixed(-724662845.0/4294967296.0,1,-nbitq), 
to_sfixed(28431496.0/4294967296.0,1,-nbitq), 
to_sfixed(126292113.0/4294967296.0,1,-nbitq), 
to_sfixed(-163554633.0/4294967296.0,1,-nbitq), 
to_sfixed(-283737252.0/4294967296.0,1,-nbitq), 
to_sfixed(-7222949.0/4294967296.0,1,-nbitq), 
to_sfixed(275152303.0/4294967296.0,1,-nbitq), 
to_sfixed(466477224.0/4294967296.0,1,-nbitq), 
to_sfixed(-573679761.0/4294967296.0,1,-nbitq), 
to_sfixed(650497917.0/4294967296.0,1,-nbitq), 
to_sfixed(-174338051.0/4294967296.0,1,-nbitq), 
to_sfixed(70034505.0/4294967296.0,1,-nbitq), 
to_sfixed(-123185140.0/4294967296.0,1,-nbitq), 
to_sfixed(253680137.0/4294967296.0,1,-nbitq), 
to_sfixed(-548462712.0/4294967296.0,1,-nbitq), 
to_sfixed(-283768546.0/4294967296.0,1,-nbitq), 
to_sfixed(-87953955.0/4294967296.0,1,-nbitq), 
to_sfixed(72974153.0/4294967296.0,1,-nbitq), 
to_sfixed(-261029927.0/4294967296.0,1,-nbitq), 
to_sfixed(-597176407.0/4294967296.0,1,-nbitq), 
to_sfixed(581417946.0/4294967296.0,1,-nbitq), 
to_sfixed(-201172403.0/4294967296.0,1,-nbitq), 
to_sfixed(-296017896.0/4294967296.0,1,-nbitq), 
to_sfixed(-61247957.0/4294967296.0,1,-nbitq), 
to_sfixed(176278214.0/4294967296.0,1,-nbitq), 
to_sfixed(-6797771.0/4294967296.0,1,-nbitq), 
to_sfixed(432062615.0/4294967296.0,1,-nbitq), 
to_sfixed(269482046.0/4294967296.0,1,-nbitq), 
to_sfixed(-670372749.0/4294967296.0,1,-nbitq), 
to_sfixed(56308388.0/4294967296.0,1,-nbitq), 
to_sfixed(298702237.0/4294967296.0,1,-nbitq), 
to_sfixed(51356037.0/4294967296.0,1,-nbitq), 
to_sfixed(-225839766.0/4294967296.0,1,-nbitq), 
to_sfixed(-612915781.0/4294967296.0,1,-nbitq), 
to_sfixed(-749231810.0/4294967296.0,1,-nbitq), 
to_sfixed(234460342.0/4294967296.0,1,-nbitq), 
to_sfixed(-496647645.0/4294967296.0,1,-nbitq), 
to_sfixed(308817098.0/4294967296.0,1,-nbitq), 
to_sfixed(79516315.0/4294967296.0,1,-nbitq), 
to_sfixed(322358718.0/4294967296.0,1,-nbitq), 
to_sfixed(145617276.0/4294967296.0,1,-nbitq), 
to_sfixed(-227636599.0/4294967296.0,1,-nbitq), 
to_sfixed(474481752.0/4294967296.0,1,-nbitq), 
to_sfixed(-981023205.0/4294967296.0,1,-nbitq), 
to_sfixed(-471419600.0/4294967296.0,1,-nbitq), 
to_sfixed(-401180487.0/4294967296.0,1,-nbitq), 
to_sfixed(-262798681.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-281627066.0/4294967296.0,1,-nbitq), 
to_sfixed(1280029978.0/4294967296.0,1,-nbitq), 
to_sfixed(133289634.0/4294967296.0,1,-nbitq), 
to_sfixed(-227246715.0/4294967296.0,1,-nbitq), 
to_sfixed(337857852.0/4294967296.0,1,-nbitq), 
to_sfixed(247298295.0/4294967296.0,1,-nbitq), 
to_sfixed(-415118584.0/4294967296.0,1,-nbitq), 
to_sfixed(332673038.0/4294967296.0,1,-nbitq), 
to_sfixed(-489598562.0/4294967296.0,1,-nbitq), 
to_sfixed(144390518.0/4294967296.0,1,-nbitq), 
to_sfixed(823384387.0/4294967296.0,1,-nbitq), 
to_sfixed(178813598.0/4294967296.0,1,-nbitq), 
to_sfixed(860745184.0/4294967296.0,1,-nbitq), 
to_sfixed(-619081211.0/4294967296.0,1,-nbitq), 
to_sfixed(-68042184.0/4294967296.0,1,-nbitq), 
to_sfixed(-342471671.0/4294967296.0,1,-nbitq), 
to_sfixed(7187470.0/4294967296.0,1,-nbitq), 
to_sfixed(-160170068.0/4294967296.0,1,-nbitq), 
to_sfixed(408458707.0/4294967296.0,1,-nbitq), 
to_sfixed(384568627.0/4294967296.0,1,-nbitq), 
to_sfixed(145144774.0/4294967296.0,1,-nbitq), 
to_sfixed(123400541.0/4294967296.0,1,-nbitq), 
to_sfixed(-300289548.0/4294967296.0,1,-nbitq), 
to_sfixed(-222853501.0/4294967296.0,1,-nbitq), 
to_sfixed(279091955.0/4294967296.0,1,-nbitq), 
to_sfixed(551597032.0/4294967296.0,1,-nbitq), 
to_sfixed(-360704904.0/4294967296.0,1,-nbitq), 
to_sfixed(773594523.0/4294967296.0,1,-nbitq), 
to_sfixed(-443542497.0/4294967296.0,1,-nbitq), 
to_sfixed(-177978903.0/4294967296.0,1,-nbitq), 
to_sfixed(288813319.0/4294967296.0,1,-nbitq), 
to_sfixed(19422251.0/4294967296.0,1,-nbitq), 
to_sfixed(437428445.0/4294967296.0,1,-nbitq), 
to_sfixed(39095994.0/4294967296.0,1,-nbitq), 
to_sfixed(1399731.0/4294967296.0,1,-nbitq), 
to_sfixed(105087432.0/4294967296.0,1,-nbitq), 
to_sfixed(-86298066.0/4294967296.0,1,-nbitq), 
to_sfixed(-1127539811.0/4294967296.0,1,-nbitq), 
to_sfixed(-105951556.0/4294967296.0,1,-nbitq), 
to_sfixed(51534746.0/4294967296.0,1,-nbitq), 
to_sfixed(286593845.0/4294967296.0,1,-nbitq), 
to_sfixed(164957708.0/4294967296.0,1,-nbitq), 
to_sfixed(-178698093.0/4294967296.0,1,-nbitq), 
to_sfixed(-282212238.0/4294967296.0,1,-nbitq), 
to_sfixed(135277145.0/4294967296.0,1,-nbitq), 
to_sfixed(-36711515.0/4294967296.0,1,-nbitq), 
to_sfixed(-330624776.0/4294967296.0,1,-nbitq), 
to_sfixed(-171458066.0/4294967296.0,1,-nbitq), 
to_sfixed(-273087464.0/4294967296.0,1,-nbitq), 
to_sfixed(-414488154.0/4294967296.0,1,-nbitq), 
to_sfixed(-261530072.0/4294967296.0,1,-nbitq), 
to_sfixed(-760839749.0/4294967296.0,1,-nbitq), 
to_sfixed(-179534641.0/4294967296.0,1,-nbitq), 
to_sfixed(619299898.0/4294967296.0,1,-nbitq), 
to_sfixed(-459444444.0/4294967296.0,1,-nbitq), 
to_sfixed(-661359323.0/4294967296.0,1,-nbitq), 
to_sfixed(-50714590.0/4294967296.0,1,-nbitq), 
to_sfixed(-404588543.0/4294967296.0,1,-nbitq), 
to_sfixed(73341070.0/4294967296.0,1,-nbitq), 
to_sfixed(164909888.0/4294967296.0,1,-nbitq), 
to_sfixed(-843036.0/4294967296.0,1,-nbitq), 
to_sfixed(-678852662.0/4294967296.0,1,-nbitq), 
to_sfixed(433639241.0/4294967296.0,1,-nbitq), 
to_sfixed(42182790.0/4294967296.0,1,-nbitq), 
to_sfixed(-200964520.0/4294967296.0,1,-nbitq), 
to_sfixed(-365073031.0/4294967296.0,1,-nbitq), 
to_sfixed(-954462157.0/4294967296.0,1,-nbitq), 
to_sfixed(-205883543.0/4294967296.0,1,-nbitq), 
to_sfixed(371365797.0/4294967296.0,1,-nbitq), 
to_sfixed(-550304608.0/4294967296.0,1,-nbitq), 
to_sfixed(699891357.0/4294967296.0,1,-nbitq), 
to_sfixed(-383061733.0/4294967296.0,1,-nbitq), 
to_sfixed(-120991182.0/4294967296.0,1,-nbitq), 
to_sfixed(-341203316.0/4294967296.0,1,-nbitq), 
to_sfixed(150485371.0/4294967296.0,1,-nbitq), 
to_sfixed(-144495163.0/4294967296.0,1,-nbitq), 
to_sfixed(-199092658.0/4294967296.0,1,-nbitq), 
to_sfixed(-371663742.0/4294967296.0,1,-nbitq), 
to_sfixed(-120495555.0/4294967296.0,1,-nbitq), 
to_sfixed(40357246.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(175353440.0/4294967296.0,1,-nbitq), 
to_sfixed(127839433.0/4294967296.0,1,-nbitq), 
to_sfixed(-322201001.0/4294967296.0,1,-nbitq), 
to_sfixed(518108840.0/4294967296.0,1,-nbitq), 
to_sfixed(319409426.0/4294967296.0,1,-nbitq), 
to_sfixed(212125142.0/4294967296.0,1,-nbitq), 
to_sfixed(-8388599.0/4294967296.0,1,-nbitq), 
to_sfixed(251238242.0/4294967296.0,1,-nbitq), 
to_sfixed(-604284743.0/4294967296.0,1,-nbitq), 
to_sfixed(326865277.0/4294967296.0,1,-nbitq), 
to_sfixed(1178442320.0/4294967296.0,1,-nbitq), 
to_sfixed(834418007.0/4294967296.0,1,-nbitq), 
to_sfixed(835415704.0/4294967296.0,1,-nbitq), 
to_sfixed(-378812765.0/4294967296.0,1,-nbitq), 
to_sfixed(161737277.0/4294967296.0,1,-nbitq), 
to_sfixed(-476133763.0/4294967296.0,1,-nbitq), 
to_sfixed(-359030778.0/4294967296.0,1,-nbitq), 
to_sfixed(112080458.0/4294967296.0,1,-nbitq), 
to_sfixed(378089231.0/4294967296.0,1,-nbitq), 
to_sfixed(136796344.0/4294967296.0,1,-nbitq), 
to_sfixed(273817903.0/4294967296.0,1,-nbitq), 
to_sfixed(617571625.0/4294967296.0,1,-nbitq), 
to_sfixed(68990495.0/4294967296.0,1,-nbitq), 
to_sfixed(-397935548.0/4294967296.0,1,-nbitq), 
to_sfixed(-243292807.0/4294967296.0,1,-nbitq), 
to_sfixed(762521859.0/4294967296.0,1,-nbitq), 
to_sfixed(-824857350.0/4294967296.0,1,-nbitq), 
to_sfixed(-45891457.0/4294967296.0,1,-nbitq), 
to_sfixed(453273889.0/4294967296.0,1,-nbitq), 
to_sfixed(-680821028.0/4294967296.0,1,-nbitq), 
to_sfixed(166838075.0/4294967296.0,1,-nbitq), 
to_sfixed(29416957.0/4294967296.0,1,-nbitq), 
to_sfixed(431276380.0/4294967296.0,1,-nbitq), 
to_sfixed(-385192.0/4294967296.0,1,-nbitq), 
to_sfixed(188855384.0/4294967296.0,1,-nbitq), 
to_sfixed(-258596014.0/4294967296.0,1,-nbitq), 
to_sfixed(-524531225.0/4294967296.0,1,-nbitq), 
to_sfixed(-1009718480.0/4294967296.0,1,-nbitq), 
to_sfixed(-77888480.0/4294967296.0,1,-nbitq), 
to_sfixed(123651158.0/4294967296.0,1,-nbitq), 
to_sfixed(154723817.0/4294967296.0,1,-nbitq), 
to_sfixed(82661660.0/4294967296.0,1,-nbitq), 
to_sfixed(223177969.0/4294967296.0,1,-nbitq), 
to_sfixed(-9469003.0/4294967296.0,1,-nbitq), 
to_sfixed(501539483.0/4294967296.0,1,-nbitq), 
to_sfixed(-241591128.0/4294967296.0,1,-nbitq), 
to_sfixed(-406209053.0/4294967296.0,1,-nbitq), 
to_sfixed(-80805413.0/4294967296.0,1,-nbitq), 
to_sfixed(-370910921.0/4294967296.0,1,-nbitq), 
to_sfixed(-278373105.0/4294967296.0,1,-nbitq), 
to_sfixed(-356410537.0/4294967296.0,1,-nbitq), 
to_sfixed(78945304.0/4294967296.0,1,-nbitq), 
to_sfixed(47277708.0/4294967296.0,1,-nbitq), 
to_sfixed(118537381.0/4294967296.0,1,-nbitq), 
to_sfixed(-245464396.0/4294967296.0,1,-nbitq), 
to_sfixed(45448688.0/4294967296.0,1,-nbitq), 
to_sfixed(-422418958.0/4294967296.0,1,-nbitq), 
to_sfixed(-25863360.0/4294967296.0,1,-nbitq), 
to_sfixed(-145845812.0/4294967296.0,1,-nbitq), 
to_sfixed(129126151.0/4294967296.0,1,-nbitq), 
to_sfixed(-70843452.0/4294967296.0,1,-nbitq), 
to_sfixed(-688119515.0/4294967296.0,1,-nbitq), 
to_sfixed(-82039970.0/4294967296.0,1,-nbitq), 
to_sfixed(-334388573.0/4294967296.0,1,-nbitq), 
to_sfixed(-203000318.0/4294967296.0,1,-nbitq), 
to_sfixed(-105889848.0/4294967296.0,1,-nbitq), 
to_sfixed(-753434383.0/4294967296.0,1,-nbitq), 
to_sfixed(-602284254.0/4294967296.0,1,-nbitq), 
to_sfixed(174103752.0/4294967296.0,1,-nbitq), 
to_sfixed(-196572711.0/4294967296.0,1,-nbitq), 
to_sfixed(168405173.0/4294967296.0,1,-nbitq), 
to_sfixed(341495849.0/4294967296.0,1,-nbitq), 
to_sfixed(-81665640.0/4294967296.0,1,-nbitq), 
to_sfixed(-123473131.0/4294967296.0,1,-nbitq), 
to_sfixed(497296263.0/4294967296.0,1,-nbitq), 
to_sfixed(38319434.0/4294967296.0,1,-nbitq), 
to_sfixed(-467736917.0/4294967296.0,1,-nbitq), 
to_sfixed(100696176.0/4294967296.0,1,-nbitq), 
to_sfixed(-646316308.0/4294967296.0,1,-nbitq), 
to_sfixed(-285158123.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(228168011.0/4294967296.0,1,-nbitq), 
to_sfixed(356923184.0/4294967296.0,1,-nbitq), 
to_sfixed(-412640433.0/4294967296.0,1,-nbitq), 
to_sfixed(187642558.0/4294967296.0,1,-nbitq), 
to_sfixed(-95730170.0/4294967296.0,1,-nbitq), 
to_sfixed(-25298493.0/4294967296.0,1,-nbitq), 
to_sfixed(-215188461.0/4294967296.0,1,-nbitq), 
to_sfixed(323995675.0/4294967296.0,1,-nbitq), 
to_sfixed(115336558.0/4294967296.0,1,-nbitq), 
to_sfixed(369744959.0/4294967296.0,1,-nbitq), 
to_sfixed(556680733.0/4294967296.0,1,-nbitq), 
to_sfixed(377532286.0/4294967296.0,1,-nbitq), 
to_sfixed(260684876.0/4294967296.0,1,-nbitq), 
to_sfixed(72972632.0/4294967296.0,1,-nbitq), 
to_sfixed(-77290574.0/4294967296.0,1,-nbitq), 
to_sfixed(-301570002.0/4294967296.0,1,-nbitq), 
to_sfixed(365602186.0/4294967296.0,1,-nbitq), 
to_sfixed(-172875527.0/4294967296.0,1,-nbitq), 
to_sfixed(133296418.0/4294967296.0,1,-nbitq), 
to_sfixed(-43284686.0/4294967296.0,1,-nbitq), 
to_sfixed(-307567930.0/4294967296.0,1,-nbitq), 
to_sfixed(-191100297.0/4294967296.0,1,-nbitq), 
to_sfixed(91328922.0/4294967296.0,1,-nbitq), 
to_sfixed(-57579732.0/4294967296.0,1,-nbitq), 
to_sfixed(286538242.0/4294967296.0,1,-nbitq), 
to_sfixed(486459548.0/4294967296.0,1,-nbitq), 
to_sfixed(11634353.0/4294967296.0,1,-nbitq), 
to_sfixed(51003129.0/4294967296.0,1,-nbitq), 
to_sfixed(75639927.0/4294967296.0,1,-nbitq), 
to_sfixed(-222728597.0/4294967296.0,1,-nbitq), 
to_sfixed(-294636200.0/4294967296.0,1,-nbitq), 
to_sfixed(318769855.0/4294967296.0,1,-nbitq), 
to_sfixed(520580558.0/4294967296.0,1,-nbitq), 
to_sfixed(-47459702.0/4294967296.0,1,-nbitq), 
to_sfixed(112412668.0/4294967296.0,1,-nbitq), 
to_sfixed(220019647.0/4294967296.0,1,-nbitq), 
to_sfixed(163859747.0/4294967296.0,1,-nbitq), 
to_sfixed(-155722206.0/4294967296.0,1,-nbitq), 
to_sfixed(214126855.0/4294967296.0,1,-nbitq), 
to_sfixed(105084408.0/4294967296.0,1,-nbitq), 
to_sfixed(253776654.0/4294967296.0,1,-nbitq), 
to_sfixed(277345902.0/4294967296.0,1,-nbitq), 
to_sfixed(-377935781.0/4294967296.0,1,-nbitq), 
to_sfixed(146991183.0/4294967296.0,1,-nbitq), 
to_sfixed(74217923.0/4294967296.0,1,-nbitq), 
to_sfixed(-324239662.0/4294967296.0,1,-nbitq), 
to_sfixed(-436700410.0/4294967296.0,1,-nbitq), 
to_sfixed(191504967.0/4294967296.0,1,-nbitq), 
to_sfixed(-332906655.0/4294967296.0,1,-nbitq), 
to_sfixed(-386973472.0/4294967296.0,1,-nbitq), 
to_sfixed(-179527058.0/4294967296.0,1,-nbitq), 
to_sfixed(10347790.0/4294967296.0,1,-nbitq), 
to_sfixed(-137560299.0/4294967296.0,1,-nbitq), 
to_sfixed(-57696005.0/4294967296.0,1,-nbitq), 
to_sfixed(-175276292.0/4294967296.0,1,-nbitq), 
to_sfixed(95947644.0/4294967296.0,1,-nbitq), 
to_sfixed(-13774048.0/4294967296.0,1,-nbitq), 
to_sfixed(138093176.0/4294967296.0,1,-nbitq), 
to_sfixed(204173564.0/4294967296.0,1,-nbitq), 
to_sfixed(-52498229.0/4294967296.0,1,-nbitq), 
to_sfixed(-132732236.0/4294967296.0,1,-nbitq), 
to_sfixed(95745601.0/4294967296.0,1,-nbitq), 
to_sfixed(-167816562.0/4294967296.0,1,-nbitq), 
to_sfixed(-197082426.0/4294967296.0,1,-nbitq), 
to_sfixed(2396305.0/4294967296.0,1,-nbitq), 
to_sfixed(27450877.0/4294967296.0,1,-nbitq), 
to_sfixed(353739751.0/4294967296.0,1,-nbitq), 
to_sfixed(-140971631.0/4294967296.0,1,-nbitq), 
to_sfixed(-351897323.0/4294967296.0,1,-nbitq), 
to_sfixed(-86180474.0/4294967296.0,1,-nbitq), 
to_sfixed(255524024.0/4294967296.0,1,-nbitq), 
to_sfixed(314313783.0/4294967296.0,1,-nbitq), 
to_sfixed(100561408.0/4294967296.0,1,-nbitq), 
to_sfixed(77050552.0/4294967296.0,1,-nbitq), 
to_sfixed(-197798589.0/4294967296.0,1,-nbitq), 
to_sfixed(-464434682.0/4294967296.0,1,-nbitq), 
to_sfixed(340257986.0/4294967296.0,1,-nbitq), 
to_sfixed(-230358174.0/4294967296.0,1,-nbitq), 
to_sfixed(-453311628.0/4294967296.0,1,-nbitq), 
to_sfixed(77898817.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(157004560.0/4294967296.0,1,-nbitq), 
to_sfixed(-270183359.0/4294967296.0,1,-nbitq), 
to_sfixed(-142804435.0/4294967296.0,1,-nbitq), 
to_sfixed(13958785.0/4294967296.0,1,-nbitq), 
to_sfixed(32576739.0/4294967296.0,1,-nbitq), 
to_sfixed(-132551064.0/4294967296.0,1,-nbitq), 
to_sfixed(-98439193.0/4294967296.0,1,-nbitq), 
to_sfixed(90773454.0/4294967296.0,1,-nbitq), 
to_sfixed(151537592.0/4294967296.0,1,-nbitq), 
to_sfixed(32094260.0/4294967296.0,1,-nbitq), 
to_sfixed(-51829322.0/4294967296.0,1,-nbitq), 
to_sfixed(1524594.0/4294967296.0,1,-nbitq), 
to_sfixed(217371937.0/4294967296.0,1,-nbitq), 
to_sfixed(162069006.0/4294967296.0,1,-nbitq), 
to_sfixed(-283061266.0/4294967296.0,1,-nbitq), 
to_sfixed(-215342023.0/4294967296.0,1,-nbitq), 
to_sfixed(286967018.0/4294967296.0,1,-nbitq), 
to_sfixed(238641625.0/4294967296.0,1,-nbitq), 
to_sfixed(57684363.0/4294967296.0,1,-nbitq), 
to_sfixed(-279687873.0/4294967296.0,1,-nbitq), 
to_sfixed(-165067045.0/4294967296.0,1,-nbitq), 
to_sfixed(439214796.0/4294967296.0,1,-nbitq), 
to_sfixed(247328365.0/4294967296.0,1,-nbitq), 
to_sfixed(-123675789.0/4294967296.0,1,-nbitq), 
to_sfixed(78800407.0/4294967296.0,1,-nbitq), 
to_sfixed(600406523.0/4294967296.0,1,-nbitq), 
to_sfixed(27818737.0/4294967296.0,1,-nbitq), 
to_sfixed(-155711017.0/4294967296.0,1,-nbitq), 
to_sfixed(47316546.0/4294967296.0,1,-nbitq), 
to_sfixed(-530716795.0/4294967296.0,1,-nbitq), 
to_sfixed(56426207.0/4294967296.0,1,-nbitq), 
to_sfixed(-340022850.0/4294967296.0,1,-nbitq), 
to_sfixed(-328609302.0/4294967296.0,1,-nbitq), 
to_sfixed(-285779959.0/4294967296.0,1,-nbitq), 
to_sfixed(108129175.0/4294967296.0,1,-nbitq), 
to_sfixed(-419612811.0/4294967296.0,1,-nbitq), 
to_sfixed(67453191.0/4294967296.0,1,-nbitq), 
to_sfixed(-233892014.0/4294967296.0,1,-nbitq), 
to_sfixed(-243908893.0/4294967296.0,1,-nbitq), 
to_sfixed(461905548.0/4294967296.0,1,-nbitq), 
to_sfixed(-109149469.0/4294967296.0,1,-nbitq), 
to_sfixed(317295476.0/4294967296.0,1,-nbitq), 
to_sfixed(277781999.0/4294967296.0,1,-nbitq), 
to_sfixed(-148212615.0/4294967296.0,1,-nbitq), 
to_sfixed(132515594.0/4294967296.0,1,-nbitq), 
to_sfixed(54487296.0/4294967296.0,1,-nbitq), 
to_sfixed(-268744450.0/4294967296.0,1,-nbitq), 
to_sfixed(118492777.0/4294967296.0,1,-nbitq), 
to_sfixed(290356617.0/4294967296.0,1,-nbitq), 
to_sfixed(128832265.0/4294967296.0,1,-nbitq), 
to_sfixed(-279573909.0/4294967296.0,1,-nbitq), 
to_sfixed(196080038.0/4294967296.0,1,-nbitq), 
to_sfixed(-40923096.0/4294967296.0,1,-nbitq), 
to_sfixed(328292963.0/4294967296.0,1,-nbitq), 
to_sfixed(210374494.0/4294967296.0,1,-nbitq), 
to_sfixed(276073966.0/4294967296.0,1,-nbitq), 
to_sfixed(-87671179.0/4294967296.0,1,-nbitq), 
to_sfixed(-282575607.0/4294967296.0,1,-nbitq), 
to_sfixed(250831490.0/4294967296.0,1,-nbitq), 
to_sfixed(-172356595.0/4294967296.0,1,-nbitq), 
to_sfixed(100691456.0/4294967296.0,1,-nbitq), 
to_sfixed(375552261.0/4294967296.0,1,-nbitq), 
to_sfixed(-316389774.0/4294967296.0,1,-nbitq), 
to_sfixed(281234829.0/4294967296.0,1,-nbitq), 
to_sfixed(263540184.0/4294967296.0,1,-nbitq), 
to_sfixed(357024618.0/4294967296.0,1,-nbitq), 
to_sfixed(880167061.0/4294967296.0,1,-nbitq), 
to_sfixed(249812307.0/4294967296.0,1,-nbitq), 
to_sfixed(-12562016.0/4294967296.0,1,-nbitq), 
to_sfixed(350895465.0/4294967296.0,1,-nbitq), 
to_sfixed(-462675138.0/4294967296.0,1,-nbitq), 
to_sfixed(115972986.0/4294967296.0,1,-nbitq), 
to_sfixed(-42084263.0/4294967296.0,1,-nbitq), 
to_sfixed(143249375.0/4294967296.0,1,-nbitq), 
to_sfixed(-44880590.0/4294967296.0,1,-nbitq), 
to_sfixed(110996479.0/4294967296.0,1,-nbitq), 
to_sfixed(-54255287.0/4294967296.0,1,-nbitq), 
to_sfixed(-142912492.0/4294967296.0,1,-nbitq), 
to_sfixed(24972144.0/4294967296.0,1,-nbitq), 
to_sfixed(374154325.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-23410215.0/4294967296.0,1,-nbitq), 
to_sfixed(-485180145.0/4294967296.0,1,-nbitq), 
to_sfixed(-261832505.0/4294967296.0,1,-nbitq), 
to_sfixed(-378489196.0/4294967296.0,1,-nbitq), 
to_sfixed(-255301361.0/4294967296.0,1,-nbitq), 
to_sfixed(-157140356.0/4294967296.0,1,-nbitq), 
to_sfixed(128867669.0/4294967296.0,1,-nbitq), 
to_sfixed(358381280.0/4294967296.0,1,-nbitq), 
to_sfixed(53570236.0/4294967296.0,1,-nbitq), 
to_sfixed(227256889.0/4294967296.0,1,-nbitq), 
to_sfixed(253965286.0/4294967296.0,1,-nbitq), 
to_sfixed(62024679.0/4294967296.0,1,-nbitq), 
to_sfixed(230464847.0/4294967296.0,1,-nbitq), 
to_sfixed(-49177351.0/4294967296.0,1,-nbitq), 
to_sfixed(-382353708.0/4294967296.0,1,-nbitq), 
to_sfixed(185595332.0/4294967296.0,1,-nbitq), 
to_sfixed(10628111.0/4294967296.0,1,-nbitq), 
to_sfixed(-101286016.0/4294967296.0,1,-nbitq), 
to_sfixed(-172033731.0/4294967296.0,1,-nbitq), 
to_sfixed(209103212.0/4294967296.0,1,-nbitq), 
to_sfixed(346049735.0/4294967296.0,1,-nbitq), 
to_sfixed(443493184.0/4294967296.0,1,-nbitq), 
to_sfixed(42619187.0/4294967296.0,1,-nbitq), 
to_sfixed(398469685.0/4294967296.0,1,-nbitq), 
to_sfixed(-336841048.0/4294967296.0,1,-nbitq), 
to_sfixed(-112798260.0/4294967296.0,1,-nbitq), 
to_sfixed(1124643.0/4294967296.0,1,-nbitq), 
to_sfixed(45402543.0/4294967296.0,1,-nbitq), 
to_sfixed(-243678269.0/4294967296.0,1,-nbitq), 
to_sfixed(-298778926.0/4294967296.0,1,-nbitq), 
to_sfixed(-251466983.0/4294967296.0,1,-nbitq), 
to_sfixed(164979175.0/4294967296.0,1,-nbitq), 
to_sfixed(-325519059.0/4294967296.0,1,-nbitq), 
to_sfixed(-192872194.0/4294967296.0,1,-nbitq), 
to_sfixed(-97243817.0/4294967296.0,1,-nbitq), 
to_sfixed(-184172500.0/4294967296.0,1,-nbitq), 
to_sfixed(53142774.0/4294967296.0,1,-nbitq), 
to_sfixed(-113181585.0/4294967296.0,1,-nbitq), 
to_sfixed(-16388906.0/4294967296.0,1,-nbitq), 
to_sfixed(354324747.0/4294967296.0,1,-nbitq), 
to_sfixed(-189541947.0/4294967296.0,1,-nbitq), 
to_sfixed(494934446.0/4294967296.0,1,-nbitq), 
to_sfixed(-136468615.0/4294967296.0,1,-nbitq), 
to_sfixed(378732883.0/4294967296.0,1,-nbitq), 
to_sfixed(-213696921.0/4294967296.0,1,-nbitq), 
to_sfixed(164610584.0/4294967296.0,1,-nbitq), 
to_sfixed(311659265.0/4294967296.0,1,-nbitq), 
to_sfixed(-339346344.0/4294967296.0,1,-nbitq), 
to_sfixed(-29715351.0/4294967296.0,1,-nbitq), 
to_sfixed(-203435632.0/4294967296.0,1,-nbitq), 
to_sfixed(-122126738.0/4294967296.0,1,-nbitq), 
to_sfixed(-224093147.0/4294967296.0,1,-nbitq), 
to_sfixed(-317213208.0/4294967296.0,1,-nbitq), 
to_sfixed(-25435003.0/4294967296.0,1,-nbitq), 
to_sfixed(462806140.0/4294967296.0,1,-nbitq), 
to_sfixed(87927435.0/4294967296.0,1,-nbitq), 
to_sfixed(336767246.0/4294967296.0,1,-nbitq), 
to_sfixed(-330797983.0/4294967296.0,1,-nbitq), 
to_sfixed(172733423.0/4294967296.0,1,-nbitq), 
to_sfixed(-231727472.0/4294967296.0,1,-nbitq), 
to_sfixed(202640113.0/4294967296.0,1,-nbitq), 
to_sfixed(177677702.0/4294967296.0,1,-nbitq), 
to_sfixed(109953105.0/4294967296.0,1,-nbitq), 
to_sfixed(371494213.0/4294967296.0,1,-nbitq), 
to_sfixed(161272532.0/4294967296.0,1,-nbitq), 
to_sfixed(-161296709.0/4294967296.0,1,-nbitq), 
to_sfixed(416763428.0/4294967296.0,1,-nbitq), 
to_sfixed(-303603502.0/4294967296.0,1,-nbitq), 
to_sfixed(-131667318.0/4294967296.0,1,-nbitq), 
to_sfixed(-149906114.0/4294967296.0,1,-nbitq), 
to_sfixed(-359400322.0/4294967296.0,1,-nbitq), 
to_sfixed(100711014.0/4294967296.0,1,-nbitq), 
to_sfixed(143904806.0/4294967296.0,1,-nbitq), 
to_sfixed(144133665.0/4294967296.0,1,-nbitq), 
to_sfixed(-218466731.0/4294967296.0,1,-nbitq), 
to_sfixed(-367193201.0/4294967296.0,1,-nbitq), 
to_sfixed(-184272434.0/4294967296.0,1,-nbitq), 
to_sfixed(-442206042.0/4294967296.0,1,-nbitq), 
to_sfixed(-428461017.0/4294967296.0,1,-nbitq), 
to_sfixed(283334019.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-108626657.0/4294967296.0,1,-nbitq), 
to_sfixed(-474952262.0/4294967296.0,1,-nbitq), 
to_sfixed(6072945.0/4294967296.0,1,-nbitq), 
to_sfixed(-396143527.0/4294967296.0,1,-nbitq), 
to_sfixed(497150703.0/4294967296.0,1,-nbitq), 
to_sfixed(278052865.0/4294967296.0,1,-nbitq), 
to_sfixed(-25572978.0/4294967296.0,1,-nbitq), 
to_sfixed(-3498390.0/4294967296.0,1,-nbitq), 
to_sfixed(-124644112.0/4294967296.0,1,-nbitq), 
to_sfixed(113453609.0/4294967296.0,1,-nbitq), 
to_sfixed(212608520.0/4294967296.0,1,-nbitq), 
to_sfixed(430862501.0/4294967296.0,1,-nbitq), 
to_sfixed(354716087.0/4294967296.0,1,-nbitq), 
to_sfixed(107814961.0/4294967296.0,1,-nbitq), 
to_sfixed(118802077.0/4294967296.0,1,-nbitq), 
to_sfixed(27519079.0/4294967296.0,1,-nbitq), 
to_sfixed(369381978.0/4294967296.0,1,-nbitq), 
to_sfixed(-63187284.0/4294967296.0,1,-nbitq), 
to_sfixed(64806408.0/4294967296.0,1,-nbitq), 
to_sfixed(-430688239.0/4294967296.0,1,-nbitq), 
to_sfixed(-241557536.0/4294967296.0,1,-nbitq), 
to_sfixed(-120481979.0/4294967296.0,1,-nbitq), 
to_sfixed(-14598524.0/4294967296.0,1,-nbitq), 
to_sfixed(217125300.0/4294967296.0,1,-nbitq), 
to_sfixed(-224229774.0/4294967296.0,1,-nbitq), 
to_sfixed(117950942.0/4294967296.0,1,-nbitq), 
to_sfixed(-165203691.0/4294967296.0,1,-nbitq), 
to_sfixed(108555387.0/4294967296.0,1,-nbitq), 
to_sfixed(463449919.0/4294967296.0,1,-nbitq), 
to_sfixed(98868232.0/4294967296.0,1,-nbitq), 
to_sfixed(-109783137.0/4294967296.0,1,-nbitq), 
to_sfixed(-206176492.0/4294967296.0,1,-nbitq), 
to_sfixed(409011621.0/4294967296.0,1,-nbitq), 
to_sfixed(-316139599.0/4294967296.0,1,-nbitq), 
to_sfixed(-156568099.0/4294967296.0,1,-nbitq), 
to_sfixed(-114007493.0/4294967296.0,1,-nbitq), 
to_sfixed(-66685238.0/4294967296.0,1,-nbitq), 
to_sfixed(473555702.0/4294967296.0,1,-nbitq), 
to_sfixed(-70252491.0/4294967296.0,1,-nbitq), 
to_sfixed(-76175085.0/4294967296.0,1,-nbitq), 
to_sfixed(-194250804.0/4294967296.0,1,-nbitq), 
to_sfixed(199674182.0/4294967296.0,1,-nbitq), 
to_sfixed(325007023.0/4294967296.0,1,-nbitq), 
to_sfixed(-202333036.0/4294967296.0,1,-nbitq), 
to_sfixed(-139157057.0/4294967296.0,1,-nbitq), 
to_sfixed(-119601019.0/4294967296.0,1,-nbitq), 
to_sfixed(326655934.0/4294967296.0,1,-nbitq), 
to_sfixed(241076425.0/4294967296.0,1,-nbitq), 
to_sfixed(-16297627.0/4294967296.0,1,-nbitq), 
to_sfixed(310509927.0/4294967296.0,1,-nbitq), 
to_sfixed(-97759386.0/4294967296.0,1,-nbitq), 
to_sfixed(-230849139.0/4294967296.0,1,-nbitq), 
to_sfixed(-425025892.0/4294967296.0,1,-nbitq), 
to_sfixed(-389248680.0/4294967296.0,1,-nbitq), 
to_sfixed(71141665.0/4294967296.0,1,-nbitq), 
to_sfixed(70533866.0/4294967296.0,1,-nbitq), 
to_sfixed(361122079.0/4294967296.0,1,-nbitq), 
to_sfixed(-218346010.0/4294967296.0,1,-nbitq), 
to_sfixed(-370368541.0/4294967296.0,1,-nbitq), 
to_sfixed(-248604699.0/4294967296.0,1,-nbitq), 
to_sfixed(-348933497.0/4294967296.0,1,-nbitq), 
to_sfixed(454494183.0/4294967296.0,1,-nbitq), 
to_sfixed(-496254809.0/4294967296.0,1,-nbitq), 
to_sfixed(-165877054.0/4294967296.0,1,-nbitq), 
to_sfixed(49342069.0/4294967296.0,1,-nbitq), 
to_sfixed(194900060.0/4294967296.0,1,-nbitq), 
to_sfixed(490936539.0/4294967296.0,1,-nbitq), 
to_sfixed(-35030397.0/4294967296.0,1,-nbitq), 
to_sfixed(-339785984.0/4294967296.0,1,-nbitq), 
to_sfixed(226282732.0/4294967296.0,1,-nbitq), 
to_sfixed(-451303231.0/4294967296.0,1,-nbitq), 
to_sfixed(-156364612.0/4294967296.0,1,-nbitq), 
to_sfixed(-105085249.0/4294967296.0,1,-nbitq), 
to_sfixed(30850433.0/4294967296.0,1,-nbitq), 
to_sfixed(353915670.0/4294967296.0,1,-nbitq), 
to_sfixed(-55195092.0/4294967296.0,1,-nbitq), 
to_sfixed(230141121.0/4294967296.0,1,-nbitq), 
to_sfixed(-145592059.0/4294967296.0,1,-nbitq), 
to_sfixed(-438979637.0/4294967296.0,1,-nbitq), 
to_sfixed(163332733.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-315770564.0/4294967296.0,1,-nbitq), 
to_sfixed(-38657191.0/4294967296.0,1,-nbitq), 
to_sfixed(-104312162.0/4294967296.0,1,-nbitq), 
to_sfixed(269722433.0/4294967296.0,1,-nbitq), 
to_sfixed(365121148.0/4294967296.0,1,-nbitq), 
to_sfixed(320138296.0/4294967296.0,1,-nbitq), 
to_sfixed(-357657334.0/4294967296.0,1,-nbitq), 
to_sfixed(-141972178.0/4294967296.0,1,-nbitq), 
to_sfixed(-79757189.0/4294967296.0,1,-nbitq), 
to_sfixed(3436960.0/4294967296.0,1,-nbitq), 
to_sfixed(-382700923.0/4294967296.0,1,-nbitq), 
to_sfixed(115540641.0/4294967296.0,1,-nbitq), 
to_sfixed(20366545.0/4294967296.0,1,-nbitq), 
to_sfixed(113626373.0/4294967296.0,1,-nbitq), 
to_sfixed(-42746242.0/4294967296.0,1,-nbitq), 
to_sfixed(-248457611.0/4294967296.0,1,-nbitq), 
to_sfixed(151964426.0/4294967296.0,1,-nbitq), 
to_sfixed(-5146402.0/4294967296.0,1,-nbitq), 
to_sfixed(315592576.0/4294967296.0,1,-nbitq), 
to_sfixed(213065017.0/4294967296.0,1,-nbitq), 
to_sfixed(63048202.0/4294967296.0,1,-nbitq), 
to_sfixed(517623912.0/4294967296.0,1,-nbitq), 
to_sfixed(354328631.0/4294967296.0,1,-nbitq), 
to_sfixed(312031859.0/4294967296.0,1,-nbitq), 
to_sfixed(-202949391.0/4294967296.0,1,-nbitq), 
to_sfixed(-19367650.0/4294967296.0,1,-nbitq), 
to_sfixed(-57382974.0/4294967296.0,1,-nbitq), 
to_sfixed(-555172889.0/4294967296.0,1,-nbitq), 
to_sfixed(-220179765.0/4294967296.0,1,-nbitq), 
to_sfixed(76165766.0/4294967296.0,1,-nbitq), 
to_sfixed(-604323270.0/4294967296.0,1,-nbitq), 
to_sfixed(91258318.0/4294967296.0,1,-nbitq), 
to_sfixed(-265097117.0/4294967296.0,1,-nbitq), 
to_sfixed(-78040569.0/4294967296.0,1,-nbitq), 
to_sfixed(71727683.0/4294967296.0,1,-nbitq), 
to_sfixed(316532508.0/4294967296.0,1,-nbitq), 
to_sfixed(99900239.0/4294967296.0,1,-nbitq), 
to_sfixed(322317063.0/4294967296.0,1,-nbitq), 
to_sfixed(32631383.0/4294967296.0,1,-nbitq), 
to_sfixed(-47568337.0/4294967296.0,1,-nbitq), 
to_sfixed(192611187.0/4294967296.0,1,-nbitq), 
to_sfixed(-211440709.0/4294967296.0,1,-nbitq), 
to_sfixed(-332014295.0/4294967296.0,1,-nbitq), 
to_sfixed(-100542821.0/4294967296.0,1,-nbitq), 
to_sfixed(-285134623.0/4294967296.0,1,-nbitq), 
to_sfixed(-145340987.0/4294967296.0,1,-nbitq), 
to_sfixed(-198142375.0/4294967296.0,1,-nbitq), 
to_sfixed(-152969991.0/4294967296.0,1,-nbitq), 
to_sfixed(-243801535.0/4294967296.0,1,-nbitq), 
to_sfixed(541405611.0/4294967296.0,1,-nbitq), 
to_sfixed(178750481.0/4294967296.0,1,-nbitq), 
to_sfixed(112722820.0/4294967296.0,1,-nbitq), 
to_sfixed(-444723393.0/4294967296.0,1,-nbitq), 
to_sfixed(-57914434.0/4294967296.0,1,-nbitq), 
to_sfixed(-1901018.0/4294967296.0,1,-nbitq), 
to_sfixed(-329369688.0/4294967296.0,1,-nbitq), 
to_sfixed(403086016.0/4294967296.0,1,-nbitq), 
to_sfixed(-609852879.0/4294967296.0,1,-nbitq), 
to_sfixed(28986544.0/4294967296.0,1,-nbitq), 
to_sfixed(123285568.0/4294967296.0,1,-nbitq), 
to_sfixed(-40912284.0/4294967296.0,1,-nbitq), 
to_sfixed(194627202.0/4294967296.0,1,-nbitq), 
to_sfixed(21404132.0/4294967296.0,1,-nbitq), 
to_sfixed(-110461126.0/4294967296.0,1,-nbitq), 
to_sfixed(279272052.0/4294967296.0,1,-nbitq), 
to_sfixed(-105601730.0/4294967296.0,1,-nbitq), 
to_sfixed(333931285.0/4294967296.0,1,-nbitq), 
to_sfixed(-371386427.0/4294967296.0,1,-nbitq), 
to_sfixed(-303603830.0/4294967296.0,1,-nbitq), 
to_sfixed(221168325.0/4294967296.0,1,-nbitq), 
to_sfixed(-364876219.0/4294967296.0,1,-nbitq), 
to_sfixed(-307643462.0/4294967296.0,1,-nbitq), 
to_sfixed(-281123565.0/4294967296.0,1,-nbitq), 
to_sfixed(78563991.0/4294967296.0,1,-nbitq), 
to_sfixed(-195676320.0/4294967296.0,1,-nbitq), 
to_sfixed(-512689154.0/4294967296.0,1,-nbitq), 
to_sfixed(14669652.0/4294967296.0,1,-nbitq), 
to_sfixed(148764599.0/4294967296.0,1,-nbitq), 
to_sfixed(85117609.0/4294967296.0,1,-nbitq), 
to_sfixed(99765348.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-46617982.0/4294967296.0,1,-nbitq), 
to_sfixed(-191534160.0/4294967296.0,1,-nbitq), 
to_sfixed(-99675632.0/4294967296.0,1,-nbitq), 
to_sfixed(-31174985.0/4294967296.0,1,-nbitq), 
to_sfixed(91752362.0/4294967296.0,1,-nbitq), 
to_sfixed(40257794.0/4294967296.0,1,-nbitq), 
to_sfixed(-243898837.0/4294967296.0,1,-nbitq), 
to_sfixed(-148671573.0/4294967296.0,1,-nbitq), 
to_sfixed(-77604974.0/4294967296.0,1,-nbitq), 
to_sfixed(-286727267.0/4294967296.0,1,-nbitq), 
to_sfixed(202274343.0/4294967296.0,1,-nbitq), 
to_sfixed(7197457.0/4294967296.0,1,-nbitq), 
to_sfixed(-104132049.0/4294967296.0,1,-nbitq), 
to_sfixed(211754974.0/4294967296.0,1,-nbitq), 
to_sfixed(-31958894.0/4294967296.0,1,-nbitq), 
to_sfixed(-268450749.0/4294967296.0,1,-nbitq), 
to_sfixed(-26333843.0/4294967296.0,1,-nbitq), 
to_sfixed(131271595.0/4294967296.0,1,-nbitq), 
to_sfixed(83894006.0/4294967296.0,1,-nbitq), 
to_sfixed(-455480366.0/4294967296.0,1,-nbitq), 
to_sfixed(-363218829.0/4294967296.0,1,-nbitq), 
to_sfixed(225947136.0/4294967296.0,1,-nbitq), 
to_sfixed(-211304656.0/4294967296.0,1,-nbitq), 
to_sfixed(152629926.0/4294967296.0,1,-nbitq), 
to_sfixed(-105229748.0/4294967296.0,1,-nbitq), 
to_sfixed(264641043.0/4294967296.0,1,-nbitq), 
to_sfixed(245326232.0/4294967296.0,1,-nbitq), 
to_sfixed(66588629.0/4294967296.0,1,-nbitq), 
to_sfixed(81205866.0/4294967296.0,1,-nbitq), 
to_sfixed(77863884.0/4294967296.0,1,-nbitq), 
to_sfixed(-494671875.0/4294967296.0,1,-nbitq), 
to_sfixed(-628083491.0/4294967296.0,1,-nbitq), 
to_sfixed(-111574956.0/4294967296.0,1,-nbitq), 
to_sfixed(171049523.0/4294967296.0,1,-nbitq), 
to_sfixed(464829457.0/4294967296.0,1,-nbitq), 
to_sfixed(331020908.0/4294967296.0,1,-nbitq), 
to_sfixed(97240615.0/4294967296.0,1,-nbitq), 
to_sfixed(-50384792.0/4294967296.0,1,-nbitq), 
to_sfixed(97273129.0/4294967296.0,1,-nbitq), 
to_sfixed(340068746.0/4294967296.0,1,-nbitq), 
to_sfixed(-220183960.0/4294967296.0,1,-nbitq), 
to_sfixed(-299656576.0/4294967296.0,1,-nbitq), 
to_sfixed(292888013.0/4294967296.0,1,-nbitq), 
to_sfixed(-190632922.0/4294967296.0,1,-nbitq), 
to_sfixed(82138508.0/4294967296.0,1,-nbitq), 
to_sfixed(-126441030.0/4294967296.0,1,-nbitq), 
to_sfixed(-135035923.0/4294967296.0,1,-nbitq), 
to_sfixed(-372527301.0/4294967296.0,1,-nbitq), 
to_sfixed(-205039674.0/4294967296.0,1,-nbitq), 
to_sfixed(-213499840.0/4294967296.0,1,-nbitq), 
to_sfixed(-351224819.0/4294967296.0,1,-nbitq), 
to_sfixed(-284574746.0/4294967296.0,1,-nbitq), 
to_sfixed(128924827.0/4294967296.0,1,-nbitq), 
to_sfixed(8523350.0/4294967296.0,1,-nbitq), 
to_sfixed(-154645271.0/4294967296.0,1,-nbitq), 
to_sfixed(311028008.0/4294967296.0,1,-nbitq), 
to_sfixed(237520028.0/4294967296.0,1,-nbitq), 
to_sfixed(-39106846.0/4294967296.0,1,-nbitq), 
to_sfixed(259415854.0/4294967296.0,1,-nbitq), 
to_sfixed(-80350549.0/4294967296.0,1,-nbitq), 
to_sfixed(236254556.0/4294967296.0,1,-nbitq), 
to_sfixed(365195276.0/4294967296.0,1,-nbitq), 
to_sfixed(83244972.0/4294967296.0,1,-nbitq), 
to_sfixed(-69069398.0/4294967296.0,1,-nbitq), 
to_sfixed(341111867.0/4294967296.0,1,-nbitq), 
to_sfixed(171409234.0/4294967296.0,1,-nbitq), 
to_sfixed(767948044.0/4294967296.0,1,-nbitq), 
to_sfixed(378099601.0/4294967296.0,1,-nbitq), 
to_sfixed(-155385938.0/4294967296.0,1,-nbitq), 
to_sfixed(-54675515.0/4294967296.0,1,-nbitq), 
to_sfixed(-161952021.0/4294967296.0,1,-nbitq), 
to_sfixed(250599885.0/4294967296.0,1,-nbitq), 
to_sfixed(-467370456.0/4294967296.0,1,-nbitq), 
to_sfixed(369084521.0/4294967296.0,1,-nbitq), 
to_sfixed(-90541518.0/4294967296.0,1,-nbitq), 
to_sfixed(95792491.0/4294967296.0,1,-nbitq), 
to_sfixed(-239042590.0/4294967296.0,1,-nbitq), 
to_sfixed(-343100949.0/4294967296.0,1,-nbitq), 
to_sfixed(-424749027.0/4294967296.0,1,-nbitq), 
to_sfixed(133815426.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-92041132.0/4294967296.0,1,-nbitq), 
to_sfixed(-164456602.0/4294967296.0,1,-nbitq), 
to_sfixed(-103716871.0/4294967296.0,1,-nbitq), 
to_sfixed(80121429.0/4294967296.0,1,-nbitq), 
to_sfixed(283781921.0/4294967296.0,1,-nbitq), 
to_sfixed(-27951385.0/4294967296.0,1,-nbitq), 
to_sfixed(74191398.0/4294967296.0,1,-nbitq), 
to_sfixed(-355512511.0/4294967296.0,1,-nbitq), 
to_sfixed(-572248889.0/4294967296.0,1,-nbitq), 
to_sfixed(420712467.0/4294967296.0,1,-nbitq), 
to_sfixed(99425997.0/4294967296.0,1,-nbitq), 
to_sfixed(-583664112.0/4294967296.0,1,-nbitq), 
to_sfixed(453296497.0/4294967296.0,1,-nbitq), 
to_sfixed(902451675.0/4294967296.0,1,-nbitq), 
to_sfixed(-398501609.0/4294967296.0,1,-nbitq), 
to_sfixed(238326304.0/4294967296.0,1,-nbitq), 
to_sfixed(221435595.0/4294967296.0,1,-nbitq), 
to_sfixed(159189955.0/4294967296.0,1,-nbitq), 
to_sfixed(508972148.0/4294967296.0,1,-nbitq), 
to_sfixed(-64058731.0/4294967296.0,1,-nbitq), 
to_sfixed(345223559.0/4294967296.0,1,-nbitq), 
to_sfixed(-82151116.0/4294967296.0,1,-nbitq), 
to_sfixed(272160738.0/4294967296.0,1,-nbitq), 
to_sfixed(391046217.0/4294967296.0,1,-nbitq), 
to_sfixed(-34237655.0/4294967296.0,1,-nbitq), 
to_sfixed(627350046.0/4294967296.0,1,-nbitq), 
to_sfixed(-258925735.0/4294967296.0,1,-nbitq), 
to_sfixed(-208980038.0/4294967296.0,1,-nbitq), 
to_sfixed(335711665.0/4294967296.0,1,-nbitq), 
to_sfixed(236253053.0/4294967296.0,1,-nbitq), 
to_sfixed(-342313324.0/4294967296.0,1,-nbitq), 
to_sfixed(50272020.0/4294967296.0,1,-nbitq), 
to_sfixed(-256958733.0/4294967296.0,1,-nbitq), 
to_sfixed(-90241349.0/4294967296.0,1,-nbitq), 
to_sfixed(176663957.0/4294967296.0,1,-nbitq), 
to_sfixed(67331477.0/4294967296.0,1,-nbitq), 
to_sfixed(45661908.0/4294967296.0,1,-nbitq), 
to_sfixed(539177199.0/4294967296.0,1,-nbitq), 
to_sfixed(-417781146.0/4294967296.0,1,-nbitq), 
to_sfixed(-223825223.0/4294967296.0,1,-nbitq), 
to_sfixed(-411460883.0/4294967296.0,1,-nbitq), 
to_sfixed(230798918.0/4294967296.0,1,-nbitq), 
to_sfixed(87230856.0/4294967296.0,1,-nbitq), 
to_sfixed(-15763582.0/4294967296.0,1,-nbitq), 
to_sfixed(-50869606.0/4294967296.0,1,-nbitq), 
to_sfixed(59774170.0/4294967296.0,1,-nbitq), 
to_sfixed(80598410.0/4294967296.0,1,-nbitq), 
to_sfixed(-277928401.0/4294967296.0,1,-nbitq), 
to_sfixed(12260625.0/4294967296.0,1,-nbitq), 
to_sfixed(-302385691.0/4294967296.0,1,-nbitq), 
to_sfixed(-2883317.0/4294967296.0,1,-nbitq), 
to_sfixed(8583118.0/4294967296.0,1,-nbitq), 
to_sfixed(-103183326.0/4294967296.0,1,-nbitq), 
to_sfixed(46419687.0/4294967296.0,1,-nbitq), 
to_sfixed(105226432.0/4294967296.0,1,-nbitq), 
to_sfixed(92304564.0/4294967296.0,1,-nbitq), 
to_sfixed(-311690016.0/4294967296.0,1,-nbitq), 
to_sfixed(296287949.0/4294967296.0,1,-nbitq), 
to_sfixed(-269531771.0/4294967296.0,1,-nbitq), 
to_sfixed(-137945444.0/4294967296.0,1,-nbitq), 
to_sfixed(318070211.0/4294967296.0,1,-nbitq), 
to_sfixed(106563802.0/4294967296.0,1,-nbitq), 
to_sfixed(-15403641.0/4294967296.0,1,-nbitq), 
to_sfixed(235300687.0/4294967296.0,1,-nbitq), 
to_sfixed(-76815135.0/4294967296.0,1,-nbitq), 
to_sfixed(175560404.0/4294967296.0,1,-nbitq), 
to_sfixed(353080690.0/4294967296.0,1,-nbitq), 
to_sfixed(208281840.0/4294967296.0,1,-nbitq), 
to_sfixed(-82043807.0/4294967296.0,1,-nbitq), 
to_sfixed(184282453.0/4294967296.0,1,-nbitq), 
to_sfixed(206943405.0/4294967296.0,1,-nbitq), 
to_sfixed(216932881.0/4294967296.0,1,-nbitq), 
to_sfixed(157917055.0/4294967296.0,1,-nbitq), 
to_sfixed(239884853.0/4294967296.0,1,-nbitq), 
to_sfixed(-42270366.0/4294967296.0,1,-nbitq), 
to_sfixed(-109014893.0/4294967296.0,1,-nbitq), 
to_sfixed(204255393.0/4294967296.0,1,-nbitq), 
to_sfixed(151615780.0/4294967296.0,1,-nbitq), 
to_sfixed(166306003.0/4294967296.0,1,-nbitq), 
to_sfixed(294720970.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(393264366.0/4294967296.0,1,-nbitq), 
to_sfixed(20017107.0/4294967296.0,1,-nbitq), 
to_sfixed(-245383032.0/4294967296.0,1,-nbitq), 
to_sfixed(1043240389.0/4294967296.0,1,-nbitq), 
to_sfixed(194694027.0/4294967296.0,1,-nbitq), 
to_sfixed(667578786.0/4294967296.0,1,-nbitq), 
to_sfixed(-305610570.0/4294967296.0,1,-nbitq), 
to_sfixed(-379998020.0/4294967296.0,1,-nbitq), 
to_sfixed(-692004494.0/4294967296.0,1,-nbitq), 
to_sfixed(42154684.0/4294967296.0,1,-nbitq), 
to_sfixed(493113089.0/4294967296.0,1,-nbitq), 
to_sfixed(-359848433.0/4294967296.0,1,-nbitq), 
to_sfixed(519779805.0/4294967296.0,1,-nbitq), 
to_sfixed(189341484.0/4294967296.0,1,-nbitq), 
to_sfixed(175013505.0/4294967296.0,1,-nbitq), 
to_sfixed(-192617172.0/4294967296.0,1,-nbitq), 
to_sfixed(358774571.0/4294967296.0,1,-nbitq), 
to_sfixed(234505785.0/4294967296.0,1,-nbitq), 
to_sfixed(272602425.0/4294967296.0,1,-nbitq), 
to_sfixed(-59233422.0/4294967296.0,1,-nbitq), 
to_sfixed(142402443.0/4294967296.0,1,-nbitq), 
to_sfixed(-466574454.0/4294967296.0,1,-nbitq), 
to_sfixed(-448225875.0/4294967296.0,1,-nbitq), 
to_sfixed(541095704.0/4294967296.0,1,-nbitq), 
to_sfixed(-238985074.0/4294967296.0,1,-nbitq), 
to_sfixed(640163061.0/4294967296.0,1,-nbitq), 
to_sfixed(285795729.0/4294967296.0,1,-nbitq), 
to_sfixed(390913705.0/4294967296.0,1,-nbitq), 
to_sfixed(562075079.0/4294967296.0,1,-nbitq), 
to_sfixed(-42227362.0/4294967296.0,1,-nbitq), 
to_sfixed(-153929292.0/4294967296.0,1,-nbitq), 
to_sfixed(-356195689.0/4294967296.0,1,-nbitq), 
to_sfixed(-65503716.0/4294967296.0,1,-nbitq), 
to_sfixed(16251176.0/4294967296.0,1,-nbitq), 
to_sfixed(-184330353.0/4294967296.0,1,-nbitq), 
to_sfixed(18598054.0/4294967296.0,1,-nbitq), 
to_sfixed(378858609.0/4294967296.0,1,-nbitq), 
to_sfixed(777039470.0/4294967296.0,1,-nbitq), 
to_sfixed(-119604746.0/4294967296.0,1,-nbitq), 
to_sfixed(29837225.0/4294967296.0,1,-nbitq), 
to_sfixed(-371999884.0/4294967296.0,1,-nbitq), 
to_sfixed(-233336287.0/4294967296.0,1,-nbitq), 
to_sfixed(634668735.0/4294967296.0,1,-nbitq), 
to_sfixed(-275920807.0/4294967296.0,1,-nbitq), 
to_sfixed(-154667054.0/4294967296.0,1,-nbitq), 
to_sfixed(581776054.0/4294967296.0,1,-nbitq), 
to_sfixed(-245198174.0/4294967296.0,1,-nbitq), 
to_sfixed(-110621752.0/4294967296.0,1,-nbitq), 
to_sfixed(-180797776.0/4294967296.0,1,-nbitq), 
to_sfixed(-628604083.0/4294967296.0,1,-nbitq), 
to_sfixed(-381534639.0/4294967296.0,1,-nbitq), 
to_sfixed(153556390.0/4294967296.0,1,-nbitq), 
to_sfixed(816502952.0/4294967296.0,1,-nbitq), 
to_sfixed(-208195268.0/4294967296.0,1,-nbitq), 
to_sfixed(1020987032.0/4294967296.0,1,-nbitq), 
to_sfixed(291969522.0/4294967296.0,1,-nbitq), 
to_sfixed(-23027616.0/4294967296.0,1,-nbitq), 
to_sfixed(-81550444.0/4294967296.0,1,-nbitq), 
to_sfixed(233393154.0/4294967296.0,1,-nbitq), 
to_sfixed(-24845222.0/4294967296.0,1,-nbitq), 
to_sfixed(-84259571.0/4294967296.0,1,-nbitq), 
to_sfixed(259054122.0/4294967296.0,1,-nbitq), 
to_sfixed(-508068093.0/4294967296.0,1,-nbitq), 
to_sfixed(439338540.0/4294967296.0,1,-nbitq), 
to_sfixed(-562999973.0/4294967296.0,1,-nbitq), 
to_sfixed(-221870081.0/4294967296.0,1,-nbitq), 
to_sfixed(-51885144.0/4294967296.0,1,-nbitq), 
to_sfixed(-71776271.0/4294967296.0,1,-nbitq), 
to_sfixed(-104294575.0/4294967296.0,1,-nbitq), 
to_sfixed(-87607443.0/4294967296.0,1,-nbitq), 
to_sfixed(143333446.0/4294967296.0,1,-nbitq), 
to_sfixed(391170676.0/4294967296.0,1,-nbitq), 
to_sfixed(192185145.0/4294967296.0,1,-nbitq), 
to_sfixed(88684372.0/4294967296.0,1,-nbitq), 
to_sfixed(35828076.0/4294967296.0,1,-nbitq), 
to_sfixed(-447193613.0/4294967296.0,1,-nbitq), 
to_sfixed(-20786527.0/4294967296.0,1,-nbitq), 
to_sfixed(-77859474.0/4294967296.0,1,-nbitq), 
to_sfixed(360526091.0/4294967296.0,1,-nbitq), 
to_sfixed(-297550688.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-129456342.0/4294967296.0,1,-nbitq), 
to_sfixed(409942564.0/4294967296.0,1,-nbitq), 
to_sfixed(249704085.0/4294967296.0,1,-nbitq), 
to_sfixed(607527140.0/4294967296.0,1,-nbitq), 
to_sfixed(878495173.0/4294967296.0,1,-nbitq), 
to_sfixed(71743306.0/4294967296.0,1,-nbitq), 
to_sfixed(167797136.0/4294967296.0,1,-nbitq), 
to_sfixed(-402777733.0/4294967296.0,1,-nbitq), 
to_sfixed(-312905661.0/4294967296.0,1,-nbitq), 
to_sfixed(11912645.0/4294967296.0,1,-nbitq), 
to_sfixed(692898541.0/4294967296.0,1,-nbitq), 
to_sfixed(-743168374.0/4294967296.0,1,-nbitq), 
to_sfixed(518919433.0/4294967296.0,1,-nbitq), 
to_sfixed(740010195.0/4294967296.0,1,-nbitq), 
to_sfixed(122767739.0/4294967296.0,1,-nbitq), 
to_sfixed(-728818145.0/4294967296.0,1,-nbitq), 
to_sfixed(-194932845.0/4294967296.0,1,-nbitq), 
to_sfixed(230628675.0/4294967296.0,1,-nbitq), 
to_sfixed(-340807133.0/4294967296.0,1,-nbitq), 
to_sfixed(345249638.0/4294967296.0,1,-nbitq), 
to_sfixed(-119760674.0/4294967296.0,1,-nbitq), 
to_sfixed(-278046422.0/4294967296.0,1,-nbitq), 
to_sfixed(-151751074.0/4294967296.0,1,-nbitq), 
to_sfixed(198145937.0/4294967296.0,1,-nbitq), 
to_sfixed(-345190503.0/4294967296.0,1,-nbitq), 
to_sfixed(-96123388.0/4294967296.0,1,-nbitq), 
to_sfixed(-185462161.0/4294967296.0,1,-nbitq), 
to_sfixed(9293450.0/4294967296.0,1,-nbitq), 
to_sfixed(358265021.0/4294967296.0,1,-nbitq), 
to_sfixed(-230051274.0/4294967296.0,1,-nbitq), 
to_sfixed(-215602094.0/4294967296.0,1,-nbitq), 
to_sfixed(-121717508.0/4294967296.0,1,-nbitq), 
to_sfixed(-217129080.0/4294967296.0,1,-nbitq), 
to_sfixed(-184831212.0/4294967296.0,1,-nbitq), 
to_sfixed(7754278.0/4294967296.0,1,-nbitq), 
to_sfixed(202314490.0/4294967296.0,1,-nbitq), 
to_sfixed(-230101536.0/4294967296.0,1,-nbitq), 
to_sfixed(892210825.0/4294967296.0,1,-nbitq), 
to_sfixed(102776394.0/4294967296.0,1,-nbitq), 
to_sfixed(266196942.0/4294967296.0,1,-nbitq), 
to_sfixed(-29572393.0/4294967296.0,1,-nbitq), 
to_sfixed(-84735564.0/4294967296.0,1,-nbitq), 
to_sfixed(215719363.0/4294967296.0,1,-nbitq), 
to_sfixed(-13786746.0/4294967296.0,1,-nbitq), 
to_sfixed(309577644.0/4294967296.0,1,-nbitq), 
to_sfixed(352544232.0/4294967296.0,1,-nbitq), 
to_sfixed(141366227.0/4294967296.0,1,-nbitq), 
to_sfixed(-420917522.0/4294967296.0,1,-nbitq), 
to_sfixed(-15989566.0/4294967296.0,1,-nbitq), 
to_sfixed(-593450538.0/4294967296.0,1,-nbitq), 
to_sfixed(345833215.0/4294967296.0,1,-nbitq), 
to_sfixed(194808899.0/4294967296.0,1,-nbitq), 
to_sfixed(1207294973.0/4294967296.0,1,-nbitq), 
to_sfixed(-509960534.0/4294967296.0,1,-nbitq), 
to_sfixed(318682363.0/4294967296.0,1,-nbitq), 
to_sfixed(540647385.0/4294967296.0,1,-nbitq), 
to_sfixed(-299815294.0/4294967296.0,1,-nbitq), 
to_sfixed(162055836.0/4294967296.0,1,-nbitq), 
to_sfixed(-90451035.0/4294967296.0,1,-nbitq), 
to_sfixed(-27994936.0/4294967296.0,1,-nbitq), 
to_sfixed(-24986381.0/4294967296.0,1,-nbitq), 
to_sfixed(-279873668.0/4294967296.0,1,-nbitq), 
to_sfixed(-1416381687.0/4294967296.0,1,-nbitq), 
to_sfixed(214419373.0/4294967296.0,1,-nbitq), 
to_sfixed(-195885215.0/4294967296.0,1,-nbitq), 
to_sfixed(-399706431.0/4294967296.0,1,-nbitq), 
to_sfixed(-543588767.0/4294967296.0,1,-nbitq), 
to_sfixed(918141936.0/4294967296.0,1,-nbitq), 
to_sfixed(295978972.0/4294967296.0,1,-nbitq), 
to_sfixed(-98395487.0/4294967296.0,1,-nbitq), 
to_sfixed(-940740.0/4294967296.0,1,-nbitq), 
to_sfixed(489138914.0/4294967296.0,1,-nbitq), 
to_sfixed(-387565956.0/4294967296.0,1,-nbitq), 
to_sfixed(-158076983.0/4294967296.0,1,-nbitq), 
to_sfixed(467225213.0/4294967296.0,1,-nbitq), 
to_sfixed(-694335592.0/4294967296.0,1,-nbitq), 
to_sfixed(528152114.0/4294967296.0,1,-nbitq), 
to_sfixed(-7957787.0/4294967296.0,1,-nbitq), 
to_sfixed(206722052.0/4294967296.0,1,-nbitq), 
to_sfixed(-44051847.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(142439648.0/4294967296.0,1,-nbitq), 
to_sfixed(-55989139.0/4294967296.0,1,-nbitq), 
to_sfixed(-173331128.0/4294967296.0,1,-nbitq), 
to_sfixed(967588921.0/4294967296.0,1,-nbitq), 
to_sfixed(1176370374.0/4294967296.0,1,-nbitq), 
to_sfixed(311293349.0/4294967296.0,1,-nbitq), 
to_sfixed(226095681.0/4294967296.0,1,-nbitq), 
to_sfixed(214566557.0/4294967296.0,1,-nbitq), 
to_sfixed(179985334.0/4294967296.0,1,-nbitq), 
to_sfixed(164610036.0/4294967296.0,1,-nbitq), 
to_sfixed(481144191.0/4294967296.0,1,-nbitq), 
to_sfixed(-371599866.0/4294967296.0,1,-nbitq), 
to_sfixed(542465096.0/4294967296.0,1,-nbitq), 
to_sfixed(-5846560.0/4294967296.0,1,-nbitq), 
to_sfixed(155074581.0/4294967296.0,1,-nbitq), 
to_sfixed(-839441077.0/4294967296.0,1,-nbitq), 
to_sfixed(-322556691.0/4294967296.0,1,-nbitq), 
to_sfixed(17307899.0/4294967296.0,1,-nbitq), 
to_sfixed(316851338.0/4294967296.0,1,-nbitq), 
to_sfixed(-40880526.0/4294967296.0,1,-nbitq), 
to_sfixed(-202200292.0/4294967296.0,1,-nbitq), 
to_sfixed(-210330653.0/4294967296.0,1,-nbitq), 
to_sfixed(-472571558.0/4294967296.0,1,-nbitq), 
to_sfixed(551663354.0/4294967296.0,1,-nbitq), 
to_sfixed(-154500925.0/4294967296.0,1,-nbitq), 
to_sfixed(-54626736.0/4294967296.0,1,-nbitq), 
to_sfixed(140806682.0/4294967296.0,1,-nbitq), 
to_sfixed(-281091720.0/4294967296.0,1,-nbitq), 
to_sfixed(380803374.0/4294967296.0,1,-nbitq), 
to_sfixed(-588144187.0/4294967296.0,1,-nbitq), 
to_sfixed(-356022573.0/4294967296.0,1,-nbitq), 
to_sfixed(-465712808.0/4294967296.0,1,-nbitq), 
to_sfixed(-224212392.0/4294967296.0,1,-nbitq), 
to_sfixed(175516957.0/4294967296.0,1,-nbitq), 
to_sfixed(116902587.0/4294967296.0,1,-nbitq), 
to_sfixed(-274415836.0/4294967296.0,1,-nbitq), 
to_sfixed(19066322.0/4294967296.0,1,-nbitq), 
to_sfixed(531843871.0/4294967296.0,1,-nbitq), 
to_sfixed(-305968797.0/4294967296.0,1,-nbitq), 
to_sfixed(503257038.0/4294967296.0,1,-nbitq), 
to_sfixed(-461715111.0/4294967296.0,1,-nbitq), 
to_sfixed(-135516577.0/4294967296.0,1,-nbitq), 
to_sfixed(-377202788.0/4294967296.0,1,-nbitq), 
to_sfixed(-547605313.0/4294967296.0,1,-nbitq), 
to_sfixed(455429163.0/4294967296.0,1,-nbitq), 
to_sfixed(433544893.0/4294967296.0,1,-nbitq), 
to_sfixed(-346784095.0/4294967296.0,1,-nbitq), 
to_sfixed(-493121564.0/4294967296.0,1,-nbitq), 
to_sfixed(149316992.0/4294967296.0,1,-nbitq), 
to_sfixed(-767840830.0/4294967296.0,1,-nbitq), 
to_sfixed(108297669.0/4294967296.0,1,-nbitq), 
to_sfixed(574143563.0/4294967296.0,1,-nbitq), 
to_sfixed(764344059.0/4294967296.0,1,-nbitq), 
to_sfixed(-384852247.0/4294967296.0,1,-nbitq), 
to_sfixed(430770683.0/4294967296.0,1,-nbitq), 
to_sfixed(1122657798.0/4294967296.0,1,-nbitq), 
to_sfixed(-233531416.0/4294967296.0,1,-nbitq), 
to_sfixed(398556048.0/4294967296.0,1,-nbitq), 
to_sfixed(-224028293.0/4294967296.0,1,-nbitq), 
to_sfixed(-143420238.0/4294967296.0,1,-nbitq), 
to_sfixed(118014254.0/4294967296.0,1,-nbitq), 
to_sfixed(126810339.0/4294967296.0,1,-nbitq), 
to_sfixed(-883526831.0/4294967296.0,1,-nbitq), 
to_sfixed(552519723.0/4294967296.0,1,-nbitq), 
to_sfixed(-435091515.0/4294967296.0,1,-nbitq), 
to_sfixed(-273014047.0/4294967296.0,1,-nbitq), 
to_sfixed(-354503474.0/4294967296.0,1,-nbitq), 
to_sfixed(689805933.0/4294967296.0,1,-nbitq), 
to_sfixed(143038579.0/4294967296.0,1,-nbitq), 
to_sfixed(-1027942090.0/4294967296.0,1,-nbitq), 
to_sfixed(213081932.0/4294967296.0,1,-nbitq), 
to_sfixed(90947082.0/4294967296.0,1,-nbitq), 
to_sfixed(-334490362.0/4294967296.0,1,-nbitq), 
to_sfixed(-303597095.0/4294967296.0,1,-nbitq), 
to_sfixed(339696650.0/4294967296.0,1,-nbitq), 
to_sfixed(350078628.0/4294967296.0,1,-nbitq), 
to_sfixed(501529887.0/4294967296.0,1,-nbitq), 
to_sfixed(388946900.0/4294967296.0,1,-nbitq), 
to_sfixed(61987554.0/4294967296.0,1,-nbitq), 
to_sfixed(283532813.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-376932559.0/4294967296.0,1,-nbitq), 
to_sfixed(-42155885.0/4294967296.0,1,-nbitq), 
to_sfixed(-295158685.0/4294967296.0,1,-nbitq), 
to_sfixed(470278571.0/4294967296.0,1,-nbitq), 
to_sfixed(1522626105.0/4294967296.0,1,-nbitq), 
to_sfixed(1132217877.0/4294967296.0,1,-nbitq), 
to_sfixed(454176821.0/4294967296.0,1,-nbitq), 
to_sfixed(272168621.0/4294967296.0,1,-nbitq), 
to_sfixed(335559739.0/4294967296.0,1,-nbitq), 
to_sfixed(81406913.0/4294967296.0,1,-nbitq), 
to_sfixed(414919286.0/4294967296.0,1,-nbitq), 
to_sfixed(-769590386.0/4294967296.0,1,-nbitq), 
to_sfixed(972058725.0/4294967296.0,1,-nbitq), 
to_sfixed(-386559397.0/4294967296.0,1,-nbitq), 
to_sfixed(-118778996.0/4294967296.0,1,-nbitq), 
to_sfixed(-822513998.0/4294967296.0,1,-nbitq), 
to_sfixed(159155203.0/4294967296.0,1,-nbitq), 
to_sfixed(-76967862.0/4294967296.0,1,-nbitq), 
to_sfixed(223282068.0/4294967296.0,1,-nbitq), 
to_sfixed(439898159.0/4294967296.0,1,-nbitq), 
to_sfixed(38393606.0/4294967296.0,1,-nbitq), 
to_sfixed(-384644098.0/4294967296.0,1,-nbitq), 
to_sfixed(-57745668.0/4294967296.0,1,-nbitq), 
to_sfixed(432939923.0/4294967296.0,1,-nbitq), 
to_sfixed(340513350.0/4294967296.0,1,-nbitq), 
to_sfixed(115878169.0/4294967296.0,1,-nbitq), 
to_sfixed(-66703279.0/4294967296.0,1,-nbitq), 
to_sfixed(-446942538.0/4294967296.0,1,-nbitq), 
to_sfixed(577265107.0/4294967296.0,1,-nbitq), 
to_sfixed(-933801732.0/4294967296.0,1,-nbitq), 
to_sfixed(-132258441.0/4294967296.0,1,-nbitq), 
to_sfixed(-174069913.0/4294967296.0,1,-nbitq), 
to_sfixed(-144721072.0/4294967296.0,1,-nbitq), 
to_sfixed(312899927.0/4294967296.0,1,-nbitq), 
to_sfixed(-110383798.0/4294967296.0,1,-nbitq), 
to_sfixed(-231669020.0/4294967296.0,1,-nbitq), 
to_sfixed(295113196.0/4294967296.0,1,-nbitq), 
to_sfixed(-144033023.0/4294967296.0,1,-nbitq), 
to_sfixed(-281094870.0/4294967296.0,1,-nbitq), 
to_sfixed(165377730.0/4294967296.0,1,-nbitq), 
to_sfixed(-433864777.0/4294967296.0,1,-nbitq), 
to_sfixed(-362925287.0/4294967296.0,1,-nbitq), 
to_sfixed(-25465861.0/4294967296.0,1,-nbitq), 
to_sfixed(-410538719.0/4294967296.0,1,-nbitq), 
to_sfixed(-112947.0/4294967296.0,1,-nbitq), 
to_sfixed(-394187080.0/4294967296.0,1,-nbitq), 
to_sfixed(-380194030.0/4294967296.0,1,-nbitq), 
to_sfixed(-455414333.0/4294967296.0,1,-nbitq), 
to_sfixed(337283017.0/4294967296.0,1,-nbitq), 
to_sfixed(-657014306.0/4294967296.0,1,-nbitq), 
to_sfixed(-36246935.0/4294967296.0,1,-nbitq), 
to_sfixed(349541754.0/4294967296.0,1,-nbitq), 
to_sfixed(611921182.0/4294967296.0,1,-nbitq), 
to_sfixed(-109943680.0/4294967296.0,1,-nbitq), 
to_sfixed(961856750.0/4294967296.0,1,-nbitq), 
to_sfixed(1670619870.0/4294967296.0,1,-nbitq), 
to_sfixed(-68648456.0/4294967296.0,1,-nbitq), 
to_sfixed(19817423.0/4294967296.0,1,-nbitq), 
to_sfixed(273609996.0/4294967296.0,1,-nbitq), 
to_sfixed(-84734565.0/4294967296.0,1,-nbitq), 
to_sfixed(-131892885.0/4294967296.0,1,-nbitq), 
to_sfixed(-246506068.0/4294967296.0,1,-nbitq), 
to_sfixed(-715752057.0/4294967296.0,1,-nbitq), 
to_sfixed(1078369863.0/4294967296.0,1,-nbitq), 
to_sfixed(-98795539.0/4294967296.0,1,-nbitq), 
to_sfixed(-193175312.0/4294967296.0,1,-nbitq), 
to_sfixed(-372913157.0/4294967296.0,1,-nbitq), 
to_sfixed(329667965.0/4294967296.0,1,-nbitq), 
to_sfixed(-173777409.0/4294967296.0,1,-nbitq), 
to_sfixed(-818520547.0/4294967296.0,1,-nbitq), 
to_sfixed(-628001634.0/4294967296.0,1,-nbitq), 
to_sfixed(283996892.0/4294967296.0,1,-nbitq), 
to_sfixed(347958004.0/4294967296.0,1,-nbitq), 
to_sfixed(379979271.0/4294967296.0,1,-nbitq), 
to_sfixed(-222609442.0/4294967296.0,1,-nbitq), 
to_sfixed(135958804.0/4294967296.0,1,-nbitq), 
to_sfixed(278624702.0/4294967296.0,1,-nbitq), 
to_sfixed(484017002.0/4294967296.0,1,-nbitq), 
to_sfixed(-62250918.0/4294967296.0,1,-nbitq), 
to_sfixed(-264189921.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-68102140.0/4294967296.0,1,-nbitq), 
to_sfixed(-1260593652.0/4294967296.0,1,-nbitq), 
to_sfixed(232620914.0/4294967296.0,1,-nbitq), 
to_sfixed(204763385.0/4294967296.0,1,-nbitq), 
to_sfixed(370072271.0/4294967296.0,1,-nbitq), 
to_sfixed(1974317852.0/4294967296.0,1,-nbitq), 
to_sfixed(-117373539.0/4294967296.0,1,-nbitq), 
to_sfixed(491758867.0/4294967296.0,1,-nbitq), 
to_sfixed(511474703.0/4294967296.0,1,-nbitq), 
to_sfixed(118488132.0/4294967296.0,1,-nbitq), 
to_sfixed(19908531.0/4294967296.0,1,-nbitq), 
to_sfixed(-611075123.0/4294967296.0,1,-nbitq), 
to_sfixed(779224236.0/4294967296.0,1,-nbitq), 
to_sfixed(-742630935.0/4294967296.0,1,-nbitq), 
to_sfixed(440940779.0/4294967296.0,1,-nbitq), 
to_sfixed(-598916597.0/4294967296.0,1,-nbitq), 
to_sfixed(-225005794.0/4294967296.0,1,-nbitq), 
to_sfixed(-47421326.0/4294967296.0,1,-nbitq), 
to_sfixed(293439969.0/4294967296.0,1,-nbitq), 
to_sfixed(723944536.0/4294967296.0,1,-nbitq), 
to_sfixed(-266741639.0/4294967296.0,1,-nbitq), 
to_sfixed(-293539696.0/4294967296.0,1,-nbitq), 
to_sfixed(-598599218.0/4294967296.0,1,-nbitq), 
to_sfixed(826815174.0/4294967296.0,1,-nbitq), 
to_sfixed(-377568117.0/4294967296.0,1,-nbitq), 
to_sfixed(210280998.0/4294967296.0,1,-nbitq), 
to_sfixed(-264427851.0/4294967296.0,1,-nbitq), 
to_sfixed(-105935431.0/4294967296.0,1,-nbitq), 
to_sfixed(-66292516.0/4294967296.0,1,-nbitq), 
to_sfixed(-233094949.0/4294967296.0,1,-nbitq), 
to_sfixed(206467009.0/4294967296.0,1,-nbitq), 
to_sfixed(-1070044264.0/4294967296.0,1,-nbitq), 
to_sfixed(568465584.0/4294967296.0,1,-nbitq), 
to_sfixed(89269154.0/4294967296.0,1,-nbitq), 
to_sfixed(-117457491.0/4294967296.0,1,-nbitq), 
to_sfixed(-223008054.0/4294967296.0,1,-nbitq), 
to_sfixed(243899472.0/4294967296.0,1,-nbitq), 
to_sfixed(-223769296.0/4294967296.0,1,-nbitq), 
to_sfixed(-97300314.0/4294967296.0,1,-nbitq), 
to_sfixed(16870320.0/4294967296.0,1,-nbitq), 
to_sfixed(-39586238.0/4294967296.0,1,-nbitq), 
to_sfixed(-549833091.0/4294967296.0,1,-nbitq), 
to_sfixed(400331864.0/4294967296.0,1,-nbitq), 
to_sfixed(-514432594.0/4294967296.0,1,-nbitq), 
to_sfixed(437607280.0/4294967296.0,1,-nbitq), 
to_sfixed(-211153053.0/4294967296.0,1,-nbitq), 
to_sfixed(36818706.0/4294967296.0,1,-nbitq), 
to_sfixed(-631002655.0/4294967296.0,1,-nbitq), 
to_sfixed(371929715.0/4294967296.0,1,-nbitq), 
to_sfixed(-653973043.0/4294967296.0,1,-nbitq), 
to_sfixed(226670780.0/4294967296.0,1,-nbitq), 
to_sfixed(-282768286.0/4294967296.0,1,-nbitq), 
to_sfixed(412381971.0/4294967296.0,1,-nbitq), 
to_sfixed(-510537475.0/4294967296.0,1,-nbitq), 
to_sfixed(-49962803.0/4294967296.0,1,-nbitq), 
to_sfixed(762862046.0/4294967296.0,1,-nbitq), 
to_sfixed(28663164.0/4294967296.0,1,-nbitq), 
to_sfixed(255298105.0/4294967296.0,1,-nbitq), 
to_sfixed(72752088.0/4294967296.0,1,-nbitq), 
to_sfixed(-307333786.0/4294967296.0,1,-nbitq), 
to_sfixed(-225102675.0/4294967296.0,1,-nbitq), 
to_sfixed(-75564154.0/4294967296.0,1,-nbitq), 
to_sfixed(-700985509.0/4294967296.0,1,-nbitq), 
to_sfixed(1128997282.0/4294967296.0,1,-nbitq), 
to_sfixed(-222819247.0/4294967296.0,1,-nbitq), 
to_sfixed(159231044.0/4294967296.0,1,-nbitq), 
to_sfixed(-1075876499.0/4294967296.0,1,-nbitq), 
to_sfixed(2549394.0/4294967296.0,1,-nbitq), 
to_sfixed(-188292524.0/4294967296.0,1,-nbitq), 
to_sfixed(-1119169864.0/4294967296.0,1,-nbitq), 
to_sfixed(-868970388.0/4294967296.0,1,-nbitq), 
to_sfixed(-17446052.0/4294967296.0,1,-nbitq), 
to_sfixed(-75500731.0/4294967296.0,1,-nbitq), 
to_sfixed(-292607937.0/4294967296.0,1,-nbitq), 
to_sfixed(88326289.0/4294967296.0,1,-nbitq), 
to_sfixed(-205996815.0/4294967296.0,1,-nbitq), 
to_sfixed(1110365674.0/4294967296.0,1,-nbitq), 
to_sfixed(685838545.0/4294967296.0,1,-nbitq), 
to_sfixed(-484292856.0/4294967296.0,1,-nbitq), 
to_sfixed(-246947792.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-155894030.0/4294967296.0,1,-nbitq), 
to_sfixed(-1034059120.0/4294967296.0,1,-nbitq), 
to_sfixed(360028001.0/4294967296.0,1,-nbitq), 
to_sfixed(-32902461.0/4294967296.0,1,-nbitq), 
to_sfixed(1235290745.0/4294967296.0,1,-nbitq), 
to_sfixed(1018285104.0/4294967296.0,1,-nbitq), 
to_sfixed(38160058.0/4294967296.0,1,-nbitq), 
to_sfixed(86847538.0/4294967296.0,1,-nbitq), 
to_sfixed(657611143.0/4294967296.0,1,-nbitq), 
to_sfixed(151598193.0/4294967296.0,1,-nbitq), 
to_sfixed(-414847510.0/4294967296.0,1,-nbitq), 
to_sfixed(-93123340.0/4294967296.0,1,-nbitq), 
to_sfixed(512391952.0/4294967296.0,1,-nbitq), 
to_sfixed(-1413895886.0/4294967296.0,1,-nbitq), 
to_sfixed(366683879.0/4294967296.0,1,-nbitq), 
to_sfixed(-667238193.0/4294967296.0,1,-nbitq), 
to_sfixed(379620531.0/4294967296.0,1,-nbitq), 
to_sfixed(-98587461.0/4294967296.0,1,-nbitq), 
to_sfixed(882194396.0/4294967296.0,1,-nbitq), 
to_sfixed(348724365.0/4294967296.0,1,-nbitq), 
to_sfixed(-385700642.0/4294967296.0,1,-nbitq), 
to_sfixed(212009063.0/4294967296.0,1,-nbitq), 
to_sfixed(-471512354.0/4294967296.0,1,-nbitq), 
to_sfixed(378131827.0/4294967296.0,1,-nbitq), 
to_sfixed(-205205717.0/4294967296.0,1,-nbitq), 
to_sfixed(101322845.0/4294967296.0,1,-nbitq), 
to_sfixed(134058669.0/4294967296.0,1,-nbitq), 
to_sfixed(382037529.0/4294967296.0,1,-nbitq), 
to_sfixed(361252524.0/4294967296.0,1,-nbitq), 
to_sfixed(-622595150.0/4294967296.0,1,-nbitq), 
to_sfixed(891762272.0/4294967296.0,1,-nbitq), 
to_sfixed(-1071907918.0/4294967296.0,1,-nbitq), 
to_sfixed(435195811.0/4294967296.0,1,-nbitq), 
to_sfixed(459416694.0/4294967296.0,1,-nbitq), 
to_sfixed(-1089178938.0/4294967296.0,1,-nbitq), 
to_sfixed(432204179.0/4294967296.0,1,-nbitq), 
to_sfixed(831503571.0/4294967296.0,1,-nbitq), 
to_sfixed(-571495641.0/4294967296.0,1,-nbitq), 
to_sfixed(91357543.0/4294967296.0,1,-nbitq), 
to_sfixed(57308730.0/4294967296.0,1,-nbitq), 
to_sfixed(-609043050.0/4294967296.0,1,-nbitq), 
to_sfixed(-421883903.0/4294967296.0,1,-nbitq), 
to_sfixed(-413850969.0/4294967296.0,1,-nbitq), 
to_sfixed(-769260578.0/4294967296.0,1,-nbitq), 
to_sfixed(203751991.0/4294967296.0,1,-nbitq), 
to_sfixed(-644914242.0/4294967296.0,1,-nbitq), 
to_sfixed(-152076420.0/4294967296.0,1,-nbitq), 
to_sfixed(-362662937.0/4294967296.0,1,-nbitq), 
to_sfixed(-298167955.0/4294967296.0,1,-nbitq), 
to_sfixed(-809493490.0/4294967296.0,1,-nbitq), 
to_sfixed(-289677446.0/4294967296.0,1,-nbitq), 
to_sfixed(489590822.0/4294967296.0,1,-nbitq), 
to_sfixed(762402282.0/4294967296.0,1,-nbitq), 
to_sfixed(273447632.0/4294967296.0,1,-nbitq), 
to_sfixed(-475654791.0/4294967296.0,1,-nbitq), 
to_sfixed(820615574.0/4294967296.0,1,-nbitq), 
to_sfixed(31586917.0/4294967296.0,1,-nbitq), 
to_sfixed(591542898.0/4294967296.0,1,-nbitq), 
to_sfixed(152878448.0/4294967296.0,1,-nbitq), 
to_sfixed(61193345.0/4294967296.0,1,-nbitq), 
to_sfixed(-197138547.0/4294967296.0,1,-nbitq), 
to_sfixed(94841748.0/4294967296.0,1,-nbitq), 
to_sfixed(-331962826.0/4294967296.0,1,-nbitq), 
to_sfixed(1535869850.0/4294967296.0,1,-nbitq), 
to_sfixed(96706892.0/4294967296.0,1,-nbitq), 
to_sfixed(-131378466.0/4294967296.0,1,-nbitq), 
to_sfixed(-442465801.0/4294967296.0,1,-nbitq), 
to_sfixed(-88647740.0/4294967296.0,1,-nbitq), 
to_sfixed(-285080265.0/4294967296.0,1,-nbitq), 
to_sfixed(-77037522.0/4294967296.0,1,-nbitq), 
to_sfixed(-1197212639.0/4294967296.0,1,-nbitq), 
to_sfixed(-4763473.0/4294967296.0,1,-nbitq), 
to_sfixed(-131629431.0/4294967296.0,1,-nbitq), 
to_sfixed(435547393.0/4294967296.0,1,-nbitq), 
to_sfixed(129861950.0/4294967296.0,1,-nbitq), 
to_sfixed(-347231063.0/4294967296.0,1,-nbitq), 
to_sfixed(1050811961.0/4294967296.0,1,-nbitq), 
to_sfixed(455599917.0/4294967296.0,1,-nbitq), 
to_sfixed(-424102058.0/4294967296.0,1,-nbitq), 
to_sfixed(137990444.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-136054953.0/4294967296.0,1,-nbitq), 
to_sfixed(-469811467.0/4294967296.0,1,-nbitq), 
to_sfixed(473059860.0/4294967296.0,1,-nbitq), 
to_sfixed(401046483.0/4294967296.0,1,-nbitq), 
to_sfixed(878070674.0/4294967296.0,1,-nbitq), 
to_sfixed(-418302175.0/4294967296.0,1,-nbitq), 
to_sfixed(-457032157.0/4294967296.0,1,-nbitq), 
to_sfixed(-1108378459.0/4294967296.0,1,-nbitq), 
to_sfixed(1073931049.0/4294967296.0,1,-nbitq), 
to_sfixed(359328415.0/4294967296.0,1,-nbitq), 
to_sfixed(-183757934.0/4294967296.0,1,-nbitq), 
to_sfixed(88548456.0/4294967296.0,1,-nbitq), 
to_sfixed(97337590.0/4294967296.0,1,-nbitq), 
to_sfixed(-1718411033.0/4294967296.0,1,-nbitq), 
to_sfixed(-198983933.0/4294967296.0,1,-nbitq), 
to_sfixed(-726736128.0/4294967296.0,1,-nbitq), 
to_sfixed(357135103.0/4294967296.0,1,-nbitq), 
to_sfixed(-309395762.0/4294967296.0,1,-nbitq), 
to_sfixed(1049916747.0/4294967296.0,1,-nbitq), 
to_sfixed(106224247.0/4294967296.0,1,-nbitq), 
to_sfixed(-192866144.0/4294967296.0,1,-nbitq), 
to_sfixed(439517539.0/4294967296.0,1,-nbitq), 
to_sfixed(-411576757.0/4294967296.0,1,-nbitq), 
to_sfixed(-392967193.0/4294967296.0,1,-nbitq), 
to_sfixed(321228360.0/4294967296.0,1,-nbitq), 
to_sfixed(-552314053.0/4294967296.0,1,-nbitq), 
to_sfixed(-48613467.0/4294967296.0,1,-nbitq), 
to_sfixed(903675332.0/4294967296.0,1,-nbitq), 
to_sfixed(868881028.0/4294967296.0,1,-nbitq), 
to_sfixed(-1335902972.0/4294967296.0,1,-nbitq), 
to_sfixed(1545181786.0/4294967296.0,1,-nbitq), 
to_sfixed(-206851679.0/4294967296.0,1,-nbitq), 
to_sfixed(702314153.0/4294967296.0,1,-nbitq), 
to_sfixed(71806483.0/4294967296.0,1,-nbitq), 
to_sfixed(-787400817.0/4294967296.0,1,-nbitq), 
to_sfixed(160330029.0/4294967296.0,1,-nbitq), 
to_sfixed(621495110.0/4294967296.0,1,-nbitq), 
to_sfixed(-66415887.0/4294967296.0,1,-nbitq), 
to_sfixed(385367567.0/4294967296.0,1,-nbitq), 
to_sfixed(269861651.0/4294967296.0,1,-nbitq), 
to_sfixed(-613508755.0/4294967296.0,1,-nbitq), 
to_sfixed(-140204058.0/4294967296.0,1,-nbitq), 
to_sfixed(475307334.0/4294967296.0,1,-nbitq), 
to_sfixed(68552328.0/4294967296.0,1,-nbitq), 
to_sfixed(-367727547.0/4294967296.0,1,-nbitq), 
to_sfixed(-1113799755.0/4294967296.0,1,-nbitq), 
to_sfixed(-141347007.0/4294967296.0,1,-nbitq), 
to_sfixed(-685771086.0/4294967296.0,1,-nbitq), 
to_sfixed(-29497669.0/4294967296.0,1,-nbitq), 
to_sfixed(-438365389.0/4294967296.0,1,-nbitq), 
to_sfixed(-132110757.0/4294967296.0,1,-nbitq), 
to_sfixed(248460088.0/4294967296.0,1,-nbitq), 
to_sfixed(409358453.0/4294967296.0,1,-nbitq), 
to_sfixed(1266914789.0/4294967296.0,1,-nbitq), 
to_sfixed(-787091250.0/4294967296.0,1,-nbitq), 
to_sfixed(-18012927.0/4294967296.0,1,-nbitq), 
to_sfixed(90983545.0/4294967296.0,1,-nbitq), 
to_sfixed(628649531.0/4294967296.0,1,-nbitq), 
to_sfixed(182648159.0/4294967296.0,1,-nbitq), 
to_sfixed(309649659.0/4294967296.0,1,-nbitq), 
to_sfixed(87997448.0/4294967296.0,1,-nbitq), 
to_sfixed(160022396.0/4294967296.0,1,-nbitq), 
to_sfixed(59621987.0/4294967296.0,1,-nbitq), 
to_sfixed(655987596.0/4294967296.0,1,-nbitq), 
to_sfixed(5125570.0/4294967296.0,1,-nbitq), 
to_sfixed(-338139789.0/4294967296.0,1,-nbitq), 
to_sfixed(121087743.0/4294967296.0,1,-nbitq), 
to_sfixed(-423207047.0/4294967296.0,1,-nbitq), 
to_sfixed(-289390897.0/4294967296.0,1,-nbitq), 
to_sfixed(438683892.0/4294967296.0,1,-nbitq), 
to_sfixed(-1139980320.0/4294967296.0,1,-nbitq), 
to_sfixed(156945024.0/4294967296.0,1,-nbitq), 
to_sfixed(-475395249.0/4294967296.0,1,-nbitq), 
to_sfixed(-238675773.0/4294967296.0,1,-nbitq), 
to_sfixed(86847675.0/4294967296.0,1,-nbitq), 
to_sfixed(377381160.0/4294967296.0,1,-nbitq), 
to_sfixed(941391474.0/4294967296.0,1,-nbitq), 
to_sfixed(851195174.0/4294967296.0,1,-nbitq), 
to_sfixed(-774277051.0/4294967296.0,1,-nbitq), 
to_sfixed(-137043390.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-493232622.0/4294967296.0,1,-nbitq), 
to_sfixed(-627146928.0/4294967296.0,1,-nbitq), 
to_sfixed(80227220.0/4294967296.0,1,-nbitq), 
to_sfixed(605505761.0/4294967296.0,1,-nbitq), 
to_sfixed(401937020.0/4294967296.0,1,-nbitq), 
to_sfixed(-677017799.0/4294967296.0,1,-nbitq), 
to_sfixed(-488897341.0/4294967296.0,1,-nbitq), 
to_sfixed(-1114893372.0/4294967296.0,1,-nbitq), 
to_sfixed(1365806393.0/4294967296.0,1,-nbitq), 
to_sfixed(228464886.0/4294967296.0,1,-nbitq), 
to_sfixed(-514030731.0/4294967296.0,1,-nbitq), 
to_sfixed(-826598234.0/4294967296.0,1,-nbitq), 
to_sfixed(-395455962.0/4294967296.0,1,-nbitq), 
to_sfixed(-831320389.0/4294967296.0,1,-nbitq), 
to_sfixed(340680426.0/4294967296.0,1,-nbitq), 
to_sfixed(-1232614611.0/4294967296.0,1,-nbitq), 
to_sfixed(133690553.0/4294967296.0,1,-nbitq), 
to_sfixed(366889077.0/4294967296.0,1,-nbitq), 
to_sfixed(918950360.0/4294967296.0,1,-nbitq), 
to_sfixed(-612024472.0/4294967296.0,1,-nbitq), 
to_sfixed(-284304927.0/4294967296.0,1,-nbitq), 
to_sfixed(520779109.0/4294967296.0,1,-nbitq), 
to_sfixed(-487380223.0/4294967296.0,1,-nbitq), 
to_sfixed(25787317.0/4294967296.0,1,-nbitq), 
to_sfixed(132653499.0/4294967296.0,1,-nbitq), 
to_sfixed(-182614565.0/4294967296.0,1,-nbitq), 
to_sfixed(-268544377.0/4294967296.0,1,-nbitq), 
to_sfixed(276379107.0/4294967296.0,1,-nbitq), 
to_sfixed(634246265.0/4294967296.0,1,-nbitq), 
to_sfixed(-1098439987.0/4294967296.0,1,-nbitq), 
to_sfixed(638382739.0/4294967296.0,1,-nbitq), 
to_sfixed(245156454.0/4294967296.0,1,-nbitq), 
to_sfixed(115886060.0/4294967296.0,1,-nbitq), 
to_sfixed(285348178.0/4294967296.0,1,-nbitq), 
to_sfixed(-285014441.0/4294967296.0,1,-nbitq), 
to_sfixed(182883596.0/4294967296.0,1,-nbitq), 
to_sfixed(-524877439.0/4294967296.0,1,-nbitq), 
to_sfixed(-932580377.0/4294967296.0,1,-nbitq), 
to_sfixed(206387484.0/4294967296.0,1,-nbitq), 
to_sfixed(602059824.0/4294967296.0,1,-nbitq), 
to_sfixed(347247660.0/4294967296.0,1,-nbitq), 
to_sfixed(-567463374.0/4294967296.0,1,-nbitq), 
to_sfixed(641791194.0/4294967296.0,1,-nbitq), 
to_sfixed(-682126724.0/4294967296.0,1,-nbitq), 
to_sfixed(187389637.0/4294967296.0,1,-nbitq), 
to_sfixed(-1131007451.0/4294967296.0,1,-nbitq), 
to_sfixed(-53068144.0/4294967296.0,1,-nbitq), 
to_sfixed(-616131759.0/4294967296.0,1,-nbitq), 
to_sfixed(-203592731.0/4294967296.0,1,-nbitq), 
to_sfixed(85310042.0/4294967296.0,1,-nbitq), 
to_sfixed(-498737956.0/4294967296.0,1,-nbitq), 
to_sfixed(-250094787.0/4294967296.0,1,-nbitq), 
to_sfixed(211006017.0/4294967296.0,1,-nbitq), 
to_sfixed(872205290.0/4294967296.0,1,-nbitq), 
to_sfixed(-1490723978.0/4294967296.0,1,-nbitq), 
to_sfixed(299109320.0/4294967296.0,1,-nbitq), 
to_sfixed(-418663510.0/4294967296.0,1,-nbitq), 
to_sfixed(176494378.0/4294967296.0,1,-nbitq), 
to_sfixed(53210017.0/4294967296.0,1,-nbitq), 
to_sfixed(290679597.0/4294967296.0,1,-nbitq), 
to_sfixed(235061040.0/4294967296.0,1,-nbitq), 
to_sfixed(381893426.0/4294967296.0,1,-nbitq), 
to_sfixed(313304126.0/4294967296.0,1,-nbitq), 
to_sfixed(558785607.0/4294967296.0,1,-nbitq), 
to_sfixed(243825370.0/4294967296.0,1,-nbitq), 
to_sfixed(-284502612.0/4294967296.0,1,-nbitq), 
to_sfixed(702217344.0/4294967296.0,1,-nbitq), 
to_sfixed(-854316411.0/4294967296.0,1,-nbitq), 
to_sfixed(100126833.0/4294967296.0,1,-nbitq), 
to_sfixed(-72345586.0/4294967296.0,1,-nbitq), 
to_sfixed(-2231417568.0/4294967296.0,1,-nbitq), 
to_sfixed(-201698737.0/4294967296.0,1,-nbitq), 
to_sfixed(418502271.0/4294967296.0,1,-nbitq), 
to_sfixed(288779803.0/4294967296.0,1,-nbitq), 
to_sfixed(-83397518.0/4294967296.0,1,-nbitq), 
to_sfixed(436323901.0/4294967296.0,1,-nbitq), 
to_sfixed(983100028.0/4294967296.0,1,-nbitq), 
to_sfixed(290531297.0/4294967296.0,1,-nbitq), 
to_sfixed(-674560238.0/4294967296.0,1,-nbitq), 
to_sfixed(-318727067.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-717454835.0/4294967296.0,1,-nbitq), 
to_sfixed(-1506566325.0/4294967296.0,1,-nbitq), 
to_sfixed(740991066.0/4294967296.0,1,-nbitq), 
to_sfixed(835649744.0/4294967296.0,1,-nbitq), 
to_sfixed(127191908.0/4294967296.0,1,-nbitq), 
to_sfixed(-304370269.0/4294967296.0,1,-nbitq), 
to_sfixed(-438582570.0/4294967296.0,1,-nbitq), 
to_sfixed(-73616114.0/4294967296.0,1,-nbitq), 
to_sfixed(977032007.0/4294967296.0,1,-nbitq), 
to_sfixed(-182630442.0/4294967296.0,1,-nbitq), 
to_sfixed(-705011141.0/4294967296.0,1,-nbitq), 
to_sfixed(-359093322.0/4294967296.0,1,-nbitq), 
to_sfixed(-197230075.0/4294967296.0,1,-nbitq), 
to_sfixed(-1029164058.0/4294967296.0,1,-nbitq), 
to_sfixed(-176294196.0/4294967296.0,1,-nbitq), 
to_sfixed(-1402812445.0/4294967296.0,1,-nbitq), 
to_sfixed(89418079.0/4294967296.0,1,-nbitq), 
to_sfixed(-219442878.0/4294967296.0,1,-nbitq), 
to_sfixed(413366657.0/4294967296.0,1,-nbitq), 
to_sfixed(-455957044.0/4294967296.0,1,-nbitq), 
to_sfixed(243493883.0/4294967296.0,1,-nbitq), 
to_sfixed(1067437105.0/4294967296.0,1,-nbitq), 
to_sfixed(-398871457.0/4294967296.0,1,-nbitq), 
to_sfixed(132603068.0/4294967296.0,1,-nbitq), 
to_sfixed(213730824.0/4294967296.0,1,-nbitq), 
to_sfixed(1015851807.0/4294967296.0,1,-nbitq), 
to_sfixed(-858385508.0/4294967296.0,1,-nbitq), 
to_sfixed(761905329.0/4294967296.0,1,-nbitq), 
to_sfixed(-710124815.0/4294967296.0,1,-nbitq), 
to_sfixed(-540847709.0/4294967296.0,1,-nbitq), 
to_sfixed(1037873789.0/4294967296.0,1,-nbitq), 
to_sfixed(691604596.0/4294967296.0,1,-nbitq), 
to_sfixed(-121462266.0/4294967296.0,1,-nbitq), 
to_sfixed(-154186785.0/4294967296.0,1,-nbitq), 
to_sfixed(589257575.0/4294967296.0,1,-nbitq), 
to_sfixed(1012832206.0/4294967296.0,1,-nbitq), 
to_sfixed(-621973952.0/4294967296.0,1,-nbitq), 
to_sfixed(-1338238265.0/4294967296.0,1,-nbitq), 
to_sfixed(535275340.0/4294967296.0,1,-nbitq), 
to_sfixed(267268177.0/4294967296.0,1,-nbitq), 
to_sfixed(39794950.0/4294967296.0,1,-nbitq), 
to_sfixed(-230708285.0/4294967296.0,1,-nbitq), 
to_sfixed(1756240506.0/4294967296.0,1,-nbitq), 
to_sfixed(-243383834.0/4294967296.0,1,-nbitq), 
to_sfixed(118197927.0/4294967296.0,1,-nbitq), 
to_sfixed(-1142748115.0/4294967296.0,1,-nbitq), 
to_sfixed(-306044041.0/4294967296.0,1,-nbitq), 
to_sfixed(-1354366698.0/4294967296.0,1,-nbitq), 
to_sfixed(-395125003.0/4294967296.0,1,-nbitq), 
to_sfixed(84261387.0/4294967296.0,1,-nbitq), 
to_sfixed(-70182790.0/4294967296.0,1,-nbitq), 
to_sfixed(628301198.0/4294967296.0,1,-nbitq), 
to_sfixed(-829530524.0/4294967296.0,1,-nbitq), 
to_sfixed(1395441381.0/4294967296.0,1,-nbitq), 
to_sfixed(-430465518.0/4294967296.0,1,-nbitq), 
to_sfixed(650360443.0/4294967296.0,1,-nbitq), 
to_sfixed(-214776955.0/4294967296.0,1,-nbitq), 
to_sfixed(-207364062.0/4294967296.0,1,-nbitq), 
to_sfixed(-355708038.0/4294967296.0,1,-nbitq), 
to_sfixed(346756479.0/4294967296.0,1,-nbitq), 
to_sfixed(-82272100.0/4294967296.0,1,-nbitq), 
to_sfixed(236910771.0/4294967296.0,1,-nbitq), 
to_sfixed(-43065341.0/4294967296.0,1,-nbitq), 
to_sfixed(968874774.0/4294967296.0,1,-nbitq), 
to_sfixed(-230710947.0/4294967296.0,1,-nbitq), 
to_sfixed(399701979.0/4294967296.0,1,-nbitq), 
to_sfixed(-28441259.0/4294967296.0,1,-nbitq), 
to_sfixed(-1174194284.0/4294967296.0,1,-nbitq), 
to_sfixed(-312631316.0/4294967296.0,1,-nbitq), 
to_sfixed(69957412.0/4294967296.0,1,-nbitq), 
to_sfixed(-921851166.0/4294967296.0,1,-nbitq), 
to_sfixed(407283904.0/4294967296.0,1,-nbitq), 
to_sfixed(70697894.0/4294967296.0,1,-nbitq), 
to_sfixed(10029893.0/4294967296.0,1,-nbitq), 
to_sfixed(-263861649.0/4294967296.0,1,-nbitq), 
to_sfixed(682471770.0/4294967296.0,1,-nbitq), 
to_sfixed(1735584454.0/4294967296.0,1,-nbitq), 
to_sfixed(536204982.0/4294967296.0,1,-nbitq), 
to_sfixed(-567944174.0/4294967296.0,1,-nbitq), 
to_sfixed(268656348.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-249874706.0/4294967296.0,1,-nbitq), 
to_sfixed(-271073181.0/4294967296.0,1,-nbitq), 
to_sfixed(512925482.0/4294967296.0,1,-nbitq), 
to_sfixed(635766290.0/4294967296.0,1,-nbitq), 
to_sfixed(460931273.0/4294967296.0,1,-nbitq), 
to_sfixed(-377945325.0/4294967296.0,1,-nbitq), 
to_sfixed(-136176710.0/4294967296.0,1,-nbitq), 
to_sfixed(500883064.0/4294967296.0,1,-nbitq), 
to_sfixed(663321505.0/4294967296.0,1,-nbitq), 
to_sfixed(-45191400.0/4294967296.0,1,-nbitq), 
to_sfixed(-328377229.0/4294967296.0,1,-nbitq), 
to_sfixed(-330578578.0/4294967296.0,1,-nbitq), 
to_sfixed(-282153870.0/4294967296.0,1,-nbitq), 
to_sfixed(-1123670482.0/4294967296.0,1,-nbitq), 
to_sfixed(-10120718.0/4294967296.0,1,-nbitq), 
to_sfixed(-409465740.0/4294967296.0,1,-nbitq), 
to_sfixed(-261265287.0/4294967296.0,1,-nbitq), 
to_sfixed(-229463569.0/4294967296.0,1,-nbitq), 
to_sfixed(384442452.0/4294967296.0,1,-nbitq), 
to_sfixed(-106461126.0/4294967296.0,1,-nbitq), 
to_sfixed(-211785584.0/4294967296.0,1,-nbitq), 
to_sfixed(900719591.0/4294967296.0,1,-nbitq), 
to_sfixed(370556247.0/4294967296.0,1,-nbitq), 
to_sfixed(-634281827.0/4294967296.0,1,-nbitq), 
to_sfixed(372719741.0/4294967296.0,1,-nbitq), 
to_sfixed(292327165.0/4294967296.0,1,-nbitq), 
to_sfixed(21552239.0/4294967296.0,1,-nbitq), 
to_sfixed(138150623.0/4294967296.0,1,-nbitq), 
to_sfixed(-765487601.0/4294967296.0,1,-nbitq), 
to_sfixed(-176066057.0/4294967296.0,1,-nbitq), 
to_sfixed(366064687.0/4294967296.0,1,-nbitq), 
to_sfixed(811029977.0/4294967296.0,1,-nbitq), 
to_sfixed(-355939168.0/4294967296.0,1,-nbitq), 
to_sfixed(176011895.0/4294967296.0,1,-nbitq), 
to_sfixed(-17218569.0/4294967296.0,1,-nbitq), 
to_sfixed(798558817.0/4294967296.0,1,-nbitq), 
to_sfixed(-999078011.0/4294967296.0,1,-nbitq), 
to_sfixed(-343326633.0/4294967296.0,1,-nbitq), 
to_sfixed(190586984.0/4294967296.0,1,-nbitq), 
to_sfixed(261734992.0/4294967296.0,1,-nbitq), 
to_sfixed(-498742101.0/4294967296.0,1,-nbitq), 
to_sfixed(143731542.0/4294967296.0,1,-nbitq), 
to_sfixed(722702056.0/4294967296.0,1,-nbitq), 
to_sfixed(-168333296.0/4294967296.0,1,-nbitq), 
to_sfixed(-398127997.0/4294967296.0,1,-nbitq), 
to_sfixed(-1557286538.0/4294967296.0,1,-nbitq), 
to_sfixed(294010749.0/4294967296.0,1,-nbitq), 
to_sfixed(-694536520.0/4294967296.0,1,-nbitq), 
to_sfixed(111108117.0/4294967296.0,1,-nbitq), 
to_sfixed(-26046154.0/4294967296.0,1,-nbitq), 
to_sfixed(208530954.0/4294967296.0,1,-nbitq), 
to_sfixed(305130479.0/4294967296.0,1,-nbitq), 
to_sfixed(-925307235.0/4294967296.0,1,-nbitq), 
to_sfixed(1414636059.0/4294967296.0,1,-nbitq), 
to_sfixed(176388317.0/4294967296.0,1,-nbitq), 
to_sfixed(1223637033.0/4294967296.0,1,-nbitq), 
to_sfixed(-178718878.0/4294967296.0,1,-nbitq), 
to_sfixed(-635216576.0/4294967296.0,1,-nbitq), 
to_sfixed(-86271658.0/4294967296.0,1,-nbitq), 
to_sfixed(99054117.0/4294967296.0,1,-nbitq), 
to_sfixed(13425476.0/4294967296.0,1,-nbitq), 
to_sfixed(-244378703.0/4294967296.0,1,-nbitq), 
to_sfixed(388727990.0/4294967296.0,1,-nbitq), 
to_sfixed(955209466.0/4294967296.0,1,-nbitq), 
to_sfixed(500815537.0/4294967296.0,1,-nbitq), 
to_sfixed(403267971.0/4294967296.0,1,-nbitq), 
to_sfixed(358232310.0/4294967296.0,1,-nbitq), 
to_sfixed(-615173666.0/4294967296.0,1,-nbitq), 
to_sfixed(-265600486.0/4294967296.0,1,-nbitq), 
to_sfixed(-772688762.0/4294967296.0,1,-nbitq), 
to_sfixed(-1107017847.0/4294967296.0,1,-nbitq), 
to_sfixed(167967369.0/4294967296.0,1,-nbitq), 
to_sfixed(655690760.0/4294967296.0,1,-nbitq), 
to_sfixed(-385765642.0/4294967296.0,1,-nbitq), 
to_sfixed(41654288.0/4294967296.0,1,-nbitq), 
to_sfixed(894214072.0/4294967296.0,1,-nbitq), 
to_sfixed(1719071822.0/4294967296.0,1,-nbitq), 
to_sfixed(458379595.0/4294967296.0,1,-nbitq), 
to_sfixed(322736087.0/4294967296.0,1,-nbitq), 
to_sfixed(-223197777.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-236567231.0/4294967296.0,1,-nbitq), 
to_sfixed(203863276.0/4294967296.0,1,-nbitq), 
to_sfixed(1139463798.0/4294967296.0,1,-nbitq), 
to_sfixed(171835056.0/4294967296.0,1,-nbitq), 
to_sfixed(370378912.0/4294967296.0,1,-nbitq), 
to_sfixed(-276823851.0/4294967296.0,1,-nbitq), 
to_sfixed(206036701.0/4294967296.0,1,-nbitq), 
to_sfixed(360722735.0/4294967296.0,1,-nbitq), 
to_sfixed(867024945.0/4294967296.0,1,-nbitq), 
to_sfixed(93231640.0/4294967296.0,1,-nbitq), 
to_sfixed(596025761.0/4294967296.0,1,-nbitq), 
to_sfixed(-308279676.0/4294967296.0,1,-nbitq), 
to_sfixed(-17888673.0/4294967296.0,1,-nbitq), 
to_sfixed(-436822734.0/4294967296.0,1,-nbitq), 
to_sfixed(118896609.0/4294967296.0,1,-nbitq), 
to_sfixed(113183671.0/4294967296.0,1,-nbitq), 
to_sfixed(-139266539.0/4294967296.0,1,-nbitq), 
to_sfixed(-232004191.0/4294967296.0,1,-nbitq), 
to_sfixed(-94225719.0/4294967296.0,1,-nbitq), 
to_sfixed(59784297.0/4294967296.0,1,-nbitq), 
to_sfixed(301046130.0/4294967296.0,1,-nbitq), 
to_sfixed(68642696.0/4294967296.0,1,-nbitq), 
to_sfixed(944518141.0/4294967296.0,1,-nbitq), 
to_sfixed(-1374568286.0/4294967296.0,1,-nbitq), 
to_sfixed(105305378.0/4294967296.0,1,-nbitq), 
to_sfixed(254636263.0/4294967296.0,1,-nbitq), 
to_sfixed(435965520.0/4294967296.0,1,-nbitq), 
to_sfixed(-207518866.0/4294967296.0,1,-nbitq), 
to_sfixed(-1516779760.0/4294967296.0,1,-nbitq), 
to_sfixed(-408591685.0/4294967296.0,1,-nbitq), 
to_sfixed(362202134.0/4294967296.0,1,-nbitq), 
to_sfixed(1137358129.0/4294967296.0,1,-nbitq), 
to_sfixed(-133647424.0/4294967296.0,1,-nbitq), 
to_sfixed(195697325.0/4294967296.0,1,-nbitq), 
to_sfixed(54058178.0/4294967296.0,1,-nbitq), 
to_sfixed(329013342.0/4294967296.0,1,-nbitq), 
to_sfixed(-808195994.0/4294967296.0,1,-nbitq), 
to_sfixed(369041962.0/4294967296.0,1,-nbitq), 
to_sfixed(-200887759.0/4294967296.0,1,-nbitq), 
to_sfixed(-128828579.0/4294967296.0,1,-nbitq), 
to_sfixed(-618900239.0/4294967296.0,1,-nbitq), 
to_sfixed(313031702.0/4294967296.0,1,-nbitq), 
to_sfixed(430738169.0/4294967296.0,1,-nbitq), 
to_sfixed(-172400772.0/4294967296.0,1,-nbitq), 
to_sfixed(-165584025.0/4294967296.0,1,-nbitq), 
to_sfixed(-1849109193.0/4294967296.0,1,-nbitq), 
to_sfixed(-273883321.0/4294967296.0,1,-nbitq), 
to_sfixed(-810643432.0/4294967296.0,1,-nbitq), 
to_sfixed(-408918360.0/4294967296.0,1,-nbitq), 
to_sfixed(751077119.0/4294967296.0,1,-nbitq), 
to_sfixed(311420242.0/4294967296.0,1,-nbitq), 
to_sfixed(195570129.0/4294967296.0,1,-nbitq), 
to_sfixed(123682098.0/4294967296.0,1,-nbitq), 
to_sfixed(509062143.0/4294967296.0,1,-nbitq), 
to_sfixed(605082426.0/4294967296.0,1,-nbitq), 
to_sfixed(410796660.0/4294967296.0,1,-nbitq), 
to_sfixed(-94512789.0/4294967296.0,1,-nbitq), 
to_sfixed(-375447061.0/4294967296.0,1,-nbitq), 
to_sfixed(234890550.0/4294967296.0,1,-nbitq), 
to_sfixed(269178390.0/4294967296.0,1,-nbitq), 
to_sfixed(205174811.0/4294967296.0,1,-nbitq), 
to_sfixed(-216956934.0/4294967296.0,1,-nbitq), 
to_sfixed(556859754.0/4294967296.0,1,-nbitq), 
to_sfixed(836662924.0/4294967296.0,1,-nbitq), 
to_sfixed(1829255.0/4294967296.0,1,-nbitq), 
to_sfixed(-446765120.0/4294967296.0,1,-nbitq), 
to_sfixed(633515422.0/4294967296.0,1,-nbitq), 
to_sfixed(-668680370.0/4294967296.0,1,-nbitq), 
to_sfixed(-224414304.0/4294967296.0,1,-nbitq), 
to_sfixed(-1033730615.0/4294967296.0,1,-nbitq), 
to_sfixed(-963852971.0/4294967296.0,1,-nbitq), 
to_sfixed(-82307272.0/4294967296.0,1,-nbitq), 
to_sfixed(247749250.0/4294967296.0,1,-nbitq), 
to_sfixed(96251297.0/4294967296.0,1,-nbitq), 
to_sfixed(-42613367.0/4294967296.0,1,-nbitq), 
to_sfixed(238838393.0/4294967296.0,1,-nbitq), 
to_sfixed(1565521178.0/4294967296.0,1,-nbitq), 
to_sfixed(-98950069.0/4294967296.0,1,-nbitq), 
to_sfixed(373620026.0/4294967296.0,1,-nbitq), 
to_sfixed(-191625886.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(11331184.0/4294967296.0,1,-nbitq), 
to_sfixed(173385505.0/4294967296.0,1,-nbitq), 
to_sfixed(856434368.0/4294967296.0,1,-nbitq), 
to_sfixed(-545382716.0/4294967296.0,1,-nbitq), 
to_sfixed(263012218.0/4294967296.0,1,-nbitq), 
to_sfixed(-809512799.0/4294967296.0,1,-nbitq), 
to_sfixed(-319903443.0/4294967296.0,1,-nbitq), 
to_sfixed(-135805867.0/4294967296.0,1,-nbitq), 
to_sfixed(321405961.0/4294967296.0,1,-nbitq), 
to_sfixed(-204403878.0/4294967296.0,1,-nbitq), 
to_sfixed(1052862523.0/4294967296.0,1,-nbitq), 
to_sfixed(60614332.0/4294967296.0,1,-nbitq), 
to_sfixed(64905934.0/4294967296.0,1,-nbitq), 
to_sfixed(1164250544.0/4294967296.0,1,-nbitq), 
to_sfixed(-242457986.0/4294967296.0,1,-nbitq), 
to_sfixed(-88302205.0/4294967296.0,1,-nbitq), 
to_sfixed(-308392848.0/4294967296.0,1,-nbitq), 
to_sfixed(141578253.0/4294967296.0,1,-nbitq), 
to_sfixed(89350673.0/4294967296.0,1,-nbitq), 
to_sfixed(-192633597.0/4294967296.0,1,-nbitq), 
to_sfixed(44084698.0/4294967296.0,1,-nbitq), 
to_sfixed(-725700590.0/4294967296.0,1,-nbitq), 
to_sfixed(325576978.0/4294967296.0,1,-nbitq), 
to_sfixed(-1547989136.0/4294967296.0,1,-nbitq), 
to_sfixed(382756295.0/4294967296.0,1,-nbitq), 
to_sfixed(-126520988.0/4294967296.0,1,-nbitq), 
to_sfixed(239929561.0/4294967296.0,1,-nbitq), 
to_sfixed(-1122697683.0/4294967296.0,1,-nbitq), 
to_sfixed(-1124211695.0/4294967296.0,1,-nbitq), 
to_sfixed(-738936714.0/4294967296.0,1,-nbitq), 
to_sfixed(-560417564.0/4294967296.0,1,-nbitq), 
to_sfixed(787492543.0/4294967296.0,1,-nbitq), 
to_sfixed(-64627245.0/4294967296.0,1,-nbitq), 
to_sfixed(-424712939.0/4294967296.0,1,-nbitq), 
to_sfixed(372187485.0/4294967296.0,1,-nbitq), 
to_sfixed(-126173631.0/4294967296.0,1,-nbitq), 
to_sfixed(-479331865.0/4294967296.0,1,-nbitq), 
to_sfixed(-327234771.0/4294967296.0,1,-nbitq), 
to_sfixed(-121547765.0/4294967296.0,1,-nbitq), 
to_sfixed(-375515123.0/4294967296.0,1,-nbitq), 
to_sfixed(-251693715.0/4294967296.0,1,-nbitq), 
to_sfixed(-145778946.0/4294967296.0,1,-nbitq), 
to_sfixed(512080017.0/4294967296.0,1,-nbitq), 
to_sfixed(-315835300.0/4294967296.0,1,-nbitq), 
to_sfixed(-396951035.0/4294967296.0,1,-nbitq), 
to_sfixed(-1664372389.0/4294967296.0,1,-nbitq), 
to_sfixed(103475861.0/4294967296.0,1,-nbitq), 
to_sfixed(-1257389727.0/4294967296.0,1,-nbitq), 
to_sfixed(373746249.0/4294967296.0,1,-nbitq), 
to_sfixed(579758607.0/4294967296.0,1,-nbitq), 
to_sfixed(116971120.0/4294967296.0,1,-nbitq), 
to_sfixed(-84751728.0/4294967296.0,1,-nbitq), 
to_sfixed(-117137542.0/4294967296.0,1,-nbitq), 
to_sfixed(188886024.0/4294967296.0,1,-nbitq), 
to_sfixed(1100419915.0/4294967296.0,1,-nbitq), 
to_sfixed(-1153481002.0/4294967296.0,1,-nbitq), 
to_sfixed(-45801595.0/4294967296.0,1,-nbitq), 
to_sfixed(-67847365.0/4294967296.0,1,-nbitq), 
to_sfixed(150093843.0/4294967296.0,1,-nbitq), 
to_sfixed(-346875744.0/4294967296.0,1,-nbitq), 
to_sfixed(-332400514.0/4294967296.0,1,-nbitq), 
to_sfixed(-146830261.0/4294967296.0,1,-nbitq), 
to_sfixed(1036159011.0/4294967296.0,1,-nbitq), 
to_sfixed(929776428.0/4294967296.0,1,-nbitq), 
to_sfixed(-94000965.0/4294967296.0,1,-nbitq), 
to_sfixed(-516098860.0/4294967296.0,1,-nbitq), 
to_sfixed(-494231557.0/4294967296.0,1,-nbitq), 
to_sfixed(-1020641951.0/4294967296.0,1,-nbitq), 
to_sfixed(32403009.0/4294967296.0,1,-nbitq), 
to_sfixed(-1420744587.0/4294967296.0,1,-nbitq), 
to_sfixed(-201175220.0/4294967296.0,1,-nbitq), 
to_sfixed(298221079.0/4294967296.0,1,-nbitq), 
to_sfixed(-178731855.0/4294967296.0,1,-nbitq), 
to_sfixed(223274763.0/4294967296.0,1,-nbitq), 
to_sfixed(-261127965.0/4294967296.0,1,-nbitq), 
to_sfixed(610621353.0/4294967296.0,1,-nbitq), 
to_sfixed(833439267.0/4294967296.0,1,-nbitq), 
to_sfixed(-126360779.0/4294967296.0,1,-nbitq), 
to_sfixed(188267881.0/4294967296.0,1,-nbitq), 
to_sfixed(118415159.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-153917700.0/4294967296.0,1,-nbitq), 
to_sfixed(260685033.0/4294967296.0,1,-nbitq), 
to_sfixed(-44780563.0/4294967296.0,1,-nbitq), 
to_sfixed(-757485659.0/4294967296.0,1,-nbitq), 
to_sfixed(-538246079.0/4294967296.0,1,-nbitq), 
to_sfixed(-1605427444.0/4294967296.0,1,-nbitq), 
to_sfixed(85571507.0/4294967296.0,1,-nbitq), 
to_sfixed(-80658109.0/4294967296.0,1,-nbitq), 
to_sfixed(626562665.0/4294967296.0,1,-nbitq), 
to_sfixed(18399204.0/4294967296.0,1,-nbitq), 
to_sfixed(546185479.0/4294967296.0,1,-nbitq), 
to_sfixed(-499860302.0/4294967296.0,1,-nbitq), 
to_sfixed(52168025.0/4294967296.0,1,-nbitq), 
to_sfixed(1537694527.0/4294967296.0,1,-nbitq), 
to_sfixed(186882641.0/4294967296.0,1,-nbitq), 
to_sfixed(-595361184.0/4294967296.0,1,-nbitq), 
to_sfixed(-177497553.0/4294967296.0,1,-nbitq), 
to_sfixed(97527039.0/4294967296.0,1,-nbitq), 
to_sfixed(-349723198.0/4294967296.0,1,-nbitq), 
to_sfixed(203117556.0/4294967296.0,1,-nbitq), 
to_sfixed(120350255.0/4294967296.0,1,-nbitq), 
to_sfixed(-44888569.0/4294967296.0,1,-nbitq), 
to_sfixed(656111101.0/4294967296.0,1,-nbitq), 
to_sfixed(-447749580.0/4294967296.0,1,-nbitq), 
to_sfixed(-241726520.0/4294967296.0,1,-nbitq), 
to_sfixed(-413288483.0/4294967296.0,1,-nbitq), 
to_sfixed(-213077173.0/4294967296.0,1,-nbitq), 
to_sfixed(-980716117.0/4294967296.0,1,-nbitq), 
to_sfixed(50389587.0/4294967296.0,1,-nbitq), 
to_sfixed(-1442619121.0/4294967296.0,1,-nbitq), 
to_sfixed(-616575595.0/4294967296.0,1,-nbitq), 
to_sfixed(313936337.0/4294967296.0,1,-nbitq), 
to_sfixed(-278284124.0/4294967296.0,1,-nbitq), 
to_sfixed(-185457839.0/4294967296.0,1,-nbitq), 
to_sfixed(497434726.0/4294967296.0,1,-nbitq), 
to_sfixed(199642948.0/4294967296.0,1,-nbitq), 
to_sfixed(59496877.0/4294967296.0,1,-nbitq), 
to_sfixed(-119282753.0/4294967296.0,1,-nbitq), 
to_sfixed(259991499.0/4294967296.0,1,-nbitq), 
to_sfixed(-174603995.0/4294967296.0,1,-nbitq), 
to_sfixed(-191478714.0/4294967296.0,1,-nbitq), 
to_sfixed(542687138.0/4294967296.0,1,-nbitq), 
to_sfixed(147967666.0/4294967296.0,1,-nbitq), 
to_sfixed(469487701.0/4294967296.0,1,-nbitq), 
to_sfixed(-613937856.0/4294967296.0,1,-nbitq), 
to_sfixed(-1353838100.0/4294967296.0,1,-nbitq), 
to_sfixed(-320146722.0/4294967296.0,1,-nbitq), 
to_sfixed(-1364264213.0/4294967296.0,1,-nbitq), 
to_sfixed(-183683015.0/4294967296.0,1,-nbitq), 
to_sfixed(378421798.0/4294967296.0,1,-nbitq), 
to_sfixed(-122292289.0/4294967296.0,1,-nbitq), 
to_sfixed(533122812.0/4294967296.0,1,-nbitq), 
to_sfixed(157275911.0/4294967296.0,1,-nbitq), 
to_sfixed(304496134.0/4294967296.0,1,-nbitq), 
to_sfixed(1077015112.0/4294967296.0,1,-nbitq), 
to_sfixed(-790493775.0/4294967296.0,1,-nbitq), 
to_sfixed(142128593.0/4294967296.0,1,-nbitq), 
to_sfixed(706332947.0/4294967296.0,1,-nbitq), 
to_sfixed(200926976.0/4294967296.0,1,-nbitq), 
to_sfixed(-281510727.0/4294967296.0,1,-nbitq), 
to_sfixed(-249974222.0/4294967296.0,1,-nbitq), 
to_sfixed(-463133361.0/4294967296.0,1,-nbitq), 
to_sfixed(601132536.0/4294967296.0,1,-nbitq), 
to_sfixed(704520016.0/4294967296.0,1,-nbitq), 
to_sfixed(-283550822.0/4294967296.0,1,-nbitq), 
to_sfixed(-30328382.0/4294967296.0,1,-nbitq), 
to_sfixed(-543847814.0/4294967296.0,1,-nbitq), 
to_sfixed(-10778515.0/4294967296.0,1,-nbitq), 
to_sfixed(244127793.0/4294967296.0,1,-nbitq), 
to_sfixed(-1316380286.0/4294967296.0,1,-nbitq), 
to_sfixed(396580639.0/4294967296.0,1,-nbitq), 
to_sfixed(555075112.0/4294967296.0,1,-nbitq), 
to_sfixed(-286390600.0/4294967296.0,1,-nbitq), 
to_sfixed(269962271.0/4294967296.0,1,-nbitq), 
to_sfixed(322108277.0/4294967296.0,1,-nbitq), 
to_sfixed(152910016.0/4294967296.0,1,-nbitq), 
to_sfixed(885082839.0/4294967296.0,1,-nbitq), 
to_sfixed(295211666.0/4294967296.0,1,-nbitq), 
to_sfixed(128533860.0/4294967296.0,1,-nbitq), 
to_sfixed(-351081162.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(166200346.0/4294967296.0,1,-nbitq), 
to_sfixed(729495253.0/4294967296.0,1,-nbitq), 
to_sfixed(-565476511.0/4294967296.0,1,-nbitq), 
to_sfixed(-1139039192.0/4294967296.0,1,-nbitq), 
to_sfixed(-492263372.0/4294967296.0,1,-nbitq), 
to_sfixed(-1260224571.0/4294967296.0,1,-nbitq), 
to_sfixed(-45491435.0/4294967296.0,1,-nbitq), 
to_sfixed(-597153691.0/4294967296.0,1,-nbitq), 
to_sfixed(680615918.0/4294967296.0,1,-nbitq), 
to_sfixed(-341413632.0/4294967296.0,1,-nbitq), 
to_sfixed(191317575.0/4294967296.0,1,-nbitq), 
to_sfixed(-910898752.0/4294967296.0,1,-nbitq), 
to_sfixed(-87408079.0/4294967296.0,1,-nbitq), 
to_sfixed(1404053967.0/4294967296.0,1,-nbitq), 
to_sfixed(-115463445.0/4294967296.0,1,-nbitq), 
to_sfixed(599468183.0/4294967296.0,1,-nbitq), 
to_sfixed(-347435492.0/4294967296.0,1,-nbitq), 
to_sfixed(324988893.0/4294967296.0,1,-nbitq), 
to_sfixed(385994042.0/4294967296.0,1,-nbitq), 
to_sfixed(508964839.0/4294967296.0,1,-nbitq), 
to_sfixed(-79900713.0/4294967296.0,1,-nbitq), 
to_sfixed(-215729239.0/4294967296.0,1,-nbitq), 
to_sfixed(239458995.0/4294967296.0,1,-nbitq), 
to_sfixed(-511632962.0/4294967296.0,1,-nbitq), 
to_sfixed(31595696.0/4294967296.0,1,-nbitq), 
to_sfixed(-365266739.0/4294967296.0,1,-nbitq), 
to_sfixed(-182891453.0/4294967296.0,1,-nbitq), 
to_sfixed(-363079986.0/4294967296.0,1,-nbitq), 
to_sfixed(544695581.0/4294967296.0,1,-nbitq), 
to_sfixed(-1308382402.0/4294967296.0,1,-nbitq), 
to_sfixed(203254970.0/4294967296.0,1,-nbitq), 
to_sfixed(804757381.0/4294967296.0,1,-nbitq), 
to_sfixed(-138569545.0/4294967296.0,1,-nbitq), 
to_sfixed(81991401.0/4294967296.0,1,-nbitq), 
to_sfixed(215917409.0/4294967296.0,1,-nbitq), 
to_sfixed(631706785.0/4294967296.0,1,-nbitq), 
to_sfixed(427104096.0/4294967296.0,1,-nbitq), 
to_sfixed(7412360.0/4294967296.0,1,-nbitq), 
to_sfixed(-5778821.0/4294967296.0,1,-nbitq), 
to_sfixed(314381911.0/4294967296.0,1,-nbitq), 
to_sfixed(-219565540.0/4294967296.0,1,-nbitq), 
to_sfixed(718522722.0/4294967296.0,1,-nbitq), 
to_sfixed(408675649.0/4294967296.0,1,-nbitq), 
to_sfixed(722536454.0/4294967296.0,1,-nbitq), 
to_sfixed(-276237305.0/4294967296.0,1,-nbitq), 
to_sfixed(-351776712.0/4294967296.0,1,-nbitq), 
to_sfixed(104476907.0/4294967296.0,1,-nbitq), 
to_sfixed(-960412754.0/4294967296.0,1,-nbitq), 
to_sfixed(-272308109.0/4294967296.0,1,-nbitq), 
to_sfixed(-54635767.0/4294967296.0,1,-nbitq), 
to_sfixed(-352262856.0/4294967296.0,1,-nbitq), 
to_sfixed(-71420487.0/4294967296.0,1,-nbitq), 
to_sfixed(-110894492.0/4294967296.0,1,-nbitq), 
to_sfixed(458588657.0/4294967296.0,1,-nbitq), 
to_sfixed(958637123.0/4294967296.0,1,-nbitq), 
to_sfixed(-759238513.0/4294967296.0,1,-nbitq), 
to_sfixed(-111290006.0/4294967296.0,1,-nbitq), 
to_sfixed(64089600.0/4294967296.0,1,-nbitq), 
to_sfixed(-293557750.0/4294967296.0,1,-nbitq), 
to_sfixed(-27926346.0/4294967296.0,1,-nbitq), 
to_sfixed(132260795.0/4294967296.0,1,-nbitq), 
to_sfixed(-717829019.0/4294967296.0,1,-nbitq), 
to_sfixed(1085574389.0/4294967296.0,1,-nbitq), 
to_sfixed(689901806.0/4294967296.0,1,-nbitq), 
to_sfixed(101232489.0/4294967296.0,1,-nbitq), 
to_sfixed(-261083612.0/4294967296.0,1,-nbitq), 
to_sfixed(-845162127.0/4294967296.0,1,-nbitq), 
to_sfixed(268530489.0/4294967296.0,1,-nbitq), 
to_sfixed(361834144.0/4294967296.0,1,-nbitq), 
to_sfixed(-337382028.0/4294967296.0,1,-nbitq), 
to_sfixed(202797811.0/4294967296.0,1,-nbitq), 
to_sfixed(-31558720.0/4294967296.0,1,-nbitq), 
to_sfixed(-232228231.0/4294967296.0,1,-nbitq), 
to_sfixed(-294840912.0/4294967296.0,1,-nbitq), 
to_sfixed(313938330.0/4294967296.0,1,-nbitq), 
to_sfixed(-211666121.0/4294967296.0,1,-nbitq), 
to_sfixed(394946722.0/4294967296.0,1,-nbitq), 
to_sfixed(-86155023.0/4294967296.0,1,-nbitq), 
to_sfixed(-453248861.0/4294967296.0,1,-nbitq), 
to_sfixed(-274452427.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-244721030.0/4294967296.0,1,-nbitq), 
to_sfixed(461314107.0/4294967296.0,1,-nbitq), 
to_sfixed(-708572074.0/4294967296.0,1,-nbitq), 
to_sfixed(-112414448.0/4294967296.0,1,-nbitq), 
to_sfixed(-288849779.0/4294967296.0,1,-nbitq), 
to_sfixed(413072341.0/4294967296.0,1,-nbitq), 
to_sfixed(-334190533.0/4294967296.0,1,-nbitq), 
to_sfixed(-105528767.0/4294967296.0,1,-nbitq), 
to_sfixed(167003552.0/4294967296.0,1,-nbitq), 
to_sfixed(172605616.0/4294967296.0,1,-nbitq), 
to_sfixed(-281512135.0/4294967296.0,1,-nbitq), 
to_sfixed(-1069704834.0/4294967296.0,1,-nbitq), 
to_sfixed(-89258232.0/4294967296.0,1,-nbitq), 
to_sfixed(959747845.0/4294967296.0,1,-nbitq), 
to_sfixed(-70931326.0/4294967296.0,1,-nbitq), 
to_sfixed(-307269239.0/4294967296.0,1,-nbitq), 
to_sfixed(24896252.0/4294967296.0,1,-nbitq), 
to_sfixed(-93948838.0/4294967296.0,1,-nbitq), 
to_sfixed(759171745.0/4294967296.0,1,-nbitq), 
to_sfixed(649474057.0/4294967296.0,1,-nbitq), 
to_sfixed(300634441.0/4294967296.0,1,-nbitq), 
to_sfixed(207442156.0/4294967296.0,1,-nbitq), 
to_sfixed(382868718.0/4294967296.0,1,-nbitq), 
to_sfixed(-661352965.0/4294967296.0,1,-nbitq), 
to_sfixed(-282928033.0/4294967296.0,1,-nbitq), 
to_sfixed(790863700.0/4294967296.0,1,-nbitq), 
to_sfixed(468845833.0/4294967296.0,1,-nbitq), 
to_sfixed(-642013943.0/4294967296.0,1,-nbitq), 
to_sfixed(732128230.0/4294967296.0,1,-nbitq), 
to_sfixed(-898222227.0/4294967296.0,1,-nbitq), 
to_sfixed(-459934133.0/4294967296.0,1,-nbitq), 
to_sfixed(115750235.0/4294967296.0,1,-nbitq), 
to_sfixed(-476376356.0/4294967296.0,1,-nbitq), 
to_sfixed(-504777931.0/4294967296.0,1,-nbitq), 
to_sfixed(703700377.0/4294967296.0,1,-nbitq), 
to_sfixed(361751342.0/4294967296.0,1,-nbitq), 
to_sfixed(24475371.0/4294967296.0,1,-nbitq), 
to_sfixed(29888058.0/4294967296.0,1,-nbitq), 
to_sfixed(256630392.0/4294967296.0,1,-nbitq), 
to_sfixed(502557561.0/4294967296.0,1,-nbitq), 
to_sfixed(-330805495.0/4294967296.0,1,-nbitq), 
to_sfixed(671122610.0/4294967296.0,1,-nbitq), 
to_sfixed(-63944071.0/4294967296.0,1,-nbitq), 
to_sfixed(760008318.0/4294967296.0,1,-nbitq), 
to_sfixed(154332437.0/4294967296.0,1,-nbitq), 
to_sfixed(-384167370.0/4294967296.0,1,-nbitq), 
to_sfixed(-104663313.0/4294967296.0,1,-nbitq), 
to_sfixed(-992706181.0/4294967296.0,1,-nbitq), 
to_sfixed(251386987.0/4294967296.0,1,-nbitq), 
to_sfixed(560490125.0/4294967296.0,1,-nbitq), 
to_sfixed(-109011877.0/4294967296.0,1,-nbitq), 
to_sfixed(-21827559.0/4294967296.0,1,-nbitq), 
to_sfixed(-359606137.0/4294967296.0,1,-nbitq), 
to_sfixed(536586836.0/4294967296.0,1,-nbitq), 
to_sfixed(548614188.0/4294967296.0,1,-nbitq), 
to_sfixed(-115252338.0/4294967296.0,1,-nbitq), 
to_sfixed(-211303979.0/4294967296.0,1,-nbitq), 
to_sfixed(-163344670.0/4294967296.0,1,-nbitq), 
to_sfixed(-78299839.0/4294967296.0,1,-nbitq), 
to_sfixed(-226446747.0/4294967296.0,1,-nbitq), 
to_sfixed(-211987238.0/4294967296.0,1,-nbitq), 
to_sfixed(-581609680.0/4294967296.0,1,-nbitq), 
to_sfixed(500946196.0/4294967296.0,1,-nbitq), 
to_sfixed(27174516.0/4294967296.0,1,-nbitq), 
to_sfixed(-267479057.0/4294967296.0,1,-nbitq), 
to_sfixed(-176186543.0/4294967296.0,1,-nbitq), 
to_sfixed(-637338419.0/4294967296.0,1,-nbitq), 
to_sfixed(53018297.0/4294967296.0,1,-nbitq), 
to_sfixed(223669002.0/4294967296.0,1,-nbitq), 
to_sfixed(-457198946.0/4294967296.0,1,-nbitq), 
to_sfixed(279197015.0/4294967296.0,1,-nbitq), 
to_sfixed(479224412.0/4294967296.0,1,-nbitq), 
to_sfixed(-507768950.0/4294967296.0,1,-nbitq), 
to_sfixed(-330777737.0/4294967296.0,1,-nbitq), 
to_sfixed(-251878828.0/4294967296.0,1,-nbitq), 
to_sfixed(-290618180.0/4294967296.0,1,-nbitq), 
to_sfixed(616862847.0/4294967296.0,1,-nbitq), 
to_sfixed(414548236.0/4294967296.0,1,-nbitq), 
to_sfixed(-846817310.0/4294967296.0,1,-nbitq), 
to_sfixed(-228367185.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(21958294.0/4294967296.0,1,-nbitq), 
to_sfixed(631033848.0/4294967296.0,1,-nbitq), 
to_sfixed(-463799552.0/4294967296.0,1,-nbitq), 
to_sfixed(-442071966.0/4294967296.0,1,-nbitq), 
to_sfixed(772168460.0/4294967296.0,1,-nbitq), 
to_sfixed(470750481.0/4294967296.0,1,-nbitq), 
to_sfixed(1915838.0/4294967296.0,1,-nbitq), 
to_sfixed(-123176891.0/4294967296.0,1,-nbitq), 
to_sfixed(81627126.0/4294967296.0,1,-nbitq), 
to_sfixed(-18012304.0/4294967296.0,1,-nbitq), 
to_sfixed(42774119.0/4294967296.0,1,-nbitq), 
to_sfixed(-573053573.0/4294967296.0,1,-nbitq), 
to_sfixed(102597410.0/4294967296.0,1,-nbitq), 
to_sfixed(-88015256.0/4294967296.0,1,-nbitq), 
to_sfixed(207688839.0/4294967296.0,1,-nbitq), 
to_sfixed(-852802593.0/4294967296.0,1,-nbitq), 
to_sfixed(293177197.0/4294967296.0,1,-nbitq), 
to_sfixed(-89484875.0/4294967296.0,1,-nbitq), 
to_sfixed(252091450.0/4294967296.0,1,-nbitq), 
to_sfixed(42056918.0/4294967296.0,1,-nbitq), 
to_sfixed(-182511387.0/4294967296.0,1,-nbitq), 
to_sfixed(-376763566.0/4294967296.0,1,-nbitq), 
to_sfixed(10911588.0/4294967296.0,1,-nbitq), 
to_sfixed(-214392598.0/4294967296.0,1,-nbitq), 
to_sfixed(98578313.0/4294967296.0,1,-nbitq), 
to_sfixed(1108772893.0/4294967296.0,1,-nbitq), 
to_sfixed(-401466047.0/4294967296.0,1,-nbitq), 
to_sfixed(269367681.0/4294967296.0,1,-nbitq), 
to_sfixed(-73082830.0/4294967296.0,1,-nbitq), 
to_sfixed(-812908087.0/4294967296.0,1,-nbitq), 
to_sfixed(-64584866.0/4294967296.0,1,-nbitq), 
to_sfixed(607189740.0/4294967296.0,1,-nbitq), 
to_sfixed(112069945.0/4294967296.0,1,-nbitq), 
to_sfixed(-844755392.0/4294967296.0,1,-nbitq), 
to_sfixed(137298077.0/4294967296.0,1,-nbitq), 
to_sfixed(658793237.0/4294967296.0,1,-nbitq), 
to_sfixed(205216527.0/4294967296.0,1,-nbitq), 
to_sfixed(-102090956.0/4294967296.0,1,-nbitq), 
to_sfixed(91862908.0/4294967296.0,1,-nbitq), 
to_sfixed(493035881.0/4294967296.0,1,-nbitq), 
to_sfixed(8863144.0/4294967296.0,1,-nbitq), 
to_sfixed(-20597294.0/4294967296.0,1,-nbitq), 
to_sfixed(494315104.0/4294967296.0,1,-nbitq), 
to_sfixed(54789593.0/4294967296.0,1,-nbitq), 
to_sfixed(-48415633.0/4294967296.0,1,-nbitq), 
to_sfixed(46692528.0/4294967296.0,1,-nbitq), 
to_sfixed(-40532111.0/4294967296.0,1,-nbitq), 
to_sfixed(-896401433.0/4294967296.0,1,-nbitq), 
to_sfixed(-66292530.0/4294967296.0,1,-nbitq), 
to_sfixed(258816213.0/4294967296.0,1,-nbitq), 
to_sfixed(-158211136.0/4294967296.0,1,-nbitq), 
to_sfixed(-853351958.0/4294967296.0,1,-nbitq), 
to_sfixed(-390846994.0/4294967296.0,1,-nbitq), 
to_sfixed(-2464511.0/4294967296.0,1,-nbitq), 
to_sfixed(760940816.0/4294967296.0,1,-nbitq), 
to_sfixed(194889714.0/4294967296.0,1,-nbitq), 
to_sfixed(-118960800.0/4294967296.0,1,-nbitq), 
to_sfixed(-70380899.0/4294967296.0,1,-nbitq), 
to_sfixed(405892417.0/4294967296.0,1,-nbitq), 
to_sfixed(-180651429.0/4294967296.0,1,-nbitq), 
to_sfixed(-83058025.0/4294967296.0,1,-nbitq), 
to_sfixed(-826883355.0/4294967296.0,1,-nbitq), 
to_sfixed(111900319.0/4294967296.0,1,-nbitq), 
to_sfixed(233125672.0/4294967296.0,1,-nbitq), 
to_sfixed(340014196.0/4294967296.0,1,-nbitq), 
to_sfixed(387606178.0/4294967296.0,1,-nbitq), 
to_sfixed(-617059183.0/4294967296.0,1,-nbitq), 
to_sfixed(-813578933.0/4294967296.0,1,-nbitq), 
to_sfixed(-261969166.0/4294967296.0,1,-nbitq), 
to_sfixed(-9442939.0/4294967296.0,1,-nbitq), 
to_sfixed(664173574.0/4294967296.0,1,-nbitq), 
to_sfixed(-307079866.0/4294967296.0,1,-nbitq), 
to_sfixed(-336645527.0/4294967296.0,1,-nbitq), 
to_sfixed(315607320.0/4294967296.0,1,-nbitq), 
to_sfixed(-101812489.0/4294967296.0,1,-nbitq), 
to_sfixed(49331877.0/4294967296.0,1,-nbitq), 
to_sfixed(-416756417.0/4294967296.0,1,-nbitq), 
to_sfixed(-399970974.0/4294967296.0,1,-nbitq), 
to_sfixed(-57953924.0/4294967296.0,1,-nbitq), 
to_sfixed(-78326149.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-121399271.0/4294967296.0,1,-nbitq), 
to_sfixed(1113485884.0/4294967296.0,1,-nbitq), 
to_sfixed(-205897819.0/4294967296.0,1,-nbitq), 
to_sfixed(-632566531.0/4294967296.0,1,-nbitq), 
to_sfixed(765185246.0/4294967296.0,1,-nbitq), 
to_sfixed(-294007444.0/4294967296.0,1,-nbitq), 
to_sfixed(249450357.0/4294967296.0,1,-nbitq), 
to_sfixed(441958856.0/4294967296.0,1,-nbitq), 
to_sfixed(-249352246.0/4294967296.0,1,-nbitq), 
to_sfixed(-56986803.0/4294967296.0,1,-nbitq), 
to_sfixed(713262078.0/4294967296.0,1,-nbitq), 
to_sfixed(-187080980.0/4294967296.0,1,-nbitq), 
to_sfixed(596888480.0/4294967296.0,1,-nbitq), 
to_sfixed(123421196.0/4294967296.0,1,-nbitq), 
to_sfixed(337992230.0/4294967296.0,1,-nbitq), 
to_sfixed(-208789519.0/4294967296.0,1,-nbitq), 
to_sfixed(166167222.0/4294967296.0,1,-nbitq), 
to_sfixed(-354477313.0/4294967296.0,1,-nbitq), 
to_sfixed(216890789.0/4294967296.0,1,-nbitq), 
to_sfixed(151331022.0/4294967296.0,1,-nbitq), 
to_sfixed(96903621.0/4294967296.0,1,-nbitq), 
to_sfixed(35956334.0/4294967296.0,1,-nbitq), 
to_sfixed(-150488826.0/4294967296.0,1,-nbitq), 
to_sfixed(-285463473.0/4294967296.0,1,-nbitq), 
to_sfixed(-187665348.0/4294967296.0,1,-nbitq), 
to_sfixed(965470112.0/4294967296.0,1,-nbitq), 
to_sfixed(-168004758.0/4294967296.0,1,-nbitq), 
to_sfixed(292807700.0/4294967296.0,1,-nbitq), 
to_sfixed(346284003.0/4294967296.0,1,-nbitq), 
to_sfixed(-851541109.0/4294967296.0,1,-nbitq), 
to_sfixed(-97394572.0/4294967296.0,1,-nbitq), 
to_sfixed(609546850.0/4294967296.0,1,-nbitq), 
to_sfixed(-41582956.0/4294967296.0,1,-nbitq), 
to_sfixed(-195301118.0/4294967296.0,1,-nbitq), 
to_sfixed(-104234067.0/4294967296.0,1,-nbitq), 
to_sfixed(548035544.0/4294967296.0,1,-nbitq), 
to_sfixed(-200201044.0/4294967296.0,1,-nbitq), 
to_sfixed(-84654418.0/4294967296.0,1,-nbitq), 
to_sfixed(189260738.0/4294967296.0,1,-nbitq), 
to_sfixed(178234208.0/4294967296.0,1,-nbitq), 
to_sfixed(385546205.0/4294967296.0,1,-nbitq), 
to_sfixed(-127799815.0/4294967296.0,1,-nbitq), 
to_sfixed(415328291.0/4294967296.0,1,-nbitq), 
to_sfixed(7072598.0/4294967296.0,1,-nbitq), 
to_sfixed(-32411659.0/4294967296.0,1,-nbitq), 
to_sfixed(431043800.0/4294967296.0,1,-nbitq), 
to_sfixed(-437666019.0/4294967296.0,1,-nbitq), 
to_sfixed(-847999687.0/4294967296.0,1,-nbitq), 
to_sfixed(-51741250.0/4294967296.0,1,-nbitq), 
to_sfixed(-536184604.0/4294967296.0,1,-nbitq), 
to_sfixed(-266077068.0/4294967296.0,1,-nbitq), 
to_sfixed(-684516724.0/4294967296.0,1,-nbitq), 
to_sfixed(270191582.0/4294967296.0,1,-nbitq), 
to_sfixed(256945938.0/4294967296.0,1,-nbitq), 
to_sfixed(519150982.0/4294967296.0,1,-nbitq), 
to_sfixed(-401127879.0/4294967296.0,1,-nbitq), 
to_sfixed(156167887.0/4294967296.0,1,-nbitq), 
to_sfixed(186293662.0/4294967296.0,1,-nbitq), 
to_sfixed(-128730546.0/4294967296.0,1,-nbitq), 
to_sfixed(250166120.0/4294967296.0,1,-nbitq), 
to_sfixed(-234902783.0/4294967296.0,1,-nbitq), 
to_sfixed(-387803087.0/4294967296.0,1,-nbitq), 
to_sfixed(872654747.0/4294967296.0,1,-nbitq), 
to_sfixed(52909918.0/4294967296.0,1,-nbitq), 
to_sfixed(293656042.0/4294967296.0,1,-nbitq), 
to_sfixed(-216641535.0/4294967296.0,1,-nbitq), 
to_sfixed(-478660095.0/4294967296.0,1,-nbitq), 
to_sfixed(-917093390.0/4294967296.0,1,-nbitq), 
to_sfixed(-100718984.0/4294967296.0,1,-nbitq), 
to_sfixed(77418591.0/4294967296.0,1,-nbitq), 
to_sfixed(1057769602.0/4294967296.0,1,-nbitq), 
to_sfixed(455832977.0/4294967296.0,1,-nbitq), 
to_sfixed(214797515.0/4294967296.0,1,-nbitq), 
to_sfixed(415435505.0/4294967296.0,1,-nbitq), 
to_sfixed(375941612.0/4294967296.0,1,-nbitq), 
to_sfixed(-260267149.0/4294967296.0,1,-nbitq), 
to_sfixed(-589353083.0/4294967296.0,1,-nbitq), 
to_sfixed(-265526409.0/4294967296.0,1,-nbitq), 
to_sfixed(-158101649.0/4294967296.0,1,-nbitq), 
to_sfixed(298771313.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(67658304.0/4294967296.0,1,-nbitq), 
to_sfixed(450639148.0/4294967296.0,1,-nbitq), 
to_sfixed(62608980.0/4294967296.0,1,-nbitq), 
to_sfixed(377267093.0/4294967296.0,1,-nbitq), 
to_sfixed(138554069.0/4294967296.0,1,-nbitq), 
to_sfixed(69854723.0/4294967296.0,1,-nbitq), 
to_sfixed(132535706.0/4294967296.0,1,-nbitq), 
to_sfixed(283372103.0/4294967296.0,1,-nbitq), 
to_sfixed(134914603.0/4294967296.0,1,-nbitq), 
to_sfixed(-123433430.0/4294967296.0,1,-nbitq), 
to_sfixed(625171013.0/4294967296.0,1,-nbitq), 
to_sfixed(-61847084.0/4294967296.0,1,-nbitq), 
to_sfixed(718305713.0/4294967296.0,1,-nbitq), 
to_sfixed(-445606448.0/4294967296.0,1,-nbitq), 
to_sfixed(-274776168.0/4294967296.0,1,-nbitq), 
to_sfixed(-360777470.0/4294967296.0,1,-nbitq), 
to_sfixed(-171981027.0/4294967296.0,1,-nbitq), 
to_sfixed(358080441.0/4294967296.0,1,-nbitq), 
to_sfixed(-72667169.0/4294967296.0,1,-nbitq), 
to_sfixed(-140813256.0/4294967296.0,1,-nbitq), 
to_sfixed(-312155361.0/4294967296.0,1,-nbitq), 
to_sfixed(272362181.0/4294967296.0,1,-nbitq), 
to_sfixed(-164913545.0/4294967296.0,1,-nbitq), 
to_sfixed(-578314634.0/4294967296.0,1,-nbitq), 
to_sfixed(254699699.0/4294967296.0,1,-nbitq), 
to_sfixed(1013503758.0/4294967296.0,1,-nbitq), 
to_sfixed(-391442620.0/4294967296.0,1,-nbitq), 
to_sfixed(204944621.0/4294967296.0,1,-nbitq), 
to_sfixed(-281457254.0/4294967296.0,1,-nbitq), 
to_sfixed(-500791808.0/4294967296.0,1,-nbitq), 
to_sfixed(341247444.0/4294967296.0,1,-nbitq), 
to_sfixed(738633180.0/4294967296.0,1,-nbitq), 
to_sfixed(408813659.0/4294967296.0,1,-nbitq), 
to_sfixed(-271655201.0/4294967296.0,1,-nbitq), 
to_sfixed(-98714232.0/4294967296.0,1,-nbitq), 
to_sfixed(-8923969.0/4294967296.0,1,-nbitq), 
to_sfixed(308109587.0/4294967296.0,1,-nbitq), 
to_sfixed(-876827275.0/4294967296.0,1,-nbitq), 
to_sfixed(170881937.0/4294967296.0,1,-nbitq), 
to_sfixed(56639604.0/4294967296.0,1,-nbitq), 
to_sfixed(705408638.0/4294967296.0,1,-nbitq), 
to_sfixed(-180170264.0/4294967296.0,1,-nbitq), 
to_sfixed(373374766.0/4294967296.0,1,-nbitq), 
to_sfixed(-59809051.0/4294967296.0,1,-nbitq), 
to_sfixed(480421580.0/4294967296.0,1,-nbitq), 
to_sfixed(537449268.0/4294967296.0,1,-nbitq), 
to_sfixed(151942312.0/4294967296.0,1,-nbitq), 
to_sfixed(-221379744.0/4294967296.0,1,-nbitq), 
to_sfixed(-479477906.0/4294967296.0,1,-nbitq), 
to_sfixed(-478654666.0/4294967296.0,1,-nbitq), 
to_sfixed(-430642950.0/4294967296.0,1,-nbitq), 
to_sfixed(-121701585.0/4294967296.0,1,-nbitq), 
to_sfixed(116968574.0/4294967296.0,1,-nbitq), 
to_sfixed(-8788692.0/4294967296.0,1,-nbitq), 
to_sfixed(217227250.0/4294967296.0,1,-nbitq), 
to_sfixed(137934953.0/4294967296.0,1,-nbitq), 
to_sfixed(-150140073.0/4294967296.0,1,-nbitq), 
to_sfixed(-304400180.0/4294967296.0,1,-nbitq), 
to_sfixed(-80476657.0/4294967296.0,1,-nbitq), 
to_sfixed(-132995376.0/4294967296.0,1,-nbitq), 
to_sfixed(-281532024.0/4294967296.0,1,-nbitq), 
to_sfixed(-273067474.0/4294967296.0,1,-nbitq), 
to_sfixed(323990330.0/4294967296.0,1,-nbitq), 
to_sfixed(-151160773.0/4294967296.0,1,-nbitq), 
to_sfixed(-5680218.0/4294967296.0,1,-nbitq), 
to_sfixed(-73149944.0/4294967296.0,1,-nbitq), 
to_sfixed(-869968109.0/4294967296.0,1,-nbitq), 
to_sfixed(-690235600.0/4294967296.0,1,-nbitq), 
to_sfixed(251733239.0/4294967296.0,1,-nbitq), 
to_sfixed(-80326904.0/4294967296.0,1,-nbitq), 
to_sfixed(768316566.0/4294967296.0,1,-nbitq), 
to_sfixed(128033720.0/4294967296.0,1,-nbitq), 
to_sfixed(-292637733.0/4294967296.0,1,-nbitq), 
to_sfixed(23321509.0/4294967296.0,1,-nbitq), 
to_sfixed(346012618.0/4294967296.0,1,-nbitq), 
to_sfixed(255122182.0/4294967296.0,1,-nbitq), 
to_sfixed(261581816.0/4294967296.0,1,-nbitq), 
to_sfixed(-231421740.0/4294967296.0,1,-nbitq), 
to_sfixed(-72730593.0/4294967296.0,1,-nbitq), 
to_sfixed(-182667760.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(299752322.0/4294967296.0,1,-nbitq), 
to_sfixed(706515335.0/4294967296.0,1,-nbitq), 
to_sfixed(-86078000.0/4294967296.0,1,-nbitq), 
to_sfixed(433567985.0/4294967296.0,1,-nbitq), 
to_sfixed(-32916862.0/4294967296.0,1,-nbitq), 
to_sfixed(9628695.0/4294967296.0,1,-nbitq), 
to_sfixed(-322411976.0/4294967296.0,1,-nbitq), 
to_sfixed(-24070996.0/4294967296.0,1,-nbitq), 
to_sfixed(-149703959.0/4294967296.0,1,-nbitq), 
to_sfixed(297674609.0/4294967296.0,1,-nbitq), 
to_sfixed(770672657.0/4294967296.0,1,-nbitq), 
to_sfixed(132232234.0/4294967296.0,1,-nbitq), 
to_sfixed(788229402.0/4294967296.0,1,-nbitq), 
to_sfixed(-850424007.0/4294967296.0,1,-nbitq), 
to_sfixed(-401560094.0/4294967296.0,1,-nbitq), 
to_sfixed(-36001268.0/4294967296.0,1,-nbitq), 
to_sfixed(-347440447.0/4294967296.0,1,-nbitq), 
to_sfixed(-349528111.0/4294967296.0,1,-nbitq), 
to_sfixed(655437052.0/4294967296.0,1,-nbitq), 
to_sfixed(-13867349.0/4294967296.0,1,-nbitq), 
to_sfixed(142450488.0/4294967296.0,1,-nbitq), 
to_sfixed(149004847.0/4294967296.0,1,-nbitq), 
to_sfixed(113528533.0/4294967296.0,1,-nbitq), 
to_sfixed(-281884221.0/4294967296.0,1,-nbitq), 
to_sfixed(318985291.0/4294967296.0,1,-nbitq), 
to_sfixed(628446042.0/4294967296.0,1,-nbitq), 
to_sfixed(-513279944.0/4294967296.0,1,-nbitq), 
to_sfixed(36835357.0/4294967296.0,1,-nbitq), 
to_sfixed(-41302681.0/4294967296.0,1,-nbitq), 
to_sfixed(-158442767.0/4294967296.0,1,-nbitq), 
to_sfixed(264572939.0/4294967296.0,1,-nbitq), 
to_sfixed(106534587.0/4294967296.0,1,-nbitq), 
to_sfixed(532057397.0/4294967296.0,1,-nbitq), 
to_sfixed(-229068609.0/4294967296.0,1,-nbitq), 
to_sfixed(-442016863.0/4294967296.0,1,-nbitq), 
to_sfixed(-146510125.0/4294967296.0,1,-nbitq), 
to_sfixed(-115509938.0/4294967296.0,1,-nbitq), 
to_sfixed(20990861.0/4294967296.0,1,-nbitq), 
to_sfixed(17915579.0/4294967296.0,1,-nbitq), 
to_sfixed(406535196.0/4294967296.0,1,-nbitq), 
to_sfixed(389923048.0/4294967296.0,1,-nbitq), 
to_sfixed(4531827.0/4294967296.0,1,-nbitq), 
to_sfixed(-271856312.0/4294967296.0,1,-nbitq), 
to_sfixed(23833974.0/4294967296.0,1,-nbitq), 
to_sfixed(365544251.0/4294967296.0,1,-nbitq), 
to_sfixed(410414590.0/4294967296.0,1,-nbitq), 
to_sfixed(-95787021.0/4294967296.0,1,-nbitq), 
to_sfixed(274022431.0/4294967296.0,1,-nbitq), 
to_sfixed(163592536.0/4294967296.0,1,-nbitq), 
to_sfixed(20393469.0/4294967296.0,1,-nbitq), 
to_sfixed(-447360836.0/4294967296.0,1,-nbitq), 
to_sfixed(-106657795.0/4294967296.0,1,-nbitq), 
to_sfixed(164829973.0/4294967296.0,1,-nbitq), 
to_sfixed(447915247.0/4294967296.0,1,-nbitq), 
to_sfixed(276572467.0/4294967296.0,1,-nbitq), 
to_sfixed(-137983694.0/4294967296.0,1,-nbitq), 
to_sfixed(-400793897.0/4294967296.0,1,-nbitq), 
to_sfixed(-36355415.0/4294967296.0,1,-nbitq), 
to_sfixed(305161178.0/4294967296.0,1,-nbitq), 
to_sfixed(147555496.0/4294967296.0,1,-nbitq), 
to_sfixed(245693884.0/4294967296.0,1,-nbitq), 
to_sfixed(-45294363.0/4294967296.0,1,-nbitq), 
to_sfixed(-19363339.0/4294967296.0,1,-nbitq), 
to_sfixed(-285244003.0/4294967296.0,1,-nbitq), 
to_sfixed(-180382713.0/4294967296.0,1,-nbitq), 
to_sfixed(-123602081.0/4294967296.0,1,-nbitq), 
to_sfixed(237940069.0/4294967296.0,1,-nbitq), 
to_sfixed(-372412810.0/4294967296.0,1,-nbitq), 
to_sfixed(-64864467.0/4294967296.0,1,-nbitq), 
to_sfixed(-349719061.0/4294967296.0,1,-nbitq), 
to_sfixed(-121829632.0/4294967296.0,1,-nbitq), 
to_sfixed(-339972243.0/4294967296.0,1,-nbitq), 
to_sfixed(-536407415.0/4294967296.0,1,-nbitq), 
to_sfixed(286107708.0/4294967296.0,1,-nbitq), 
to_sfixed(106971051.0/4294967296.0,1,-nbitq), 
to_sfixed(-20899715.0/4294967296.0,1,-nbitq), 
to_sfixed(493060017.0/4294967296.0,1,-nbitq), 
to_sfixed(262989187.0/4294967296.0,1,-nbitq), 
to_sfixed(-254767117.0/4294967296.0,1,-nbitq), 
to_sfixed(-327361044.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-280028024.0/4294967296.0,1,-nbitq), 
to_sfixed(-146777548.0/4294967296.0,1,-nbitq), 
to_sfixed(-192807934.0/4294967296.0,1,-nbitq), 
to_sfixed(41233651.0/4294967296.0,1,-nbitq), 
to_sfixed(151134090.0/4294967296.0,1,-nbitq), 
to_sfixed(-234540882.0/4294967296.0,1,-nbitq), 
to_sfixed(143325920.0/4294967296.0,1,-nbitq), 
to_sfixed(382991852.0/4294967296.0,1,-nbitq), 
to_sfixed(-233594673.0/4294967296.0,1,-nbitq), 
to_sfixed(-346035885.0/4294967296.0,1,-nbitq), 
to_sfixed(-63593941.0/4294967296.0,1,-nbitq), 
to_sfixed(237110751.0/4294967296.0,1,-nbitq), 
to_sfixed(115462369.0/4294967296.0,1,-nbitq), 
to_sfixed(285620383.0/4294967296.0,1,-nbitq), 
to_sfixed(212558220.0/4294967296.0,1,-nbitq), 
to_sfixed(-297796594.0/4294967296.0,1,-nbitq), 
to_sfixed(-155899151.0/4294967296.0,1,-nbitq), 
to_sfixed(94773442.0/4294967296.0,1,-nbitq), 
to_sfixed(113751941.0/4294967296.0,1,-nbitq), 
to_sfixed(-59093376.0/4294967296.0,1,-nbitq), 
to_sfixed(-148146706.0/4294967296.0,1,-nbitq), 
to_sfixed(-237219938.0/4294967296.0,1,-nbitq), 
to_sfixed(-45820510.0/4294967296.0,1,-nbitq), 
to_sfixed(231042817.0/4294967296.0,1,-nbitq), 
to_sfixed(-41143220.0/4294967296.0,1,-nbitq), 
to_sfixed(584936674.0/4294967296.0,1,-nbitq), 
to_sfixed(-509716043.0/4294967296.0,1,-nbitq), 
to_sfixed(-475641202.0/4294967296.0,1,-nbitq), 
to_sfixed(512237144.0/4294967296.0,1,-nbitq), 
to_sfixed(-6459190.0/4294967296.0,1,-nbitq), 
to_sfixed(202187758.0/4294967296.0,1,-nbitq), 
to_sfixed(-274457357.0/4294967296.0,1,-nbitq), 
to_sfixed(-50396289.0/4294967296.0,1,-nbitq), 
to_sfixed(-671972172.0/4294967296.0,1,-nbitq), 
to_sfixed(-205670344.0/4294967296.0,1,-nbitq), 
to_sfixed(68010229.0/4294967296.0,1,-nbitq), 
to_sfixed(-135258816.0/4294967296.0,1,-nbitq), 
to_sfixed(-164893840.0/4294967296.0,1,-nbitq), 
to_sfixed(51294639.0/4294967296.0,1,-nbitq), 
to_sfixed(-30263889.0/4294967296.0,1,-nbitq), 
to_sfixed(1288512.0/4294967296.0,1,-nbitq), 
to_sfixed(205163650.0/4294967296.0,1,-nbitq), 
to_sfixed(-406621301.0/4294967296.0,1,-nbitq), 
to_sfixed(191502162.0/4294967296.0,1,-nbitq), 
to_sfixed(547556303.0/4294967296.0,1,-nbitq), 
to_sfixed(-195105413.0/4294967296.0,1,-nbitq), 
to_sfixed(-197756350.0/4294967296.0,1,-nbitq), 
to_sfixed(193562962.0/4294967296.0,1,-nbitq), 
to_sfixed(170647607.0/4294967296.0,1,-nbitq), 
to_sfixed(288632492.0/4294967296.0,1,-nbitq), 
to_sfixed(86890568.0/4294967296.0,1,-nbitq), 
to_sfixed(-11974346.0/4294967296.0,1,-nbitq), 
to_sfixed(-64145893.0/4294967296.0,1,-nbitq), 
to_sfixed(228628093.0/4294967296.0,1,-nbitq), 
to_sfixed(501670431.0/4294967296.0,1,-nbitq), 
to_sfixed(106107270.0/4294967296.0,1,-nbitq), 
to_sfixed(-37181534.0/4294967296.0,1,-nbitq), 
to_sfixed(-409276893.0/4294967296.0,1,-nbitq), 
to_sfixed(87150656.0/4294967296.0,1,-nbitq), 
to_sfixed(-350543113.0/4294967296.0,1,-nbitq), 
to_sfixed(6609358.0/4294967296.0,1,-nbitq), 
to_sfixed(-282121778.0/4294967296.0,1,-nbitq), 
to_sfixed(191847288.0/4294967296.0,1,-nbitq), 
to_sfixed(164261616.0/4294967296.0,1,-nbitq), 
to_sfixed(-60745988.0/4294967296.0,1,-nbitq), 
to_sfixed(-152898888.0/4294967296.0,1,-nbitq), 
to_sfixed(58761728.0/4294967296.0,1,-nbitq), 
to_sfixed(-244402203.0/4294967296.0,1,-nbitq), 
to_sfixed(-15880742.0/4294967296.0,1,-nbitq), 
to_sfixed(-125320134.0/4294967296.0,1,-nbitq), 
to_sfixed(78633571.0/4294967296.0,1,-nbitq), 
to_sfixed(-287704744.0/4294967296.0,1,-nbitq), 
to_sfixed(-88858047.0/4294967296.0,1,-nbitq), 
to_sfixed(-184503128.0/4294967296.0,1,-nbitq), 
to_sfixed(370343263.0/4294967296.0,1,-nbitq), 
to_sfixed(-559523875.0/4294967296.0,1,-nbitq), 
to_sfixed(245551622.0/4294967296.0,1,-nbitq), 
to_sfixed(-210378221.0/4294967296.0,1,-nbitq), 
to_sfixed(-659090216.0/4294967296.0,1,-nbitq), 
to_sfixed(-33050957.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(295277357.0/4294967296.0,1,-nbitq), 
to_sfixed(-47248540.0/4294967296.0,1,-nbitq), 
to_sfixed(217963602.0/4294967296.0,1,-nbitq), 
to_sfixed(-294876516.0/4294967296.0,1,-nbitq), 
to_sfixed(238414872.0/4294967296.0,1,-nbitq), 
to_sfixed(-244038998.0/4294967296.0,1,-nbitq), 
to_sfixed(318498550.0/4294967296.0,1,-nbitq), 
to_sfixed(353945677.0/4294967296.0,1,-nbitq), 
to_sfixed(-224136657.0/4294967296.0,1,-nbitq), 
to_sfixed(-175313055.0/4294967296.0,1,-nbitq), 
to_sfixed(206540014.0/4294967296.0,1,-nbitq), 
to_sfixed(418813072.0/4294967296.0,1,-nbitq), 
to_sfixed(-263899186.0/4294967296.0,1,-nbitq), 
to_sfixed(252205399.0/4294967296.0,1,-nbitq), 
to_sfixed(245519213.0/4294967296.0,1,-nbitq), 
to_sfixed(-492641797.0/4294967296.0,1,-nbitq), 
to_sfixed(351540553.0/4294967296.0,1,-nbitq), 
to_sfixed(262064772.0/4294967296.0,1,-nbitq), 
to_sfixed(497832052.0/4294967296.0,1,-nbitq), 
to_sfixed(-334019827.0/4294967296.0,1,-nbitq), 
to_sfixed(-329398631.0/4294967296.0,1,-nbitq), 
to_sfixed(-228261591.0/4294967296.0,1,-nbitq), 
to_sfixed(507215227.0/4294967296.0,1,-nbitq), 
to_sfixed(-354690105.0/4294967296.0,1,-nbitq), 
to_sfixed(-42829416.0/4294967296.0,1,-nbitq), 
to_sfixed(302974130.0/4294967296.0,1,-nbitq), 
to_sfixed(336178471.0/4294967296.0,1,-nbitq), 
to_sfixed(-87841210.0/4294967296.0,1,-nbitq), 
to_sfixed(-42841389.0/4294967296.0,1,-nbitq), 
to_sfixed(-40607869.0/4294967296.0,1,-nbitq), 
to_sfixed(-554086545.0/4294967296.0,1,-nbitq), 
to_sfixed(-374174646.0/4294967296.0,1,-nbitq), 
to_sfixed(185122902.0/4294967296.0,1,-nbitq), 
to_sfixed(-520190921.0/4294967296.0,1,-nbitq), 
to_sfixed(-218688225.0/4294967296.0,1,-nbitq), 
to_sfixed(-327884910.0/4294967296.0,1,-nbitq), 
to_sfixed(179485792.0/4294967296.0,1,-nbitq), 
to_sfixed(420207724.0/4294967296.0,1,-nbitq), 
to_sfixed(-296293488.0/4294967296.0,1,-nbitq), 
to_sfixed(175173972.0/4294967296.0,1,-nbitq), 
to_sfixed(-353434068.0/4294967296.0,1,-nbitq), 
to_sfixed(-26020989.0/4294967296.0,1,-nbitq), 
to_sfixed(-309292831.0/4294967296.0,1,-nbitq), 
to_sfixed(372564033.0/4294967296.0,1,-nbitq), 
to_sfixed(-10850039.0/4294967296.0,1,-nbitq), 
to_sfixed(118314321.0/4294967296.0,1,-nbitq), 
to_sfixed(-195944536.0/4294967296.0,1,-nbitq), 
to_sfixed(-61859504.0/4294967296.0,1,-nbitq), 
to_sfixed(-18771434.0/4294967296.0,1,-nbitq), 
to_sfixed(-58607473.0/4294967296.0,1,-nbitq), 
to_sfixed(230868605.0/4294967296.0,1,-nbitq), 
to_sfixed(-329599377.0/4294967296.0,1,-nbitq), 
to_sfixed(-290744445.0/4294967296.0,1,-nbitq), 
to_sfixed(161857831.0/4294967296.0,1,-nbitq), 
to_sfixed(44789418.0/4294967296.0,1,-nbitq), 
to_sfixed(247509217.0/4294967296.0,1,-nbitq), 
to_sfixed(200057181.0/4294967296.0,1,-nbitq), 
to_sfixed(-461156911.0/4294967296.0,1,-nbitq), 
to_sfixed(-168185962.0/4294967296.0,1,-nbitq), 
to_sfixed(-262235347.0/4294967296.0,1,-nbitq), 
to_sfixed(299824026.0/4294967296.0,1,-nbitq), 
to_sfixed(244576889.0/4294967296.0,1,-nbitq), 
to_sfixed(-380209030.0/4294967296.0,1,-nbitq), 
to_sfixed(-89835993.0/4294967296.0,1,-nbitq), 
to_sfixed(14998811.0/4294967296.0,1,-nbitq), 
to_sfixed(28331845.0/4294967296.0,1,-nbitq), 
to_sfixed(297626325.0/4294967296.0,1,-nbitq), 
to_sfixed(-119663954.0/4294967296.0,1,-nbitq), 
to_sfixed(437138321.0/4294967296.0,1,-nbitq), 
to_sfixed(272301646.0/4294967296.0,1,-nbitq), 
to_sfixed(-31907387.0/4294967296.0,1,-nbitq), 
to_sfixed(327138102.0/4294967296.0,1,-nbitq), 
to_sfixed(-16318147.0/4294967296.0,1,-nbitq), 
to_sfixed(-110716969.0/4294967296.0,1,-nbitq), 
to_sfixed(393842586.0/4294967296.0,1,-nbitq), 
to_sfixed(74432485.0/4294967296.0,1,-nbitq), 
to_sfixed(72140306.0/4294967296.0,1,-nbitq), 
to_sfixed(-253201695.0/4294967296.0,1,-nbitq), 
to_sfixed(-129229172.0/4294967296.0,1,-nbitq), 
to_sfixed(325471812.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(385777964.0/4294967296.0,1,-nbitq), 
to_sfixed(-426407656.0/4294967296.0,1,-nbitq), 
to_sfixed(-83718437.0/4294967296.0,1,-nbitq), 
to_sfixed(159893916.0/4294967296.0,1,-nbitq), 
to_sfixed(229109577.0/4294967296.0,1,-nbitq), 
to_sfixed(-54688503.0/4294967296.0,1,-nbitq), 
to_sfixed(170059945.0/4294967296.0,1,-nbitq), 
to_sfixed(-163534869.0/4294967296.0,1,-nbitq), 
to_sfixed(302901436.0/4294967296.0,1,-nbitq), 
to_sfixed(-348248489.0/4294967296.0,1,-nbitq), 
to_sfixed(-212459523.0/4294967296.0,1,-nbitq), 
to_sfixed(-190403777.0/4294967296.0,1,-nbitq), 
to_sfixed(-253998380.0/4294967296.0,1,-nbitq), 
to_sfixed(41090663.0/4294967296.0,1,-nbitq), 
to_sfixed(23108805.0/4294967296.0,1,-nbitq), 
to_sfixed(-389942032.0/4294967296.0,1,-nbitq), 
to_sfixed(-295592923.0/4294967296.0,1,-nbitq), 
to_sfixed(-119034468.0/4294967296.0,1,-nbitq), 
to_sfixed(414541751.0/4294967296.0,1,-nbitq), 
to_sfixed(184885409.0/4294967296.0,1,-nbitq), 
to_sfixed(-410169791.0/4294967296.0,1,-nbitq), 
to_sfixed(265998370.0/4294967296.0,1,-nbitq), 
to_sfixed(-49781714.0/4294967296.0,1,-nbitq), 
to_sfixed(141572882.0/4294967296.0,1,-nbitq), 
to_sfixed(-273783167.0/4294967296.0,1,-nbitq), 
to_sfixed(220189321.0/4294967296.0,1,-nbitq), 
to_sfixed(133891156.0/4294967296.0,1,-nbitq), 
to_sfixed(-194580430.0/4294967296.0,1,-nbitq), 
to_sfixed(68070950.0/4294967296.0,1,-nbitq), 
to_sfixed(207621151.0/4294967296.0,1,-nbitq), 
to_sfixed(-459541962.0/4294967296.0,1,-nbitq), 
to_sfixed(4147738.0/4294967296.0,1,-nbitq), 
to_sfixed(-6674675.0/4294967296.0,1,-nbitq), 
to_sfixed(201112615.0/4294967296.0,1,-nbitq), 
to_sfixed(482960688.0/4294967296.0,1,-nbitq), 
to_sfixed(217703078.0/4294967296.0,1,-nbitq), 
to_sfixed(-103748346.0/4294967296.0,1,-nbitq), 
to_sfixed(317760936.0/4294967296.0,1,-nbitq), 
to_sfixed(204667726.0/4294967296.0,1,-nbitq), 
to_sfixed(-216095132.0/4294967296.0,1,-nbitq), 
to_sfixed(-247968048.0/4294967296.0,1,-nbitq), 
to_sfixed(-273070908.0/4294967296.0,1,-nbitq), 
to_sfixed(-335796061.0/4294967296.0,1,-nbitq), 
to_sfixed(71185053.0/4294967296.0,1,-nbitq), 
to_sfixed(-78320459.0/4294967296.0,1,-nbitq), 
to_sfixed(-220258747.0/4294967296.0,1,-nbitq), 
to_sfixed(95657545.0/4294967296.0,1,-nbitq), 
to_sfixed(89185331.0/4294967296.0,1,-nbitq), 
to_sfixed(362528115.0/4294967296.0,1,-nbitq), 
to_sfixed(120058340.0/4294967296.0,1,-nbitq), 
to_sfixed(353064763.0/4294967296.0,1,-nbitq), 
to_sfixed(-198966405.0/4294967296.0,1,-nbitq), 
to_sfixed(-105094202.0/4294967296.0,1,-nbitq), 
to_sfixed(-27488977.0/4294967296.0,1,-nbitq), 
to_sfixed(-201077982.0/4294967296.0,1,-nbitq), 
to_sfixed(-287948218.0/4294967296.0,1,-nbitq), 
to_sfixed(380930102.0/4294967296.0,1,-nbitq), 
to_sfixed(-126937889.0/4294967296.0,1,-nbitq), 
to_sfixed(-25243972.0/4294967296.0,1,-nbitq), 
to_sfixed(37273923.0/4294967296.0,1,-nbitq), 
to_sfixed(115038698.0/4294967296.0,1,-nbitq), 
to_sfixed(397384374.0/4294967296.0,1,-nbitq), 
to_sfixed(-222391910.0/4294967296.0,1,-nbitq), 
to_sfixed(340109253.0/4294967296.0,1,-nbitq), 
to_sfixed(101301863.0/4294967296.0,1,-nbitq), 
to_sfixed(117905198.0/4294967296.0,1,-nbitq), 
to_sfixed(472620999.0/4294967296.0,1,-nbitq), 
to_sfixed(79064742.0/4294967296.0,1,-nbitq), 
to_sfixed(99132819.0/4294967296.0,1,-nbitq), 
to_sfixed(475479220.0/4294967296.0,1,-nbitq), 
to_sfixed(10545594.0/4294967296.0,1,-nbitq), 
to_sfixed(-374239949.0/4294967296.0,1,-nbitq), 
to_sfixed(131702150.0/4294967296.0,1,-nbitq), 
to_sfixed(-125789959.0/4294967296.0,1,-nbitq), 
to_sfixed(210371713.0/4294967296.0,1,-nbitq), 
to_sfixed(-17714081.0/4294967296.0,1,-nbitq), 
to_sfixed(128844102.0/4294967296.0,1,-nbitq), 
to_sfixed(319779492.0/4294967296.0,1,-nbitq), 
to_sfixed(-430721017.0/4294967296.0,1,-nbitq), 
to_sfixed(29961124.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(246978907.0/4294967296.0,1,-nbitq), 
to_sfixed(-60799171.0/4294967296.0,1,-nbitq), 
to_sfixed(-412551672.0/4294967296.0,1,-nbitq), 
to_sfixed(17837159.0/4294967296.0,1,-nbitq), 
to_sfixed(-191936904.0/4294967296.0,1,-nbitq), 
to_sfixed(56135957.0/4294967296.0,1,-nbitq), 
to_sfixed(244513113.0/4294967296.0,1,-nbitq), 
to_sfixed(-31489393.0/4294967296.0,1,-nbitq), 
to_sfixed(-206117772.0/4294967296.0,1,-nbitq), 
to_sfixed(-46206521.0/4294967296.0,1,-nbitq), 
to_sfixed(313025261.0/4294967296.0,1,-nbitq), 
to_sfixed(-116267947.0/4294967296.0,1,-nbitq), 
to_sfixed(-278499507.0/4294967296.0,1,-nbitq), 
to_sfixed(508391030.0/4294967296.0,1,-nbitq), 
to_sfixed(303156035.0/4294967296.0,1,-nbitq), 
to_sfixed(-155067175.0/4294967296.0,1,-nbitq), 
to_sfixed(-308060680.0/4294967296.0,1,-nbitq), 
to_sfixed(203217767.0/4294967296.0,1,-nbitq), 
to_sfixed(-6451953.0/4294967296.0,1,-nbitq), 
to_sfixed(152374255.0/4294967296.0,1,-nbitq), 
to_sfixed(-239855348.0/4294967296.0,1,-nbitq), 
to_sfixed(346690908.0/4294967296.0,1,-nbitq), 
to_sfixed(157204466.0/4294967296.0,1,-nbitq), 
to_sfixed(389219470.0/4294967296.0,1,-nbitq), 
to_sfixed(-141703100.0/4294967296.0,1,-nbitq), 
to_sfixed(296411906.0/4294967296.0,1,-nbitq), 
to_sfixed(141161554.0/4294967296.0,1,-nbitq), 
to_sfixed(-210938055.0/4294967296.0,1,-nbitq), 
to_sfixed(-199804888.0/4294967296.0,1,-nbitq), 
to_sfixed(379571747.0/4294967296.0,1,-nbitq), 
to_sfixed(-244356732.0/4294967296.0,1,-nbitq), 
to_sfixed(115085126.0/4294967296.0,1,-nbitq), 
to_sfixed(368007263.0/4294967296.0,1,-nbitq), 
to_sfixed(8883455.0/4294967296.0,1,-nbitq), 
to_sfixed(-178829043.0/4294967296.0,1,-nbitq), 
to_sfixed(59299334.0/4294967296.0,1,-nbitq), 
to_sfixed(429691014.0/4294967296.0,1,-nbitq), 
to_sfixed(159841431.0/4294967296.0,1,-nbitq), 
to_sfixed(-278252712.0/4294967296.0,1,-nbitq), 
to_sfixed(364695840.0/4294967296.0,1,-nbitq), 
to_sfixed(93979660.0/4294967296.0,1,-nbitq), 
to_sfixed(215094895.0/4294967296.0,1,-nbitq), 
to_sfixed(267087295.0/4294967296.0,1,-nbitq), 
to_sfixed(11813188.0/4294967296.0,1,-nbitq), 
to_sfixed(-141514341.0/4294967296.0,1,-nbitq), 
to_sfixed(57925261.0/4294967296.0,1,-nbitq), 
to_sfixed(208760018.0/4294967296.0,1,-nbitq), 
to_sfixed(-290391204.0/4294967296.0,1,-nbitq), 
to_sfixed(-388019803.0/4294967296.0,1,-nbitq), 
to_sfixed(355868784.0/4294967296.0,1,-nbitq), 
to_sfixed(388729794.0/4294967296.0,1,-nbitq), 
to_sfixed(112789761.0/4294967296.0,1,-nbitq), 
to_sfixed(188588842.0/4294967296.0,1,-nbitq), 
to_sfixed(-194490455.0/4294967296.0,1,-nbitq), 
to_sfixed(-193978878.0/4294967296.0,1,-nbitq), 
to_sfixed(-137784236.0/4294967296.0,1,-nbitq), 
to_sfixed(286775693.0/4294967296.0,1,-nbitq), 
to_sfixed(-276471071.0/4294967296.0,1,-nbitq), 
to_sfixed(411284808.0/4294967296.0,1,-nbitq), 
to_sfixed(198982029.0/4294967296.0,1,-nbitq), 
to_sfixed(-254583416.0/4294967296.0,1,-nbitq), 
to_sfixed(-76453990.0/4294967296.0,1,-nbitq), 
to_sfixed(-198475586.0/4294967296.0,1,-nbitq), 
to_sfixed(-124369848.0/4294967296.0,1,-nbitq), 
to_sfixed(-182421103.0/4294967296.0,1,-nbitq), 
to_sfixed(-430092835.0/4294967296.0,1,-nbitq), 
to_sfixed(152409880.0/4294967296.0,1,-nbitq), 
to_sfixed(-73498974.0/4294967296.0,1,-nbitq), 
to_sfixed(25571956.0/4294967296.0,1,-nbitq), 
to_sfixed(-189612200.0/4294967296.0,1,-nbitq), 
to_sfixed(-86070169.0/4294967296.0,1,-nbitq), 
to_sfixed(-238084715.0/4294967296.0,1,-nbitq), 
to_sfixed(-384811995.0/4294967296.0,1,-nbitq), 
to_sfixed(-157002684.0/4294967296.0,1,-nbitq), 
to_sfixed(116954440.0/4294967296.0,1,-nbitq), 
to_sfixed(32788278.0/4294967296.0,1,-nbitq), 
to_sfixed(-56750140.0/4294967296.0,1,-nbitq), 
to_sfixed(-191108573.0/4294967296.0,1,-nbitq), 
to_sfixed(-124537820.0/4294967296.0,1,-nbitq), 
to_sfixed(-144473746.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(177506092.0/4294967296.0,1,-nbitq), 
to_sfixed(-213967485.0/4294967296.0,1,-nbitq), 
to_sfixed(144780333.0/4294967296.0,1,-nbitq), 
to_sfixed(276317058.0/4294967296.0,1,-nbitq), 
to_sfixed(401986837.0/4294967296.0,1,-nbitq), 
to_sfixed(114733277.0/4294967296.0,1,-nbitq), 
to_sfixed(-138788702.0/4294967296.0,1,-nbitq), 
to_sfixed(-302699865.0/4294967296.0,1,-nbitq), 
to_sfixed(-646430234.0/4294967296.0,1,-nbitq), 
to_sfixed(312022019.0/4294967296.0,1,-nbitq), 
to_sfixed(27182234.0/4294967296.0,1,-nbitq), 
to_sfixed(316280827.0/4294967296.0,1,-nbitq), 
to_sfixed(267739509.0/4294967296.0,1,-nbitq), 
to_sfixed(-246826585.0/4294967296.0,1,-nbitq), 
to_sfixed(350480845.0/4294967296.0,1,-nbitq), 
to_sfixed(-480436339.0/4294967296.0,1,-nbitq), 
to_sfixed(-198775376.0/4294967296.0,1,-nbitq), 
to_sfixed(29928131.0/4294967296.0,1,-nbitq), 
to_sfixed(32698805.0/4294967296.0,1,-nbitq), 
to_sfixed(320404419.0/4294967296.0,1,-nbitq), 
to_sfixed(-26311162.0/4294967296.0,1,-nbitq), 
to_sfixed(425239176.0/4294967296.0,1,-nbitq), 
to_sfixed(556902655.0/4294967296.0,1,-nbitq), 
to_sfixed(-12211479.0/4294967296.0,1,-nbitq), 
to_sfixed(-305605311.0/4294967296.0,1,-nbitq), 
to_sfixed(351971331.0/4294967296.0,1,-nbitq), 
to_sfixed(394906223.0/4294967296.0,1,-nbitq), 
to_sfixed(-268804714.0/4294967296.0,1,-nbitq), 
to_sfixed(-3355793.0/4294967296.0,1,-nbitq), 
to_sfixed(-99263273.0/4294967296.0,1,-nbitq), 
to_sfixed(-451479919.0/4294967296.0,1,-nbitq), 
to_sfixed(-230321554.0/4294967296.0,1,-nbitq), 
to_sfixed(-338958155.0/4294967296.0,1,-nbitq), 
to_sfixed(193725221.0/4294967296.0,1,-nbitq), 
to_sfixed(39661786.0/4294967296.0,1,-nbitq), 
to_sfixed(-140081674.0/4294967296.0,1,-nbitq), 
to_sfixed(88683829.0/4294967296.0,1,-nbitq), 
to_sfixed(-333483882.0/4294967296.0,1,-nbitq), 
to_sfixed(-60622574.0/4294967296.0,1,-nbitq), 
to_sfixed(247080702.0/4294967296.0,1,-nbitq), 
to_sfixed(236621614.0/4294967296.0,1,-nbitq), 
to_sfixed(347661740.0/4294967296.0,1,-nbitq), 
to_sfixed(88414521.0/4294967296.0,1,-nbitq), 
to_sfixed(-30200976.0/4294967296.0,1,-nbitq), 
to_sfixed(-318673030.0/4294967296.0,1,-nbitq), 
to_sfixed(362800249.0/4294967296.0,1,-nbitq), 
to_sfixed(138216561.0/4294967296.0,1,-nbitq), 
to_sfixed(-472778790.0/4294967296.0,1,-nbitq), 
to_sfixed(-140895895.0/4294967296.0,1,-nbitq), 
to_sfixed(372906149.0/4294967296.0,1,-nbitq), 
to_sfixed(23982194.0/4294967296.0,1,-nbitq), 
to_sfixed(-408003606.0/4294967296.0,1,-nbitq), 
to_sfixed(-366944613.0/4294967296.0,1,-nbitq), 
to_sfixed(-120934844.0/4294967296.0,1,-nbitq), 
to_sfixed(-125065445.0/4294967296.0,1,-nbitq), 
to_sfixed(5960523.0/4294967296.0,1,-nbitq), 
to_sfixed(-173460222.0/4294967296.0,1,-nbitq), 
to_sfixed(-133731160.0/4294967296.0,1,-nbitq), 
to_sfixed(431939425.0/4294967296.0,1,-nbitq), 
to_sfixed(-83440047.0/4294967296.0,1,-nbitq), 
to_sfixed(-182186833.0/4294967296.0,1,-nbitq), 
to_sfixed(439062245.0/4294967296.0,1,-nbitq), 
to_sfixed(-145638779.0/4294967296.0,1,-nbitq), 
to_sfixed(487964771.0/4294967296.0,1,-nbitq), 
to_sfixed(-341811810.0/4294967296.0,1,-nbitq), 
to_sfixed(-387489029.0/4294967296.0,1,-nbitq), 
to_sfixed(560374088.0/4294967296.0,1,-nbitq), 
to_sfixed(-26018402.0/4294967296.0,1,-nbitq), 
to_sfixed(-317719284.0/4294967296.0,1,-nbitq), 
to_sfixed(-239916481.0/4294967296.0,1,-nbitq), 
to_sfixed(-180238593.0/4294967296.0,1,-nbitq), 
to_sfixed(-366919886.0/4294967296.0,1,-nbitq), 
to_sfixed(-350256906.0/4294967296.0,1,-nbitq), 
to_sfixed(94350631.0/4294967296.0,1,-nbitq), 
to_sfixed(392254722.0/4294967296.0,1,-nbitq), 
to_sfixed(-246260031.0/4294967296.0,1,-nbitq), 
to_sfixed(104353319.0/4294967296.0,1,-nbitq), 
to_sfixed(308019646.0/4294967296.0,1,-nbitq), 
to_sfixed(-57163922.0/4294967296.0,1,-nbitq), 
to_sfixed(-29717448.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-350223935.0/4294967296.0,1,-nbitq), 
to_sfixed(-283459574.0/4294967296.0,1,-nbitq), 
to_sfixed(-166606049.0/4294967296.0,1,-nbitq), 
to_sfixed(298575187.0/4294967296.0,1,-nbitq), 
to_sfixed(64474450.0/4294967296.0,1,-nbitq), 
to_sfixed(193304663.0/4294967296.0,1,-nbitq), 
to_sfixed(-15755324.0/4294967296.0,1,-nbitq), 
to_sfixed(244381200.0/4294967296.0,1,-nbitq), 
to_sfixed(233484219.0/4294967296.0,1,-nbitq), 
to_sfixed(158926939.0/4294967296.0,1,-nbitq), 
to_sfixed(-24440750.0/4294967296.0,1,-nbitq), 
to_sfixed(-93569522.0/4294967296.0,1,-nbitq), 
to_sfixed(-203951246.0/4294967296.0,1,-nbitq), 
to_sfixed(449759375.0/4294967296.0,1,-nbitq), 
to_sfixed(135972693.0/4294967296.0,1,-nbitq), 
to_sfixed(165168150.0/4294967296.0,1,-nbitq), 
to_sfixed(-289661938.0/4294967296.0,1,-nbitq), 
to_sfixed(255984030.0/4294967296.0,1,-nbitq), 
to_sfixed(-21167493.0/4294967296.0,1,-nbitq), 
to_sfixed(29255337.0/4294967296.0,1,-nbitq), 
to_sfixed(-378105854.0/4294967296.0,1,-nbitq), 
to_sfixed(101933117.0/4294967296.0,1,-nbitq), 
to_sfixed(478830755.0/4294967296.0,1,-nbitq), 
to_sfixed(-77921610.0/4294967296.0,1,-nbitq), 
to_sfixed(294933001.0/4294967296.0,1,-nbitq), 
to_sfixed(540864903.0/4294967296.0,1,-nbitq), 
to_sfixed(440234661.0/4294967296.0,1,-nbitq), 
to_sfixed(-74940233.0/4294967296.0,1,-nbitq), 
to_sfixed(257652759.0/4294967296.0,1,-nbitq), 
to_sfixed(217100639.0/4294967296.0,1,-nbitq), 
to_sfixed(-296982339.0/4294967296.0,1,-nbitq), 
to_sfixed(-334570062.0/4294967296.0,1,-nbitq), 
to_sfixed(-47198326.0/4294967296.0,1,-nbitq), 
to_sfixed(-142514257.0/4294967296.0,1,-nbitq), 
to_sfixed(-92793184.0/4294967296.0,1,-nbitq), 
to_sfixed(-220644775.0/4294967296.0,1,-nbitq), 
to_sfixed(264892953.0/4294967296.0,1,-nbitq), 
to_sfixed(243538431.0/4294967296.0,1,-nbitq), 
to_sfixed(-241304271.0/4294967296.0,1,-nbitq), 
to_sfixed(166602691.0/4294967296.0,1,-nbitq), 
to_sfixed(-353461087.0/4294967296.0,1,-nbitq), 
to_sfixed(289139557.0/4294967296.0,1,-nbitq), 
to_sfixed(-269466477.0/4294967296.0,1,-nbitq), 
to_sfixed(222892087.0/4294967296.0,1,-nbitq), 
to_sfixed(301932065.0/4294967296.0,1,-nbitq), 
to_sfixed(350147888.0/4294967296.0,1,-nbitq), 
to_sfixed(-41253245.0/4294967296.0,1,-nbitq), 
to_sfixed(-297525351.0/4294967296.0,1,-nbitq), 
to_sfixed(83150647.0/4294967296.0,1,-nbitq), 
to_sfixed(543172605.0/4294967296.0,1,-nbitq), 
to_sfixed(369346131.0/4294967296.0,1,-nbitq), 
to_sfixed(368402269.0/4294967296.0,1,-nbitq), 
to_sfixed(271066330.0/4294967296.0,1,-nbitq), 
to_sfixed(-115570539.0/4294967296.0,1,-nbitq), 
to_sfixed(-155558376.0/4294967296.0,1,-nbitq), 
to_sfixed(-186818300.0/4294967296.0,1,-nbitq), 
to_sfixed(-210368438.0/4294967296.0,1,-nbitq), 
to_sfixed(201086213.0/4294967296.0,1,-nbitq), 
to_sfixed(-219564963.0/4294967296.0,1,-nbitq), 
to_sfixed(28999445.0/4294967296.0,1,-nbitq), 
to_sfixed(-305885714.0/4294967296.0,1,-nbitq), 
to_sfixed(-206915944.0/4294967296.0,1,-nbitq), 
to_sfixed(-154719065.0/4294967296.0,1,-nbitq), 
to_sfixed(175802441.0/4294967296.0,1,-nbitq), 
to_sfixed(348346518.0/4294967296.0,1,-nbitq), 
to_sfixed(32123262.0/4294967296.0,1,-nbitq), 
to_sfixed(557295309.0/4294967296.0,1,-nbitq), 
to_sfixed(-235111578.0/4294967296.0,1,-nbitq), 
to_sfixed(-100289412.0/4294967296.0,1,-nbitq), 
to_sfixed(-134176462.0/4294967296.0,1,-nbitq), 
to_sfixed(-13653252.0/4294967296.0,1,-nbitq), 
to_sfixed(-14579485.0/4294967296.0,1,-nbitq), 
to_sfixed(48433203.0/4294967296.0,1,-nbitq), 
to_sfixed(288230066.0/4294967296.0,1,-nbitq), 
to_sfixed(452457912.0/4294967296.0,1,-nbitq), 
to_sfixed(-257088541.0/4294967296.0,1,-nbitq), 
to_sfixed(-41714842.0/4294967296.0,1,-nbitq), 
to_sfixed(-344113466.0/4294967296.0,1,-nbitq), 
to_sfixed(238898033.0/4294967296.0,1,-nbitq), 
to_sfixed(-344416227.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-328785493.0/4294967296.0,1,-nbitq), 
to_sfixed(-729353417.0/4294967296.0,1,-nbitq), 
to_sfixed(214923670.0/4294967296.0,1,-nbitq), 
to_sfixed(-184883587.0/4294967296.0,1,-nbitq), 
to_sfixed(283986102.0/4294967296.0,1,-nbitq), 
to_sfixed(7863451.0/4294967296.0,1,-nbitq), 
to_sfixed(-186059854.0/4294967296.0,1,-nbitq), 
to_sfixed(-268586312.0/4294967296.0,1,-nbitq), 
to_sfixed(243561327.0/4294967296.0,1,-nbitq), 
to_sfixed(-57324064.0/4294967296.0,1,-nbitq), 
to_sfixed(-422162557.0/4294967296.0,1,-nbitq), 
to_sfixed(-179624653.0/4294967296.0,1,-nbitq), 
to_sfixed(-330920497.0/4294967296.0,1,-nbitq), 
to_sfixed(136690832.0/4294967296.0,1,-nbitq), 
to_sfixed(87903056.0/4294967296.0,1,-nbitq), 
to_sfixed(-387228289.0/4294967296.0,1,-nbitq), 
to_sfixed(-29306719.0/4294967296.0,1,-nbitq), 
to_sfixed(255523334.0/4294967296.0,1,-nbitq), 
to_sfixed(81409173.0/4294967296.0,1,-nbitq), 
to_sfixed(-593568058.0/4294967296.0,1,-nbitq), 
to_sfixed(-239410821.0/4294967296.0,1,-nbitq), 
to_sfixed(16542648.0/4294967296.0,1,-nbitq), 
to_sfixed(-141577769.0/4294967296.0,1,-nbitq), 
to_sfixed(56719895.0/4294967296.0,1,-nbitq), 
to_sfixed(-298340175.0/4294967296.0,1,-nbitq), 
to_sfixed(506629283.0/4294967296.0,1,-nbitq), 
to_sfixed(56098021.0/4294967296.0,1,-nbitq), 
to_sfixed(133792193.0/4294967296.0,1,-nbitq), 
to_sfixed(-43651317.0/4294967296.0,1,-nbitq), 
to_sfixed(160500084.0/4294967296.0,1,-nbitq), 
to_sfixed(18388463.0/4294967296.0,1,-nbitq), 
to_sfixed(-296439739.0/4294967296.0,1,-nbitq), 
to_sfixed(193777337.0/4294967296.0,1,-nbitq), 
to_sfixed(274807027.0/4294967296.0,1,-nbitq), 
to_sfixed(-18022903.0/4294967296.0,1,-nbitq), 
to_sfixed(353210685.0/4294967296.0,1,-nbitq), 
to_sfixed(84971343.0/4294967296.0,1,-nbitq), 
to_sfixed(528940015.0/4294967296.0,1,-nbitq), 
to_sfixed(364071895.0/4294967296.0,1,-nbitq), 
to_sfixed(457232546.0/4294967296.0,1,-nbitq), 
to_sfixed(-60387551.0/4294967296.0,1,-nbitq), 
to_sfixed(212594834.0/4294967296.0,1,-nbitq), 
to_sfixed(186363415.0/4294967296.0,1,-nbitq), 
to_sfixed(149255078.0/4294967296.0,1,-nbitq), 
to_sfixed(-130250052.0/4294967296.0,1,-nbitq), 
to_sfixed(-160314214.0/4294967296.0,1,-nbitq), 
to_sfixed(311065842.0/4294967296.0,1,-nbitq), 
to_sfixed(-599505664.0/4294967296.0,1,-nbitq), 
to_sfixed(-326700383.0/4294967296.0,1,-nbitq), 
to_sfixed(326342749.0/4294967296.0,1,-nbitq), 
to_sfixed(-293128423.0/4294967296.0,1,-nbitq), 
to_sfixed(-62763837.0/4294967296.0,1,-nbitq), 
to_sfixed(309000347.0/4294967296.0,1,-nbitq), 
to_sfixed(-600844878.0/4294967296.0,1,-nbitq), 
to_sfixed(131414171.0/4294967296.0,1,-nbitq), 
to_sfixed(-66687623.0/4294967296.0,1,-nbitq), 
to_sfixed(207088057.0/4294967296.0,1,-nbitq), 
to_sfixed(177820338.0/4294967296.0,1,-nbitq), 
to_sfixed(344738858.0/4294967296.0,1,-nbitq), 
to_sfixed(385878700.0/4294967296.0,1,-nbitq), 
to_sfixed(197109608.0/4294967296.0,1,-nbitq), 
to_sfixed(556967489.0/4294967296.0,1,-nbitq), 
to_sfixed(-219305303.0/4294967296.0,1,-nbitq), 
to_sfixed(265771672.0/4294967296.0,1,-nbitq), 
to_sfixed(-147384132.0/4294967296.0,1,-nbitq), 
to_sfixed(-475489371.0/4294967296.0,1,-nbitq), 
to_sfixed(5582164.0/4294967296.0,1,-nbitq), 
to_sfixed(455732221.0/4294967296.0,1,-nbitq), 
to_sfixed(-230827193.0/4294967296.0,1,-nbitq), 
to_sfixed(-14588410.0/4294967296.0,1,-nbitq), 
to_sfixed(116727693.0/4294967296.0,1,-nbitq), 
to_sfixed(149238735.0/4294967296.0,1,-nbitq), 
to_sfixed(-429863396.0/4294967296.0,1,-nbitq), 
to_sfixed(-218578540.0/4294967296.0,1,-nbitq), 
to_sfixed(-129519754.0/4294967296.0,1,-nbitq), 
to_sfixed(-411472466.0/4294967296.0,1,-nbitq), 
to_sfixed(-309002052.0/4294967296.0,1,-nbitq), 
to_sfixed(176328577.0/4294967296.0,1,-nbitq), 
to_sfixed(-223261857.0/4294967296.0,1,-nbitq), 
to_sfixed(56450432.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-130750050.0/4294967296.0,1,-nbitq), 
to_sfixed(-700138213.0/4294967296.0,1,-nbitq), 
to_sfixed(561837829.0/4294967296.0,1,-nbitq), 
to_sfixed(542968535.0/4294967296.0,1,-nbitq), 
to_sfixed(258166951.0/4294967296.0,1,-nbitq), 
to_sfixed(313864531.0/4294967296.0,1,-nbitq), 
to_sfixed(254922002.0/4294967296.0,1,-nbitq), 
to_sfixed(121588859.0/4294967296.0,1,-nbitq), 
to_sfixed(207039692.0/4294967296.0,1,-nbitq), 
to_sfixed(102085725.0/4294967296.0,1,-nbitq), 
to_sfixed(6239710.0/4294967296.0,1,-nbitq), 
to_sfixed(-270895800.0/4294967296.0,1,-nbitq), 
to_sfixed(118178169.0/4294967296.0,1,-nbitq), 
to_sfixed(169397193.0/4294967296.0,1,-nbitq), 
to_sfixed(168892150.0/4294967296.0,1,-nbitq), 
to_sfixed(-16578470.0/4294967296.0,1,-nbitq), 
to_sfixed(-84612674.0/4294967296.0,1,-nbitq), 
to_sfixed(-230771461.0/4294967296.0,1,-nbitq), 
to_sfixed(-221727842.0/4294967296.0,1,-nbitq), 
to_sfixed(-239416996.0/4294967296.0,1,-nbitq), 
to_sfixed(11334098.0/4294967296.0,1,-nbitq), 
to_sfixed(-53111848.0/4294967296.0,1,-nbitq), 
to_sfixed(-493958473.0/4294967296.0,1,-nbitq), 
to_sfixed(-181529929.0/4294967296.0,1,-nbitq), 
to_sfixed(-118956789.0/4294967296.0,1,-nbitq), 
to_sfixed(307386615.0/4294967296.0,1,-nbitq), 
to_sfixed(354333201.0/4294967296.0,1,-nbitq), 
to_sfixed(250633445.0/4294967296.0,1,-nbitq), 
to_sfixed(313998647.0/4294967296.0,1,-nbitq), 
to_sfixed(121963578.0/4294967296.0,1,-nbitq), 
to_sfixed(273831671.0/4294967296.0,1,-nbitq), 
to_sfixed(-288380532.0/4294967296.0,1,-nbitq), 
to_sfixed(101517411.0/4294967296.0,1,-nbitq), 
to_sfixed(207894634.0/4294967296.0,1,-nbitq), 
to_sfixed(194794618.0/4294967296.0,1,-nbitq), 
to_sfixed(154599939.0/4294967296.0,1,-nbitq), 
to_sfixed(211411977.0/4294967296.0,1,-nbitq), 
to_sfixed(577361774.0/4294967296.0,1,-nbitq), 
to_sfixed(-216580375.0/4294967296.0,1,-nbitq), 
to_sfixed(-258836063.0/4294967296.0,1,-nbitq), 
to_sfixed(9459465.0/4294967296.0,1,-nbitq), 
to_sfixed(33859279.0/4294967296.0,1,-nbitq), 
to_sfixed(427211667.0/4294967296.0,1,-nbitq), 
to_sfixed(-16760719.0/4294967296.0,1,-nbitq), 
to_sfixed(-423123486.0/4294967296.0,1,-nbitq), 
to_sfixed(163320978.0/4294967296.0,1,-nbitq), 
to_sfixed(-425407312.0/4294967296.0,1,-nbitq), 
to_sfixed(18845783.0/4294967296.0,1,-nbitq), 
to_sfixed(52458370.0/4294967296.0,1,-nbitq), 
to_sfixed(-237965376.0/4294967296.0,1,-nbitq), 
to_sfixed(208521792.0/4294967296.0,1,-nbitq), 
to_sfixed(-244390942.0/4294967296.0,1,-nbitq), 
to_sfixed(530340655.0/4294967296.0,1,-nbitq), 
to_sfixed(-235257542.0/4294967296.0,1,-nbitq), 
to_sfixed(257586628.0/4294967296.0,1,-nbitq), 
to_sfixed(20896624.0/4294967296.0,1,-nbitq), 
to_sfixed(119065373.0/4294967296.0,1,-nbitq), 
to_sfixed(3617051.0/4294967296.0,1,-nbitq), 
to_sfixed(136574405.0/4294967296.0,1,-nbitq), 
to_sfixed(325329913.0/4294967296.0,1,-nbitq), 
to_sfixed(-275039974.0/4294967296.0,1,-nbitq), 
to_sfixed(250845554.0/4294967296.0,1,-nbitq), 
to_sfixed(-470799848.0/4294967296.0,1,-nbitq), 
to_sfixed(73714393.0/4294967296.0,1,-nbitq), 
to_sfixed(-328214216.0/4294967296.0,1,-nbitq), 
to_sfixed(-194793000.0/4294967296.0,1,-nbitq), 
to_sfixed(178707923.0/4294967296.0,1,-nbitq), 
to_sfixed(636083503.0/4294967296.0,1,-nbitq), 
to_sfixed(11865887.0/4294967296.0,1,-nbitq), 
to_sfixed(258272885.0/4294967296.0,1,-nbitq), 
to_sfixed(87799069.0/4294967296.0,1,-nbitq), 
to_sfixed(357259576.0/4294967296.0,1,-nbitq), 
to_sfixed(187379798.0/4294967296.0,1,-nbitq), 
to_sfixed(-295588986.0/4294967296.0,1,-nbitq), 
to_sfixed(75238843.0/4294967296.0,1,-nbitq), 
to_sfixed(-245868219.0/4294967296.0,1,-nbitq), 
to_sfixed(188223374.0/4294967296.0,1,-nbitq), 
to_sfixed(-17482522.0/4294967296.0,1,-nbitq), 
to_sfixed(397878504.0/4294967296.0,1,-nbitq), 
to_sfixed(-114751833.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-64915730.0/4294967296.0,1,-nbitq), 
to_sfixed(456916599.0/4294967296.0,1,-nbitq), 
to_sfixed(320920094.0/4294967296.0,1,-nbitq), 
to_sfixed(974761832.0/4294967296.0,1,-nbitq), 
to_sfixed(288870656.0/4294967296.0,1,-nbitq), 
to_sfixed(426187497.0/4294967296.0,1,-nbitq), 
to_sfixed(14857582.0/4294967296.0,1,-nbitq), 
to_sfixed(123934587.0/4294967296.0,1,-nbitq), 
to_sfixed(-269060449.0/4294967296.0,1,-nbitq), 
to_sfixed(374620749.0/4294967296.0,1,-nbitq), 
to_sfixed(150243949.0/4294967296.0,1,-nbitq), 
to_sfixed(-169622225.0/4294967296.0,1,-nbitq), 
to_sfixed(702968664.0/4294967296.0,1,-nbitq), 
to_sfixed(-526682526.0/4294967296.0,1,-nbitq), 
to_sfixed(-212542599.0/4294967296.0,1,-nbitq), 
to_sfixed(-407575143.0/4294967296.0,1,-nbitq), 
to_sfixed(36584030.0/4294967296.0,1,-nbitq), 
to_sfixed(31873306.0/4294967296.0,1,-nbitq), 
to_sfixed(236539082.0/4294967296.0,1,-nbitq), 
to_sfixed(-87502125.0/4294967296.0,1,-nbitq), 
to_sfixed(-349681089.0/4294967296.0,1,-nbitq), 
to_sfixed(59228560.0/4294967296.0,1,-nbitq), 
to_sfixed(-232120909.0/4294967296.0,1,-nbitq), 
to_sfixed(115636998.0/4294967296.0,1,-nbitq), 
to_sfixed(-136193734.0/4294967296.0,1,-nbitq), 
to_sfixed(105771261.0/4294967296.0,1,-nbitq), 
to_sfixed(226220517.0/4294967296.0,1,-nbitq), 
to_sfixed(-52367094.0/4294967296.0,1,-nbitq), 
to_sfixed(-157930739.0/4294967296.0,1,-nbitq), 
to_sfixed(-59299024.0/4294967296.0,1,-nbitq), 
to_sfixed(6690270.0/4294967296.0,1,-nbitq), 
to_sfixed(-904560215.0/4294967296.0,1,-nbitq), 
to_sfixed(-90006030.0/4294967296.0,1,-nbitq), 
to_sfixed(-90875092.0/4294967296.0,1,-nbitq), 
to_sfixed(-472652572.0/4294967296.0,1,-nbitq), 
to_sfixed(566870990.0/4294967296.0,1,-nbitq), 
to_sfixed(-215965344.0/4294967296.0,1,-nbitq), 
to_sfixed(548002721.0/4294967296.0,1,-nbitq), 
to_sfixed(-104193471.0/4294967296.0,1,-nbitq), 
to_sfixed(59302959.0/4294967296.0,1,-nbitq), 
to_sfixed(80639593.0/4294967296.0,1,-nbitq), 
to_sfixed(-111750888.0/4294967296.0,1,-nbitq), 
to_sfixed(108490420.0/4294967296.0,1,-nbitq), 
to_sfixed(-731806840.0/4294967296.0,1,-nbitq), 
to_sfixed(107756149.0/4294967296.0,1,-nbitq), 
to_sfixed(-34417507.0/4294967296.0,1,-nbitq), 
to_sfixed(-244293753.0/4294967296.0,1,-nbitq), 
to_sfixed(-93898547.0/4294967296.0,1,-nbitq), 
to_sfixed(456047582.0/4294967296.0,1,-nbitq), 
to_sfixed(64490418.0/4294967296.0,1,-nbitq), 
to_sfixed(64683375.0/4294967296.0,1,-nbitq), 
to_sfixed(319595843.0/4294967296.0,1,-nbitq), 
to_sfixed(923931740.0/4294967296.0,1,-nbitq), 
to_sfixed(-907357905.0/4294967296.0,1,-nbitq), 
to_sfixed(118847851.0/4294967296.0,1,-nbitq), 
to_sfixed(616576874.0/4294967296.0,1,-nbitq), 
to_sfixed(15696869.0/4294967296.0,1,-nbitq), 
to_sfixed(629557616.0/4294967296.0,1,-nbitq), 
to_sfixed(429024289.0/4294967296.0,1,-nbitq), 
to_sfixed(-292653234.0/4294967296.0,1,-nbitq), 
to_sfixed(190370255.0/4294967296.0,1,-nbitq), 
to_sfixed(-19647683.0/4294967296.0,1,-nbitq), 
to_sfixed(-589354912.0/4294967296.0,1,-nbitq), 
to_sfixed(840433171.0/4294967296.0,1,-nbitq), 
to_sfixed(47519763.0/4294967296.0,1,-nbitq), 
to_sfixed(204665963.0/4294967296.0,1,-nbitq), 
to_sfixed(-199605655.0/4294967296.0,1,-nbitq), 
to_sfixed(663351462.0/4294967296.0,1,-nbitq), 
to_sfixed(79346288.0/4294967296.0,1,-nbitq), 
to_sfixed(-102223229.0/4294967296.0,1,-nbitq), 
to_sfixed(-341196497.0/4294967296.0,1,-nbitq), 
to_sfixed(-162963001.0/4294967296.0,1,-nbitq), 
to_sfixed(-284461170.0/4294967296.0,1,-nbitq), 
to_sfixed(360126259.0/4294967296.0,1,-nbitq), 
to_sfixed(232049106.0/4294967296.0,1,-nbitq), 
to_sfixed(-1305669478.0/4294967296.0,1,-nbitq), 
to_sfixed(265685443.0/4294967296.0,1,-nbitq), 
to_sfixed(-295920869.0/4294967296.0,1,-nbitq), 
to_sfixed(50385945.0/4294967296.0,1,-nbitq), 
to_sfixed(-120428719.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(58401166.0/4294967296.0,1,-nbitq), 
to_sfixed(555318923.0/4294967296.0,1,-nbitq), 
to_sfixed(381266498.0/4294967296.0,1,-nbitq), 
to_sfixed(942108468.0/4294967296.0,1,-nbitq), 
to_sfixed(546992862.0/4294967296.0,1,-nbitq), 
to_sfixed(613870905.0/4294967296.0,1,-nbitq), 
to_sfixed(333743610.0/4294967296.0,1,-nbitq), 
to_sfixed(61137269.0/4294967296.0,1,-nbitq), 
to_sfixed(92324105.0/4294967296.0,1,-nbitq), 
to_sfixed(48844299.0/4294967296.0,1,-nbitq), 
to_sfixed(570290238.0/4294967296.0,1,-nbitq), 
to_sfixed(-671199995.0/4294967296.0,1,-nbitq), 
to_sfixed(195779483.0/4294967296.0,1,-nbitq), 
to_sfixed(-325395965.0/4294967296.0,1,-nbitq), 
to_sfixed(-346541272.0/4294967296.0,1,-nbitq), 
to_sfixed(-477141624.0/4294967296.0,1,-nbitq), 
to_sfixed(56366912.0/4294967296.0,1,-nbitq), 
to_sfixed(-140341293.0/4294967296.0,1,-nbitq), 
to_sfixed(141875943.0/4294967296.0,1,-nbitq), 
to_sfixed(414390883.0/4294967296.0,1,-nbitq), 
to_sfixed(101225090.0/4294967296.0,1,-nbitq), 
to_sfixed(-472642900.0/4294967296.0,1,-nbitq), 
to_sfixed(305266220.0/4294967296.0,1,-nbitq), 
to_sfixed(-2401180.0/4294967296.0,1,-nbitq), 
to_sfixed(265660454.0/4294967296.0,1,-nbitq), 
to_sfixed(-356209921.0/4294967296.0,1,-nbitq), 
to_sfixed(-167759102.0/4294967296.0,1,-nbitq), 
to_sfixed(-229874461.0/4294967296.0,1,-nbitq), 
to_sfixed(382363412.0/4294967296.0,1,-nbitq), 
to_sfixed(-840232796.0/4294967296.0,1,-nbitq), 
to_sfixed(27498569.0/4294967296.0,1,-nbitq), 
to_sfixed(-674072895.0/4294967296.0,1,-nbitq), 
to_sfixed(-189163031.0/4294967296.0,1,-nbitq), 
to_sfixed(-254926800.0/4294967296.0,1,-nbitq), 
to_sfixed(-445465960.0/4294967296.0,1,-nbitq), 
to_sfixed(-271659984.0/4294967296.0,1,-nbitq), 
to_sfixed(-403979679.0/4294967296.0,1,-nbitq), 
to_sfixed(248281484.0/4294967296.0,1,-nbitq), 
to_sfixed(-173865485.0/4294967296.0,1,-nbitq), 
to_sfixed(417099061.0/4294967296.0,1,-nbitq), 
to_sfixed(-333740060.0/4294967296.0,1,-nbitq), 
to_sfixed(-566827071.0/4294967296.0,1,-nbitq), 
to_sfixed(-466143415.0/4294967296.0,1,-nbitq), 
to_sfixed(-792642952.0/4294967296.0,1,-nbitq), 
to_sfixed(555683204.0/4294967296.0,1,-nbitq), 
to_sfixed(-158362500.0/4294967296.0,1,-nbitq), 
to_sfixed(-74409849.0/4294967296.0,1,-nbitq), 
to_sfixed(28683000.0/4294967296.0,1,-nbitq), 
to_sfixed(-183173118.0/4294967296.0,1,-nbitq), 
to_sfixed(-122861406.0/4294967296.0,1,-nbitq), 
to_sfixed(182717572.0/4294967296.0,1,-nbitq), 
to_sfixed(223059602.0/4294967296.0,1,-nbitq), 
to_sfixed(951325331.0/4294967296.0,1,-nbitq), 
to_sfixed(-15722313.0/4294967296.0,1,-nbitq), 
to_sfixed(131104433.0/4294967296.0,1,-nbitq), 
to_sfixed(1055578496.0/4294967296.0,1,-nbitq), 
to_sfixed(-84393998.0/4294967296.0,1,-nbitq), 
to_sfixed(430385317.0/4294967296.0,1,-nbitq), 
to_sfixed(405665575.0/4294967296.0,1,-nbitq), 
to_sfixed(222758658.0/4294967296.0,1,-nbitq), 
to_sfixed(-356933453.0/4294967296.0,1,-nbitq), 
to_sfixed(206914228.0/4294967296.0,1,-nbitq), 
to_sfixed(-716685321.0/4294967296.0,1,-nbitq), 
to_sfixed(894255059.0/4294967296.0,1,-nbitq), 
to_sfixed(52303244.0/4294967296.0,1,-nbitq), 
to_sfixed(-161075084.0/4294967296.0,1,-nbitq), 
to_sfixed(-208217747.0/4294967296.0,1,-nbitq), 
to_sfixed(586760768.0/4294967296.0,1,-nbitq), 
to_sfixed(225283902.0/4294967296.0,1,-nbitq), 
to_sfixed(-289440790.0/4294967296.0,1,-nbitq), 
to_sfixed(-934478547.0/4294967296.0,1,-nbitq), 
to_sfixed(129915520.0/4294967296.0,1,-nbitq), 
to_sfixed(-20355204.0/4294967296.0,1,-nbitq), 
to_sfixed(51194272.0/4294967296.0,1,-nbitq), 
to_sfixed(184200487.0/4294967296.0,1,-nbitq), 
to_sfixed(-446065322.0/4294967296.0,1,-nbitq), 
to_sfixed(172706065.0/4294967296.0,1,-nbitq), 
to_sfixed(-113286766.0/4294967296.0,1,-nbitq), 
to_sfixed(118385272.0/4294967296.0,1,-nbitq), 
to_sfixed(4863473.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(539977774.0/4294967296.0,1,-nbitq), 
to_sfixed(299596498.0/4294967296.0,1,-nbitq), 
to_sfixed(354363017.0/4294967296.0,1,-nbitq), 
to_sfixed(711820403.0/4294967296.0,1,-nbitq), 
to_sfixed(987116650.0/4294967296.0,1,-nbitq), 
to_sfixed(479023330.0/4294967296.0,1,-nbitq), 
to_sfixed(53901138.0/4294967296.0,1,-nbitq), 
to_sfixed(-120096624.0/4294967296.0,1,-nbitq), 
to_sfixed(520933987.0/4294967296.0,1,-nbitq), 
to_sfixed(351852898.0/4294967296.0,1,-nbitq), 
to_sfixed(-194061685.0/4294967296.0,1,-nbitq), 
to_sfixed(-713786224.0/4294967296.0,1,-nbitq), 
to_sfixed(198895849.0/4294967296.0,1,-nbitq), 
to_sfixed(-516909010.0/4294967296.0,1,-nbitq), 
to_sfixed(-228476839.0/4294967296.0,1,-nbitq), 
to_sfixed(-680152395.0/4294967296.0,1,-nbitq), 
to_sfixed(119026872.0/4294967296.0,1,-nbitq), 
to_sfixed(90978088.0/4294967296.0,1,-nbitq), 
to_sfixed(387082320.0/4294967296.0,1,-nbitq), 
to_sfixed(454566882.0/4294967296.0,1,-nbitq), 
to_sfixed(-152628961.0/4294967296.0,1,-nbitq), 
to_sfixed(-126015977.0/4294967296.0,1,-nbitq), 
to_sfixed(76083041.0/4294967296.0,1,-nbitq), 
to_sfixed(610080645.0/4294967296.0,1,-nbitq), 
to_sfixed(-151697617.0/4294967296.0,1,-nbitq), 
to_sfixed(-922453333.0/4294967296.0,1,-nbitq), 
to_sfixed(-80129695.0/4294967296.0,1,-nbitq), 
to_sfixed(111258918.0/4294967296.0,1,-nbitq), 
to_sfixed(356385667.0/4294967296.0,1,-nbitq), 
to_sfixed(-1129111032.0/4294967296.0,1,-nbitq), 
to_sfixed(130309843.0/4294967296.0,1,-nbitq), 
to_sfixed(-211296329.0/4294967296.0,1,-nbitq), 
to_sfixed(-116477081.0/4294967296.0,1,-nbitq), 
to_sfixed(-179721043.0/4294967296.0,1,-nbitq), 
to_sfixed(212304850.0/4294967296.0,1,-nbitq), 
to_sfixed(-160895588.0/4294967296.0,1,-nbitq), 
to_sfixed(-48259146.0/4294967296.0,1,-nbitq), 
to_sfixed(595633304.0/4294967296.0,1,-nbitq), 
to_sfixed(-596933926.0/4294967296.0,1,-nbitq), 
to_sfixed(534083949.0/4294967296.0,1,-nbitq), 
to_sfixed(101258447.0/4294967296.0,1,-nbitq), 
to_sfixed(-583591336.0/4294967296.0,1,-nbitq), 
to_sfixed(334342447.0/4294967296.0,1,-nbitq), 
to_sfixed(-205499337.0/4294967296.0,1,-nbitq), 
to_sfixed(154002677.0/4294967296.0,1,-nbitq), 
to_sfixed(-310765355.0/4294967296.0,1,-nbitq), 
to_sfixed(132791590.0/4294967296.0,1,-nbitq), 
to_sfixed(-134573822.0/4294967296.0,1,-nbitq), 
to_sfixed(-225067500.0/4294967296.0,1,-nbitq), 
to_sfixed(-44717440.0/4294967296.0,1,-nbitq), 
to_sfixed(-42964115.0/4294967296.0,1,-nbitq), 
to_sfixed(126368560.0/4294967296.0,1,-nbitq), 
to_sfixed(1365470085.0/4294967296.0,1,-nbitq), 
to_sfixed(-289711485.0/4294967296.0,1,-nbitq), 
to_sfixed(441253536.0/4294967296.0,1,-nbitq), 
to_sfixed(1158049072.0/4294967296.0,1,-nbitq), 
to_sfixed(-349924946.0/4294967296.0,1,-nbitq), 
to_sfixed(-111163601.0/4294967296.0,1,-nbitq), 
to_sfixed(24582703.0/4294967296.0,1,-nbitq), 
to_sfixed(-279322372.0/4294967296.0,1,-nbitq), 
to_sfixed(101628722.0/4294967296.0,1,-nbitq), 
to_sfixed(-358185913.0/4294967296.0,1,-nbitq), 
to_sfixed(-1097494801.0/4294967296.0,1,-nbitq), 
to_sfixed(1389608850.0/4294967296.0,1,-nbitq), 
to_sfixed(-472297985.0/4294967296.0,1,-nbitq), 
to_sfixed(-290811746.0/4294967296.0,1,-nbitq), 
to_sfixed(-338454868.0/4294967296.0,1,-nbitq), 
to_sfixed(684064281.0/4294967296.0,1,-nbitq), 
to_sfixed(87290116.0/4294967296.0,1,-nbitq), 
to_sfixed(-1404678108.0/4294967296.0,1,-nbitq), 
to_sfixed(-910514987.0/4294967296.0,1,-nbitq), 
to_sfixed(15258279.0/4294967296.0,1,-nbitq), 
to_sfixed(-183692463.0/4294967296.0,1,-nbitq), 
to_sfixed(-318316807.0/4294967296.0,1,-nbitq), 
to_sfixed(8024048.0/4294967296.0,1,-nbitq), 
to_sfixed(-174991266.0/4294967296.0,1,-nbitq), 
to_sfixed(586685406.0/4294967296.0,1,-nbitq), 
to_sfixed(48099757.0/4294967296.0,1,-nbitq), 
to_sfixed(-187456949.0/4294967296.0,1,-nbitq), 
to_sfixed(-291315613.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(261241901.0/4294967296.0,1,-nbitq), 
to_sfixed(-47081534.0/4294967296.0,1,-nbitq), 
to_sfixed(929617926.0/4294967296.0,1,-nbitq), 
to_sfixed(44097300.0/4294967296.0,1,-nbitq), 
to_sfixed(1395339264.0/4294967296.0,1,-nbitq), 
to_sfixed(807227819.0/4294967296.0,1,-nbitq), 
to_sfixed(112284519.0/4294967296.0,1,-nbitq), 
to_sfixed(-104687830.0/4294967296.0,1,-nbitq), 
to_sfixed(322968526.0/4294967296.0,1,-nbitq), 
to_sfixed(-278224205.0/4294967296.0,1,-nbitq), 
to_sfixed(522875441.0/4294967296.0,1,-nbitq), 
to_sfixed(-260264717.0/4294967296.0,1,-nbitq), 
to_sfixed(14251642.0/4294967296.0,1,-nbitq), 
to_sfixed(-1132062874.0/4294967296.0,1,-nbitq), 
to_sfixed(29423876.0/4294967296.0,1,-nbitq), 
to_sfixed(-426990519.0/4294967296.0,1,-nbitq), 
to_sfixed(-392422831.0/4294967296.0,1,-nbitq), 
to_sfixed(96627119.0/4294967296.0,1,-nbitq), 
to_sfixed(751406246.0/4294967296.0,1,-nbitq), 
to_sfixed(1003335830.0/4294967296.0,1,-nbitq), 
to_sfixed(-206338464.0/4294967296.0,1,-nbitq), 
to_sfixed(98853605.0/4294967296.0,1,-nbitq), 
to_sfixed(-234637740.0/4294967296.0,1,-nbitq), 
to_sfixed(9591072.0/4294967296.0,1,-nbitq), 
to_sfixed(-149971419.0/4294967296.0,1,-nbitq), 
to_sfixed(-547793263.0/4294967296.0,1,-nbitq), 
to_sfixed(-188883684.0/4294967296.0,1,-nbitq), 
to_sfixed(141145642.0/4294967296.0,1,-nbitq), 
to_sfixed(-14088909.0/4294967296.0,1,-nbitq), 
to_sfixed(-847040723.0/4294967296.0,1,-nbitq), 
to_sfixed(291290384.0/4294967296.0,1,-nbitq), 
to_sfixed(-307879961.0/4294967296.0,1,-nbitq), 
to_sfixed(-26136938.0/4294967296.0,1,-nbitq), 
to_sfixed(-31556200.0/4294967296.0,1,-nbitq), 
to_sfixed(-157522757.0/4294967296.0,1,-nbitq), 
to_sfixed(207358824.0/4294967296.0,1,-nbitq), 
to_sfixed(127237997.0/4294967296.0,1,-nbitq), 
to_sfixed(572354690.0/4294967296.0,1,-nbitq), 
to_sfixed(151040387.0/4294967296.0,1,-nbitq), 
to_sfixed(569721481.0/4294967296.0,1,-nbitq), 
to_sfixed(-523404256.0/4294967296.0,1,-nbitq), 
to_sfixed(-593343885.0/4294967296.0,1,-nbitq), 
to_sfixed(-60354040.0/4294967296.0,1,-nbitq), 
to_sfixed(-341443821.0/4294967296.0,1,-nbitq), 
to_sfixed(73481010.0/4294967296.0,1,-nbitq), 
to_sfixed(730166184.0/4294967296.0,1,-nbitq), 
to_sfixed(-418088953.0/4294967296.0,1,-nbitq), 
to_sfixed(-225465684.0/4294967296.0,1,-nbitq), 
to_sfixed(-241165321.0/4294967296.0,1,-nbitq), 
to_sfixed(359298277.0/4294967296.0,1,-nbitq), 
to_sfixed(299975736.0/4294967296.0,1,-nbitq), 
to_sfixed(24699378.0/4294967296.0,1,-nbitq), 
to_sfixed(847100676.0/4294967296.0,1,-nbitq), 
to_sfixed(-9955243.0/4294967296.0,1,-nbitq), 
to_sfixed(113984138.0/4294967296.0,1,-nbitq), 
to_sfixed(774571280.0/4294967296.0,1,-nbitq), 
to_sfixed(31669981.0/4294967296.0,1,-nbitq), 
to_sfixed(150464298.0/4294967296.0,1,-nbitq), 
to_sfixed(142814282.0/4294967296.0,1,-nbitq), 
to_sfixed(310010364.0/4294967296.0,1,-nbitq), 
to_sfixed(-117287637.0/4294967296.0,1,-nbitq), 
to_sfixed(-14650818.0/4294967296.0,1,-nbitq), 
to_sfixed(-398740785.0/4294967296.0,1,-nbitq), 
to_sfixed(1167470585.0/4294967296.0,1,-nbitq), 
to_sfixed(282825370.0/4294967296.0,1,-nbitq), 
to_sfixed(-312992007.0/4294967296.0,1,-nbitq), 
to_sfixed(-1137811489.0/4294967296.0,1,-nbitq), 
to_sfixed(-744738735.0/4294967296.0,1,-nbitq), 
to_sfixed(-139035301.0/4294967296.0,1,-nbitq), 
to_sfixed(-347376033.0/4294967296.0,1,-nbitq), 
to_sfixed(-1084583966.0/4294967296.0,1,-nbitq), 
to_sfixed(57324973.0/4294967296.0,1,-nbitq), 
to_sfixed(416420384.0/4294967296.0,1,-nbitq), 
to_sfixed(318346516.0/4294967296.0,1,-nbitq), 
to_sfixed(-172592036.0/4294967296.0,1,-nbitq), 
to_sfixed(70228159.0/4294967296.0,1,-nbitq), 
to_sfixed(1122767794.0/4294967296.0,1,-nbitq), 
to_sfixed(109578911.0/4294967296.0,1,-nbitq), 
to_sfixed(-174272849.0/4294967296.0,1,-nbitq), 
to_sfixed(-32976609.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-143912236.0/4294967296.0,1,-nbitq), 
to_sfixed(-962354101.0/4294967296.0,1,-nbitq), 
to_sfixed(797744767.0/4294967296.0,1,-nbitq), 
to_sfixed(-359424197.0/4294967296.0,1,-nbitq), 
to_sfixed(593824435.0/4294967296.0,1,-nbitq), 
to_sfixed(464368611.0/4294967296.0,1,-nbitq), 
to_sfixed(133074655.0/4294967296.0,1,-nbitq), 
to_sfixed(-103368460.0/4294967296.0,1,-nbitq), 
to_sfixed(930661361.0/4294967296.0,1,-nbitq), 
to_sfixed(383874906.0/4294967296.0,1,-nbitq), 
to_sfixed(-40809809.0/4294967296.0,1,-nbitq), 
to_sfixed(-573690128.0/4294967296.0,1,-nbitq), 
to_sfixed(-174442037.0/4294967296.0,1,-nbitq), 
to_sfixed(-843971720.0/4294967296.0,1,-nbitq), 
to_sfixed(446108305.0/4294967296.0,1,-nbitq), 
to_sfixed(-1103398453.0/4294967296.0,1,-nbitq), 
to_sfixed(-151734570.0/4294967296.0,1,-nbitq), 
to_sfixed(-151216896.0/4294967296.0,1,-nbitq), 
to_sfixed(349831726.0/4294967296.0,1,-nbitq), 
to_sfixed(620477200.0/4294967296.0,1,-nbitq), 
to_sfixed(343016997.0/4294967296.0,1,-nbitq), 
to_sfixed(391202523.0/4294967296.0,1,-nbitq), 
to_sfixed(273978676.0/4294967296.0,1,-nbitq), 
to_sfixed(-269834854.0/4294967296.0,1,-nbitq), 
to_sfixed(117489135.0/4294967296.0,1,-nbitq), 
to_sfixed(-1055053540.0/4294967296.0,1,-nbitq), 
to_sfixed(191508692.0/4294967296.0,1,-nbitq), 
to_sfixed(295892849.0/4294967296.0,1,-nbitq), 
to_sfixed(197941457.0/4294967296.0,1,-nbitq), 
to_sfixed(-562855000.0/4294967296.0,1,-nbitq), 
to_sfixed(254471136.0/4294967296.0,1,-nbitq), 
to_sfixed(-345087157.0/4294967296.0,1,-nbitq), 
to_sfixed(143178116.0/4294967296.0,1,-nbitq), 
to_sfixed(272341790.0/4294967296.0,1,-nbitq), 
to_sfixed(-611318682.0/4294967296.0,1,-nbitq), 
to_sfixed(68277653.0/4294967296.0,1,-nbitq), 
to_sfixed(78480822.0/4294967296.0,1,-nbitq), 
to_sfixed(590457349.0/4294967296.0,1,-nbitq), 
to_sfixed(156038300.0/4294967296.0,1,-nbitq), 
to_sfixed(-44054020.0/4294967296.0,1,-nbitq), 
to_sfixed(223269994.0/4294967296.0,1,-nbitq), 
to_sfixed(89758174.0/4294967296.0,1,-nbitq), 
to_sfixed(9992136.0/4294967296.0,1,-nbitq), 
to_sfixed(-1050727121.0/4294967296.0,1,-nbitq), 
to_sfixed(694298534.0/4294967296.0,1,-nbitq), 
to_sfixed(256956.0/4294967296.0,1,-nbitq), 
to_sfixed(-12469650.0/4294967296.0,1,-nbitq), 
to_sfixed(-247106580.0/4294967296.0,1,-nbitq), 
to_sfixed(19589921.0/4294967296.0,1,-nbitq), 
to_sfixed(671415611.0/4294967296.0,1,-nbitq), 
to_sfixed(226577750.0/4294967296.0,1,-nbitq), 
to_sfixed(331728384.0/4294967296.0,1,-nbitq), 
to_sfixed(639316815.0/4294967296.0,1,-nbitq), 
to_sfixed(-1197001903.0/4294967296.0,1,-nbitq), 
to_sfixed(-288479203.0/4294967296.0,1,-nbitq), 
to_sfixed(478400924.0/4294967296.0,1,-nbitq), 
to_sfixed(171267801.0/4294967296.0,1,-nbitq), 
to_sfixed(1106743004.0/4294967296.0,1,-nbitq), 
to_sfixed(-158464298.0/4294967296.0,1,-nbitq), 
to_sfixed(360023616.0/4294967296.0,1,-nbitq), 
to_sfixed(-39385564.0/4294967296.0,1,-nbitq), 
to_sfixed(242191564.0/4294967296.0,1,-nbitq), 
to_sfixed(85480923.0/4294967296.0,1,-nbitq), 
to_sfixed(1431654361.0/4294967296.0,1,-nbitq), 
to_sfixed(81683729.0/4294967296.0,1,-nbitq), 
to_sfixed(134438566.0/4294967296.0,1,-nbitq), 
to_sfixed(-561940935.0/4294967296.0,1,-nbitq), 
to_sfixed(-191392186.0/4294967296.0,1,-nbitq), 
to_sfixed(-277376044.0/4294967296.0,1,-nbitq), 
to_sfixed(-625036140.0/4294967296.0,1,-nbitq), 
to_sfixed(-1179359891.0/4294967296.0,1,-nbitq), 
to_sfixed(401365703.0/4294967296.0,1,-nbitq), 
to_sfixed(19150532.0/4294967296.0,1,-nbitq), 
to_sfixed(173573270.0/4294967296.0,1,-nbitq), 
to_sfixed(493527427.0/4294967296.0,1,-nbitq), 
to_sfixed(295749127.0/4294967296.0,1,-nbitq), 
to_sfixed(871859790.0/4294967296.0,1,-nbitq), 
to_sfixed(214581919.0/4294967296.0,1,-nbitq), 
to_sfixed(-53071132.0/4294967296.0,1,-nbitq), 
to_sfixed(-235850034.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-465168978.0/4294967296.0,1,-nbitq), 
to_sfixed(-641647074.0/4294967296.0,1,-nbitq), 
to_sfixed(636821644.0/4294967296.0,1,-nbitq), 
to_sfixed(325109519.0/4294967296.0,1,-nbitq), 
to_sfixed(1216783598.0/4294967296.0,1,-nbitq), 
to_sfixed(223157859.0/4294967296.0,1,-nbitq), 
to_sfixed(-348409857.0/4294967296.0,1,-nbitq), 
to_sfixed(-387816368.0/4294967296.0,1,-nbitq), 
to_sfixed(1075460668.0/4294967296.0,1,-nbitq), 
to_sfixed(-165076071.0/4294967296.0,1,-nbitq), 
to_sfixed(-300100379.0/4294967296.0,1,-nbitq), 
to_sfixed(-336426333.0/4294967296.0,1,-nbitq), 
to_sfixed(-727787661.0/4294967296.0,1,-nbitq), 
to_sfixed(-1982146840.0/4294967296.0,1,-nbitq), 
to_sfixed(198423322.0/4294967296.0,1,-nbitq), 
to_sfixed(-760509331.0/4294967296.0,1,-nbitq), 
to_sfixed(392358707.0/4294967296.0,1,-nbitq), 
to_sfixed(253091773.0/4294967296.0,1,-nbitq), 
to_sfixed(565787140.0/4294967296.0,1,-nbitq), 
to_sfixed(252345152.0/4294967296.0,1,-nbitq), 
to_sfixed(-98298054.0/4294967296.0,1,-nbitq), 
to_sfixed(982802093.0/4294967296.0,1,-nbitq), 
to_sfixed(-515025217.0/4294967296.0,1,-nbitq), 
to_sfixed(-999939776.0/4294967296.0,1,-nbitq), 
to_sfixed(187030476.0/4294967296.0,1,-nbitq), 
to_sfixed(-998613273.0/4294967296.0,1,-nbitq), 
to_sfixed(-184436190.0/4294967296.0,1,-nbitq), 
to_sfixed(794575374.0/4294967296.0,1,-nbitq), 
to_sfixed(188577990.0/4294967296.0,1,-nbitq), 
to_sfixed(-470723045.0/4294967296.0,1,-nbitq), 
to_sfixed(890395655.0/4294967296.0,1,-nbitq), 
to_sfixed(345560599.0/4294967296.0,1,-nbitq), 
to_sfixed(542095349.0/4294967296.0,1,-nbitq), 
to_sfixed(78199364.0/4294967296.0,1,-nbitq), 
to_sfixed(-248312351.0/4294967296.0,1,-nbitq), 
to_sfixed(822461772.0/4294967296.0,1,-nbitq), 
to_sfixed(3535330.0/4294967296.0,1,-nbitq), 
to_sfixed(-401798013.0/4294967296.0,1,-nbitq), 
to_sfixed(449117396.0/4294967296.0,1,-nbitq), 
to_sfixed(606491457.0/4294967296.0,1,-nbitq), 
to_sfixed(-79864214.0/4294967296.0,1,-nbitq), 
to_sfixed(-470278143.0/4294967296.0,1,-nbitq), 
to_sfixed(261685319.0/4294967296.0,1,-nbitq), 
to_sfixed(-1280066378.0/4294967296.0,1,-nbitq), 
to_sfixed(205109157.0/4294967296.0,1,-nbitq), 
to_sfixed(-111192832.0/4294967296.0,1,-nbitq), 
to_sfixed(143011982.0/4294967296.0,1,-nbitq), 
to_sfixed(-757292027.0/4294967296.0,1,-nbitq), 
to_sfixed(125903190.0/4294967296.0,1,-nbitq), 
to_sfixed(645741187.0/4294967296.0,1,-nbitq), 
to_sfixed(183803232.0/4294967296.0,1,-nbitq), 
to_sfixed(91856945.0/4294967296.0,1,-nbitq), 
to_sfixed(893004398.0/4294967296.0,1,-nbitq), 
to_sfixed(-426352838.0/4294967296.0,1,-nbitq), 
to_sfixed(-780860257.0/4294967296.0,1,-nbitq), 
to_sfixed(-311679601.0/4294967296.0,1,-nbitq), 
to_sfixed(-133055278.0/4294967296.0,1,-nbitq), 
to_sfixed(724535308.0/4294967296.0,1,-nbitq), 
to_sfixed(214261930.0/4294967296.0,1,-nbitq), 
to_sfixed(-169121824.0/4294967296.0,1,-nbitq), 
to_sfixed(-233218461.0/4294967296.0,1,-nbitq), 
to_sfixed(1119807.0/4294967296.0,1,-nbitq), 
to_sfixed(581391313.0/4294967296.0,1,-nbitq), 
to_sfixed(420971137.0/4294967296.0,1,-nbitq), 
to_sfixed(-2311810.0/4294967296.0,1,-nbitq), 
to_sfixed(244951385.0/4294967296.0,1,-nbitq), 
to_sfixed(-516125156.0/4294967296.0,1,-nbitq), 
to_sfixed(-262976094.0/4294967296.0,1,-nbitq), 
to_sfixed(384303034.0/4294967296.0,1,-nbitq), 
to_sfixed(523599711.0/4294967296.0,1,-nbitq), 
to_sfixed(-1064777967.0/4294967296.0,1,-nbitq), 
to_sfixed(472133766.0/4294967296.0,1,-nbitq), 
to_sfixed(434098328.0/4294967296.0,1,-nbitq), 
to_sfixed(264004772.0/4294967296.0,1,-nbitq), 
to_sfixed(-81028959.0/4294967296.0,1,-nbitq), 
to_sfixed(443069951.0/4294967296.0,1,-nbitq), 
to_sfixed(1291491839.0/4294967296.0,1,-nbitq), 
to_sfixed(206832505.0/4294967296.0,1,-nbitq), 
to_sfixed(-55565581.0/4294967296.0,1,-nbitq), 
to_sfixed(-267668086.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(89836649.0/4294967296.0,1,-nbitq), 
to_sfixed(-558458349.0/4294967296.0,1,-nbitq), 
to_sfixed(1024658108.0/4294967296.0,1,-nbitq), 
to_sfixed(210751710.0/4294967296.0,1,-nbitq), 
to_sfixed(880012822.0/4294967296.0,1,-nbitq), 
to_sfixed(-252306363.0/4294967296.0,1,-nbitq), 
to_sfixed(-98237842.0/4294967296.0,1,-nbitq), 
to_sfixed(-42560432.0/4294967296.0,1,-nbitq), 
to_sfixed(699502801.0/4294967296.0,1,-nbitq), 
to_sfixed(-111899293.0/4294967296.0,1,-nbitq), 
to_sfixed(-847098686.0/4294967296.0,1,-nbitq), 
to_sfixed(-680175172.0/4294967296.0,1,-nbitq), 
to_sfixed(-455650676.0/4294967296.0,1,-nbitq), 
to_sfixed(-1243687819.0/4294967296.0,1,-nbitq), 
to_sfixed(231803856.0/4294967296.0,1,-nbitq), 
to_sfixed(-903402248.0/4294967296.0,1,-nbitq), 
to_sfixed(296233135.0/4294967296.0,1,-nbitq), 
to_sfixed(-95051773.0/4294967296.0,1,-nbitq), 
to_sfixed(391520813.0/4294967296.0,1,-nbitq), 
to_sfixed(-158807362.0/4294967296.0,1,-nbitq), 
to_sfixed(-114964198.0/4294967296.0,1,-nbitq), 
to_sfixed(650186492.0/4294967296.0,1,-nbitq), 
to_sfixed(-384462986.0/4294967296.0,1,-nbitq), 
to_sfixed(-658245718.0/4294967296.0,1,-nbitq), 
to_sfixed(325004551.0/4294967296.0,1,-nbitq), 
to_sfixed(-296006158.0/4294967296.0,1,-nbitq), 
to_sfixed(-437968055.0/4294967296.0,1,-nbitq), 
to_sfixed(971516557.0/4294967296.0,1,-nbitq), 
to_sfixed(-232602265.0/4294967296.0,1,-nbitq), 
to_sfixed(-1054760733.0/4294967296.0,1,-nbitq), 
to_sfixed(1148764343.0/4294967296.0,1,-nbitq), 
to_sfixed(206242018.0/4294967296.0,1,-nbitq), 
to_sfixed(-33962817.0/4294967296.0,1,-nbitq), 
to_sfixed(-136199307.0/4294967296.0,1,-nbitq), 
to_sfixed(-463875427.0/4294967296.0,1,-nbitq), 
to_sfixed(181226911.0/4294967296.0,1,-nbitq), 
to_sfixed(-164218194.0/4294967296.0,1,-nbitq), 
to_sfixed(-745502373.0/4294967296.0,1,-nbitq), 
to_sfixed(-188553038.0/4294967296.0,1,-nbitq), 
to_sfixed(-164361672.0/4294967296.0,1,-nbitq), 
to_sfixed(30890178.0/4294967296.0,1,-nbitq), 
to_sfixed(-94183096.0/4294967296.0,1,-nbitq), 
to_sfixed(547695550.0/4294967296.0,1,-nbitq), 
to_sfixed(-855698932.0/4294967296.0,1,-nbitq), 
to_sfixed(266284167.0/4294967296.0,1,-nbitq), 
to_sfixed(2206434.0/4294967296.0,1,-nbitq), 
to_sfixed(132700813.0/4294967296.0,1,-nbitq), 
to_sfixed(-958855712.0/4294967296.0,1,-nbitq), 
to_sfixed(252283863.0/4294967296.0,1,-nbitq), 
to_sfixed(507711467.0/4294967296.0,1,-nbitq), 
to_sfixed(-439176359.0/4294967296.0,1,-nbitq), 
to_sfixed(195749005.0/4294967296.0,1,-nbitq), 
to_sfixed(-58569602.0/4294967296.0,1,-nbitq), 
to_sfixed(-900220668.0/4294967296.0,1,-nbitq), 
to_sfixed(-1146246805.0/4294967296.0,1,-nbitq), 
to_sfixed(-253871475.0/4294967296.0,1,-nbitq), 
to_sfixed(-21455283.0/4294967296.0,1,-nbitq), 
to_sfixed(347368560.0/4294967296.0,1,-nbitq), 
to_sfixed(139802158.0/4294967296.0,1,-nbitq), 
to_sfixed(62620930.0/4294967296.0,1,-nbitq), 
to_sfixed(-264686096.0/4294967296.0,1,-nbitq), 
to_sfixed(272525550.0/4294967296.0,1,-nbitq), 
to_sfixed(973368364.0/4294967296.0,1,-nbitq), 
to_sfixed(113974640.0/4294967296.0,1,-nbitq), 
to_sfixed(356758431.0/4294967296.0,1,-nbitq), 
to_sfixed(309354759.0/4294967296.0,1,-nbitq), 
to_sfixed(-70226579.0/4294967296.0,1,-nbitq), 
to_sfixed(-100246277.0/4294967296.0,1,-nbitq), 
to_sfixed(231363321.0/4294967296.0,1,-nbitq), 
to_sfixed(-546058296.0/4294967296.0,1,-nbitq), 
to_sfixed(-1341790523.0/4294967296.0,1,-nbitq), 
to_sfixed(376195190.0/4294967296.0,1,-nbitq), 
to_sfixed(220403877.0/4294967296.0,1,-nbitq), 
to_sfixed(-257812555.0/4294967296.0,1,-nbitq), 
to_sfixed(-53109857.0/4294967296.0,1,-nbitq), 
to_sfixed(-89310907.0/4294967296.0,1,-nbitq), 
to_sfixed(1650126398.0/4294967296.0,1,-nbitq), 
to_sfixed(669070775.0/4294967296.0,1,-nbitq), 
to_sfixed(-215026125.0/4294967296.0,1,-nbitq), 
to_sfixed(-152643322.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-59014174.0/4294967296.0,1,-nbitq), 
to_sfixed(-957299460.0/4294967296.0,1,-nbitq), 
to_sfixed(741364722.0/4294967296.0,1,-nbitq), 
to_sfixed(1123811386.0/4294967296.0,1,-nbitq), 
to_sfixed(307208626.0/4294967296.0,1,-nbitq), 
to_sfixed(-471492205.0/4294967296.0,1,-nbitq), 
to_sfixed(-180794327.0/4294967296.0,1,-nbitq), 
to_sfixed(166131470.0/4294967296.0,1,-nbitq), 
to_sfixed(936562811.0/4294967296.0,1,-nbitq), 
to_sfixed(-63619271.0/4294967296.0,1,-nbitq), 
to_sfixed(-1175706637.0/4294967296.0,1,-nbitq), 
to_sfixed(-475307920.0/4294967296.0,1,-nbitq), 
to_sfixed(-226518255.0/4294967296.0,1,-nbitq), 
to_sfixed(-721965037.0/4294967296.0,1,-nbitq), 
to_sfixed(148538710.0/4294967296.0,1,-nbitq), 
to_sfixed(-630815030.0/4294967296.0,1,-nbitq), 
to_sfixed(8433023.0/4294967296.0,1,-nbitq), 
to_sfixed(-218702112.0/4294967296.0,1,-nbitq), 
to_sfixed(-361052307.0/4294967296.0,1,-nbitq), 
to_sfixed(-590755542.0/4294967296.0,1,-nbitq), 
to_sfixed(-180493932.0/4294967296.0,1,-nbitq), 
to_sfixed(225820730.0/4294967296.0,1,-nbitq), 
to_sfixed(-368715468.0/4294967296.0,1,-nbitq), 
to_sfixed(-542848625.0/4294967296.0,1,-nbitq), 
to_sfixed(244683826.0/4294967296.0,1,-nbitq), 
to_sfixed(-344210035.0/4294967296.0,1,-nbitq), 
to_sfixed(-728397776.0/4294967296.0,1,-nbitq), 
to_sfixed(895762711.0/4294967296.0,1,-nbitq), 
to_sfixed(-214878335.0/4294967296.0,1,-nbitq), 
to_sfixed(-204430848.0/4294967296.0,1,-nbitq), 
to_sfixed(687080357.0/4294967296.0,1,-nbitq), 
to_sfixed(908439826.0/4294967296.0,1,-nbitq), 
to_sfixed(-102313115.0/4294967296.0,1,-nbitq), 
to_sfixed(479206601.0/4294967296.0,1,-nbitq), 
to_sfixed(-322004777.0/4294967296.0,1,-nbitq), 
to_sfixed(476200113.0/4294967296.0,1,-nbitq), 
to_sfixed(89012005.0/4294967296.0,1,-nbitq), 
to_sfixed(-481543365.0/4294967296.0,1,-nbitq), 
to_sfixed(189096018.0/4294967296.0,1,-nbitq), 
to_sfixed(-243870211.0/4294967296.0,1,-nbitq), 
to_sfixed(125939751.0/4294967296.0,1,-nbitq), 
to_sfixed(-264302408.0/4294967296.0,1,-nbitq), 
to_sfixed(507587072.0/4294967296.0,1,-nbitq), 
to_sfixed(-710999813.0/4294967296.0,1,-nbitq), 
to_sfixed(155659361.0/4294967296.0,1,-nbitq), 
to_sfixed(-865176986.0/4294967296.0,1,-nbitq), 
to_sfixed(49003113.0/4294967296.0,1,-nbitq), 
to_sfixed(-744854437.0/4294967296.0,1,-nbitq), 
to_sfixed(-282593912.0/4294967296.0,1,-nbitq), 
to_sfixed(922434595.0/4294967296.0,1,-nbitq), 
to_sfixed(-360582041.0/4294967296.0,1,-nbitq), 
to_sfixed(513614601.0/4294967296.0,1,-nbitq), 
to_sfixed(-446168573.0/4294967296.0,1,-nbitq), 
to_sfixed(-1205583648.0/4294967296.0,1,-nbitq), 
to_sfixed(-546576608.0/4294967296.0,1,-nbitq), 
to_sfixed(237775654.0/4294967296.0,1,-nbitq), 
to_sfixed(105251239.0/4294967296.0,1,-nbitq), 
to_sfixed(-333656939.0/4294967296.0,1,-nbitq), 
to_sfixed(107691140.0/4294967296.0,1,-nbitq), 
to_sfixed(224371935.0/4294967296.0,1,-nbitq), 
to_sfixed(-174144471.0/4294967296.0,1,-nbitq), 
to_sfixed(392873207.0/4294967296.0,1,-nbitq), 
to_sfixed(1638412371.0/4294967296.0,1,-nbitq), 
to_sfixed(290138526.0/4294967296.0,1,-nbitq), 
to_sfixed(-141096584.0/4294967296.0,1,-nbitq), 
to_sfixed(277041372.0/4294967296.0,1,-nbitq), 
to_sfixed(229112077.0/4294967296.0,1,-nbitq), 
to_sfixed(-945598890.0/4294967296.0,1,-nbitq), 
to_sfixed(253487759.0/4294967296.0,1,-nbitq), 
to_sfixed(-365024662.0/4294967296.0,1,-nbitq), 
to_sfixed(-621239768.0/4294967296.0,1,-nbitq), 
to_sfixed(286711880.0/4294967296.0,1,-nbitq), 
to_sfixed(398034154.0/4294967296.0,1,-nbitq), 
to_sfixed(141294912.0/4294967296.0,1,-nbitq), 
to_sfixed(-486618511.0/4294967296.0,1,-nbitq), 
to_sfixed(408347110.0/4294967296.0,1,-nbitq), 
to_sfixed(1786487002.0/4294967296.0,1,-nbitq), 
to_sfixed(139034231.0/4294967296.0,1,-nbitq), 
to_sfixed(-266969388.0/4294967296.0,1,-nbitq), 
to_sfixed(-264710301.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-333484645.0/4294967296.0,1,-nbitq), 
to_sfixed(-12379993.0/4294967296.0,1,-nbitq), 
to_sfixed(505204891.0/4294967296.0,1,-nbitq), 
to_sfixed(-198904446.0/4294967296.0,1,-nbitq), 
to_sfixed(402328664.0/4294967296.0,1,-nbitq), 
to_sfixed(-316852457.0/4294967296.0,1,-nbitq), 
to_sfixed(69017803.0/4294967296.0,1,-nbitq), 
to_sfixed(117001517.0/4294967296.0,1,-nbitq), 
to_sfixed(363276426.0/4294967296.0,1,-nbitq), 
to_sfixed(-225232815.0/4294967296.0,1,-nbitq), 
to_sfixed(-288767089.0/4294967296.0,1,-nbitq), 
to_sfixed(-395083872.0/4294967296.0,1,-nbitq), 
to_sfixed(201566672.0/4294967296.0,1,-nbitq), 
to_sfixed(-652562481.0/4294967296.0,1,-nbitq), 
to_sfixed(114105328.0/4294967296.0,1,-nbitq), 
to_sfixed(-3145493.0/4294967296.0,1,-nbitq), 
to_sfixed(176484199.0/4294967296.0,1,-nbitq), 
to_sfixed(149531540.0/4294967296.0,1,-nbitq), 
to_sfixed(301693785.0/4294967296.0,1,-nbitq), 
to_sfixed(-100719059.0/4294967296.0,1,-nbitq), 
to_sfixed(135679053.0/4294967296.0,1,-nbitq), 
to_sfixed(275291866.0/4294967296.0,1,-nbitq), 
to_sfixed(467167400.0/4294967296.0,1,-nbitq), 
to_sfixed(-940294199.0/4294967296.0,1,-nbitq), 
to_sfixed(27366333.0/4294967296.0,1,-nbitq), 
to_sfixed(-425793205.0/4294967296.0,1,-nbitq), 
to_sfixed(156237833.0/4294967296.0,1,-nbitq), 
to_sfixed(105632278.0/4294967296.0,1,-nbitq), 
to_sfixed(-718768856.0/4294967296.0,1,-nbitq), 
to_sfixed(-742317560.0/4294967296.0,1,-nbitq), 
to_sfixed(517644123.0/4294967296.0,1,-nbitq), 
to_sfixed(1372233999.0/4294967296.0,1,-nbitq), 
to_sfixed(-322513334.0/4294967296.0,1,-nbitq), 
to_sfixed(380088288.0/4294967296.0,1,-nbitq), 
to_sfixed(-463779950.0/4294967296.0,1,-nbitq), 
to_sfixed(666140684.0/4294967296.0,1,-nbitq), 
to_sfixed(-621019809.0/4294967296.0,1,-nbitq), 
to_sfixed(-635863424.0/4294967296.0,1,-nbitq), 
to_sfixed(-38272966.0/4294967296.0,1,-nbitq), 
to_sfixed(-46852082.0/4294967296.0,1,-nbitq), 
to_sfixed(-801775456.0/4294967296.0,1,-nbitq), 
to_sfixed(150269469.0/4294967296.0,1,-nbitq), 
to_sfixed(729060194.0/4294967296.0,1,-nbitq), 
to_sfixed(-378457661.0/4294967296.0,1,-nbitq), 
to_sfixed(176358688.0/4294967296.0,1,-nbitq), 
to_sfixed(-1619418353.0/4294967296.0,1,-nbitq), 
to_sfixed(239210618.0/4294967296.0,1,-nbitq), 
to_sfixed(-545886796.0/4294967296.0,1,-nbitq), 
to_sfixed(137852439.0/4294967296.0,1,-nbitq), 
to_sfixed(440485241.0/4294967296.0,1,-nbitq), 
to_sfixed(-337875649.0/4294967296.0,1,-nbitq), 
to_sfixed(199054958.0/4294967296.0,1,-nbitq), 
to_sfixed(-8882773.0/4294967296.0,1,-nbitq), 
to_sfixed(-295357734.0/4294967296.0,1,-nbitq), 
to_sfixed(-221004164.0/4294967296.0,1,-nbitq), 
to_sfixed(646936961.0/4294967296.0,1,-nbitq), 
to_sfixed(365940080.0/4294967296.0,1,-nbitq), 
to_sfixed(-442547684.0/4294967296.0,1,-nbitq), 
to_sfixed(159767215.0/4294967296.0,1,-nbitq), 
to_sfixed(-150494525.0/4294967296.0,1,-nbitq), 
to_sfixed(192134597.0/4294967296.0,1,-nbitq), 
to_sfixed(116176869.0/4294967296.0,1,-nbitq), 
to_sfixed(1455798741.0/4294967296.0,1,-nbitq), 
to_sfixed(751927158.0/4294967296.0,1,-nbitq), 
to_sfixed(216321694.0/4294967296.0,1,-nbitq), 
to_sfixed(14785041.0/4294967296.0,1,-nbitq), 
to_sfixed(322598602.0/4294967296.0,1,-nbitq), 
to_sfixed(-964480610.0/4294967296.0,1,-nbitq), 
to_sfixed(-117433795.0/4294967296.0,1,-nbitq), 
to_sfixed(-800117639.0/4294967296.0,1,-nbitq), 
to_sfixed(-200843784.0/4294967296.0,1,-nbitq), 
to_sfixed(344167097.0/4294967296.0,1,-nbitq), 
to_sfixed(437789243.0/4294967296.0,1,-nbitq), 
to_sfixed(-201450887.0/4294967296.0,1,-nbitq), 
to_sfixed(184169629.0/4294967296.0,1,-nbitq), 
to_sfixed(463401379.0/4294967296.0,1,-nbitq), 
to_sfixed(1629550037.0/4294967296.0,1,-nbitq), 
to_sfixed(149472862.0/4294967296.0,1,-nbitq), 
to_sfixed(255892658.0/4294967296.0,1,-nbitq), 
to_sfixed(-146991155.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-105390755.0/4294967296.0,1,-nbitq), 
to_sfixed(-201005384.0/4294967296.0,1,-nbitq), 
to_sfixed(542056783.0/4294967296.0,1,-nbitq), 
to_sfixed(-180025171.0/4294967296.0,1,-nbitq), 
to_sfixed(315503019.0/4294967296.0,1,-nbitq), 
to_sfixed(-411359847.0/4294967296.0,1,-nbitq), 
to_sfixed(-499909185.0/4294967296.0,1,-nbitq), 
to_sfixed(-218907405.0/4294967296.0,1,-nbitq), 
to_sfixed(-1582050.0/4294967296.0,1,-nbitq), 
to_sfixed(159791249.0/4294967296.0,1,-nbitq), 
to_sfixed(785454655.0/4294967296.0,1,-nbitq), 
to_sfixed(-66112694.0/4294967296.0,1,-nbitq), 
to_sfixed(59132054.0/4294967296.0,1,-nbitq), 
to_sfixed(-1219751482.0/4294967296.0,1,-nbitq), 
to_sfixed(-166718829.0/4294967296.0,1,-nbitq), 
to_sfixed(-143647288.0/4294967296.0,1,-nbitq), 
to_sfixed(89487321.0/4294967296.0,1,-nbitq), 
to_sfixed(-248670922.0/4294967296.0,1,-nbitq), 
to_sfixed(-276420249.0/4294967296.0,1,-nbitq), 
to_sfixed(-139418007.0/4294967296.0,1,-nbitq), 
to_sfixed(-281189904.0/4294967296.0,1,-nbitq), 
to_sfixed(-126776016.0/4294967296.0,1,-nbitq), 
to_sfixed(659866902.0/4294967296.0,1,-nbitq), 
to_sfixed(-1151803601.0/4294967296.0,1,-nbitq), 
to_sfixed(-54630823.0/4294967296.0,1,-nbitq), 
to_sfixed(-294980003.0/4294967296.0,1,-nbitq), 
to_sfixed(-16701595.0/4294967296.0,1,-nbitq), 
to_sfixed(-755450492.0/4294967296.0,1,-nbitq), 
to_sfixed(-1024818951.0/4294967296.0,1,-nbitq), 
to_sfixed(-1024186291.0/4294967296.0,1,-nbitq), 
to_sfixed(397533394.0/4294967296.0,1,-nbitq), 
to_sfixed(717979851.0/4294967296.0,1,-nbitq), 
to_sfixed(94011037.0/4294967296.0,1,-nbitq), 
to_sfixed(-79598478.0/4294967296.0,1,-nbitq), 
to_sfixed(-165812949.0/4294967296.0,1,-nbitq), 
to_sfixed(201265665.0/4294967296.0,1,-nbitq), 
to_sfixed(-356075771.0/4294967296.0,1,-nbitq), 
to_sfixed(-439880913.0/4294967296.0,1,-nbitq), 
to_sfixed(-129548086.0/4294967296.0,1,-nbitq), 
to_sfixed(-305276396.0/4294967296.0,1,-nbitq), 
to_sfixed(-554623486.0/4294967296.0,1,-nbitq), 
to_sfixed(21243865.0/4294967296.0,1,-nbitq), 
to_sfixed(1053962375.0/4294967296.0,1,-nbitq), 
to_sfixed(-746245155.0/4294967296.0,1,-nbitq), 
to_sfixed(17689389.0/4294967296.0,1,-nbitq), 
to_sfixed(-1022461858.0/4294967296.0,1,-nbitq), 
to_sfixed(-143070376.0/4294967296.0,1,-nbitq), 
to_sfixed(-681953648.0/4294967296.0,1,-nbitq), 
to_sfixed(172182412.0/4294967296.0,1,-nbitq), 
to_sfixed(668571819.0/4294967296.0,1,-nbitq), 
to_sfixed(-85262004.0/4294967296.0,1,-nbitq), 
to_sfixed(510496394.0/4294967296.0,1,-nbitq), 
to_sfixed(301551492.0/4294967296.0,1,-nbitq), 
to_sfixed(-1217714145.0/4294967296.0,1,-nbitq), 
to_sfixed(635634315.0/4294967296.0,1,-nbitq), 
to_sfixed(-706618018.0/4294967296.0,1,-nbitq), 
to_sfixed(-21475026.0/4294967296.0,1,-nbitq), 
to_sfixed(-2138637.0/4294967296.0,1,-nbitq), 
to_sfixed(58491406.0/4294967296.0,1,-nbitq), 
to_sfixed(-367099999.0/4294967296.0,1,-nbitq), 
to_sfixed(-281769911.0/4294967296.0,1,-nbitq), 
to_sfixed(-27191894.0/4294967296.0,1,-nbitq), 
to_sfixed(610345962.0/4294967296.0,1,-nbitq), 
to_sfixed(368194000.0/4294967296.0,1,-nbitq), 
to_sfixed(71708837.0/4294967296.0,1,-nbitq), 
to_sfixed(-498495855.0/4294967296.0,1,-nbitq), 
to_sfixed(-84620326.0/4294967296.0,1,-nbitq), 
to_sfixed(-187925388.0/4294967296.0,1,-nbitq), 
to_sfixed(210963731.0/4294967296.0,1,-nbitq), 
to_sfixed(-1232403702.0/4294967296.0,1,-nbitq), 
to_sfixed(-129217273.0/4294967296.0,1,-nbitq), 
to_sfixed(186563118.0/4294967296.0,1,-nbitq), 
to_sfixed(431935629.0/4294967296.0,1,-nbitq), 
to_sfixed(346653964.0/4294967296.0,1,-nbitq), 
to_sfixed(-408404842.0/4294967296.0,1,-nbitq), 
to_sfixed(540820100.0/4294967296.0,1,-nbitq), 
to_sfixed(1105782361.0/4294967296.0,1,-nbitq), 
to_sfixed(323065948.0/4294967296.0,1,-nbitq), 
to_sfixed(181199671.0/4294967296.0,1,-nbitq), 
to_sfixed(187902045.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-62876648.0/4294967296.0,1,-nbitq), 
to_sfixed(-745542323.0/4294967296.0,1,-nbitq), 
to_sfixed(501214655.0/4294967296.0,1,-nbitq), 
to_sfixed(-489318529.0/4294967296.0,1,-nbitq), 
to_sfixed(-767229315.0/4294967296.0,1,-nbitq), 
to_sfixed(-1002559118.0/4294967296.0,1,-nbitq), 
to_sfixed(-262827516.0/4294967296.0,1,-nbitq), 
to_sfixed(-122368798.0/4294967296.0,1,-nbitq), 
to_sfixed(188346474.0/4294967296.0,1,-nbitq), 
to_sfixed(269698246.0/4294967296.0,1,-nbitq), 
to_sfixed(419987092.0/4294967296.0,1,-nbitq), 
to_sfixed(231155347.0/4294967296.0,1,-nbitq), 
to_sfixed(333047120.0/4294967296.0,1,-nbitq), 
to_sfixed(-349755549.0/4294967296.0,1,-nbitq), 
to_sfixed(88231366.0/4294967296.0,1,-nbitq), 
to_sfixed(-620204848.0/4294967296.0,1,-nbitq), 
to_sfixed(-891899.0/4294967296.0,1,-nbitq), 
to_sfixed(227499609.0/4294967296.0,1,-nbitq), 
to_sfixed(127275152.0/4294967296.0,1,-nbitq), 
to_sfixed(-10463509.0/4294967296.0,1,-nbitq), 
to_sfixed(197638162.0/4294967296.0,1,-nbitq), 
to_sfixed(-556782550.0/4294967296.0,1,-nbitq), 
to_sfixed(-52467104.0/4294967296.0,1,-nbitq), 
to_sfixed(-85654026.0/4294967296.0,1,-nbitq), 
to_sfixed(-28256614.0/4294967296.0,1,-nbitq), 
to_sfixed(250440497.0/4294967296.0,1,-nbitq), 
to_sfixed(300291369.0/4294967296.0,1,-nbitq), 
to_sfixed(-469726732.0/4294967296.0,1,-nbitq), 
to_sfixed(-694021755.0/4294967296.0,1,-nbitq), 
to_sfixed(-1241225919.0/4294967296.0,1,-nbitq), 
to_sfixed(500490326.0/4294967296.0,1,-nbitq), 
to_sfixed(683826408.0/4294967296.0,1,-nbitq), 
to_sfixed(91135385.0/4294967296.0,1,-nbitq), 
to_sfixed(-184557061.0/4294967296.0,1,-nbitq), 
to_sfixed(143160009.0/4294967296.0,1,-nbitq), 
to_sfixed(-15120012.0/4294967296.0,1,-nbitq), 
to_sfixed(80132221.0/4294967296.0,1,-nbitq), 
to_sfixed(-622602644.0/4294967296.0,1,-nbitq), 
to_sfixed(260976559.0/4294967296.0,1,-nbitq), 
to_sfixed(31244056.0/4294967296.0,1,-nbitq), 
to_sfixed(-227686139.0/4294967296.0,1,-nbitq), 
to_sfixed(451661685.0/4294967296.0,1,-nbitq), 
to_sfixed(953805039.0/4294967296.0,1,-nbitq), 
to_sfixed(91586240.0/4294967296.0,1,-nbitq), 
to_sfixed(114871058.0/4294967296.0,1,-nbitq), 
to_sfixed(-809001726.0/4294967296.0,1,-nbitq), 
to_sfixed(-52739394.0/4294967296.0,1,-nbitq), 
to_sfixed(-818511223.0/4294967296.0,1,-nbitq), 
to_sfixed(-179169467.0/4294967296.0,1,-nbitq), 
to_sfixed(293623549.0/4294967296.0,1,-nbitq), 
to_sfixed(86613407.0/4294967296.0,1,-nbitq), 
to_sfixed(498518735.0/4294967296.0,1,-nbitq), 
to_sfixed(99156303.0/4294967296.0,1,-nbitq), 
to_sfixed(-1228645115.0/4294967296.0,1,-nbitq), 
to_sfixed(845238516.0/4294967296.0,1,-nbitq), 
to_sfixed(-883932192.0/4294967296.0,1,-nbitq), 
to_sfixed(161370849.0/4294967296.0,1,-nbitq), 
to_sfixed(886242024.0/4294967296.0,1,-nbitq), 
to_sfixed(131054094.0/4294967296.0,1,-nbitq), 
to_sfixed(89604526.0/4294967296.0,1,-nbitq), 
to_sfixed(186940534.0/4294967296.0,1,-nbitq), 
to_sfixed(17034430.0/4294967296.0,1,-nbitq), 
to_sfixed(1084850961.0/4294967296.0,1,-nbitq), 
to_sfixed(-54166656.0/4294967296.0,1,-nbitq), 
to_sfixed(-230303562.0/4294967296.0,1,-nbitq), 
to_sfixed(-483398977.0/4294967296.0,1,-nbitq), 
to_sfixed(-370009226.0/4294967296.0,1,-nbitq), 
to_sfixed(-60261224.0/4294967296.0,1,-nbitq), 
to_sfixed(151397915.0/4294967296.0,1,-nbitq), 
to_sfixed(-1291755716.0/4294967296.0,1,-nbitq), 
to_sfixed(936505150.0/4294967296.0,1,-nbitq), 
to_sfixed(-141115104.0/4294967296.0,1,-nbitq), 
to_sfixed(7719291.0/4294967296.0,1,-nbitq), 
to_sfixed(88606645.0/4294967296.0,1,-nbitq), 
to_sfixed(-138957916.0/4294967296.0,1,-nbitq), 
to_sfixed(311242861.0/4294967296.0,1,-nbitq), 
to_sfixed(1368133354.0/4294967296.0,1,-nbitq), 
to_sfixed(256125728.0/4294967296.0,1,-nbitq), 
to_sfixed(440443140.0/4294967296.0,1,-nbitq), 
to_sfixed(105792235.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(218511130.0/4294967296.0,1,-nbitq), 
to_sfixed(388392920.0/4294967296.0,1,-nbitq), 
to_sfixed(-111471401.0/4294967296.0,1,-nbitq), 
to_sfixed(343636784.0/4294967296.0,1,-nbitq), 
to_sfixed(-402606785.0/4294967296.0,1,-nbitq), 
to_sfixed(-1037407731.0/4294967296.0,1,-nbitq), 
to_sfixed(-131870171.0/4294967296.0,1,-nbitq), 
to_sfixed(-536686764.0/4294967296.0,1,-nbitq), 
to_sfixed(940246163.0/4294967296.0,1,-nbitq), 
to_sfixed(-329646093.0/4294967296.0,1,-nbitq), 
to_sfixed(-18378357.0/4294967296.0,1,-nbitq), 
to_sfixed(-224205009.0/4294967296.0,1,-nbitq), 
to_sfixed(-383341461.0/4294967296.0,1,-nbitq), 
to_sfixed(710969740.0/4294967296.0,1,-nbitq), 
to_sfixed(-280003812.0/4294967296.0,1,-nbitq), 
to_sfixed(23204696.0/4294967296.0,1,-nbitq), 
to_sfixed(-317170888.0/4294967296.0,1,-nbitq), 
to_sfixed(149369692.0/4294967296.0,1,-nbitq), 
to_sfixed(-523310797.0/4294967296.0,1,-nbitq), 
to_sfixed(-36241542.0/4294967296.0,1,-nbitq), 
to_sfixed(225187790.0/4294967296.0,1,-nbitq), 
to_sfixed(443849242.0/4294967296.0,1,-nbitq), 
to_sfixed(298769121.0/4294967296.0,1,-nbitq), 
to_sfixed(-491910996.0/4294967296.0,1,-nbitq), 
to_sfixed(291013636.0/4294967296.0,1,-nbitq), 
to_sfixed(230218200.0/4294967296.0,1,-nbitq), 
to_sfixed(-81684098.0/4294967296.0,1,-nbitq), 
to_sfixed(30178392.0/4294967296.0,1,-nbitq), 
to_sfixed(3257464.0/4294967296.0,1,-nbitq), 
to_sfixed(-1973943994.0/4294967296.0,1,-nbitq), 
to_sfixed(-404709756.0/4294967296.0,1,-nbitq), 
to_sfixed(640330528.0/4294967296.0,1,-nbitq), 
to_sfixed(-482907575.0/4294967296.0,1,-nbitq), 
to_sfixed(201567623.0/4294967296.0,1,-nbitq), 
to_sfixed(-64043986.0/4294967296.0,1,-nbitq), 
to_sfixed(595113295.0/4294967296.0,1,-nbitq), 
to_sfixed(251415585.0/4294967296.0,1,-nbitq), 
to_sfixed(299806969.0/4294967296.0,1,-nbitq), 
to_sfixed(-475945014.0/4294967296.0,1,-nbitq), 
to_sfixed(396812005.0/4294967296.0,1,-nbitq), 
to_sfixed(-371782167.0/4294967296.0,1,-nbitq), 
to_sfixed(736145464.0/4294967296.0,1,-nbitq), 
to_sfixed(319419759.0/4294967296.0,1,-nbitq), 
to_sfixed(1346833460.0/4294967296.0,1,-nbitq), 
to_sfixed(-130420043.0/4294967296.0,1,-nbitq), 
to_sfixed(-316170302.0/4294967296.0,1,-nbitq), 
to_sfixed(-268948862.0/4294967296.0,1,-nbitq), 
to_sfixed(-591799155.0/4294967296.0,1,-nbitq), 
to_sfixed(247395495.0/4294967296.0,1,-nbitq), 
to_sfixed(-469850160.0/4294967296.0,1,-nbitq), 
to_sfixed(-42075924.0/4294967296.0,1,-nbitq), 
to_sfixed(842938127.0/4294967296.0,1,-nbitq), 
to_sfixed(-86861310.0/4294967296.0,1,-nbitq), 
to_sfixed(-80686892.0/4294967296.0,1,-nbitq), 
to_sfixed(370450490.0/4294967296.0,1,-nbitq), 
to_sfixed(-955585754.0/4294967296.0,1,-nbitq), 
to_sfixed(19658504.0/4294967296.0,1,-nbitq), 
to_sfixed(594207152.0/4294967296.0,1,-nbitq), 
to_sfixed(493371017.0/4294967296.0,1,-nbitq), 
to_sfixed(247690302.0/4294967296.0,1,-nbitq), 
to_sfixed(-194428824.0/4294967296.0,1,-nbitq), 
to_sfixed(-405007923.0/4294967296.0,1,-nbitq), 
to_sfixed(1095354297.0/4294967296.0,1,-nbitq), 
to_sfixed(-127175059.0/4294967296.0,1,-nbitq), 
to_sfixed(-159496451.0/4294967296.0,1,-nbitq), 
to_sfixed(-206072148.0/4294967296.0,1,-nbitq), 
to_sfixed(-525081896.0/4294967296.0,1,-nbitq), 
to_sfixed(36896587.0/4294967296.0,1,-nbitq), 
to_sfixed(219388245.0/4294967296.0,1,-nbitq), 
to_sfixed(-817524842.0/4294967296.0,1,-nbitq), 
to_sfixed(664662708.0/4294967296.0,1,-nbitq), 
to_sfixed(10136907.0/4294967296.0,1,-nbitq), 
to_sfixed(-222391927.0/4294967296.0,1,-nbitq), 
to_sfixed(73588223.0/4294967296.0,1,-nbitq), 
to_sfixed(41346697.0/4294967296.0,1,-nbitq), 
to_sfixed(156317502.0/4294967296.0,1,-nbitq), 
to_sfixed(926327475.0/4294967296.0,1,-nbitq), 
to_sfixed(-291350591.0/4294967296.0,1,-nbitq), 
to_sfixed(437148977.0/4294967296.0,1,-nbitq), 
to_sfixed(218054346.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(4325005.0/4294967296.0,1,-nbitq), 
to_sfixed(590269614.0/4294967296.0,1,-nbitq), 
to_sfixed(147775047.0/4294967296.0,1,-nbitq), 
to_sfixed(251752053.0/4294967296.0,1,-nbitq), 
to_sfixed(-757430076.0/4294967296.0,1,-nbitq), 
to_sfixed(-667351455.0/4294967296.0,1,-nbitq), 
to_sfixed(-517309607.0/4294967296.0,1,-nbitq), 
to_sfixed(-534575588.0/4294967296.0,1,-nbitq), 
to_sfixed(529787580.0/4294967296.0,1,-nbitq), 
to_sfixed(-290285290.0/4294967296.0,1,-nbitq), 
to_sfixed(-418469360.0/4294967296.0,1,-nbitq), 
to_sfixed(-385903951.0/4294967296.0,1,-nbitq), 
to_sfixed(-783499937.0/4294967296.0,1,-nbitq), 
to_sfixed(481214842.0/4294967296.0,1,-nbitq), 
to_sfixed(-53697658.0/4294967296.0,1,-nbitq), 
to_sfixed(-599858199.0/4294967296.0,1,-nbitq), 
to_sfixed(-332793528.0/4294967296.0,1,-nbitq), 
to_sfixed(188831951.0/4294967296.0,1,-nbitq), 
to_sfixed(-453405687.0/4294967296.0,1,-nbitq), 
to_sfixed(338647432.0/4294967296.0,1,-nbitq), 
to_sfixed(158777702.0/4294967296.0,1,-nbitq), 
to_sfixed(23835216.0/4294967296.0,1,-nbitq), 
to_sfixed(-140939213.0/4294967296.0,1,-nbitq), 
to_sfixed(-676494455.0/4294967296.0,1,-nbitq), 
to_sfixed(-5956755.0/4294967296.0,1,-nbitq), 
to_sfixed(-41798707.0/4294967296.0,1,-nbitq), 
to_sfixed(600515459.0/4294967296.0,1,-nbitq), 
to_sfixed(-327864818.0/4294967296.0,1,-nbitq), 
to_sfixed(756975376.0/4294967296.0,1,-nbitq), 
to_sfixed(-701755239.0/4294967296.0,1,-nbitq), 
to_sfixed(-405879100.0/4294967296.0,1,-nbitq), 
to_sfixed(602157163.0/4294967296.0,1,-nbitq), 
to_sfixed(-125172221.0/4294967296.0,1,-nbitq), 
to_sfixed(-148820902.0/4294967296.0,1,-nbitq), 
to_sfixed(220751372.0/4294967296.0,1,-nbitq), 
to_sfixed(312686606.0/4294967296.0,1,-nbitq), 
to_sfixed(447447452.0/4294967296.0,1,-nbitq), 
to_sfixed(395031787.0/4294967296.0,1,-nbitq), 
to_sfixed(-412775998.0/4294967296.0,1,-nbitq), 
to_sfixed(217329468.0/4294967296.0,1,-nbitq), 
to_sfixed(-112780255.0/4294967296.0,1,-nbitq), 
to_sfixed(538301135.0/4294967296.0,1,-nbitq), 
to_sfixed(555484484.0/4294967296.0,1,-nbitq), 
to_sfixed(387762467.0/4294967296.0,1,-nbitq), 
to_sfixed(80440168.0/4294967296.0,1,-nbitq), 
to_sfixed(248841394.0/4294967296.0,1,-nbitq), 
to_sfixed(62972439.0/4294967296.0,1,-nbitq), 
to_sfixed(-684979480.0/4294967296.0,1,-nbitq), 
to_sfixed(-176333497.0/4294967296.0,1,-nbitq), 
to_sfixed(773363995.0/4294967296.0,1,-nbitq), 
to_sfixed(-359550645.0/4294967296.0,1,-nbitq), 
to_sfixed(288643212.0/4294967296.0,1,-nbitq), 
to_sfixed(156477071.0/4294967296.0,1,-nbitq), 
to_sfixed(-729378209.0/4294967296.0,1,-nbitq), 
to_sfixed(621389693.0/4294967296.0,1,-nbitq), 
to_sfixed(-395745493.0/4294967296.0,1,-nbitq), 
to_sfixed(-44692676.0/4294967296.0,1,-nbitq), 
to_sfixed(186365036.0/4294967296.0,1,-nbitq), 
to_sfixed(-58219253.0/4294967296.0,1,-nbitq), 
to_sfixed(392657172.0/4294967296.0,1,-nbitq), 
to_sfixed(210231467.0/4294967296.0,1,-nbitq), 
to_sfixed(291825922.0/4294967296.0,1,-nbitq), 
to_sfixed(445998684.0/4294967296.0,1,-nbitq), 
to_sfixed(193032040.0/4294967296.0,1,-nbitq), 
to_sfixed(28876531.0/4294967296.0,1,-nbitq), 
to_sfixed(-358610441.0/4294967296.0,1,-nbitq), 
to_sfixed(-575425505.0/4294967296.0,1,-nbitq), 
to_sfixed(357367449.0/4294967296.0,1,-nbitq), 
to_sfixed(214658362.0/4294967296.0,1,-nbitq), 
to_sfixed(-356328300.0/4294967296.0,1,-nbitq), 
to_sfixed(87809743.0/4294967296.0,1,-nbitq), 
to_sfixed(98058264.0/4294967296.0,1,-nbitq), 
to_sfixed(-4287578.0/4294967296.0,1,-nbitq), 
to_sfixed(-158366723.0/4294967296.0,1,-nbitq), 
to_sfixed(271872255.0/4294967296.0,1,-nbitq), 
to_sfixed(-567448815.0/4294967296.0,1,-nbitq), 
to_sfixed(709525172.0/4294967296.0,1,-nbitq), 
to_sfixed(-139670481.0/4294967296.0,1,-nbitq), 
to_sfixed(-79401303.0/4294967296.0,1,-nbitq), 
to_sfixed(-18969028.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-205179218.0/4294967296.0,1,-nbitq), 
to_sfixed(517273723.0/4294967296.0,1,-nbitq), 
to_sfixed(-406812204.0/4294967296.0,1,-nbitq), 
to_sfixed(-116946309.0/4294967296.0,1,-nbitq), 
to_sfixed(-10125609.0/4294967296.0,1,-nbitq), 
to_sfixed(-346517269.0/4294967296.0,1,-nbitq), 
to_sfixed(279139964.0/4294967296.0,1,-nbitq), 
to_sfixed(-134792966.0/4294967296.0,1,-nbitq), 
to_sfixed(387245762.0/4294967296.0,1,-nbitq), 
to_sfixed(-217607704.0/4294967296.0,1,-nbitq), 
to_sfixed(-188681528.0/4294967296.0,1,-nbitq), 
to_sfixed(-387524521.0/4294967296.0,1,-nbitq), 
to_sfixed(-887439.0/4294967296.0,1,-nbitq), 
to_sfixed(-98452070.0/4294967296.0,1,-nbitq), 
to_sfixed(140849455.0/4294967296.0,1,-nbitq), 
to_sfixed(-768802367.0/4294967296.0,1,-nbitq), 
to_sfixed(20800716.0/4294967296.0,1,-nbitq), 
to_sfixed(-101285930.0/4294967296.0,1,-nbitq), 
to_sfixed(-7530210.0/4294967296.0,1,-nbitq), 
to_sfixed(-69177893.0/4294967296.0,1,-nbitq), 
to_sfixed(-83495727.0/4294967296.0,1,-nbitq), 
to_sfixed(319887500.0/4294967296.0,1,-nbitq), 
to_sfixed(-10312196.0/4294967296.0,1,-nbitq), 
to_sfixed(44035249.0/4294967296.0,1,-nbitq), 
to_sfixed(399671005.0/4294967296.0,1,-nbitq), 
to_sfixed(633629198.0/4294967296.0,1,-nbitq), 
to_sfixed(55945272.0/4294967296.0,1,-nbitq), 
to_sfixed(-685654171.0/4294967296.0,1,-nbitq), 
to_sfixed(230468161.0/4294967296.0,1,-nbitq), 
to_sfixed(-858267843.0/4294967296.0,1,-nbitq), 
to_sfixed(195280979.0/4294967296.0,1,-nbitq), 
to_sfixed(693240910.0/4294967296.0,1,-nbitq), 
to_sfixed(64459365.0/4294967296.0,1,-nbitq), 
to_sfixed(29301071.0/4294967296.0,1,-nbitq), 
to_sfixed(-23137923.0/4294967296.0,1,-nbitq), 
to_sfixed(660680859.0/4294967296.0,1,-nbitq), 
to_sfixed(445117348.0/4294967296.0,1,-nbitq), 
to_sfixed(349225062.0/4294967296.0,1,-nbitq), 
to_sfixed(259827553.0/4294967296.0,1,-nbitq), 
to_sfixed(105759743.0/4294967296.0,1,-nbitq), 
to_sfixed(113772614.0/4294967296.0,1,-nbitq), 
to_sfixed(813898762.0/4294967296.0,1,-nbitq), 
to_sfixed(268344340.0/4294967296.0,1,-nbitq), 
to_sfixed(699566994.0/4294967296.0,1,-nbitq), 
to_sfixed(-494833795.0/4294967296.0,1,-nbitq), 
to_sfixed(-387511835.0/4294967296.0,1,-nbitq), 
to_sfixed(-374873896.0/4294967296.0,1,-nbitq), 
to_sfixed(-1196576047.0/4294967296.0,1,-nbitq), 
to_sfixed(-213489675.0/4294967296.0,1,-nbitq), 
to_sfixed(300624229.0/4294967296.0,1,-nbitq), 
to_sfixed(169327035.0/4294967296.0,1,-nbitq), 
to_sfixed(171620580.0/4294967296.0,1,-nbitq), 
to_sfixed(289671913.0/4294967296.0,1,-nbitq), 
to_sfixed(-26783915.0/4294967296.0,1,-nbitq), 
to_sfixed(214817121.0/4294967296.0,1,-nbitq), 
to_sfixed(-453296995.0/4294967296.0,1,-nbitq), 
to_sfixed(147019489.0/4294967296.0,1,-nbitq), 
to_sfixed(506108493.0/4294967296.0,1,-nbitq), 
to_sfixed(-264674831.0/4294967296.0,1,-nbitq), 
to_sfixed(-37014886.0/4294967296.0,1,-nbitq), 
to_sfixed(-255626790.0/4294967296.0,1,-nbitq), 
to_sfixed(-273721865.0/4294967296.0,1,-nbitq), 
to_sfixed(262892025.0/4294967296.0,1,-nbitq), 
to_sfixed(531477397.0/4294967296.0,1,-nbitq), 
to_sfixed(61462035.0/4294967296.0,1,-nbitq), 
to_sfixed(355038301.0/4294967296.0,1,-nbitq), 
to_sfixed(-170000306.0/4294967296.0,1,-nbitq), 
to_sfixed(-632781971.0/4294967296.0,1,-nbitq), 
to_sfixed(141880437.0/4294967296.0,1,-nbitq), 
to_sfixed(-390236270.0/4294967296.0,1,-nbitq), 
to_sfixed(523236530.0/4294967296.0,1,-nbitq), 
to_sfixed(108401805.0/4294967296.0,1,-nbitq), 
to_sfixed(218000218.0/4294967296.0,1,-nbitq), 
to_sfixed(408516266.0/4294967296.0,1,-nbitq), 
to_sfixed(189533099.0/4294967296.0,1,-nbitq), 
to_sfixed(-112167174.0/4294967296.0,1,-nbitq), 
to_sfixed(572458172.0/4294967296.0,1,-nbitq), 
to_sfixed(-195276553.0/4294967296.0,1,-nbitq), 
to_sfixed(-672199513.0/4294967296.0,1,-nbitq), 
to_sfixed(-62498579.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-114193575.0/4294967296.0,1,-nbitq), 
to_sfixed(544342309.0/4294967296.0,1,-nbitq), 
to_sfixed(-30531762.0/4294967296.0,1,-nbitq), 
to_sfixed(-434321922.0/4294967296.0,1,-nbitq), 
to_sfixed(614411982.0/4294967296.0,1,-nbitq), 
to_sfixed(233875016.0/4294967296.0,1,-nbitq), 
to_sfixed(-410337428.0/4294967296.0,1,-nbitq), 
to_sfixed(401992403.0/4294967296.0,1,-nbitq), 
to_sfixed(903570952.0/4294967296.0,1,-nbitq), 
to_sfixed(-159992461.0/4294967296.0,1,-nbitq), 
to_sfixed(5824514.0/4294967296.0,1,-nbitq), 
to_sfixed(-529068990.0/4294967296.0,1,-nbitq), 
to_sfixed(363263589.0/4294967296.0,1,-nbitq), 
to_sfixed(-71066641.0/4294967296.0,1,-nbitq), 
to_sfixed(-258663355.0/4294967296.0,1,-nbitq), 
to_sfixed(-601415529.0/4294967296.0,1,-nbitq), 
to_sfixed(-328511343.0/4294967296.0,1,-nbitq), 
to_sfixed(134208618.0/4294967296.0,1,-nbitq), 
to_sfixed(-187828868.0/4294967296.0,1,-nbitq), 
to_sfixed(103516717.0/4294967296.0,1,-nbitq), 
to_sfixed(60911347.0/4294967296.0,1,-nbitq), 
to_sfixed(-371381670.0/4294967296.0,1,-nbitq), 
to_sfixed(373875870.0/4294967296.0,1,-nbitq), 
to_sfixed(381848973.0/4294967296.0,1,-nbitq), 
to_sfixed(-144768807.0/4294967296.0,1,-nbitq), 
to_sfixed(725352572.0/4294967296.0,1,-nbitq), 
to_sfixed(-486822813.0/4294967296.0,1,-nbitq), 
to_sfixed(211624063.0/4294967296.0,1,-nbitq), 
to_sfixed(615399430.0/4294967296.0,1,-nbitq), 
to_sfixed(-872413208.0/4294967296.0,1,-nbitq), 
to_sfixed(163375575.0/4294967296.0,1,-nbitq), 
to_sfixed(-38465810.0/4294967296.0,1,-nbitq), 
to_sfixed(147664905.0/4294967296.0,1,-nbitq), 
to_sfixed(-792055148.0/4294967296.0,1,-nbitq), 
to_sfixed(427134713.0/4294967296.0,1,-nbitq), 
to_sfixed(102576875.0/4294967296.0,1,-nbitq), 
to_sfixed(156972848.0/4294967296.0,1,-nbitq), 
to_sfixed(396494758.0/4294967296.0,1,-nbitq), 
to_sfixed(415265705.0/4294967296.0,1,-nbitq), 
to_sfixed(-46198864.0/4294967296.0,1,-nbitq), 
to_sfixed(499657244.0/4294967296.0,1,-nbitq), 
to_sfixed(-274272211.0/4294967296.0,1,-nbitq), 
to_sfixed(589857862.0/4294967296.0,1,-nbitq), 
to_sfixed(105297440.0/4294967296.0,1,-nbitq), 
to_sfixed(-130092075.0/4294967296.0,1,-nbitq), 
to_sfixed(247013813.0/4294967296.0,1,-nbitq), 
to_sfixed(-429616691.0/4294967296.0,1,-nbitq), 
to_sfixed(-650763367.0/4294967296.0,1,-nbitq), 
to_sfixed(-254563082.0/4294967296.0,1,-nbitq), 
to_sfixed(302520038.0/4294967296.0,1,-nbitq), 
to_sfixed(-47170207.0/4294967296.0,1,-nbitq), 
to_sfixed(-530110814.0/4294967296.0,1,-nbitq), 
to_sfixed(270194711.0/4294967296.0,1,-nbitq), 
to_sfixed(-441137164.0/4294967296.0,1,-nbitq), 
to_sfixed(225416341.0/4294967296.0,1,-nbitq), 
to_sfixed(173986800.0/4294967296.0,1,-nbitq), 
to_sfixed(322678239.0/4294967296.0,1,-nbitq), 
to_sfixed(-269651767.0/4294967296.0,1,-nbitq), 
to_sfixed(-209286368.0/4294967296.0,1,-nbitq), 
to_sfixed(357397494.0/4294967296.0,1,-nbitq), 
to_sfixed(174343756.0/4294967296.0,1,-nbitq), 
to_sfixed(89568089.0/4294967296.0,1,-nbitq), 
to_sfixed(528109245.0/4294967296.0,1,-nbitq), 
to_sfixed(10077184.0/4294967296.0,1,-nbitq), 
to_sfixed(-224893791.0/4294967296.0,1,-nbitq), 
to_sfixed(-253146453.0/4294967296.0,1,-nbitq), 
to_sfixed(231294676.0/4294967296.0,1,-nbitq), 
to_sfixed(-74633726.0/4294967296.0,1,-nbitq), 
to_sfixed(385581270.0/4294967296.0,1,-nbitq), 
to_sfixed(-333081958.0/4294967296.0,1,-nbitq), 
to_sfixed(1128924743.0/4294967296.0,1,-nbitq), 
to_sfixed(-121803935.0/4294967296.0,1,-nbitq), 
to_sfixed(-559502626.0/4294967296.0,1,-nbitq), 
to_sfixed(-345721528.0/4294967296.0,1,-nbitq), 
to_sfixed(486986584.0/4294967296.0,1,-nbitq), 
to_sfixed(108447440.0/4294967296.0,1,-nbitq), 
to_sfixed(-14177672.0/4294967296.0,1,-nbitq), 
to_sfixed(263393583.0/4294967296.0,1,-nbitq), 
to_sfixed(-505872523.0/4294967296.0,1,-nbitq), 
to_sfixed(216438862.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(329252102.0/4294967296.0,1,-nbitq), 
to_sfixed(330085922.0/4294967296.0,1,-nbitq), 
to_sfixed(-215941362.0/4294967296.0,1,-nbitq), 
to_sfixed(499788421.0/4294967296.0,1,-nbitq), 
to_sfixed(1007262643.0/4294967296.0,1,-nbitq), 
to_sfixed(88084342.0/4294967296.0,1,-nbitq), 
to_sfixed(279485668.0/4294967296.0,1,-nbitq), 
to_sfixed(-100323004.0/4294967296.0,1,-nbitq), 
to_sfixed(746383874.0/4294967296.0,1,-nbitq), 
to_sfixed(-33279053.0/4294967296.0,1,-nbitq), 
to_sfixed(411003810.0/4294967296.0,1,-nbitq), 
to_sfixed(-128145947.0/4294967296.0,1,-nbitq), 
to_sfixed(1056271636.0/4294967296.0,1,-nbitq), 
to_sfixed(-135252816.0/4294967296.0,1,-nbitq), 
to_sfixed(-203207613.0/4294967296.0,1,-nbitq), 
to_sfixed(-524403162.0/4294967296.0,1,-nbitq), 
to_sfixed(328865254.0/4294967296.0,1,-nbitq), 
to_sfixed(-105084399.0/4294967296.0,1,-nbitq), 
to_sfixed(-76206014.0/4294967296.0,1,-nbitq), 
to_sfixed(121062985.0/4294967296.0,1,-nbitq), 
to_sfixed(-95348590.0/4294967296.0,1,-nbitq), 
to_sfixed(240496085.0/4294967296.0,1,-nbitq), 
to_sfixed(-252569174.0/4294967296.0,1,-nbitq), 
to_sfixed(-30078173.0/4294967296.0,1,-nbitq), 
to_sfixed(-9478283.0/4294967296.0,1,-nbitq), 
to_sfixed(584370477.0/4294967296.0,1,-nbitq), 
to_sfixed(-366655915.0/4294967296.0,1,-nbitq), 
to_sfixed(-334744497.0/4294967296.0,1,-nbitq), 
to_sfixed(107307983.0/4294967296.0,1,-nbitq), 
to_sfixed(-528553483.0/4294967296.0,1,-nbitq), 
to_sfixed(118078382.0/4294967296.0,1,-nbitq), 
to_sfixed(155068571.0/4294967296.0,1,-nbitq), 
to_sfixed(503154052.0/4294967296.0,1,-nbitq), 
to_sfixed(-403152509.0/4294967296.0,1,-nbitq), 
to_sfixed(-191027199.0/4294967296.0,1,-nbitq), 
to_sfixed(-13727921.0/4294967296.0,1,-nbitq), 
to_sfixed(-20804583.0/4294967296.0,1,-nbitq), 
to_sfixed(-113032605.0/4294967296.0,1,-nbitq), 
to_sfixed(-102387635.0/4294967296.0,1,-nbitq), 
to_sfixed(263836923.0/4294967296.0,1,-nbitq), 
to_sfixed(668456752.0/4294967296.0,1,-nbitq), 
to_sfixed(330659800.0/4294967296.0,1,-nbitq), 
to_sfixed(379033680.0/4294967296.0,1,-nbitq), 
to_sfixed(-200837229.0/4294967296.0,1,-nbitq), 
to_sfixed(-200399494.0/4294967296.0,1,-nbitq), 
to_sfixed(187332539.0/4294967296.0,1,-nbitq), 
to_sfixed(-319766574.0/4294967296.0,1,-nbitq), 
to_sfixed(-27329096.0/4294967296.0,1,-nbitq), 
to_sfixed(197284385.0/4294967296.0,1,-nbitq), 
to_sfixed(115842264.0/4294967296.0,1,-nbitq), 
to_sfixed(152414468.0/4294967296.0,1,-nbitq), 
to_sfixed(-774680613.0/4294967296.0,1,-nbitq), 
to_sfixed(26621487.0/4294967296.0,1,-nbitq), 
to_sfixed(-193229056.0/4294967296.0,1,-nbitq), 
to_sfixed(-125334774.0/4294967296.0,1,-nbitq), 
to_sfixed(-178951600.0/4294967296.0,1,-nbitq), 
to_sfixed(355521839.0/4294967296.0,1,-nbitq), 
to_sfixed(-514359678.0/4294967296.0,1,-nbitq), 
to_sfixed(250164354.0/4294967296.0,1,-nbitq), 
to_sfixed(-95663787.0/4294967296.0,1,-nbitq), 
to_sfixed(-400989111.0/4294967296.0,1,-nbitq), 
to_sfixed(-741586885.0/4294967296.0,1,-nbitq), 
to_sfixed(506539362.0/4294967296.0,1,-nbitq), 
to_sfixed(-477220910.0/4294967296.0,1,-nbitq), 
to_sfixed(261714902.0/4294967296.0,1,-nbitq), 
to_sfixed(-340895373.0/4294967296.0,1,-nbitq), 
to_sfixed(-290362973.0/4294967296.0,1,-nbitq), 
to_sfixed(-113087128.0/4294967296.0,1,-nbitq), 
to_sfixed(108835633.0/4294967296.0,1,-nbitq), 
to_sfixed(502530537.0/4294967296.0,1,-nbitq), 
to_sfixed(1328440904.0/4294967296.0,1,-nbitq), 
to_sfixed(-203187579.0/4294967296.0,1,-nbitq), 
to_sfixed(-160522324.0/4294967296.0,1,-nbitq), 
to_sfixed(246996955.0/4294967296.0,1,-nbitq), 
to_sfixed(-43193977.0/4294967296.0,1,-nbitq), 
to_sfixed(-399993703.0/4294967296.0,1,-nbitq), 
to_sfixed(-164277154.0/4294967296.0,1,-nbitq), 
to_sfixed(139943243.0/4294967296.0,1,-nbitq), 
to_sfixed(-317408450.0/4294967296.0,1,-nbitq), 
to_sfixed(-392856938.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(39352021.0/4294967296.0,1,-nbitq), 
to_sfixed(624637704.0/4294967296.0,1,-nbitq), 
to_sfixed(717438.0/4294967296.0,1,-nbitq), 
to_sfixed(432624476.0/4294967296.0,1,-nbitq), 
to_sfixed(641267901.0/4294967296.0,1,-nbitq), 
to_sfixed(79446517.0/4294967296.0,1,-nbitq), 
to_sfixed(-468892488.0/4294967296.0,1,-nbitq), 
to_sfixed(18550523.0/4294967296.0,1,-nbitq), 
to_sfixed(203839455.0/4294967296.0,1,-nbitq), 
to_sfixed(140034398.0/4294967296.0,1,-nbitq), 
to_sfixed(-150843974.0/4294967296.0,1,-nbitq), 
to_sfixed(179384939.0/4294967296.0,1,-nbitq), 
to_sfixed(585293182.0/4294967296.0,1,-nbitq), 
to_sfixed(-681246887.0/4294967296.0,1,-nbitq), 
to_sfixed(318846169.0/4294967296.0,1,-nbitq), 
to_sfixed(-589852920.0/4294967296.0,1,-nbitq), 
to_sfixed(374273232.0/4294967296.0,1,-nbitq), 
to_sfixed(-205908720.0/4294967296.0,1,-nbitq), 
to_sfixed(343635122.0/4294967296.0,1,-nbitq), 
to_sfixed(-38670584.0/4294967296.0,1,-nbitq), 
to_sfixed(-350413400.0/4294967296.0,1,-nbitq), 
to_sfixed(267803629.0/4294967296.0,1,-nbitq), 
to_sfixed(-115903649.0/4294967296.0,1,-nbitq), 
to_sfixed(-424008355.0/4294967296.0,1,-nbitq), 
to_sfixed(314278870.0/4294967296.0,1,-nbitq), 
to_sfixed(481008643.0/4294967296.0,1,-nbitq), 
to_sfixed(-324154451.0/4294967296.0,1,-nbitq), 
to_sfixed(227391246.0/4294967296.0,1,-nbitq), 
to_sfixed(89603559.0/4294967296.0,1,-nbitq), 
to_sfixed(-527324048.0/4294967296.0,1,-nbitq), 
to_sfixed(232169388.0/4294967296.0,1,-nbitq), 
to_sfixed(273856693.0/4294967296.0,1,-nbitq), 
to_sfixed(-53045007.0/4294967296.0,1,-nbitq), 
to_sfixed(317430561.0/4294967296.0,1,-nbitq), 
to_sfixed(35115877.0/4294967296.0,1,-nbitq), 
to_sfixed(257456900.0/4294967296.0,1,-nbitq), 
to_sfixed(-282234903.0/4294967296.0,1,-nbitq), 
to_sfixed(-886304076.0/4294967296.0,1,-nbitq), 
to_sfixed(318605334.0/4294967296.0,1,-nbitq), 
to_sfixed(300792931.0/4294967296.0,1,-nbitq), 
to_sfixed(147537653.0/4294967296.0,1,-nbitq), 
to_sfixed(218753883.0/4294967296.0,1,-nbitq), 
to_sfixed(-223562454.0/4294967296.0,1,-nbitq), 
to_sfixed(-157730860.0/4294967296.0,1,-nbitq), 
to_sfixed(91003223.0/4294967296.0,1,-nbitq), 
to_sfixed(30552948.0/4294967296.0,1,-nbitq), 
to_sfixed(-422221865.0/4294967296.0,1,-nbitq), 
to_sfixed(-5029714.0/4294967296.0,1,-nbitq), 
to_sfixed(-504856349.0/4294967296.0,1,-nbitq), 
to_sfixed(-64362282.0/4294967296.0,1,-nbitq), 
to_sfixed(151516244.0/4294967296.0,1,-nbitq), 
to_sfixed(101639910.0/4294967296.0,1,-nbitq), 
to_sfixed(157463777.0/4294967296.0,1,-nbitq), 
to_sfixed(171091363.0/4294967296.0,1,-nbitq), 
to_sfixed(-228784708.0/4294967296.0,1,-nbitq), 
to_sfixed(69542690.0/4294967296.0,1,-nbitq), 
to_sfixed(-499395039.0/4294967296.0,1,-nbitq), 
to_sfixed(-503293332.0/4294967296.0,1,-nbitq), 
to_sfixed(130176917.0/4294967296.0,1,-nbitq), 
to_sfixed(45448684.0/4294967296.0,1,-nbitq), 
to_sfixed(-358829979.0/4294967296.0,1,-nbitq), 
to_sfixed(-325691796.0/4294967296.0,1,-nbitq), 
to_sfixed(422602250.0/4294967296.0,1,-nbitq), 
to_sfixed(16939790.0/4294967296.0,1,-nbitq), 
to_sfixed(-226919189.0/4294967296.0,1,-nbitq), 
to_sfixed(177430777.0/4294967296.0,1,-nbitq), 
to_sfixed(-334735770.0/4294967296.0,1,-nbitq), 
to_sfixed(-333724978.0/4294967296.0,1,-nbitq), 
to_sfixed(-49535345.0/4294967296.0,1,-nbitq), 
to_sfixed(65515661.0/4294967296.0,1,-nbitq), 
to_sfixed(461936151.0/4294967296.0,1,-nbitq), 
to_sfixed(392994119.0/4294967296.0,1,-nbitq), 
to_sfixed(12615337.0/4294967296.0,1,-nbitq), 
to_sfixed(-165589125.0/4294967296.0,1,-nbitq), 
to_sfixed(227950018.0/4294967296.0,1,-nbitq), 
to_sfixed(56086227.0/4294967296.0,1,-nbitq), 
to_sfixed(127779796.0/4294967296.0,1,-nbitq), 
to_sfixed(-318124572.0/4294967296.0,1,-nbitq), 
to_sfixed(12314755.0/4294967296.0,1,-nbitq), 
to_sfixed(-147205709.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-114077195.0/4294967296.0,1,-nbitq), 
to_sfixed(293278707.0/4294967296.0,1,-nbitq), 
to_sfixed(-341726958.0/4294967296.0,1,-nbitq), 
to_sfixed(235170893.0/4294967296.0,1,-nbitq), 
to_sfixed(126570383.0/4294967296.0,1,-nbitq), 
to_sfixed(-285175706.0/4294967296.0,1,-nbitq), 
to_sfixed(-32209944.0/4294967296.0,1,-nbitq), 
to_sfixed(-342598799.0/4294967296.0,1,-nbitq), 
to_sfixed(-39980098.0/4294967296.0,1,-nbitq), 
to_sfixed(323109772.0/4294967296.0,1,-nbitq), 
to_sfixed(-43068859.0/4294967296.0,1,-nbitq), 
to_sfixed(246741625.0/4294967296.0,1,-nbitq), 
to_sfixed(823503543.0/4294967296.0,1,-nbitq), 
to_sfixed(-429140803.0/4294967296.0,1,-nbitq), 
to_sfixed(359086419.0/4294967296.0,1,-nbitq), 
to_sfixed(-503955992.0/4294967296.0,1,-nbitq), 
to_sfixed(-83411921.0/4294967296.0,1,-nbitq), 
to_sfixed(-298461.0/4294967296.0,1,-nbitq), 
to_sfixed(103253193.0/4294967296.0,1,-nbitq), 
to_sfixed(139243037.0/4294967296.0,1,-nbitq), 
to_sfixed(-14755864.0/4294967296.0,1,-nbitq), 
to_sfixed(401960036.0/4294967296.0,1,-nbitq), 
to_sfixed(205520413.0/4294967296.0,1,-nbitq), 
to_sfixed(-287768033.0/4294967296.0,1,-nbitq), 
to_sfixed(185719102.0/4294967296.0,1,-nbitq), 
to_sfixed(869891723.0/4294967296.0,1,-nbitq), 
to_sfixed(123404679.0/4294967296.0,1,-nbitq), 
to_sfixed(-463117117.0/4294967296.0,1,-nbitq), 
to_sfixed(51286218.0/4294967296.0,1,-nbitq), 
to_sfixed(-35417712.0/4294967296.0,1,-nbitq), 
to_sfixed(-70622228.0/4294967296.0,1,-nbitq), 
to_sfixed(342501980.0/4294967296.0,1,-nbitq), 
to_sfixed(-184805604.0/4294967296.0,1,-nbitq), 
to_sfixed(-36333697.0/4294967296.0,1,-nbitq), 
to_sfixed(163816756.0/4294967296.0,1,-nbitq), 
to_sfixed(-335982745.0/4294967296.0,1,-nbitq), 
to_sfixed(170389487.0/4294967296.0,1,-nbitq), 
to_sfixed(73867139.0/4294967296.0,1,-nbitq), 
to_sfixed(-173966462.0/4294967296.0,1,-nbitq), 
to_sfixed(-12395471.0/4294967296.0,1,-nbitq), 
to_sfixed(667845317.0/4294967296.0,1,-nbitq), 
to_sfixed(240129714.0/4294967296.0,1,-nbitq), 
to_sfixed(191377787.0/4294967296.0,1,-nbitq), 
to_sfixed(-186952724.0/4294967296.0,1,-nbitq), 
to_sfixed(538510338.0/4294967296.0,1,-nbitq), 
to_sfixed(-93927883.0/4294967296.0,1,-nbitq), 
to_sfixed(262196776.0/4294967296.0,1,-nbitq), 
to_sfixed(-303637337.0/4294967296.0,1,-nbitq), 
to_sfixed(-185397307.0/4294967296.0,1,-nbitq), 
to_sfixed(-252768346.0/4294967296.0,1,-nbitq), 
to_sfixed(-419023490.0/4294967296.0,1,-nbitq), 
to_sfixed(289366484.0/4294967296.0,1,-nbitq), 
to_sfixed(-173375939.0/4294967296.0,1,-nbitq), 
to_sfixed(471691754.0/4294967296.0,1,-nbitq), 
to_sfixed(49089234.0/4294967296.0,1,-nbitq), 
to_sfixed(16206246.0/4294967296.0,1,-nbitq), 
to_sfixed(-382302310.0/4294967296.0,1,-nbitq), 
to_sfixed(259405437.0/4294967296.0,1,-nbitq), 
to_sfixed(112574190.0/4294967296.0,1,-nbitq), 
to_sfixed(141752339.0/4294967296.0,1,-nbitq), 
to_sfixed(-430195707.0/4294967296.0,1,-nbitq), 
to_sfixed(151491114.0/4294967296.0,1,-nbitq), 
to_sfixed(182084720.0/4294967296.0,1,-nbitq), 
to_sfixed(186509008.0/4294967296.0,1,-nbitq), 
to_sfixed(-17420775.0/4294967296.0,1,-nbitq), 
to_sfixed(-390139374.0/4294967296.0,1,-nbitq), 
to_sfixed(291039912.0/4294967296.0,1,-nbitq), 
to_sfixed(332382043.0/4294967296.0,1,-nbitq), 
to_sfixed(-238306709.0/4294967296.0,1,-nbitq), 
to_sfixed(110701177.0/4294967296.0,1,-nbitq), 
to_sfixed(-248764166.0/4294967296.0,1,-nbitq), 
to_sfixed(-125569245.0/4294967296.0,1,-nbitq), 
to_sfixed(-82466520.0/4294967296.0,1,-nbitq), 
to_sfixed(-90634527.0/4294967296.0,1,-nbitq), 
to_sfixed(150326380.0/4294967296.0,1,-nbitq), 
to_sfixed(38468032.0/4294967296.0,1,-nbitq), 
to_sfixed(265846244.0/4294967296.0,1,-nbitq), 
to_sfixed(200204185.0/4294967296.0,1,-nbitq), 
to_sfixed(-207257319.0/4294967296.0,1,-nbitq), 
to_sfixed(-208148398.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(177674771.0/4294967296.0,1,-nbitq), 
to_sfixed(-81195323.0/4294967296.0,1,-nbitq), 
to_sfixed(-132765480.0/4294967296.0,1,-nbitq), 
to_sfixed(255800823.0/4294967296.0,1,-nbitq), 
to_sfixed(-13308467.0/4294967296.0,1,-nbitq), 
to_sfixed(-428144508.0/4294967296.0,1,-nbitq), 
to_sfixed(-363569214.0/4294967296.0,1,-nbitq), 
to_sfixed(41193434.0/4294967296.0,1,-nbitq), 
to_sfixed(161957849.0/4294967296.0,1,-nbitq), 
to_sfixed(126805076.0/4294967296.0,1,-nbitq), 
to_sfixed(128675555.0/4294967296.0,1,-nbitq), 
to_sfixed(111998440.0/4294967296.0,1,-nbitq), 
to_sfixed(-29893449.0/4294967296.0,1,-nbitq), 
to_sfixed(173816915.0/4294967296.0,1,-nbitq), 
to_sfixed(-321159139.0/4294967296.0,1,-nbitq), 
to_sfixed(-409055309.0/4294967296.0,1,-nbitq), 
to_sfixed(-117689868.0/4294967296.0,1,-nbitq), 
to_sfixed(64451400.0/4294967296.0,1,-nbitq), 
to_sfixed(465789608.0/4294967296.0,1,-nbitq), 
to_sfixed(-188431403.0/4294967296.0,1,-nbitq), 
to_sfixed(-159409150.0/4294967296.0,1,-nbitq), 
to_sfixed(464487992.0/4294967296.0,1,-nbitq), 
to_sfixed(5792280.0/4294967296.0,1,-nbitq), 
to_sfixed(-23672429.0/4294967296.0,1,-nbitq), 
to_sfixed(247084845.0/4294967296.0,1,-nbitq), 
to_sfixed(703579423.0/4294967296.0,1,-nbitq), 
to_sfixed(-400566659.0/4294967296.0,1,-nbitq), 
to_sfixed(-549390562.0/4294967296.0,1,-nbitq), 
to_sfixed(227865066.0/4294967296.0,1,-nbitq), 
to_sfixed(66318744.0/4294967296.0,1,-nbitq), 
to_sfixed(-109868004.0/4294967296.0,1,-nbitq), 
to_sfixed(-208093496.0/4294967296.0,1,-nbitq), 
to_sfixed(127450125.0/4294967296.0,1,-nbitq), 
to_sfixed(-19113535.0/4294967296.0,1,-nbitq), 
to_sfixed(-115552958.0/4294967296.0,1,-nbitq), 
to_sfixed(-257589307.0/4294967296.0,1,-nbitq), 
to_sfixed(-215142028.0/4294967296.0,1,-nbitq), 
to_sfixed(-351343320.0/4294967296.0,1,-nbitq), 
to_sfixed(314835327.0/4294967296.0,1,-nbitq), 
to_sfixed(151096824.0/4294967296.0,1,-nbitq), 
to_sfixed(-212832376.0/4294967296.0,1,-nbitq), 
to_sfixed(286589583.0/4294967296.0,1,-nbitq), 
to_sfixed(-119294490.0/4294967296.0,1,-nbitq), 
to_sfixed(-59769187.0/4294967296.0,1,-nbitq), 
to_sfixed(-52060390.0/4294967296.0,1,-nbitq), 
to_sfixed(301688455.0/4294967296.0,1,-nbitq), 
to_sfixed(304818929.0/4294967296.0,1,-nbitq), 
to_sfixed(188883041.0/4294967296.0,1,-nbitq), 
to_sfixed(-143423690.0/4294967296.0,1,-nbitq), 
to_sfixed(-126206937.0/4294967296.0,1,-nbitq), 
to_sfixed(-257526129.0/4294967296.0,1,-nbitq), 
to_sfixed(145698766.0/4294967296.0,1,-nbitq), 
to_sfixed(-223130789.0/4294967296.0,1,-nbitq), 
to_sfixed(-153623217.0/4294967296.0,1,-nbitq), 
to_sfixed(-114021922.0/4294967296.0,1,-nbitq), 
to_sfixed(283801930.0/4294967296.0,1,-nbitq), 
to_sfixed(238841750.0/4294967296.0,1,-nbitq), 
to_sfixed(-136582404.0/4294967296.0,1,-nbitq), 
to_sfixed(-234370423.0/4294967296.0,1,-nbitq), 
to_sfixed(-298005491.0/4294967296.0,1,-nbitq), 
to_sfixed(-27886854.0/4294967296.0,1,-nbitq), 
to_sfixed(124709786.0/4294967296.0,1,-nbitq), 
to_sfixed(-118504709.0/4294967296.0,1,-nbitq), 
to_sfixed(14068293.0/4294967296.0,1,-nbitq), 
to_sfixed(-75821147.0/4294967296.0,1,-nbitq), 
to_sfixed(-283264742.0/4294967296.0,1,-nbitq), 
to_sfixed(660738058.0/4294967296.0,1,-nbitq), 
to_sfixed(-70680979.0/4294967296.0,1,-nbitq), 
to_sfixed(434369484.0/4294967296.0,1,-nbitq), 
to_sfixed(-86508101.0/4294967296.0,1,-nbitq), 
to_sfixed(58719076.0/4294967296.0,1,-nbitq), 
to_sfixed(48743722.0/4294967296.0,1,-nbitq), 
to_sfixed(-250771429.0/4294967296.0,1,-nbitq), 
to_sfixed(-84180521.0/4294967296.0,1,-nbitq), 
to_sfixed(405977633.0/4294967296.0,1,-nbitq), 
to_sfixed(23935555.0/4294967296.0,1,-nbitq), 
to_sfixed(-187979470.0/4294967296.0,1,-nbitq), 
to_sfixed(11224308.0/4294967296.0,1,-nbitq), 
to_sfixed(113740588.0/4294967296.0,1,-nbitq), 
to_sfixed(355856193.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-176201269.0/4294967296.0,1,-nbitq), 
to_sfixed(-279803702.0/4294967296.0,1,-nbitq), 
to_sfixed(124184373.0/4294967296.0,1,-nbitq), 
to_sfixed(-247460709.0/4294967296.0,1,-nbitq), 
to_sfixed(-56520535.0/4294967296.0,1,-nbitq), 
to_sfixed(-224320443.0/4294967296.0,1,-nbitq), 
to_sfixed(162452478.0/4294967296.0,1,-nbitq), 
to_sfixed(-41446712.0/4294967296.0,1,-nbitq), 
to_sfixed(-278285691.0/4294967296.0,1,-nbitq), 
to_sfixed(407988079.0/4294967296.0,1,-nbitq), 
to_sfixed(-381221185.0/4294967296.0,1,-nbitq), 
to_sfixed(74242570.0/4294967296.0,1,-nbitq), 
to_sfixed(-160748372.0/4294967296.0,1,-nbitq), 
to_sfixed(-248974470.0/4294967296.0,1,-nbitq), 
to_sfixed(38933851.0/4294967296.0,1,-nbitq), 
to_sfixed(135879791.0/4294967296.0,1,-nbitq), 
to_sfixed(-47277183.0/4294967296.0,1,-nbitq), 
to_sfixed(316282491.0/4294967296.0,1,-nbitq), 
to_sfixed(606489612.0/4294967296.0,1,-nbitq), 
to_sfixed(276583270.0/4294967296.0,1,-nbitq), 
to_sfixed(-174185181.0/4294967296.0,1,-nbitq), 
to_sfixed(359909225.0/4294967296.0,1,-nbitq), 
to_sfixed(67010328.0/4294967296.0,1,-nbitq), 
to_sfixed(266400680.0/4294967296.0,1,-nbitq), 
to_sfixed(350124159.0/4294967296.0,1,-nbitq), 
to_sfixed(165069010.0/4294967296.0,1,-nbitq), 
to_sfixed(55965941.0/4294967296.0,1,-nbitq), 
to_sfixed(-302562802.0/4294967296.0,1,-nbitq), 
to_sfixed(136226580.0/4294967296.0,1,-nbitq), 
to_sfixed(157448852.0/4294967296.0,1,-nbitq), 
to_sfixed(-508255286.0/4294967296.0,1,-nbitq), 
to_sfixed(-500431511.0/4294967296.0,1,-nbitq), 
to_sfixed(24693467.0/4294967296.0,1,-nbitq), 
to_sfixed(107944894.0/4294967296.0,1,-nbitq), 
to_sfixed(362658118.0/4294967296.0,1,-nbitq), 
to_sfixed(237246877.0/4294967296.0,1,-nbitq), 
to_sfixed(-248239524.0/4294967296.0,1,-nbitq), 
to_sfixed(234640122.0/4294967296.0,1,-nbitq), 
to_sfixed(354927638.0/4294967296.0,1,-nbitq), 
to_sfixed(-257038050.0/4294967296.0,1,-nbitq), 
to_sfixed(12650097.0/4294967296.0,1,-nbitq), 
to_sfixed(-237021924.0/4294967296.0,1,-nbitq), 
to_sfixed(391559042.0/4294967296.0,1,-nbitq), 
to_sfixed(348762941.0/4294967296.0,1,-nbitq), 
to_sfixed(362337449.0/4294967296.0,1,-nbitq), 
to_sfixed(241627449.0/4294967296.0,1,-nbitq), 
to_sfixed(-327072950.0/4294967296.0,1,-nbitq), 
to_sfixed(-401311818.0/4294967296.0,1,-nbitq), 
to_sfixed(154914287.0/4294967296.0,1,-nbitq), 
to_sfixed(528520723.0/4294967296.0,1,-nbitq), 
to_sfixed(-153427315.0/4294967296.0,1,-nbitq), 
to_sfixed(225353197.0/4294967296.0,1,-nbitq), 
to_sfixed(-529778968.0/4294967296.0,1,-nbitq), 
to_sfixed(-293825481.0/4294967296.0,1,-nbitq), 
to_sfixed(40441430.0/4294967296.0,1,-nbitq), 
to_sfixed(239489033.0/4294967296.0,1,-nbitq), 
to_sfixed(-291808939.0/4294967296.0,1,-nbitq), 
to_sfixed(-427201097.0/4294967296.0,1,-nbitq), 
to_sfixed(325091943.0/4294967296.0,1,-nbitq), 
to_sfixed(282764097.0/4294967296.0,1,-nbitq), 
to_sfixed(128596657.0/4294967296.0,1,-nbitq), 
to_sfixed(368408752.0/4294967296.0,1,-nbitq), 
to_sfixed(-376897653.0/4294967296.0,1,-nbitq), 
to_sfixed(245194022.0/4294967296.0,1,-nbitq), 
to_sfixed(-17535786.0/4294967296.0,1,-nbitq), 
to_sfixed(-68910398.0/4294967296.0,1,-nbitq), 
to_sfixed(-20692223.0/4294967296.0,1,-nbitq), 
to_sfixed(344879665.0/4294967296.0,1,-nbitq), 
to_sfixed(-295444322.0/4294967296.0,1,-nbitq), 
to_sfixed(-50164244.0/4294967296.0,1,-nbitq), 
to_sfixed(-330531953.0/4294967296.0,1,-nbitq), 
to_sfixed(-401598140.0/4294967296.0,1,-nbitq), 
to_sfixed(-281212179.0/4294967296.0,1,-nbitq), 
to_sfixed(-136298093.0/4294967296.0,1,-nbitq), 
to_sfixed(-108838977.0/4294967296.0,1,-nbitq), 
to_sfixed(-445093373.0/4294967296.0,1,-nbitq), 
to_sfixed(242483287.0/4294967296.0,1,-nbitq), 
to_sfixed(-350444350.0/4294967296.0,1,-nbitq), 
to_sfixed(-551628400.0/4294967296.0,1,-nbitq), 
to_sfixed(96362069.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(38340767.0/4294967296.0,1,-nbitq), 
to_sfixed(-131619221.0/4294967296.0,1,-nbitq), 
to_sfixed(295241144.0/4294967296.0,1,-nbitq), 
to_sfixed(-152186603.0/4294967296.0,1,-nbitq), 
to_sfixed(470305842.0/4294967296.0,1,-nbitq), 
to_sfixed(-459598497.0/4294967296.0,1,-nbitq), 
to_sfixed(-149000785.0/4294967296.0,1,-nbitq), 
to_sfixed(-77418327.0/4294967296.0,1,-nbitq), 
to_sfixed(261987884.0/4294967296.0,1,-nbitq), 
to_sfixed(-79197843.0/4294967296.0,1,-nbitq), 
to_sfixed(-359424055.0/4294967296.0,1,-nbitq), 
to_sfixed(492860893.0/4294967296.0,1,-nbitq), 
to_sfixed(-277341020.0/4294967296.0,1,-nbitq), 
to_sfixed(-145183654.0/4294967296.0,1,-nbitq), 
to_sfixed(321992950.0/4294967296.0,1,-nbitq), 
to_sfixed(215025790.0/4294967296.0,1,-nbitq), 
to_sfixed(338352509.0/4294967296.0,1,-nbitq), 
to_sfixed(184698683.0/4294967296.0,1,-nbitq), 
to_sfixed(-215691005.0/4294967296.0,1,-nbitq), 
to_sfixed(-322616993.0/4294967296.0,1,-nbitq), 
to_sfixed(-145727751.0/4294967296.0,1,-nbitq), 
to_sfixed(416824756.0/4294967296.0,1,-nbitq), 
to_sfixed(394952029.0/4294967296.0,1,-nbitq), 
to_sfixed(-272159618.0/4294967296.0,1,-nbitq), 
to_sfixed(271996934.0/4294967296.0,1,-nbitq), 
to_sfixed(-126403781.0/4294967296.0,1,-nbitq), 
to_sfixed(-19040518.0/4294967296.0,1,-nbitq), 
to_sfixed(-125228584.0/4294967296.0,1,-nbitq), 
to_sfixed(380639372.0/4294967296.0,1,-nbitq), 
to_sfixed(437040559.0/4294967296.0,1,-nbitq), 
to_sfixed(-14831594.0/4294967296.0,1,-nbitq), 
to_sfixed(-350904002.0/4294967296.0,1,-nbitq), 
to_sfixed(338404048.0/4294967296.0,1,-nbitq), 
to_sfixed(66269085.0/4294967296.0,1,-nbitq), 
to_sfixed(539177947.0/4294967296.0,1,-nbitq), 
to_sfixed(426554863.0/4294967296.0,1,-nbitq), 
to_sfixed(41108106.0/4294967296.0,1,-nbitq), 
to_sfixed(-344421353.0/4294967296.0,1,-nbitq), 
to_sfixed(319580096.0/4294967296.0,1,-nbitq), 
to_sfixed(45142758.0/4294967296.0,1,-nbitq), 
to_sfixed(-413416115.0/4294967296.0,1,-nbitq), 
to_sfixed(255259863.0/4294967296.0,1,-nbitq), 
to_sfixed(-109042664.0/4294967296.0,1,-nbitq), 
to_sfixed(-327968323.0/4294967296.0,1,-nbitq), 
to_sfixed(31094220.0/4294967296.0,1,-nbitq), 
to_sfixed(292871428.0/4294967296.0,1,-nbitq), 
to_sfixed(-364574923.0/4294967296.0,1,-nbitq), 
to_sfixed(134216219.0/4294967296.0,1,-nbitq), 
to_sfixed(146333152.0/4294967296.0,1,-nbitq), 
to_sfixed(-140896949.0/4294967296.0,1,-nbitq), 
to_sfixed(249511273.0/4294967296.0,1,-nbitq), 
to_sfixed(-29758502.0/4294967296.0,1,-nbitq), 
to_sfixed(-49523244.0/4294967296.0,1,-nbitq), 
to_sfixed(319998639.0/4294967296.0,1,-nbitq), 
to_sfixed(-189497119.0/4294967296.0,1,-nbitq), 
to_sfixed(-237530771.0/4294967296.0,1,-nbitq), 
to_sfixed(447407821.0/4294967296.0,1,-nbitq), 
to_sfixed(-380758930.0/4294967296.0,1,-nbitq), 
to_sfixed(179574182.0/4294967296.0,1,-nbitq), 
to_sfixed(-240607384.0/4294967296.0,1,-nbitq), 
to_sfixed(82329984.0/4294967296.0,1,-nbitq), 
to_sfixed(66826575.0/4294967296.0,1,-nbitq), 
to_sfixed(159676520.0/4294967296.0,1,-nbitq), 
to_sfixed(24460121.0/4294967296.0,1,-nbitq), 
to_sfixed(-251577010.0/4294967296.0,1,-nbitq), 
to_sfixed(-174718526.0/4294967296.0,1,-nbitq), 
to_sfixed(483489723.0/4294967296.0,1,-nbitq), 
to_sfixed(76947503.0/4294967296.0,1,-nbitq), 
to_sfixed(-223109315.0/4294967296.0,1,-nbitq), 
to_sfixed(447299333.0/4294967296.0,1,-nbitq), 
to_sfixed(114284831.0/4294967296.0,1,-nbitq), 
to_sfixed(-366069532.0/4294967296.0,1,-nbitq), 
to_sfixed(-356594582.0/4294967296.0,1,-nbitq), 
to_sfixed(191415622.0/4294967296.0,1,-nbitq), 
to_sfixed(-145420430.0/4294967296.0,1,-nbitq), 
to_sfixed(101574002.0/4294967296.0,1,-nbitq), 
to_sfixed(-66529298.0/4294967296.0,1,-nbitq), 
to_sfixed(-270434912.0/4294967296.0,1,-nbitq), 
to_sfixed(18454099.0/4294967296.0,1,-nbitq), 
to_sfixed(162200829.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-290391334.0/4294967296.0,1,-nbitq), 
to_sfixed(230545026.0/4294967296.0,1,-nbitq), 
to_sfixed(372375037.0/4294967296.0,1,-nbitq), 
to_sfixed(-121494490.0/4294967296.0,1,-nbitq), 
to_sfixed(143716268.0/4294967296.0,1,-nbitq), 
to_sfixed(-121848310.0/4294967296.0,1,-nbitq), 
to_sfixed(155463230.0/4294967296.0,1,-nbitq), 
to_sfixed(-257016909.0/4294967296.0,1,-nbitq), 
to_sfixed(69282078.0/4294967296.0,1,-nbitq), 
to_sfixed(280860972.0/4294967296.0,1,-nbitq), 
to_sfixed(-47199972.0/4294967296.0,1,-nbitq), 
to_sfixed(194132728.0/4294967296.0,1,-nbitq), 
to_sfixed(-88221657.0/4294967296.0,1,-nbitq), 
to_sfixed(18821558.0/4294967296.0,1,-nbitq), 
to_sfixed(344669208.0/4294967296.0,1,-nbitq), 
to_sfixed(101166185.0/4294967296.0,1,-nbitq), 
to_sfixed(-162716253.0/4294967296.0,1,-nbitq), 
to_sfixed(-49824505.0/4294967296.0,1,-nbitq), 
to_sfixed(231616770.0/4294967296.0,1,-nbitq), 
to_sfixed(-16510504.0/4294967296.0,1,-nbitq), 
to_sfixed(-359825677.0/4294967296.0,1,-nbitq), 
to_sfixed(135618545.0/4294967296.0,1,-nbitq), 
to_sfixed(21646106.0/4294967296.0,1,-nbitq), 
to_sfixed(110609531.0/4294967296.0,1,-nbitq), 
to_sfixed(-315477021.0/4294967296.0,1,-nbitq), 
to_sfixed(383410552.0/4294967296.0,1,-nbitq), 
to_sfixed(410441970.0/4294967296.0,1,-nbitq), 
to_sfixed(-228194294.0/4294967296.0,1,-nbitq), 
to_sfixed(180766371.0/4294967296.0,1,-nbitq), 
to_sfixed(434075005.0/4294967296.0,1,-nbitq), 
to_sfixed(-26621862.0/4294967296.0,1,-nbitq), 
to_sfixed(-56495106.0/4294967296.0,1,-nbitq), 
to_sfixed(35528789.0/4294967296.0,1,-nbitq), 
to_sfixed(111888038.0/4294967296.0,1,-nbitq), 
to_sfixed(510795775.0/4294967296.0,1,-nbitq), 
to_sfixed(253803245.0/4294967296.0,1,-nbitq), 
to_sfixed(-89589659.0/4294967296.0,1,-nbitq), 
to_sfixed(250689439.0/4294967296.0,1,-nbitq), 
to_sfixed(-318770962.0/4294967296.0,1,-nbitq), 
to_sfixed(267989714.0/4294967296.0,1,-nbitq), 
to_sfixed(-479090439.0/4294967296.0,1,-nbitq), 
to_sfixed(190551488.0/4294967296.0,1,-nbitq), 
to_sfixed(5889129.0/4294967296.0,1,-nbitq), 
to_sfixed(-331407440.0/4294967296.0,1,-nbitq), 
to_sfixed(-210538339.0/4294967296.0,1,-nbitq), 
to_sfixed(407546100.0/4294967296.0,1,-nbitq), 
to_sfixed(-54155111.0/4294967296.0,1,-nbitq), 
to_sfixed(-297266805.0/4294967296.0,1,-nbitq), 
to_sfixed(343819322.0/4294967296.0,1,-nbitq), 
to_sfixed(429703727.0/4294967296.0,1,-nbitq), 
to_sfixed(176777087.0/4294967296.0,1,-nbitq), 
to_sfixed(241358226.0/4294967296.0,1,-nbitq), 
to_sfixed(49496895.0/4294967296.0,1,-nbitq), 
to_sfixed(-268802236.0/4294967296.0,1,-nbitq), 
to_sfixed(-138893237.0/4294967296.0,1,-nbitq), 
to_sfixed(-88467394.0/4294967296.0,1,-nbitq), 
to_sfixed(-310238679.0/4294967296.0,1,-nbitq), 
to_sfixed(-248680355.0/4294967296.0,1,-nbitq), 
to_sfixed(-216656270.0/4294967296.0,1,-nbitq), 
to_sfixed(-52170693.0/4294967296.0,1,-nbitq), 
to_sfixed(353929561.0/4294967296.0,1,-nbitq), 
to_sfixed(-57038214.0/4294967296.0,1,-nbitq), 
to_sfixed(157624512.0/4294967296.0,1,-nbitq), 
to_sfixed(-268118938.0/4294967296.0,1,-nbitq), 
to_sfixed(-198474121.0/4294967296.0,1,-nbitq), 
to_sfixed(-4449325.0/4294967296.0,1,-nbitq), 
to_sfixed(528827501.0/4294967296.0,1,-nbitq), 
to_sfixed(-10061978.0/4294967296.0,1,-nbitq), 
to_sfixed(345079450.0/4294967296.0,1,-nbitq), 
to_sfixed(-5631856.0/4294967296.0,1,-nbitq), 
to_sfixed(277694449.0/4294967296.0,1,-nbitq), 
to_sfixed(242791822.0/4294967296.0,1,-nbitq), 
to_sfixed(-349848202.0/4294967296.0,1,-nbitq), 
to_sfixed(235353127.0/4294967296.0,1,-nbitq), 
to_sfixed(393223845.0/4294967296.0,1,-nbitq), 
to_sfixed(-439400620.0/4294967296.0,1,-nbitq), 
to_sfixed(78809966.0/4294967296.0,1,-nbitq), 
to_sfixed(-11838582.0/4294967296.0,1,-nbitq), 
to_sfixed(-449988106.0/4294967296.0,1,-nbitq), 
to_sfixed(354502134.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-173056746.0/4294967296.0,1,-nbitq), 
to_sfixed(54121310.0/4294967296.0,1,-nbitq), 
to_sfixed(541271512.0/4294967296.0,1,-nbitq), 
to_sfixed(-362147321.0/4294967296.0,1,-nbitq), 
to_sfixed(-150847917.0/4294967296.0,1,-nbitq), 
to_sfixed(-173724932.0/4294967296.0,1,-nbitq), 
to_sfixed(94643635.0/4294967296.0,1,-nbitq), 
to_sfixed(-352035537.0/4294967296.0,1,-nbitq), 
to_sfixed(-74002806.0/4294967296.0,1,-nbitq), 
to_sfixed(-109206085.0/4294967296.0,1,-nbitq), 
to_sfixed(-224602490.0/4294967296.0,1,-nbitq), 
to_sfixed(-67862163.0/4294967296.0,1,-nbitq), 
to_sfixed(-269491485.0/4294967296.0,1,-nbitq), 
to_sfixed(227739847.0/4294967296.0,1,-nbitq), 
to_sfixed(-218788988.0/4294967296.0,1,-nbitq), 
to_sfixed(29117215.0/4294967296.0,1,-nbitq), 
to_sfixed(-207835832.0/4294967296.0,1,-nbitq), 
to_sfixed(-312602924.0/4294967296.0,1,-nbitq), 
to_sfixed(-206855868.0/4294967296.0,1,-nbitq), 
to_sfixed(275816903.0/4294967296.0,1,-nbitq), 
to_sfixed(-319220419.0/4294967296.0,1,-nbitq), 
to_sfixed(-239800106.0/4294967296.0,1,-nbitq), 
to_sfixed(288229234.0/4294967296.0,1,-nbitq), 
to_sfixed(-62828085.0/4294967296.0,1,-nbitq), 
to_sfixed(-274332930.0/4294967296.0,1,-nbitq), 
to_sfixed(-113460983.0/4294967296.0,1,-nbitq), 
to_sfixed(36160939.0/4294967296.0,1,-nbitq), 
to_sfixed(-331802769.0/4294967296.0,1,-nbitq), 
to_sfixed(194982050.0/4294967296.0,1,-nbitq), 
to_sfixed(52850008.0/4294967296.0,1,-nbitq), 
to_sfixed(-2504772.0/4294967296.0,1,-nbitq), 
to_sfixed(-66255669.0/4294967296.0,1,-nbitq), 
to_sfixed(161723952.0/4294967296.0,1,-nbitq), 
to_sfixed(-401958819.0/4294967296.0,1,-nbitq), 
to_sfixed(40060991.0/4294967296.0,1,-nbitq), 
to_sfixed(-214289227.0/4294967296.0,1,-nbitq), 
to_sfixed(147552448.0/4294967296.0,1,-nbitq), 
to_sfixed(-91331774.0/4294967296.0,1,-nbitq), 
to_sfixed(279879382.0/4294967296.0,1,-nbitq), 
to_sfixed(-27038540.0/4294967296.0,1,-nbitq), 
to_sfixed(245040185.0/4294967296.0,1,-nbitq), 
to_sfixed(-145351690.0/4294967296.0,1,-nbitq), 
to_sfixed(378023808.0/4294967296.0,1,-nbitq), 
to_sfixed(392196157.0/4294967296.0,1,-nbitq), 
to_sfixed(15921967.0/4294967296.0,1,-nbitq), 
to_sfixed(-172353610.0/4294967296.0,1,-nbitq), 
to_sfixed(-93179169.0/4294967296.0,1,-nbitq), 
to_sfixed(762928.0/4294967296.0,1,-nbitq), 
to_sfixed(-157135329.0/4294967296.0,1,-nbitq), 
to_sfixed(267059057.0/4294967296.0,1,-nbitq), 
to_sfixed(-265254128.0/4294967296.0,1,-nbitq), 
to_sfixed(-2285927.0/4294967296.0,1,-nbitq), 
to_sfixed(-376019521.0/4294967296.0,1,-nbitq), 
to_sfixed(-75530163.0/4294967296.0,1,-nbitq), 
to_sfixed(207388222.0/4294967296.0,1,-nbitq), 
to_sfixed(-89991851.0/4294967296.0,1,-nbitq), 
to_sfixed(-17205711.0/4294967296.0,1,-nbitq), 
to_sfixed(-152135315.0/4294967296.0,1,-nbitq), 
to_sfixed(62692178.0/4294967296.0,1,-nbitq), 
to_sfixed(414709048.0/4294967296.0,1,-nbitq), 
to_sfixed(-114238291.0/4294967296.0,1,-nbitq), 
to_sfixed(-45135636.0/4294967296.0,1,-nbitq), 
to_sfixed(-151348423.0/4294967296.0,1,-nbitq), 
to_sfixed(402178780.0/4294967296.0,1,-nbitq), 
to_sfixed(-288435836.0/4294967296.0,1,-nbitq), 
to_sfixed(147548364.0/4294967296.0,1,-nbitq), 
to_sfixed(755729673.0/4294967296.0,1,-nbitq), 
to_sfixed(-125559928.0/4294967296.0,1,-nbitq), 
to_sfixed(-193650339.0/4294967296.0,1,-nbitq), 
to_sfixed(90469460.0/4294967296.0,1,-nbitq), 
to_sfixed(147854623.0/4294967296.0,1,-nbitq), 
to_sfixed(-99175568.0/4294967296.0,1,-nbitq), 
to_sfixed(-328640786.0/4294967296.0,1,-nbitq), 
to_sfixed(-216323739.0/4294967296.0,1,-nbitq), 
to_sfixed(-161682669.0/4294967296.0,1,-nbitq), 
to_sfixed(-613393657.0/4294967296.0,1,-nbitq), 
to_sfixed(-363074457.0/4294967296.0,1,-nbitq), 
to_sfixed(62968770.0/4294967296.0,1,-nbitq), 
to_sfixed(36832294.0/4294967296.0,1,-nbitq), 
to_sfixed(-232587694.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-153278424.0/4294967296.0,1,-nbitq), 
to_sfixed(-409880071.0/4294967296.0,1,-nbitq), 
to_sfixed(154002014.0/4294967296.0,1,-nbitq), 
to_sfixed(-95439777.0/4294967296.0,1,-nbitq), 
to_sfixed(-320764924.0/4294967296.0,1,-nbitq), 
to_sfixed(-54997276.0/4294967296.0,1,-nbitq), 
to_sfixed(-123984860.0/4294967296.0,1,-nbitq), 
to_sfixed(-300307995.0/4294967296.0,1,-nbitq), 
to_sfixed(-453176818.0/4294967296.0,1,-nbitq), 
to_sfixed(-266073320.0/4294967296.0,1,-nbitq), 
to_sfixed(16849408.0/4294967296.0,1,-nbitq), 
to_sfixed(288471606.0/4294967296.0,1,-nbitq), 
to_sfixed(154771385.0/4294967296.0,1,-nbitq), 
to_sfixed(401426161.0/4294967296.0,1,-nbitq), 
to_sfixed(-205411651.0/4294967296.0,1,-nbitq), 
to_sfixed(-141824641.0/4294967296.0,1,-nbitq), 
to_sfixed(7054209.0/4294967296.0,1,-nbitq), 
to_sfixed(-191690534.0/4294967296.0,1,-nbitq), 
to_sfixed(307267331.0/4294967296.0,1,-nbitq), 
to_sfixed(137973794.0/4294967296.0,1,-nbitq), 
to_sfixed(36791403.0/4294967296.0,1,-nbitq), 
to_sfixed(496462769.0/4294967296.0,1,-nbitq), 
to_sfixed(444752366.0/4294967296.0,1,-nbitq), 
to_sfixed(334173167.0/4294967296.0,1,-nbitq), 
to_sfixed(289376270.0/4294967296.0,1,-nbitq), 
to_sfixed(-87849005.0/4294967296.0,1,-nbitq), 
to_sfixed(325512729.0/4294967296.0,1,-nbitq), 
to_sfixed(-496093474.0/4294967296.0,1,-nbitq), 
to_sfixed(127790222.0/4294967296.0,1,-nbitq), 
to_sfixed(301770242.0/4294967296.0,1,-nbitq), 
to_sfixed(-465003721.0/4294967296.0,1,-nbitq), 
to_sfixed(-622287123.0/4294967296.0,1,-nbitq), 
to_sfixed(176940368.0/4294967296.0,1,-nbitq), 
to_sfixed(-33868089.0/4294967296.0,1,-nbitq), 
to_sfixed(-202780770.0/4294967296.0,1,-nbitq), 
to_sfixed(388515007.0/4294967296.0,1,-nbitq), 
to_sfixed(289292909.0/4294967296.0,1,-nbitq), 
to_sfixed(300387361.0/4294967296.0,1,-nbitq), 
to_sfixed(328563477.0/4294967296.0,1,-nbitq), 
to_sfixed(1519261.0/4294967296.0,1,-nbitq), 
to_sfixed(41456406.0/4294967296.0,1,-nbitq), 
to_sfixed(272353019.0/4294967296.0,1,-nbitq), 
to_sfixed(321102629.0/4294967296.0,1,-nbitq), 
to_sfixed(171950032.0/4294967296.0,1,-nbitq), 
to_sfixed(363492752.0/4294967296.0,1,-nbitq), 
to_sfixed(688769420.0/4294967296.0,1,-nbitq), 
to_sfixed(775010.0/4294967296.0,1,-nbitq), 
to_sfixed(-239380472.0/4294967296.0,1,-nbitq), 
to_sfixed(-331922337.0/4294967296.0,1,-nbitq), 
to_sfixed(-148950604.0/4294967296.0,1,-nbitq), 
to_sfixed(-244254986.0/4294967296.0,1,-nbitq), 
to_sfixed(-315746543.0/4294967296.0,1,-nbitq), 
to_sfixed(-163876751.0/4294967296.0,1,-nbitq), 
to_sfixed(-352720677.0/4294967296.0,1,-nbitq), 
to_sfixed(315002621.0/4294967296.0,1,-nbitq), 
to_sfixed(-220852165.0/4294967296.0,1,-nbitq), 
to_sfixed(-310982435.0/4294967296.0,1,-nbitq), 
to_sfixed(-348199276.0/4294967296.0,1,-nbitq), 
to_sfixed(447251755.0/4294967296.0,1,-nbitq), 
to_sfixed(-307854394.0/4294967296.0,1,-nbitq), 
to_sfixed(133854999.0/4294967296.0,1,-nbitq), 
to_sfixed(77557592.0/4294967296.0,1,-nbitq), 
to_sfixed(-432651342.0/4294967296.0,1,-nbitq), 
to_sfixed(473390102.0/4294967296.0,1,-nbitq), 
to_sfixed(318052359.0/4294967296.0,1,-nbitq), 
to_sfixed(-426834154.0/4294967296.0,1,-nbitq), 
to_sfixed(216741838.0/4294967296.0,1,-nbitq), 
to_sfixed(289281240.0/4294967296.0,1,-nbitq), 
to_sfixed(203167482.0/4294967296.0,1,-nbitq), 
to_sfixed(-482402996.0/4294967296.0,1,-nbitq), 
to_sfixed(144124397.0/4294967296.0,1,-nbitq), 
to_sfixed(404090515.0/4294967296.0,1,-nbitq), 
to_sfixed(53128594.0/4294967296.0,1,-nbitq), 
to_sfixed(-283720499.0/4294967296.0,1,-nbitq), 
to_sfixed(-62854710.0/4294967296.0,1,-nbitq), 
to_sfixed(-543357784.0/4294967296.0,1,-nbitq), 
to_sfixed(113136475.0/4294967296.0,1,-nbitq), 
to_sfixed(106897623.0/4294967296.0,1,-nbitq), 
to_sfixed(-222935628.0/4294967296.0,1,-nbitq), 
to_sfixed(321157767.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(296129199.0/4294967296.0,1,-nbitq), 
to_sfixed(-567090358.0/4294967296.0,1,-nbitq), 
to_sfixed(441029889.0/4294967296.0,1,-nbitq), 
to_sfixed(431676776.0/4294967296.0,1,-nbitq), 
to_sfixed(-165432572.0/4294967296.0,1,-nbitq), 
to_sfixed(-393915327.0/4294967296.0,1,-nbitq), 
to_sfixed(155488158.0/4294967296.0,1,-nbitq), 
to_sfixed(-306113715.0/4294967296.0,1,-nbitq), 
to_sfixed(-368457221.0/4294967296.0,1,-nbitq), 
to_sfixed(262467537.0/4294967296.0,1,-nbitq), 
to_sfixed(-266086188.0/4294967296.0,1,-nbitq), 
to_sfixed(160717105.0/4294967296.0,1,-nbitq), 
to_sfixed(83134467.0/4294967296.0,1,-nbitq), 
to_sfixed(78724077.0/4294967296.0,1,-nbitq), 
to_sfixed(169635887.0/4294967296.0,1,-nbitq), 
to_sfixed(28026611.0/4294967296.0,1,-nbitq), 
to_sfixed(-417751952.0/4294967296.0,1,-nbitq), 
to_sfixed(-233161901.0/4294967296.0,1,-nbitq), 
to_sfixed(-171266977.0/4294967296.0,1,-nbitq), 
to_sfixed(266500968.0/4294967296.0,1,-nbitq), 
to_sfixed(-136216070.0/4294967296.0,1,-nbitq), 
to_sfixed(87098872.0/4294967296.0,1,-nbitq), 
to_sfixed(-261853447.0/4294967296.0,1,-nbitq), 
to_sfixed(203862309.0/4294967296.0,1,-nbitq), 
to_sfixed(13250611.0/4294967296.0,1,-nbitq), 
to_sfixed(-130729729.0/4294967296.0,1,-nbitq), 
to_sfixed(-188047577.0/4294967296.0,1,-nbitq), 
to_sfixed(336659549.0/4294967296.0,1,-nbitq), 
to_sfixed(293510947.0/4294967296.0,1,-nbitq), 
to_sfixed(-279920411.0/4294967296.0,1,-nbitq), 
to_sfixed(106356608.0/4294967296.0,1,-nbitq), 
to_sfixed(-201212356.0/4294967296.0,1,-nbitq), 
to_sfixed(-103549297.0/4294967296.0,1,-nbitq), 
to_sfixed(71219325.0/4294967296.0,1,-nbitq), 
to_sfixed(-312892545.0/4294967296.0,1,-nbitq), 
to_sfixed(97205948.0/4294967296.0,1,-nbitq), 
to_sfixed(-53720799.0/4294967296.0,1,-nbitq), 
to_sfixed(-427056283.0/4294967296.0,1,-nbitq), 
to_sfixed(308313750.0/4294967296.0,1,-nbitq), 
to_sfixed(-220877214.0/4294967296.0,1,-nbitq), 
to_sfixed(119481069.0/4294967296.0,1,-nbitq), 
to_sfixed(305755023.0/4294967296.0,1,-nbitq), 
to_sfixed(411975640.0/4294967296.0,1,-nbitq), 
to_sfixed(51797135.0/4294967296.0,1,-nbitq), 
to_sfixed(-208951534.0/4294967296.0,1,-nbitq), 
to_sfixed(24776782.0/4294967296.0,1,-nbitq), 
to_sfixed(158953887.0/4294967296.0,1,-nbitq), 
to_sfixed(-84087276.0/4294967296.0,1,-nbitq), 
to_sfixed(-29000936.0/4294967296.0,1,-nbitq), 
to_sfixed(-4799718.0/4294967296.0,1,-nbitq), 
to_sfixed(2775251.0/4294967296.0,1,-nbitq), 
to_sfixed(-230372699.0/4294967296.0,1,-nbitq), 
to_sfixed(134252346.0/4294967296.0,1,-nbitq), 
to_sfixed(-688218961.0/4294967296.0,1,-nbitq), 
to_sfixed(-120807827.0/4294967296.0,1,-nbitq), 
to_sfixed(199628626.0/4294967296.0,1,-nbitq), 
to_sfixed(-72651987.0/4294967296.0,1,-nbitq), 
to_sfixed(377641467.0/4294967296.0,1,-nbitq), 
to_sfixed(274795531.0/4294967296.0,1,-nbitq), 
to_sfixed(-193916948.0/4294967296.0,1,-nbitq), 
to_sfixed(-57572115.0/4294967296.0,1,-nbitq), 
to_sfixed(225920385.0/4294967296.0,1,-nbitq), 
to_sfixed(-93426056.0/4294967296.0,1,-nbitq), 
to_sfixed(135999743.0/4294967296.0,1,-nbitq), 
to_sfixed(-472030366.0/4294967296.0,1,-nbitq), 
to_sfixed(-243672484.0/4294967296.0,1,-nbitq), 
to_sfixed(-337464514.0/4294967296.0,1,-nbitq), 
to_sfixed(-22780116.0/4294967296.0,1,-nbitq), 
to_sfixed(352530295.0/4294967296.0,1,-nbitq), 
to_sfixed(114668148.0/4294967296.0,1,-nbitq), 
to_sfixed(196053071.0/4294967296.0,1,-nbitq), 
to_sfixed(74788598.0/4294967296.0,1,-nbitq), 
to_sfixed(-371706528.0/4294967296.0,1,-nbitq), 
to_sfixed(-32341517.0/4294967296.0,1,-nbitq), 
to_sfixed(28580716.0/4294967296.0,1,-nbitq), 
to_sfixed(-641008891.0/4294967296.0,1,-nbitq), 
to_sfixed(-96822672.0/4294967296.0,1,-nbitq), 
to_sfixed(267158863.0/4294967296.0,1,-nbitq), 
to_sfixed(464087896.0/4294967296.0,1,-nbitq), 
to_sfixed(211891131.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(450997286.0/4294967296.0,1,-nbitq), 
to_sfixed(-157138600.0/4294967296.0,1,-nbitq), 
to_sfixed(-59129910.0/4294967296.0,1,-nbitq), 
to_sfixed(1063070023.0/4294967296.0,1,-nbitq), 
to_sfixed(-220774382.0/4294967296.0,1,-nbitq), 
to_sfixed(283998831.0/4294967296.0,1,-nbitq), 
to_sfixed(-142622577.0/4294967296.0,1,-nbitq), 
to_sfixed(-159450458.0/4294967296.0,1,-nbitq), 
to_sfixed(-83670082.0/4294967296.0,1,-nbitq), 
to_sfixed(-302622787.0/4294967296.0,1,-nbitq), 
to_sfixed(9175748.0/4294967296.0,1,-nbitq), 
to_sfixed(-289108657.0/4294967296.0,1,-nbitq), 
to_sfixed(163003331.0/4294967296.0,1,-nbitq), 
to_sfixed(-230081441.0/4294967296.0,1,-nbitq), 
to_sfixed(7490754.0/4294967296.0,1,-nbitq), 
to_sfixed(77917314.0/4294967296.0,1,-nbitq), 
to_sfixed(384506078.0/4294967296.0,1,-nbitq), 
to_sfixed(203959054.0/4294967296.0,1,-nbitq), 
to_sfixed(-261382812.0/4294967296.0,1,-nbitq), 
to_sfixed(-59432867.0/4294967296.0,1,-nbitq), 
to_sfixed(-33476382.0/4294967296.0,1,-nbitq), 
to_sfixed(147103914.0/4294967296.0,1,-nbitq), 
to_sfixed(-607548280.0/4294967296.0,1,-nbitq), 
to_sfixed(-105684632.0/4294967296.0,1,-nbitq), 
to_sfixed(158949274.0/4294967296.0,1,-nbitq), 
to_sfixed(-88353185.0/4294967296.0,1,-nbitq), 
to_sfixed(87060936.0/4294967296.0,1,-nbitq), 
to_sfixed(48172781.0/4294967296.0,1,-nbitq), 
to_sfixed(103457294.0/4294967296.0,1,-nbitq), 
to_sfixed(-261370202.0/4294967296.0,1,-nbitq), 
to_sfixed(199830413.0/4294967296.0,1,-nbitq), 
to_sfixed(-536852476.0/4294967296.0,1,-nbitq), 
to_sfixed(-21063749.0/4294967296.0,1,-nbitq), 
to_sfixed(346670862.0/4294967296.0,1,-nbitq), 
to_sfixed(-375711757.0/4294967296.0,1,-nbitq), 
to_sfixed(-103388887.0/4294967296.0,1,-nbitq), 
to_sfixed(395983995.0/4294967296.0,1,-nbitq), 
to_sfixed(-60224849.0/4294967296.0,1,-nbitq), 
to_sfixed(-207469994.0/4294967296.0,1,-nbitq), 
to_sfixed(83857433.0/4294967296.0,1,-nbitq), 
to_sfixed(-154644264.0/4294967296.0,1,-nbitq), 
to_sfixed(211841024.0/4294967296.0,1,-nbitq), 
to_sfixed(91328817.0/4294967296.0,1,-nbitq), 
to_sfixed(-884415475.0/4294967296.0,1,-nbitq), 
to_sfixed(25727244.0/4294967296.0,1,-nbitq), 
to_sfixed(235231978.0/4294967296.0,1,-nbitq), 
to_sfixed(-269644576.0/4294967296.0,1,-nbitq), 
to_sfixed(103724691.0/4294967296.0,1,-nbitq), 
to_sfixed(313717931.0/4294967296.0,1,-nbitq), 
to_sfixed(227143543.0/4294967296.0,1,-nbitq), 
to_sfixed(34464670.0/4294967296.0,1,-nbitq), 
to_sfixed(155145809.0/4294967296.0,1,-nbitq), 
to_sfixed(811472849.0/4294967296.0,1,-nbitq), 
to_sfixed(-253773230.0/4294967296.0,1,-nbitq), 
to_sfixed(394427903.0/4294967296.0,1,-nbitq), 
to_sfixed(327779012.0/4294967296.0,1,-nbitq), 
to_sfixed(108298772.0/4294967296.0,1,-nbitq), 
to_sfixed(564939822.0/4294967296.0,1,-nbitq), 
to_sfixed(133026137.0/4294967296.0,1,-nbitq), 
to_sfixed(-244525984.0/4294967296.0,1,-nbitq), 
to_sfixed(170143504.0/4294967296.0,1,-nbitq), 
to_sfixed(191023106.0/4294967296.0,1,-nbitq), 
to_sfixed(-446209932.0/4294967296.0,1,-nbitq), 
to_sfixed(259120101.0/4294967296.0,1,-nbitq), 
to_sfixed(-523218745.0/4294967296.0,1,-nbitq), 
to_sfixed(-300408354.0/4294967296.0,1,-nbitq), 
to_sfixed(-321779230.0/4294967296.0,1,-nbitq), 
to_sfixed(138409078.0/4294967296.0,1,-nbitq), 
to_sfixed(76621580.0/4294967296.0,1,-nbitq), 
to_sfixed(-144412239.0/4294967296.0,1,-nbitq), 
to_sfixed(-313455445.0/4294967296.0,1,-nbitq), 
to_sfixed(-37445683.0/4294967296.0,1,-nbitq), 
to_sfixed(-333768786.0/4294967296.0,1,-nbitq), 
to_sfixed(42486463.0/4294967296.0,1,-nbitq), 
to_sfixed(520519717.0/4294967296.0,1,-nbitq), 
to_sfixed(-234876401.0/4294967296.0,1,-nbitq), 
to_sfixed(210010184.0/4294967296.0,1,-nbitq), 
to_sfixed(-404326605.0/4294967296.0,1,-nbitq), 
to_sfixed(-146603844.0/4294967296.0,1,-nbitq), 
to_sfixed(-194638149.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(135405475.0/4294967296.0,1,-nbitq), 
to_sfixed(-450036471.0/4294967296.0,1,-nbitq), 
to_sfixed(-216592511.0/4294967296.0,1,-nbitq), 
to_sfixed(944864100.0/4294967296.0,1,-nbitq), 
to_sfixed(292787757.0/4294967296.0,1,-nbitq), 
to_sfixed(108283509.0/4294967296.0,1,-nbitq), 
to_sfixed(-272299084.0/4294967296.0,1,-nbitq), 
to_sfixed(-118397699.0/4294967296.0,1,-nbitq), 
to_sfixed(145868954.0/4294967296.0,1,-nbitq), 
to_sfixed(-275338811.0/4294967296.0,1,-nbitq), 
to_sfixed(277484366.0/4294967296.0,1,-nbitq), 
to_sfixed(-163213614.0/4294967296.0,1,-nbitq), 
to_sfixed(81512128.0/4294967296.0,1,-nbitq), 
to_sfixed(-403448814.0/4294967296.0,1,-nbitq), 
to_sfixed(-112812813.0/4294967296.0,1,-nbitq), 
to_sfixed(-335112743.0/4294967296.0,1,-nbitq), 
to_sfixed(204231767.0/4294967296.0,1,-nbitq), 
to_sfixed(234376834.0/4294967296.0,1,-nbitq), 
to_sfixed(484913837.0/4294967296.0,1,-nbitq), 
to_sfixed(36975432.0/4294967296.0,1,-nbitq), 
to_sfixed(160998753.0/4294967296.0,1,-nbitq), 
to_sfixed(169896121.0/4294967296.0,1,-nbitq), 
to_sfixed(310188153.0/4294967296.0,1,-nbitq), 
to_sfixed(-742815169.0/4294967296.0,1,-nbitq), 
to_sfixed(-273360156.0/4294967296.0,1,-nbitq), 
to_sfixed(271425600.0/4294967296.0,1,-nbitq), 
to_sfixed(331725105.0/4294967296.0,1,-nbitq), 
to_sfixed(326998532.0/4294967296.0,1,-nbitq), 
to_sfixed(-362687017.0/4294967296.0,1,-nbitq), 
to_sfixed(-1040738590.0/4294967296.0,1,-nbitq), 
to_sfixed(484600359.0/4294967296.0,1,-nbitq), 
to_sfixed(-214422353.0/4294967296.0,1,-nbitq), 
to_sfixed(-440638912.0/4294967296.0,1,-nbitq), 
to_sfixed(-175607911.0/4294967296.0,1,-nbitq), 
to_sfixed(-305081404.0/4294967296.0,1,-nbitq), 
to_sfixed(35138314.0/4294967296.0,1,-nbitq), 
to_sfixed(382657788.0/4294967296.0,1,-nbitq), 
to_sfixed(183620305.0/4294967296.0,1,-nbitq), 
to_sfixed(-344589293.0/4294967296.0,1,-nbitq), 
to_sfixed(-43534526.0/4294967296.0,1,-nbitq), 
to_sfixed(382662817.0/4294967296.0,1,-nbitq), 
to_sfixed(-424642462.0/4294967296.0,1,-nbitq), 
to_sfixed(143046954.0/4294967296.0,1,-nbitq), 
to_sfixed(-779039430.0/4294967296.0,1,-nbitq), 
to_sfixed(693441779.0/4294967296.0,1,-nbitq), 
to_sfixed(-274962338.0/4294967296.0,1,-nbitq), 
to_sfixed(330154653.0/4294967296.0,1,-nbitq), 
to_sfixed(818760363.0/4294967296.0,1,-nbitq), 
to_sfixed(215828950.0/4294967296.0,1,-nbitq), 
to_sfixed(508787562.0/4294967296.0,1,-nbitq), 
to_sfixed(-365936807.0/4294967296.0,1,-nbitq), 
to_sfixed(-121507199.0/4294967296.0,1,-nbitq), 
to_sfixed(761151050.0/4294967296.0,1,-nbitq), 
to_sfixed(-523241255.0/4294967296.0,1,-nbitq), 
to_sfixed(602886649.0/4294967296.0,1,-nbitq), 
to_sfixed(763688532.0/4294967296.0,1,-nbitq), 
to_sfixed(112017258.0/4294967296.0,1,-nbitq), 
to_sfixed(-143482960.0/4294967296.0,1,-nbitq), 
to_sfixed(68002044.0/4294967296.0,1,-nbitq), 
to_sfixed(418748604.0/4294967296.0,1,-nbitq), 
to_sfixed(-204262063.0/4294967296.0,1,-nbitq), 
to_sfixed(81372615.0/4294967296.0,1,-nbitq), 
to_sfixed(-272877219.0/4294967296.0,1,-nbitq), 
to_sfixed(963713034.0/4294967296.0,1,-nbitq), 
to_sfixed(-485965561.0/4294967296.0,1,-nbitq), 
to_sfixed(-255745468.0/4294967296.0,1,-nbitq), 
to_sfixed(-516406637.0/4294967296.0,1,-nbitq), 
to_sfixed(358845115.0/4294967296.0,1,-nbitq), 
to_sfixed(173625861.0/4294967296.0,1,-nbitq), 
to_sfixed(-328112420.0/4294967296.0,1,-nbitq), 
to_sfixed(-961689772.0/4294967296.0,1,-nbitq), 
to_sfixed(235216627.0/4294967296.0,1,-nbitq), 
to_sfixed(-295780756.0/4294967296.0,1,-nbitq), 
to_sfixed(246283088.0/4294967296.0,1,-nbitq), 
to_sfixed(177708651.0/4294967296.0,1,-nbitq), 
to_sfixed(-876369009.0/4294967296.0,1,-nbitq), 
to_sfixed(-89023727.0/4294967296.0,1,-nbitq), 
to_sfixed(217045780.0/4294967296.0,1,-nbitq), 
to_sfixed(-164672294.0/4294967296.0,1,-nbitq), 
to_sfixed(223425712.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(296820623.0/4294967296.0,1,-nbitq), 
to_sfixed(-216500946.0/4294967296.0,1,-nbitq), 
to_sfixed(19288893.0/4294967296.0,1,-nbitq), 
to_sfixed(1125168186.0/4294967296.0,1,-nbitq), 
to_sfixed(562451069.0/4294967296.0,1,-nbitq), 
to_sfixed(-207369716.0/4294967296.0,1,-nbitq), 
to_sfixed(-196420479.0/4294967296.0,1,-nbitq), 
to_sfixed(233082544.0/4294967296.0,1,-nbitq), 
to_sfixed(844754714.0/4294967296.0,1,-nbitq), 
to_sfixed(368273130.0/4294967296.0,1,-nbitq), 
to_sfixed(756262163.0/4294967296.0,1,-nbitq), 
to_sfixed(125615434.0/4294967296.0,1,-nbitq), 
to_sfixed(95430629.0/4294967296.0,1,-nbitq), 
to_sfixed(-379966988.0/4294967296.0,1,-nbitq), 
to_sfixed(98073194.0/4294967296.0,1,-nbitq), 
to_sfixed(-232372124.0/4294967296.0,1,-nbitq), 
to_sfixed(88925009.0/4294967296.0,1,-nbitq), 
to_sfixed(372571034.0/4294967296.0,1,-nbitq), 
to_sfixed(627768396.0/4294967296.0,1,-nbitq), 
to_sfixed(697974299.0/4294967296.0,1,-nbitq), 
to_sfixed(-154214088.0/4294967296.0,1,-nbitq), 
to_sfixed(109059963.0/4294967296.0,1,-nbitq), 
to_sfixed(-49373860.0/4294967296.0,1,-nbitq), 
to_sfixed(-625031183.0/4294967296.0,1,-nbitq), 
to_sfixed(263064274.0/4294967296.0,1,-nbitq), 
to_sfixed(-133725884.0/4294967296.0,1,-nbitq), 
to_sfixed(195211068.0/4294967296.0,1,-nbitq), 
to_sfixed(395844538.0/4294967296.0,1,-nbitq), 
to_sfixed(15962905.0/4294967296.0,1,-nbitq), 
to_sfixed(-1304491837.0/4294967296.0,1,-nbitq), 
to_sfixed(41160613.0/4294967296.0,1,-nbitq), 
to_sfixed(47572738.0/4294967296.0,1,-nbitq), 
to_sfixed(128153335.0/4294967296.0,1,-nbitq), 
to_sfixed(467498310.0/4294967296.0,1,-nbitq), 
to_sfixed(-494724232.0/4294967296.0,1,-nbitq), 
to_sfixed(-344868043.0/4294967296.0,1,-nbitq), 
to_sfixed(-36351071.0/4294967296.0,1,-nbitq), 
to_sfixed(129835609.0/4294967296.0,1,-nbitq), 
to_sfixed(-620814895.0/4294967296.0,1,-nbitq), 
to_sfixed(236908048.0/4294967296.0,1,-nbitq), 
to_sfixed(-264021145.0/4294967296.0,1,-nbitq), 
to_sfixed(70167890.0/4294967296.0,1,-nbitq), 
to_sfixed(272732366.0/4294967296.0,1,-nbitq), 
to_sfixed(-753112373.0/4294967296.0,1,-nbitq), 
to_sfixed(1021398683.0/4294967296.0,1,-nbitq), 
to_sfixed(32096992.0/4294967296.0,1,-nbitq), 
to_sfixed(-223242556.0/4294967296.0,1,-nbitq), 
to_sfixed(779314241.0/4294967296.0,1,-nbitq), 
to_sfixed(-240565835.0/4294967296.0,1,-nbitq), 
to_sfixed(147850051.0/4294967296.0,1,-nbitq), 
to_sfixed(-389524683.0/4294967296.0,1,-nbitq), 
to_sfixed(453124748.0/4294967296.0,1,-nbitq), 
to_sfixed(899615500.0/4294967296.0,1,-nbitq), 
to_sfixed(-607952808.0/4294967296.0,1,-nbitq), 
to_sfixed(751430067.0/4294967296.0,1,-nbitq), 
to_sfixed(921227750.0/4294967296.0,1,-nbitq), 
to_sfixed(590580641.0/4294967296.0,1,-nbitq), 
to_sfixed(348360496.0/4294967296.0,1,-nbitq), 
to_sfixed(-312543802.0/4294967296.0,1,-nbitq), 
to_sfixed(-265562695.0/4294967296.0,1,-nbitq), 
to_sfixed(230367608.0/4294967296.0,1,-nbitq), 
to_sfixed(-336184914.0/4294967296.0,1,-nbitq), 
to_sfixed(291672106.0/4294967296.0,1,-nbitq), 
to_sfixed(1257040205.0/4294967296.0,1,-nbitq), 
to_sfixed(-209947602.0/4294967296.0,1,-nbitq), 
to_sfixed(225383095.0/4294967296.0,1,-nbitq), 
to_sfixed(-493554620.0/4294967296.0,1,-nbitq), 
to_sfixed(-273356865.0/4294967296.0,1,-nbitq), 
to_sfixed(218616603.0/4294967296.0,1,-nbitq), 
to_sfixed(-397752024.0/4294967296.0,1,-nbitq), 
to_sfixed(-903882074.0/4294967296.0,1,-nbitq), 
to_sfixed(-36655282.0/4294967296.0,1,-nbitq), 
to_sfixed(340935466.0/4294967296.0,1,-nbitq), 
to_sfixed(17897733.0/4294967296.0,1,-nbitq), 
to_sfixed(-155966816.0/4294967296.0,1,-nbitq), 
to_sfixed(-168493727.0/4294967296.0,1,-nbitq), 
to_sfixed(412059972.0/4294967296.0,1,-nbitq), 
to_sfixed(-203300338.0/4294967296.0,1,-nbitq), 
to_sfixed(-302170933.0/4294967296.0,1,-nbitq), 
to_sfixed(131979147.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(398307273.0/4294967296.0,1,-nbitq), 
to_sfixed(-516205616.0/4294967296.0,1,-nbitq), 
to_sfixed(316206882.0/4294967296.0,1,-nbitq), 
to_sfixed(581479265.0/4294967296.0,1,-nbitq), 
to_sfixed(730885974.0/4294967296.0,1,-nbitq), 
to_sfixed(131508489.0/4294967296.0,1,-nbitq), 
to_sfixed(-128257523.0/4294967296.0,1,-nbitq), 
to_sfixed(-286470674.0/4294967296.0,1,-nbitq), 
to_sfixed(893344496.0/4294967296.0,1,-nbitq), 
to_sfixed(282096566.0/4294967296.0,1,-nbitq), 
to_sfixed(738661607.0/4294967296.0,1,-nbitq), 
to_sfixed(-85578521.0/4294967296.0,1,-nbitq), 
to_sfixed(-386150882.0/4294967296.0,1,-nbitq), 
to_sfixed(-1068051775.0/4294967296.0,1,-nbitq), 
to_sfixed(166755627.0/4294967296.0,1,-nbitq), 
to_sfixed(-384301081.0/4294967296.0,1,-nbitq), 
to_sfixed(59346498.0/4294967296.0,1,-nbitq), 
to_sfixed(183877597.0/4294967296.0,1,-nbitq), 
to_sfixed(647268540.0/4294967296.0,1,-nbitq), 
to_sfixed(763200981.0/4294967296.0,1,-nbitq), 
to_sfixed(-327710505.0/4294967296.0,1,-nbitq), 
to_sfixed(-281918796.0/4294967296.0,1,-nbitq), 
to_sfixed(266727291.0/4294967296.0,1,-nbitq), 
to_sfixed(-384166354.0/4294967296.0,1,-nbitq), 
to_sfixed(298308454.0/4294967296.0,1,-nbitq), 
to_sfixed(-1006195462.0/4294967296.0,1,-nbitq), 
to_sfixed(-236299503.0/4294967296.0,1,-nbitq), 
to_sfixed(201504313.0/4294967296.0,1,-nbitq), 
to_sfixed(-260075960.0/4294967296.0,1,-nbitq), 
to_sfixed(-678027600.0/4294967296.0,1,-nbitq), 
to_sfixed(161355962.0/4294967296.0,1,-nbitq), 
to_sfixed(94834970.0/4294967296.0,1,-nbitq), 
to_sfixed(-413028735.0/4294967296.0,1,-nbitq), 
to_sfixed(383127535.0/4294967296.0,1,-nbitq), 
to_sfixed(-696330373.0/4294967296.0,1,-nbitq), 
to_sfixed(-171108945.0/4294967296.0,1,-nbitq), 
to_sfixed(-20078619.0/4294967296.0,1,-nbitq), 
to_sfixed(569512858.0/4294967296.0,1,-nbitq), 
to_sfixed(-15667999.0/4294967296.0,1,-nbitq), 
to_sfixed(621327252.0/4294967296.0,1,-nbitq), 
to_sfixed(-23795618.0/4294967296.0,1,-nbitq), 
to_sfixed(43775663.0/4294967296.0,1,-nbitq), 
to_sfixed(206185914.0/4294967296.0,1,-nbitq), 
to_sfixed(-703988439.0/4294967296.0,1,-nbitq), 
to_sfixed(663343452.0/4294967296.0,1,-nbitq), 
to_sfixed(278544569.0/4294967296.0,1,-nbitq), 
to_sfixed(235728771.0/4294967296.0,1,-nbitq), 
to_sfixed(531771076.0/4294967296.0,1,-nbitq), 
to_sfixed(-304568482.0/4294967296.0,1,-nbitq), 
to_sfixed(595374436.0/4294967296.0,1,-nbitq), 
to_sfixed(-127872413.0/4294967296.0,1,-nbitq), 
to_sfixed(-11448057.0/4294967296.0,1,-nbitq), 
to_sfixed(875669741.0/4294967296.0,1,-nbitq), 
to_sfixed(-576545695.0/4294967296.0,1,-nbitq), 
to_sfixed(268773649.0/4294967296.0,1,-nbitq), 
to_sfixed(40333704.0/4294967296.0,1,-nbitq), 
to_sfixed(-44884659.0/4294967296.0,1,-nbitq), 
to_sfixed(98368942.0/4294967296.0,1,-nbitq), 
to_sfixed(-117315940.0/4294967296.0,1,-nbitq), 
to_sfixed(-181089843.0/4294967296.0,1,-nbitq), 
to_sfixed(-43587375.0/4294967296.0,1,-nbitq), 
to_sfixed(-289185088.0/4294967296.0,1,-nbitq), 
to_sfixed(32005531.0/4294967296.0,1,-nbitq), 
to_sfixed(331747286.0/4294967296.0,1,-nbitq), 
to_sfixed(-556039582.0/4294967296.0,1,-nbitq), 
to_sfixed(-135428723.0/4294967296.0,1,-nbitq), 
to_sfixed(-119246042.0/4294967296.0,1,-nbitq), 
to_sfixed(-1254197852.0/4294967296.0,1,-nbitq), 
to_sfixed(202382560.0/4294967296.0,1,-nbitq), 
to_sfixed(-215691215.0/4294967296.0,1,-nbitq), 
to_sfixed(-1494281542.0/4294967296.0,1,-nbitq), 
to_sfixed(-117715506.0/4294967296.0,1,-nbitq), 
to_sfixed(540685806.0/4294967296.0,1,-nbitq), 
to_sfixed(383157277.0/4294967296.0,1,-nbitq), 
to_sfixed(2306773.0/4294967296.0,1,-nbitq), 
to_sfixed(166802422.0/4294967296.0,1,-nbitq), 
to_sfixed(608437412.0/4294967296.0,1,-nbitq), 
to_sfixed(260875026.0/4294967296.0,1,-nbitq), 
to_sfixed(145611075.0/4294967296.0,1,-nbitq), 
to_sfixed(-10551224.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-43441114.0/4294967296.0,1,-nbitq), 
to_sfixed(-916130089.0/4294967296.0,1,-nbitq), 
to_sfixed(232570417.0/4294967296.0,1,-nbitq), 
to_sfixed(-445821152.0/4294967296.0,1,-nbitq), 
to_sfixed(181657682.0/4294967296.0,1,-nbitq), 
to_sfixed(680969711.0/4294967296.0,1,-nbitq), 
to_sfixed(-342749706.0/4294967296.0,1,-nbitq), 
to_sfixed(-329970040.0/4294967296.0,1,-nbitq), 
to_sfixed(991218461.0/4294967296.0,1,-nbitq), 
to_sfixed(223741197.0/4294967296.0,1,-nbitq), 
to_sfixed(680123773.0/4294967296.0,1,-nbitq), 
to_sfixed(-462805087.0/4294967296.0,1,-nbitq), 
to_sfixed(-635424404.0/4294967296.0,1,-nbitq), 
to_sfixed(-1009027845.0/4294967296.0,1,-nbitq), 
to_sfixed(-117011765.0/4294967296.0,1,-nbitq), 
to_sfixed(-45965644.0/4294967296.0,1,-nbitq), 
to_sfixed(120108787.0/4294967296.0,1,-nbitq), 
to_sfixed(-328034257.0/4294967296.0,1,-nbitq), 
to_sfixed(1071551171.0/4294967296.0,1,-nbitq), 
to_sfixed(501357492.0/4294967296.0,1,-nbitq), 
to_sfixed(128460949.0/4294967296.0,1,-nbitq), 
to_sfixed(635054204.0/4294967296.0,1,-nbitq), 
to_sfixed(272237107.0/4294967296.0,1,-nbitq), 
to_sfixed(-713486377.0/4294967296.0,1,-nbitq), 
to_sfixed(-46037691.0/4294967296.0,1,-nbitq), 
to_sfixed(-936099914.0/4294967296.0,1,-nbitq), 
to_sfixed(-29804940.0/4294967296.0,1,-nbitq), 
to_sfixed(-171240546.0/4294967296.0,1,-nbitq), 
to_sfixed(-122120343.0/4294967296.0,1,-nbitq), 
to_sfixed(-897782860.0/4294967296.0,1,-nbitq), 
to_sfixed(345159113.0/4294967296.0,1,-nbitq), 
to_sfixed(424676512.0/4294967296.0,1,-nbitq), 
to_sfixed(119616403.0/4294967296.0,1,-nbitq), 
to_sfixed(646903287.0/4294967296.0,1,-nbitq), 
to_sfixed(-329267392.0/4294967296.0,1,-nbitq), 
to_sfixed(-203062010.0/4294967296.0,1,-nbitq), 
to_sfixed(-300672232.0/4294967296.0,1,-nbitq), 
to_sfixed(-12489811.0/4294967296.0,1,-nbitq), 
to_sfixed(-98857291.0/4294967296.0,1,-nbitq), 
to_sfixed(806925237.0/4294967296.0,1,-nbitq), 
to_sfixed(269146620.0/4294967296.0,1,-nbitq), 
to_sfixed(-309875650.0/4294967296.0,1,-nbitq), 
to_sfixed(-34631192.0/4294967296.0,1,-nbitq), 
to_sfixed(-1390741798.0/4294967296.0,1,-nbitq), 
to_sfixed(-37533409.0/4294967296.0,1,-nbitq), 
to_sfixed(1066150996.0/4294967296.0,1,-nbitq), 
to_sfixed(-265679101.0/4294967296.0,1,-nbitq), 
to_sfixed(499393828.0/4294967296.0,1,-nbitq), 
to_sfixed(-275951711.0/4294967296.0,1,-nbitq), 
to_sfixed(474480471.0/4294967296.0,1,-nbitq), 
to_sfixed(233064352.0/4294967296.0,1,-nbitq), 
to_sfixed(1006525347.0/4294967296.0,1,-nbitq), 
to_sfixed(637315503.0/4294967296.0,1,-nbitq), 
to_sfixed(-1396514487.0/4294967296.0,1,-nbitq), 
to_sfixed(-33237262.0/4294967296.0,1,-nbitq), 
to_sfixed(63892840.0/4294967296.0,1,-nbitq), 
to_sfixed(435794775.0/4294967296.0,1,-nbitq), 
to_sfixed(987999067.0/4294967296.0,1,-nbitq), 
to_sfixed(-295092655.0/4294967296.0,1,-nbitq), 
to_sfixed(232891899.0/4294967296.0,1,-nbitq), 
to_sfixed(33867639.0/4294967296.0,1,-nbitq), 
to_sfixed(-271421635.0/4294967296.0,1,-nbitq), 
to_sfixed(908371226.0/4294967296.0,1,-nbitq), 
to_sfixed(504328828.0/4294967296.0,1,-nbitq), 
to_sfixed(30047953.0/4294967296.0,1,-nbitq), 
to_sfixed(197970036.0/4294967296.0,1,-nbitq), 
to_sfixed(-1281824010.0/4294967296.0,1,-nbitq), 
to_sfixed(-1548709220.0/4294967296.0,1,-nbitq), 
to_sfixed(71943721.0/4294967296.0,1,-nbitq), 
to_sfixed(-988626003.0/4294967296.0,1,-nbitq), 
to_sfixed(-1021806594.0/4294967296.0,1,-nbitq), 
to_sfixed(115110116.0/4294967296.0,1,-nbitq), 
to_sfixed(318090780.0/4294967296.0,1,-nbitq), 
to_sfixed(380856986.0/4294967296.0,1,-nbitq), 
to_sfixed(353492996.0/4294967296.0,1,-nbitq), 
to_sfixed(-324190285.0/4294967296.0,1,-nbitq), 
to_sfixed(1114548568.0/4294967296.0,1,-nbitq), 
to_sfixed(-72366712.0/4294967296.0,1,-nbitq), 
to_sfixed(43089856.0/4294967296.0,1,-nbitq), 
to_sfixed(-36975262.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(706381812.0/4294967296.0,1,-nbitq), 
to_sfixed(-406539590.0/4294967296.0,1,-nbitq), 
to_sfixed(346309973.0/4294967296.0,1,-nbitq), 
to_sfixed(-52144748.0/4294967296.0,1,-nbitq), 
to_sfixed(531786388.0/4294967296.0,1,-nbitq), 
to_sfixed(-232671757.0/4294967296.0,1,-nbitq), 
to_sfixed(186443318.0/4294967296.0,1,-nbitq), 
to_sfixed(-749534359.0/4294967296.0,1,-nbitq), 
to_sfixed(1406804726.0/4294967296.0,1,-nbitq), 
to_sfixed(-94809859.0/4294967296.0,1,-nbitq), 
to_sfixed(364876313.0/4294967296.0,1,-nbitq), 
to_sfixed(-511105956.0/4294967296.0,1,-nbitq), 
to_sfixed(-459737231.0/4294967296.0,1,-nbitq), 
to_sfixed(-213877180.0/4294967296.0,1,-nbitq), 
to_sfixed(84894190.0/4294967296.0,1,-nbitq), 
to_sfixed(-118716857.0/4294967296.0,1,-nbitq), 
to_sfixed(-50790966.0/4294967296.0,1,-nbitq), 
to_sfixed(314831555.0/4294967296.0,1,-nbitq), 
to_sfixed(759131932.0/4294967296.0,1,-nbitq), 
to_sfixed(25564889.0/4294967296.0,1,-nbitq), 
to_sfixed(182372544.0/4294967296.0,1,-nbitq), 
to_sfixed(585123715.0/4294967296.0,1,-nbitq), 
to_sfixed(-57604410.0/4294967296.0,1,-nbitq), 
to_sfixed(-961075818.0/4294967296.0,1,-nbitq), 
to_sfixed(302130840.0/4294967296.0,1,-nbitq), 
to_sfixed(-959633061.0/4294967296.0,1,-nbitq), 
to_sfixed(-18703308.0/4294967296.0,1,-nbitq), 
to_sfixed(758561199.0/4294967296.0,1,-nbitq), 
to_sfixed(199519653.0/4294967296.0,1,-nbitq), 
to_sfixed(-735938161.0/4294967296.0,1,-nbitq), 
to_sfixed(637210818.0/4294967296.0,1,-nbitq), 
to_sfixed(289656650.0/4294967296.0,1,-nbitq), 
to_sfixed(-371815259.0/4294967296.0,1,-nbitq), 
to_sfixed(105638267.0/4294967296.0,1,-nbitq), 
to_sfixed(-141143297.0/4294967296.0,1,-nbitq), 
to_sfixed(465563206.0/4294967296.0,1,-nbitq), 
to_sfixed(114243907.0/4294967296.0,1,-nbitq), 
to_sfixed(-821249836.0/4294967296.0,1,-nbitq), 
to_sfixed(210159307.0/4294967296.0,1,-nbitq), 
to_sfixed(794106462.0/4294967296.0,1,-nbitq), 
to_sfixed(266757164.0/4294967296.0,1,-nbitq), 
to_sfixed(-188409951.0/4294967296.0,1,-nbitq), 
to_sfixed(628622821.0/4294967296.0,1,-nbitq), 
to_sfixed(-695360875.0/4294967296.0,1,-nbitq), 
to_sfixed(303404497.0/4294967296.0,1,-nbitq), 
to_sfixed(1202897697.0/4294967296.0,1,-nbitq), 
to_sfixed(-5091032.0/4294967296.0,1,-nbitq), 
to_sfixed(139427470.0/4294967296.0,1,-nbitq), 
to_sfixed(20720899.0/4294967296.0,1,-nbitq), 
to_sfixed(1234134912.0/4294967296.0,1,-nbitq), 
to_sfixed(19824407.0/4294967296.0,1,-nbitq), 
to_sfixed(658672620.0/4294967296.0,1,-nbitq), 
to_sfixed(235079883.0/4294967296.0,1,-nbitq), 
to_sfixed(-1046445853.0/4294967296.0,1,-nbitq), 
to_sfixed(-467094931.0/4294967296.0,1,-nbitq), 
to_sfixed(168110091.0/4294967296.0,1,-nbitq), 
to_sfixed(415116459.0/4294967296.0,1,-nbitq), 
to_sfixed(682334726.0/4294967296.0,1,-nbitq), 
to_sfixed(342841719.0/4294967296.0,1,-nbitq), 
to_sfixed(-218570183.0/4294967296.0,1,-nbitq), 
to_sfixed(-358857918.0/4294967296.0,1,-nbitq), 
to_sfixed(-363851994.0/4294967296.0,1,-nbitq), 
to_sfixed(776951674.0/4294967296.0,1,-nbitq), 
to_sfixed(781513111.0/4294967296.0,1,-nbitq), 
to_sfixed(164474772.0/4294967296.0,1,-nbitq), 
to_sfixed(-173205299.0/4294967296.0,1,-nbitq), 
to_sfixed(-848904529.0/4294967296.0,1,-nbitq), 
to_sfixed(-1201182980.0/4294967296.0,1,-nbitq), 
to_sfixed(-365783879.0/4294967296.0,1,-nbitq), 
to_sfixed(-225626988.0/4294967296.0,1,-nbitq), 
to_sfixed(-1394828958.0/4294967296.0,1,-nbitq), 
to_sfixed(13094849.0/4294967296.0,1,-nbitq), 
to_sfixed(272217.0/4294967296.0,1,-nbitq), 
to_sfixed(274363828.0/4294967296.0,1,-nbitq), 
to_sfixed(495805428.0/4294967296.0,1,-nbitq), 
to_sfixed(-469913106.0/4294967296.0,1,-nbitq), 
to_sfixed(1467819471.0/4294967296.0,1,-nbitq), 
to_sfixed(-170544466.0/4294967296.0,1,-nbitq), 
to_sfixed(-31316108.0/4294967296.0,1,-nbitq), 
to_sfixed(-44237388.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(381168843.0/4294967296.0,1,-nbitq), 
to_sfixed(-214452080.0/4294967296.0,1,-nbitq), 
to_sfixed(552360894.0/4294967296.0,1,-nbitq), 
to_sfixed(179420845.0/4294967296.0,1,-nbitq), 
to_sfixed(796840490.0/4294967296.0,1,-nbitq), 
to_sfixed(-153147069.0/4294967296.0,1,-nbitq), 
to_sfixed(163393257.0/4294967296.0,1,-nbitq), 
to_sfixed(-435218166.0/4294967296.0,1,-nbitq), 
to_sfixed(399031412.0/4294967296.0,1,-nbitq), 
to_sfixed(-7117126.0/4294967296.0,1,-nbitq), 
to_sfixed(-113383841.0/4294967296.0,1,-nbitq), 
to_sfixed(-924789256.0/4294967296.0,1,-nbitq), 
to_sfixed(-1076756179.0/4294967296.0,1,-nbitq), 
to_sfixed(-609431606.0/4294967296.0,1,-nbitq), 
to_sfixed(387966875.0/4294967296.0,1,-nbitq), 
to_sfixed(-428362446.0/4294967296.0,1,-nbitq), 
to_sfixed(-149604248.0/4294967296.0,1,-nbitq), 
to_sfixed(-318201994.0/4294967296.0,1,-nbitq), 
to_sfixed(286442568.0/4294967296.0,1,-nbitq), 
to_sfixed(-70295707.0/4294967296.0,1,-nbitq), 
to_sfixed(55793897.0/4294967296.0,1,-nbitq), 
to_sfixed(317203599.0/4294967296.0,1,-nbitq), 
to_sfixed(-145186979.0/4294967296.0,1,-nbitq), 
to_sfixed(-1193908220.0/4294967296.0,1,-nbitq), 
to_sfixed(280460172.0/4294967296.0,1,-nbitq), 
to_sfixed(-276006160.0/4294967296.0,1,-nbitq), 
to_sfixed(-24738759.0/4294967296.0,1,-nbitq), 
to_sfixed(789769125.0/4294967296.0,1,-nbitq), 
to_sfixed(160906213.0/4294967296.0,1,-nbitq), 
to_sfixed(-1087981312.0/4294967296.0,1,-nbitq), 
to_sfixed(622339219.0/4294967296.0,1,-nbitq), 
to_sfixed(1382090177.0/4294967296.0,1,-nbitq), 
to_sfixed(-38242942.0/4294967296.0,1,-nbitq), 
to_sfixed(469681841.0/4294967296.0,1,-nbitq), 
to_sfixed(38791636.0/4294967296.0,1,-nbitq), 
to_sfixed(-87216955.0/4294967296.0,1,-nbitq), 
to_sfixed(126777159.0/4294967296.0,1,-nbitq), 
to_sfixed(-498756027.0/4294967296.0,1,-nbitq), 
to_sfixed(-154623505.0/4294967296.0,1,-nbitq), 
to_sfixed(570908886.0/4294967296.0,1,-nbitq), 
to_sfixed(380440737.0/4294967296.0,1,-nbitq), 
to_sfixed(-601131615.0/4294967296.0,1,-nbitq), 
to_sfixed(379798843.0/4294967296.0,1,-nbitq), 
to_sfixed(-322674824.0/4294967296.0,1,-nbitq), 
to_sfixed(435547371.0/4294967296.0,1,-nbitq), 
to_sfixed(412909830.0/4294967296.0,1,-nbitq), 
to_sfixed(-139145919.0/4294967296.0,1,-nbitq), 
to_sfixed(-475485526.0/4294967296.0,1,-nbitq), 
to_sfixed(182202870.0/4294967296.0,1,-nbitq), 
to_sfixed(742831956.0/4294967296.0,1,-nbitq), 
to_sfixed(124788226.0/4294967296.0,1,-nbitq), 
to_sfixed(667916186.0/4294967296.0,1,-nbitq), 
to_sfixed(262357407.0/4294967296.0,1,-nbitq), 
to_sfixed(-402174774.0/4294967296.0,1,-nbitq), 
to_sfixed(-478972041.0/4294967296.0,1,-nbitq), 
to_sfixed(-444017147.0/4294967296.0,1,-nbitq), 
to_sfixed(65820894.0/4294967296.0,1,-nbitq), 
to_sfixed(-165935128.0/4294967296.0,1,-nbitq), 
to_sfixed(350371209.0/4294967296.0,1,-nbitq), 
to_sfixed(-63024030.0/4294967296.0,1,-nbitq), 
to_sfixed(152105901.0/4294967296.0,1,-nbitq), 
to_sfixed(35331854.0/4294967296.0,1,-nbitq), 
to_sfixed(1590062226.0/4294967296.0,1,-nbitq), 
to_sfixed(-103367044.0/4294967296.0,1,-nbitq), 
to_sfixed(-530308500.0/4294967296.0,1,-nbitq), 
to_sfixed(-443215964.0/4294967296.0,1,-nbitq), 
to_sfixed(86349343.0/4294967296.0,1,-nbitq), 
to_sfixed(-1347605467.0/4294967296.0,1,-nbitq), 
to_sfixed(234921340.0/4294967296.0,1,-nbitq), 
to_sfixed(19384700.0/4294967296.0,1,-nbitq), 
to_sfixed(-1088592785.0/4294967296.0,1,-nbitq), 
to_sfixed(209135451.0/4294967296.0,1,-nbitq), 
to_sfixed(783638924.0/4294967296.0,1,-nbitq), 
to_sfixed(-200798675.0/4294967296.0,1,-nbitq), 
to_sfixed(223765904.0/4294967296.0,1,-nbitq), 
to_sfixed(190245007.0/4294967296.0,1,-nbitq), 
to_sfixed(1945844847.0/4294967296.0,1,-nbitq), 
to_sfixed(-67827161.0/4294967296.0,1,-nbitq), 
to_sfixed(-201923336.0/4294967296.0,1,-nbitq), 
to_sfixed(125417135.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(73053806.0/4294967296.0,1,-nbitq), 
to_sfixed(-94231542.0/4294967296.0,1,-nbitq), 
to_sfixed(266336678.0/4294967296.0,1,-nbitq), 
to_sfixed(430689670.0/4294967296.0,1,-nbitq), 
to_sfixed(882073075.0/4294967296.0,1,-nbitq), 
to_sfixed(-654654023.0/4294967296.0,1,-nbitq), 
to_sfixed(-179424756.0/4294967296.0,1,-nbitq), 
to_sfixed(-312547899.0/4294967296.0,1,-nbitq), 
to_sfixed(616403415.0/4294967296.0,1,-nbitq), 
to_sfixed(210064104.0/4294967296.0,1,-nbitq), 
to_sfixed(3164771.0/4294967296.0,1,-nbitq), 
to_sfixed(-667920078.0/4294967296.0,1,-nbitq), 
to_sfixed(-622137258.0/4294967296.0,1,-nbitq), 
to_sfixed(71844766.0/4294967296.0,1,-nbitq), 
to_sfixed(-144775791.0/4294967296.0,1,-nbitq), 
to_sfixed(-395158664.0/4294967296.0,1,-nbitq), 
to_sfixed(228448924.0/4294967296.0,1,-nbitq), 
to_sfixed(113273702.0/4294967296.0,1,-nbitq), 
to_sfixed(-69234791.0/4294967296.0,1,-nbitq), 
to_sfixed(311073250.0/4294967296.0,1,-nbitq), 
to_sfixed(-353730220.0/4294967296.0,1,-nbitq), 
to_sfixed(371496830.0/4294967296.0,1,-nbitq), 
to_sfixed(355809241.0/4294967296.0,1,-nbitq), 
to_sfixed(-954617637.0/4294967296.0,1,-nbitq), 
to_sfixed(99337666.0/4294967296.0,1,-nbitq), 
to_sfixed(358832824.0/4294967296.0,1,-nbitq), 
to_sfixed(228416098.0/4294967296.0,1,-nbitq), 
to_sfixed(667084288.0/4294967296.0,1,-nbitq), 
to_sfixed(-212611468.0/4294967296.0,1,-nbitq), 
to_sfixed(-952757275.0/4294967296.0,1,-nbitq), 
to_sfixed(845195389.0/4294967296.0,1,-nbitq), 
to_sfixed(1264424981.0/4294967296.0,1,-nbitq), 
to_sfixed(99135915.0/4294967296.0,1,-nbitq), 
to_sfixed(759542687.0/4294967296.0,1,-nbitq), 
to_sfixed(119559278.0/4294967296.0,1,-nbitq), 
to_sfixed(275691285.0/4294967296.0,1,-nbitq), 
to_sfixed(-162735274.0/4294967296.0,1,-nbitq), 
to_sfixed(-249763647.0/4294967296.0,1,-nbitq), 
to_sfixed(-350183310.0/4294967296.0,1,-nbitq), 
to_sfixed(105964112.0/4294967296.0,1,-nbitq), 
to_sfixed(234107089.0/4294967296.0,1,-nbitq), 
to_sfixed(96738197.0/4294967296.0,1,-nbitq), 
to_sfixed(30449692.0/4294967296.0,1,-nbitq), 
to_sfixed(-178829788.0/4294967296.0,1,-nbitq), 
to_sfixed(-167888207.0/4294967296.0,1,-nbitq), 
to_sfixed(-352385011.0/4294967296.0,1,-nbitq), 
to_sfixed(130544195.0/4294967296.0,1,-nbitq), 
to_sfixed(-169088237.0/4294967296.0,1,-nbitq), 
to_sfixed(-397323079.0/4294967296.0,1,-nbitq), 
to_sfixed(207743593.0/4294967296.0,1,-nbitq), 
to_sfixed(163015980.0/4294967296.0,1,-nbitq), 
to_sfixed(616280692.0/4294967296.0,1,-nbitq), 
to_sfixed(-362371211.0/4294967296.0,1,-nbitq), 
to_sfixed(-548392170.0/4294967296.0,1,-nbitq), 
to_sfixed(-489791281.0/4294967296.0,1,-nbitq), 
to_sfixed(18174026.0/4294967296.0,1,-nbitq), 
to_sfixed(-286511679.0/4294967296.0,1,-nbitq), 
to_sfixed(-305267778.0/4294967296.0,1,-nbitq), 
to_sfixed(42564226.0/4294967296.0,1,-nbitq), 
to_sfixed(-96212457.0/4294967296.0,1,-nbitq), 
to_sfixed(-93337331.0/4294967296.0,1,-nbitq), 
to_sfixed(442091360.0/4294967296.0,1,-nbitq), 
to_sfixed(1498905809.0/4294967296.0,1,-nbitq), 
to_sfixed(452152842.0/4294967296.0,1,-nbitq), 
to_sfixed(-260065216.0/4294967296.0,1,-nbitq), 
to_sfixed(-380313326.0/4294967296.0,1,-nbitq), 
to_sfixed(833295787.0/4294967296.0,1,-nbitq), 
to_sfixed(-1173590440.0/4294967296.0,1,-nbitq), 
to_sfixed(74435368.0/4294967296.0,1,-nbitq), 
to_sfixed(-717901366.0/4294967296.0,1,-nbitq), 
to_sfixed(-1168298141.0/4294967296.0,1,-nbitq), 
to_sfixed(140713665.0/4294967296.0,1,-nbitq), 
to_sfixed(712709851.0/4294967296.0,1,-nbitq), 
to_sfixed(-306705916.0/4294967296.0,1,-nbitq), 
to_sfixed(-133239392.0/4294967296.0,1,-nbitq), 
to_sfixed(584619124.0/4294967296.0,1,-nbitq), 
to_sfixed(1741889827.0/4294967296.0,1,-nbitq), 
to_sfixed(185202746.0/4294967296.0,1,-nbitq), 
to_sfixed(-44126564.0/4294967296.0,1,-nbitq), 
to_sfixed(361449399.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-83200338.0/4294967296.0,1,-nbitq), 
to_sfixed(-561538032.0/4294967296.0,1,-nbitq), 
to_sfixed(-164517852.0/4294967296.0,1,-nbitq), 
to_sfixed(305103207.0/4294967296.0,1,-nbitq), 
to_sfixed(662784050.0/4294967296.0,1,-nbitq), 
to_sfixed(-111376490.0/4294967296.0,1,-nbitq), 
to_sfixed(-53368977.0/4294967296.0,1,-nbitq), 
to_sfixed(-558756064.0/4294967296.0,1,-nbitq), 
to_sfixed(376878719.0/4294967296.0,1,-nbitq), 
to_sfixed(405615298.0/4294967296.0,1,-nbitq), 
to_sfixed(-362883934.0/4294967296.0,1,-nbitq), 
to_sfixed(-531113579.0/4294967296.0,1,-nbitq), 
to_sfixed(-192799135.0/4294967296.0,1,-nbitq), 
to_sfixed(-167757186.0/4294967296.0,1,-nbitq), 
to_sfixed(216557236.0/4294967296.0,1,-nbitq), 
to_sfixed(86234314.0/4294967296.0,1,-nbitq), 
to_sfixed(-37849917.0/4294967296.0,1,-nbitq), 
to_sfixed(30230491.0/4294967296.0,1,-nbitq), 
to_sfixed(-155490707.0/4294967296.0,1,-nbitq), 
to_sfixed(148184163.0/4294967296.0,1,-nbitq), 
to_sfixed(78094218.0/4294967296.0,1,-nbitq), 
to_sfixed(-280272391.0/4294967296.0,1,-nbitq), 
to_sfixed(719092403.0/4294967296.0,1,-nbitq), 
to_sfixed(-537119589.0/4294967296.0,1,-nbitq), 
to_sfixed(272107775.0/4294967296.0,1,-nbitq), 
to_sfixed(666624226.0/4294967296.0,1,-nbitq), 
to_sfixed(-357004989.0/4294967296.0,1,-nbitq), 
to_sfixed(65875879.0/4294967296.0,1,-nbitq), 
to_sfixed(-403421467.0/4294967296.0,1,-nbitq), 
to_sfixed(-988216298.0/4294967296.0,1,-nbitq), 
to_sfixed(753693087.0/4294967296.0,1,-nbitq), 
to_sfixed(1320651533.0/4294967296.0,1,-nbitq), 
to_sfixed(55934285.0/4294967296.0,1,-nbitq), 
to_sfixed(63352558.0/4294967296.0,1,-nbitq), 
to_sfixed(165106832.0/4294967296.0,1,-nbitq), 
to_sfixed(479725350.0/4294967296.0,1,-nbitq), 
to_sfixed(334509740.0/4294967296.0,1,-nbitq), 
to_sfixed(-545368760.0/4294967296.0,1,-nbitq), 
to_sfixed(-33584094.0/4294967296.0,1,-nbitq), 
to_sfixed(286214597.0/4294967296.0,1,-nbitq), 
to_sfixed(384188751.0/4294967296.0,1,-nbitq), 
to_sfixed(367195370.0/4294967296.0,1,-nbitq), 
to_sfixed(1033529941.0/4294967296.0,1,-nbitq), 
to_sfixed(-195396658.0/4294967296.0,1,-nbitq), 
to_sfixed(-205244226.0/4294967296.0,1,-nbitq), 
to_sfixed(-580139528.0/4294967296.0,1,-nbitq), 
to_sfixed(-299551.0/4294967296.0,1,-nbitq), 
to_sfixed(-208832324.0/4294967296.0,1,-nbitq), 
to_sfixed(103045893.0/4294967296.0,1,-nbitq), 
to_sfixed(122567428.0/4294967296.0,1,-nbitq), 
to_sfixed(-348868831.0/4294967296.0,1,-nbitq), 
to_sfixed(749749902.0/4294967296.0,1,-nbitq), 
to_sfixed(96841592.0/4294967296.0,1,-nbitq), 
to_sfixed(-378541901.0/4294967296.0,1,-nbitq), 
to_sfixed(-322442305.0/4294967296.0,1,-nbitq), 
to_sfixed(-244014048.0/4294967296.0,1,-nbitq), 
to_sfixed(119881702.0/4294967296.0,1,-nbitq), 
to_sfixed(89398118.0/4294967296.0,1,-nbitq), 
to_sfixed(-5928034.0/4294967296.0,1,-nbitq), 
to_sfixed(-165073132.0/4294967296.0,1,-nbitq), 
to_sfixed(-291754898.0/4294967296.0,1,-nbitq), 
to_sfixed(621953331.0/4294967296.0,1,-nbitq), 
to_sfixed(524148196.0/4294967296.0,1,-nbitq), 
to_sfixed(301059647.0/4294967296.0,1,-nbitq), 
to_sfixed(-21289037.0/4294967296.0,1,-nbitq), 
to_sfixed(190850160.0/4294967296.0,1,-nbitq), 
to_sfixed(885271282.0/4294967296.0,1,-nbitq), 
to_sfixed(-1216666705.0/4294967296.0,1,-nbitq), 
to_sfixed(7774902.0/4294967296.0,1,-nbitq), 
to_sfixed(-1202416509.0/4294967296.0,1,-nbitq), 
to_sfixed(-736320133.0/4294967296.0,1,-nbitq), 
to_sfixed(-58440371.0/4294967296.0,1,-nbitq), 
to_sfixed(602690906.0/4294967296.0,1,-nbitq), 
to_sfixed(344819642.0/4294967296.0,1,-nbitq), 
to_sfixed(-15408523.0/4294967296.0,1,-nbitq), 
to_sfixed(494994222.0/4294967296.0,1,-nbitq), 
to_sfixed(1226955309.0/4294967296.0,1,-nbitq), 
to_sfixed(-105094174.0/4294967296.0,1,-nbitq), 
to_sfixed(177376819.0/4294967296.0,1,-nbitq), 
to_sfixed(-41180980.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-239758967.0/4294967296.0,1,-nbitq), 
to_sfixed(-575902669.0/4294967296.0,1,-nbitq), 
to_sfixed(546393837.0/4294967296.0,1,-nbitq), 
to_sfixed(14646564.0/4294967296.0,1,-nbitq), 
to_sfixed(-491716900.0/4294967296.0,1,-nbitq), 
to_sfixed(-252703527.0/4294967296.0,1,-nbitq), 
to_sfixed(-309181911.0/4294967296.0,1,-nbitq), 
to_sfixed(-757233764.0/4294967296.0,1,-nbitq), 
to_sfixed(313325118.0/4294967296.0,1,-nbitq), 
to_sfixed(-116442720.0/4294967296.0,1,-nbitq), 
to_sfixed(-649950158.0/4294967296.0,1,-nbitq), 
to_sfixed(-43730781.0/4294967296.0,1,-nbitq), 
to_sfixed(-161087854.0/4294967296.0,1,-nbitq), 
to_sfixed(-134206056.0/4294967296.0,1,-nbitq), 
to_sfixed(-228817801.0/4294967296.0,1,-nbitq), 
to_sfixed(274014722.0/4294967296.0,1,-nbitq), 
to_sfixed(61751064.0/4294967296.0,1,-nbitq), 
to_sfixed(328938302.0/4294967296.0,1,-nbitq), 
to_sfixed(500096832.0/4294967296.0,1,-nbitq), 
to_sfixed(123479257.0/4294967296.0,1,-nbitq), 
to_sfixed(-312487486.0/4294967296.0,1,-nbitq), 
to_sfixed(-292612816.0/4294967296.0,1,-nbitq), 
to_sfixed(729295570.0/4294967296.0,1,-nbitq), 
to_sfixed(-222166013.0/4294967296.0,1,-nbitq), 
to_sfixed(325961812.0/4294967296.0,1,-nbitq), 
to_sfixed(1142600915.0/4294967296.0,1,-nbitq), 
to_sfixed(-145734326.0/4294967296.0,1,-nbitq), 
to_sfixed(367898039.0/4294967296.0,1,-nbitq), 
to_sfixed(-483098083.0/4294967296.0,1,-nbitq), 
to_sfixed(-890586209.0/4294967296.0,1,-nbitq), 
to_sfixed(615355793.0/4294967296.0,1,-nbitq), 
to_sfixed(833704557.0/4294967296.0,1,-nbitq), 
to_sfixed(149453524.0/4294967296.0,1,-nbitq), 
to_sfixed(110837132.0/4294967296.0,1,-nbitq), 
to_sfixed(164985299.0/4294967296.0,1,-nbitq), 
to_sfixed(140085629.0/4294967296.0,1,-nbitq), 
to_sfixed(228315668.0/4294967296.0,1,-nbitq), 
to_sfixed(-865945549.0/4294967296.0,1,-nbitq), 
to_sfixed(-356129072.0/4294967296.0,1,-nbitq), 
to_sfixed(336702362.0/4294967296.0,1,-nbitq), 
to_sfixed(158409628.0/4294967296.0,1,-nbitq), 
to_sfixed(-219117315.0/4294967296.0,1,-nbitq), 
to_sfixed(375906747.0/4294967296.0,1,-nbitq), 
to_sfixed(-101808329.0/4294967296.0,1,-nbitq), 
to_sfixed(194612789.0/4294967296.0,1,-nbitq), 
to_sfixed(-596295535.0/4294967296.0,1,-nbitq), 
to_sfixed(153584762.0/4294967296.0,1,-nbitq), 
to_sfixed(-210006428.0/4294967296.0,1,-nbitq), 
to_sfixed(-366252937.0/4294967296.0,1,-nbitq), 
to_sfixed(-178343606.0/4294967296.0,1,-nbitq), 
to_sfixed(134911640.0/4294967296.0,1,-nbitq), 
to_sfixed(932198411.0/4294967296.0,1,-nbitq), 
to_sfixed(79033838.0/4294967296.0,1,-nbitq), 
to_sfixed(-899336868.0/4294967296.0,1,-nbitq), 
to_sfixed(306879720.0/4294967296.0,1,-nbitq), 
to_sfixed(-405091675.0/4294967296.0,1,-nbitq), 
to_sfixed(527944873.0/4294967296.0,1,-nbitq), 
to_sfixed(113616183.0/4294967296.0,1,-nbitq), 
to_sfixed(-330948108.0/4294967296.0,1,-nbitq), 
to_sfixed(-5304687.0/4294967296.0,1,-nbitq), 
to_sfixed(27724791.0/4294967296.0,1,-nbitq), 
to_sfixed(23223195.0/4294967296.0,1,-nbitq), 
to_sfixed(179762766.0/4294967296.0,1,-nbitq), 
to_sfixed(423484304.0/4294967296.0,1,-nbitq), 
to_sfixed(-125342997.0/4294967296.0,1,-nbitq), 
to_sfixed(-164922705.0/4294967296.0,1,-nbitq), 
to_sfixed(401560582.0/4294967296.0,1,-nbitq), 
to_sfixed(-831315327.0/4294967296.0,1,-nbitq), 
to_sfixed(-106123052.0/4294967296.0,1,-nbitq), 
to_sfixed(-785746575.0/4294967296.0,1,-nbitq), 
to_sfixed(-37245666.0/4294967296.0,1,-nbitq), 
to_sfixed(-46581043.0/4294967296.0,1,-nbitq), 
to_sfixed(358560072.0/4294967296.0,1,-nbitq), 
to_sfixed(229908758.0/4294967296.0,1,-nbitq), 
to_sfixed(-315424308.0/4294967296.0,1,-nbitq), 
to_sfixed(-96085164.0/4294967296.0,1,-nbitq), 
to_sfixed(439496615.0/4294967296.0,1,-nbitq), 
to_sfixed(112952170.0/4294967296.0,1,-nbitq), 
to_sfixed(-43971742.0/4294967296.0,1,-nbitq), 
to_sfixed(213547792.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(127926639.0/4294967296.0,1,-nbitq), 
to_sfixed(-877550616.0/4294967296.0,1,-nbitq), 
to_sfixed(1135134262.0/4294967296.0,1,-nbitq), 
to_sfixed(-285107558.0/4294967296.0,1,-nbitq), 
to_sfixed(-545957513.0/4294967296.0,1,-nbitq), 
to_sfixed(-1248269144.0/4294967296.0,1,-nbitq), 
to_sfixed(195504191.0/4294967296.0,1,-nbitq), 
to_sfixed(-255209096.0/4294967296.0,1,-nbitq), 
to_sfixed(760270303.0/4294967296.0,1,-nbitq), 
to_sfixed(116042122.0/4294967296.0,1,-nbitq), 
to_sfixed(-863812045.0/4294967296.0,1,-nbitq), 
to_sfixed(-215161584.0/4294967296.0,1,-nbitq), 
to_sfixed(-784958654.0/4294967296.0,1,-nbitq), 
to_sfixed(619512633.0/4294967296.0,1,-nbitq), 
to_sfixed(464851233.0/4294967296.0,1,-nbitq), 
to_sfixed(285361378.0/4294967296.0,1,-nbitq), 
to_sfixed(138057064.0/4294967296.0,1,-nbitq), 
to_sfixed(185415896.0/4294967296.0,1,-nbitq), 
to_sfixed(77833283.0/4294967296.0,1,-nbitq), 
to_sfixed(-48830881.0/4294967296.0,1,-nbitq), 
to_sfixed(-407525079.0/4294967296.0,1,-nbitq), 
to_sfixed(195232345.0/4294967296.0,1,-nbitq), 
to_sfixed(175820284.0/4294967296.0,1,-nbitq), 
to_sfixed(86993417.0/4294967296.0,1,-nbitq), 
to_sfixed(-271831239.0/4294967296.0,1,-nbitq), 
to_sfixed(878443478.0/4294967296.0,1,-nbitq), 
to_sfixed(177154312.0/4294967296.0,1,-nbitq), 
to_sfixed(-131101182.0/4294967296.0,1,-nbitq), 
to_sfixed(-244676919.0/4294967296.0,1,-nbitq), 
to_sfixed(-1760165741.0/4294967296.0,1,-nbitq), 
to_sfixed(-62777475.0/4294967296.0,1,-nbitq), 
to_sfixed(913296130.0/4294967296.0,1,-nbitq), 
to_sfixed(-469665894.0/4294967296.0,1,-nbitq), 
to_sfixed(-43277673.0/4294967296.0,1,-nbitq), 
to_sfixed(219678830.0/4294967296.0,1,-nbitq), 
to_sfixed(323218256.0/4294967296.0,1,-nbitq), 
to_sfixed(474486462.0/4294967296.0,1,-nbitq), 
to_sfixed(-850240896.0/4294967296.0,1,-nbitq), 
to_sfixed(-77785849.0/4294967296.0,1,-nbitq), 
to_sfixed(303543199.0/4294967296.0,1,-nbitq), 
to_sfixed(138761572.0/4294967296.0,1,-nbitq), 
to_sfixed(306663159.0/4294967296.0,1,-nbitq), 
to_sfixed(750406215.0/4294967296.0,1,-nbitq), 
to_sfixed(552066752.0/4294967296.0,1,-nbitq), 
to_sfixed(-359923383.0/4294967296.0,1,-nbitq), 
to_sfixed(-154710654.0/4294967296.0,1,-nbitq), 
to_sfixed(-224969404.0/4294967296.0,1,-nbitq), 
to_sfixed(-779912922.0/4294967296.0,1,-nbitq), 
to_sfixed(307673335.0/4294967296.0,1,-nbitq), 
to_sfixed(-604358464.0/4294967296.0,1,-nbitq), 
to_sfixed(-334974832.0/4294967296.0,1,-nbitq), 
to_sfixed(730027871.0/4294967296.0,1,-nbitq), 
to_sfixed(-10245247.0/4294967296.0,1,-nbitq), 
to_sfixed(-158972768.0/4294967296.0,1,-nbitq), 
to_sfixed(-198315045.0/4294967296.0,1,-nbitq), 
to_sfixed(-321532876.0/4294967296.0,1,-nbitq), 
to_sfixed(-111151103.0/4294967296.0,1,-nbitq), 
to_sfixed(612148378.0/4294967296.0,1,-nbitq), 
to_sfixed(248226467.0/4294967296.0,1,-nbitq), 
to_sfixed(380218059.0/4294967296.0,1,-nbitq), 
to_sfixed(-356758800.0/4294967296.0,1,-nbitq), 
to_sfixed(-276514004.0/4294967296.0,1,-nbitq), 
to_sfixed(695006678.0/4294967296.0,1,-nbitq), 
to_sfixed(592463346.0/4294967296.0,1,-nbitq), 
to_sfixed(361080100.0/4294967296.0,1,-nbitq), 
to_sfixed(35497148.0/4294967296.0,1,-nbitq), 
to_sfixed(-460510996.0/4294967296.0,1,-nbitq), 
to_sfixed(-377927951.0/4294967296.0,1,-nbitq), 
to_sfixed(323671649.0/4294967296.0,1,-nbitq), 
to_sfixed(-796756604.0/4294967296.0,1,-nbitq), 
to_sfixed(211257043.0/4294967296.0,1,-nbitq), 
to_sfixed(318855084.0/4294967296.0,1,-nbitq), 
to_sfixed(-141643900.0/4294967296.0,1,-nbitq), 
to_sfixed(-255811354.0/4294967296.0,1,-nbitq), 
to_sfixed(158178554.0/4294967296.0,1,-nbitq), 
to_sfixed(-187442478.0/4294967296.0,1,-nbitq), 
to_sfixed(930162307.0/4294967296.0,1,-nbitq), 
to_sfixed(425451815.0/4294967296.0,1,-nbitq), 
to_sfixed(-365115923.0/4294967296.0,1,-nbitq), 
to_sfixed(-237964104.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(323537835.0/4294967296.0,1,-nbitq), 
to_sfixed(-249200034.0/4294967296.0,1,-nbitq), 
to_sfixed(1037890700.0/4294967296.0,1,-nbitq), 
to_sfixed(263983407.0/4294967296.0,1,-nbitq), 
to_sfixed(-721965504.0/4294967296.0,1,-nbitq), 
to_sfixed(-832531475.0/4294967296.0,1,-nbitq), 
to_sfixed(-164835862.0/4294967296.0,1,-nbitq), 
to_sfixed(-474282471.0/4294967296.0,1,-nbitq), 
to_sfixed(965802360.0/4294967296.0,1,-nbitq), 
to_sfixed(346112748.0/4294967296.0,1,-nbitq), 
to_sfixed(-236001056.0/4294967296.0,1,-nbitq), 
to_sfixed(-323308888.0/4294967296.0,1,-nbitq), 
to_sfixed(-758303647.0/4294967296.0,1,-nbitq), 
to_sfixed(294759947.0/4294967296.0,1,-nbitq), 
to_sfixed(-241202757.0/4294967296.0,1,-nbitq), 
to_sfixed(728254576.0/4294967296.0,1,-nbitq), 
to_sfixed(168325879.0/4294967296.0,1,-nbitq), 
to_sfixed(451771596.0/4294967296.0,1,-nbitq), 
to_sfixed(-133710404.0/4294967296.0,1,-nbitq), 
to_sfixed(25941975.0/4294967296.0,1,-nbitq), 
to_sfixed(-149686542.0/4294967296.0,1,-nbitq), 
to_sfixed(261209657.0/4294967296.0,1,-nbitq), 
to_sfixed(-125797841.0/4294967296.0,1,-nbitq), 
to_sfixed(-354883808.0/4294967296.0,1,-nbitq), 
to_sfixed(-319069177.0/4294967296.0,1,-nbitq), 
to_sfixed(19839505.0/4294967296.0,1,-nbitq), 
to_sfixed(6654044.0/4294967296.0,1,-nbitq), 
to_sfixed(-93475088.0/4294967296.0,1,-nbitq), 
to_sfixed(-426123291.0/4294967296.0,1,-nbitq), 
to_sfixed(-1803712735.0/4294967296.0,1,-nbitq), 
to_sfixed(-2043508.0/4294967296.0,1,-nbitq), 
to_sfixed(204886999.0/4294967296.0,1,-nbitq), 
to_sfixed(-491794688.0/4294967296.0,1,-nbitq), 
to_sfixed(604545235.0/4294967296.0,1,-nbitq), 
to_sfixed(464491348.0/4294967296.0,1,-nbitq), 
to_sfixed(448353525.0/4294967296.0,1,-nbitq), 
to_sfixed(705873198.0/4294967296.0,1,-nbitq), 
to_sfixed(-40832469.0/4294967296.0,1,-nbitq), 
to_sfixed(-218464905.0/4294967296.0,1,-nbitq), 
to_sfixed(560042463.0/4294967296.0,1,-nbitq), 
to_sfixed(-422902675.0/4294967296.0,1,-nbitq), 
to_sfixed(827689429.0/4294967296.0,1,-nbitq), 
to_sfixed(93673210.0/4294967296.0,1,-nbitq), 
to_sfixed(888653829.0/4294967296.0,1,-nbitq), 
to_sfixed(-547982404.0/4294967296.0,1,-nbitq), 
to_sfixed(-462505804.0/4294967296.0,1,-nbitq), 
to_sfixed(-296521525.0/4294967296.0,1,-nbitq), 
to_sfixed(-789500582.0/4294967296.0,1,-nbitq), 
to_sfixed(-433954853.0/4294967296.0,1,-nbitq), 
to_sfixed(-486876319.0/4294967296.0,1,-nbitq), 
to_sfixed(173938144.0/4294967296.0,1,-nbitq), 
to_sfixed(633500228.0/4294967296.0,1,-nbitq), 
to_sfixed(-85614902.0/4294967296.0,1,-nbitq), 
to_sfixed(-4778283.0/4294967296.0,1,-nbitq), 
to_sfixed(197505829.0/4294967296.0,1,-nbitq), 
to_sfixed(-220804301.0/4294967296.0,1,-nbitq), 
to_sfixed(26838153.0/4294967296.0,1,-nbitq), 
to_sfixed(387019068.0/4294967296.0,1,-nbitq), 
to_sfixed(306877365.0/4294967296.0,1,-nbitq), 
to_sfixed(259581964.0/4294967296.0,1,-nbitq), 
to_sfixed(278812365.0/4294967296.0,1,-nbitq), 
to_sfixed(284804055.0/4294967296.0,1,-nbitq), 
to_sfixed(941042779.0/4294967296.0,1,-nbitq), 
to_sfixed(520025049.0/4294967296.0,1,-nbitq), 
to_sfixed(275351361.0/4294967296.0,1,-nbitq), 
to_sfixed(-414955482.0/4294967296.0,1,-nbitq), 
to_sfixed(-367803080.0/4294967296.0,1,-nbitq), 
to_sfixed(35801977.0/4294967296.0,1,-nbitq), 
to_sfixed(331038672.0/4294967296.0,1,-nbitq), 
to_sfixed(-363447974.0/4294967296.0,1,-nbitq), 
to_sfixed(1342721289.0/4294967296.0,1,-nbitq), 
to_sfixed(-49127666.0/4294967296.0,1,-nbitq), 
to_sfixed(14873640.0/4294967296.0,1,-nbitq), 
to_sfixed(-121559424.0/4294967296.0,1,-nbitq), 
to_sfixed(-81064833.0/4294967296.0,1,-nbitq), 
to_sfixed(85874037.0/4294967296.0,1,-nbitq), 
to_sfixed(926219911.0/4294967296.0,1,-nbitq), 
to_sfixed(348673040.0/4294967296.0,1,-nbitq), 
to_sfixed(179925847.0/4294967296.0,1,-nbitq), 
to_sfixed(414288156.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(47214655.0/4294967296.0,1,-nbitq), 
to_sfixed(614266542.0/4294967296.0,1,-nbitq), 
to_sfixed(123598716.0/4294967296.0,1,-nbitq), 
to_sfixed(-178890987.0/4294967296.0,1,-nbitq), 
to_sfixed(-351469028.0/4294967296.0,1,-nbitq), 
to_sfixed(-308499746.0/4294967296.0,1,-nbitq), 
to_sfixed(-91376785.0/4294967296.0,1,-nbitq), 
to_sfixed(12672961.0/4294967296.0,1,-nbitq), 
to_sfixed(309564901.0/4294967296.0,1,-nbitq), 
to_sfixed(147855414.0/4294967296.0,1,-nbitq), 
to_sfixed(-474577902.0/4294967296.0,1,-nbitq), 
to_sfixed(-938692725.0/4294967296.0,1,-nbitq), 
to_sfixed(-198182964.0/4294967296.0,1,-nbitq), 
to_sfixed(466969851.0/4294967296.0,1,-nbitq), 
to_sfixed(-232488072.0/4294967296.0,1,-nbitq), 
to_sfixed(-348482424.0/4294967296.0,1,-nbitq), 
to_sfixed(-54708038.0/4294967296.0,1,-nbitq), 
to_sfixed(361799050.0/4294967296.0,1,-nbitq), 
to_sfixed(-373558015.0/4294967296.0,1,-nbitq), 
to_sfixed(195604525.0/4294967296.0,1,-nbitq), 
to_sfixed(89071644.0/4294967296.0,1,-nbitq), 
to_sfixed(351163933.0/4294967296.0,1,-nbitq), 
to_sfixed(124401222.0/4294967296.0,1,-nbitq), 
to_sfixed(231107882.0/4294967296.0,1,-nbitq), 
to_sfixed(-304460140.0/4294967296.0,1,-nbitq), 
to_sfixed(362571737.0/4294967296.0,1,-nbitq), 
to_sfixed(150616698.0/4294967296.0,1,-nbitq), 
to_sfixed(-326188331.0/4294967296.0,1,-nbitq), 
to_sfixed(56075373.0/4294967296.0,1,-nbitq), 
to_sfixed(-764013540.0/4294967296.0,1,-nbitq), 
to_sfixed(-184654706.0/4294967296.0,1,-nbitq), 
to_sfixed(125414489.0/4294967296.0,1,-nbitq), 
to_sfixed(-469566884.0/4294967296.0,1,-nbitq), 
to_sfixed(400708508.0/4294967296.0,1,-nbitq), 
to_sfixed(194868631.0/4294967296.0,1,-nbitq), 
to_sfixed(563924554.0/4294967296.0,1,-nbitq), 
to_sfixed(-42824323.0/4294967296.0,1,-nbitq), 
to_sfixed(-239807463.0/4294967296.0,1,-nbitq), 
to_sfixed(41086967.0/4294967296.0,1,-nbitq), 
to_sfixed(739729083.0/4294967296.0,1,-nbitq), 
to_sfixed(-339757780.0/4294967296.0,1,-nbitq), 
to_sfixed(195476239.0/4294967296.0,1,-nbitq), 
to_sfixed(286822462.0/4294967296.0,1,-nbitq), 
to_sfixed(1253173546.0/4294967296.0,1,-nbitq), 
to_sfixed(-303485938.0/4294967296.0,1,-nbitq), 
to_sfixed(-377578706.0/4294967296.0,1,-nbitq), 
to_sfixed(-69861802.0/4294967296.0,1,-nbitq), 
to_sfixed(-1021300896.0/4294967296.0,1,-nbitq), 
to_sfixed(-210011309.0/4294967296.0,1,-nbitq), 
to_sfixed(-237138368.0/4294967296.0,1,-nbitq), 
to_sfixed(-411434113.0/4294967296.0,1,-nbitq), 
to_sfixed(-174396900.0/4294967296.0,1,-nbitq), 
to_sfixed(-13426151.0/4294967296.0,1,-nbitq), 
to_sfixed(-371396251.0/4294967296.0,1,-nbitq), 
to_sfixed(575362128.0/4294967296.0,1,-nbitq), 
to_sfixed(-509881453.0/4294967296.0,1,-nbitq), 
to_sfixed(-84808590.0/4294967296.0,1,-nbitq), 
to_sfixed(890887654.0/4294967296.0,1,-nbitq), 
to_sfixed(224088418.0/4294967296.0,1,-nbitq), 
to_sfixed(-164634243.0/4294967296.0,1,-nbitq), 
to_sfixed(244335386.0/4294967296.0,1,-nbitq), 
to_sfixed(437621517.0/4294967296.0,1,-nbitq), 
to_sfixed(532644344.0/4294967296.0,1,-nbitq), 
to_sfixed(323697124.0/4294967296.0,1,-nbitq), 
to_sfixed(-231099468.0/4294967296.0,1,-nbitq), 
to_sfixed(-345920190.0/4294967296.0,1,-nbitq), 
to_sfixed(-63011218.0/4294967296.0,1,-nbitq), 
to_sfixed(106847174.0/4294967296.0,1,-nbitq), 
to_sfixed(168417318.0/4294967296.0,1,-nbitq), 
to_sfixed(-425190510.0/4294967296.0,1,-nbitq), 
to_sfixed(1186349407.0/4294967296.0,1,-nbitq), 
to_sfixed(-33813655.0/4294967296.0,1,-nbitq), 
to_sfixed(-219309200.0/4294967296.0,1,-nbitq), 
to_sfixed(222097181.0/4294967296.0,1,-nbitq), 
to_sfixed(11530349.0/4294967296.0,1,-nbitq), 
to_sfixed(-440357971.0/4294967296.0,1,-nbitq), 
to_sfixed(845441823.0/4294967296.0,1,-nbitq), 
to_sfixed(371965042.0/4294967296.0,1,-nbitq), 
to_sfixed(-153498777.0/4294967296.0,1,-nbitq), 
to_sfixed(-352414383.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(404935610.0/4294967296.0,1,-nbitq), 
to_sfixed(546360421.0/4294967296.0,1,-nbitq), 
to_sfixed(208317401.0/4294967296.0,1,-nbitq), 
to_sfixed(-178054936.0/4294967296.0,1,-nbitq), 
to_sfixed(170968446.0/4294967296.0,1,-nbitq), 
to_sfixed(-638134399.0/4294967296.0,1,-nbitq), 
to_sfixed(-402466913.0/4294967296.0,1,-nbitq), 
to_sfixed(129751028.0/4294967296.0,1,-nbitq), 
to_sfixed(739039516.0/4294967296.0,1,-nbitq), 
to_sfixed(402806498.0/4294967296.0,1,-nbitq), 
to_sfixed(99755370.0/4294967296.0,1,-nbitq), 
to_sfixed(-492044639.0/4294967296.0,1,-nbitq), 
to_sfixed(115659585.0/4294967296.0,1,-nbitq), 
to_sfixed(284049983.0/4294967296.0,1,-nbitq), 
to_sfixed(159702166.0/4294967296.0,1,-nbitq), 
to_sfixed(-75313161.0/4294967296.0,1,-nbitq), 
to_sfixed(146033421.0/4294967296.0,1,-nbitq), 
to_sfixed(426744660.0/4294967296.0,1,-nbitq), 
to_sfixed(-369940481.0/4294967296.0,1,-nbitq), 
to_sfixed(220408060.0/4294967296.0,1,-nbitq), 
to_sfixed(325867897.0/4294967296.0,1,-nbitq), 
to_sfixed(-187191032.0/4294967296.0,1,-nbitq), 
to_sfixed(245074378.0/4294967296.0,1,-nbitq), 
to_sfixed(-195363611.0/4294967296.0,1,-nbitq), 
to_sfixed(340591466.0/4294967296.0,1,-nbitq), 
to_sfixed(773313330.0/4294967296.0,1,-nbitq), 
to_sfixed(-211848499.0/4294967296.0,1,-nbitq), 
to_sfixed(-55272203.0/4294967296.0,1,-nbitq), 
to_sfixed(792171398.0/4294967296.0,1,-nbitq), 
to_sfixed(-400553060.0/4294967296.0,1,-nbitq), 
to_sfixed(-364764461.0/4294967296.0,1,-nbitq), 
to_sfixed(53001798.0/4294967296.0,1,-nbitq), 
to_sfixed(-70287141.0/4294967296.0,1,-nbitq), 
to_sfixed(-442103083.0/4294967296.0,1,-nbitq), 
to_sfixed(464274639.0/4294967296.0,1,-nbitq), 
to_sfixed(-148696981.0/4294967296.0,1,-nbitq), 
to_sfixed(-153946988.0/4294967296.0,1,-nbitq), 
to_sfixed(35523045.0/4294967296.0,1,-nbitq), 
to_sfixed(-191737271.0/4294967296.0,1,-nbitq), 
to_sfixed(-42944006.0/4294967296.0,1,-nbitq), 
to_sfixed(410103244.0/4294967296.0,1,-nbitq), 
to_sfixed(369449575.0/4294967296.0,1,-nbitq), 
to_sfixed(605369799.0/4294967296.0,1,-nbitq), 
to_sfixed(903986388.0/4294967296.0,1,-nbitq), 
to_sfixed(-77263140.0/4294967296.0,1,-nbitq), 
to_sfixed(-22229635.0/4294967296.0,1,-nbitq), 
to_sfixed(-241937240.0/4294967296.0,1,-nbitq), 
to_sfixed(-1281562201.0/4294967296.0,1,-nbitq), 
to_sfixed(-196756704.0/4294967296.0,1,-nbitq), 
to_sfixed(-137342432.0/4294967296.0,1,-nbitq), 
to_sfixed(77068009.0/4294967296.0,1,-nbitq), 
to_sfixed(-763047090.0/4294967296.0,1,-nbitq), 
to_sfixed(91500156.0/4294967296.0,1,-nbitq), 
to_sfixed(-261143421.0/4294967296.0,1,-nbitq), 
to_sfixed(493165772.0/4294967296.0,1,-nbitq), 
to_sfixed(-547921605.0/4294967296.0,1,-nbitq), 
to_sfixed(177742970.0/4294967296.0,1,-nbitq), 
to_sfixed(433136437.0/4294967296.0,1,-nbitq), 
to_sfixed(-81621081.0/4294967296.0,1,-nbitq), 
to_sfixed(-348030111.0/4294967296.0,1,-nbitq), 
to_sfixed(52525310.0/4294967296.0,1,-nbitq), 
to_sfixed(179023282.0/4294967296.0,1,-nbitq), 
to_sfixed(570378062.0/4294967296.0,1,-nbitq), 
to_sfixed(56753184.0/4294967296.0,1,-nbitq), 
to_sfixed(-33023460.0/4294967296.0,1,-nbitq), 
to_sfixed(49749691.0/4294967296.0,1,-nbitq), 
to_sfixed(95979919.0/4294967296.0,1,-nbitq), 
to_sfixed(322814996.0/4294967296.0,1,-nbitq), 
to_sfixed(-185690916.0/4294967296.0,1,-nbitq), 
to_sfixed(-551392831.0/4294967296.0,1,-nbitq), 
to_sfixed(742969025.0/4294967296.0,1,-nbitq), 
to_sfixed(-172499983.0/4294967296.0,1,-nbitq), 
to_sfixed(-109880201.0/4294967296.0,1,-nbitq), 
to_sfixed(99898062.0/4294967296.0,1,-nbitq), 
to_sfixed(-149478496.0/4294967296.0,1,-nbitq), 
to_sfixed(-47651436.0/4294967296.0,1,-nbitq), 
to_sfixed(466270564.0/4294967296.0,1,-nbitq), 
to_sfixed(429073212.0/4294967296.0,1,-nbitq), 
to_sfixed(123949180.0/4294967296.0,1,-nbitq), 
to_sfixed(393242747.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-347614484.0/4294967296.0,1,-nbitq), 
to_sfixed(564975630.0/4294967296.0,1,-nbitq), 
to_sfixed(233325688.0/4294967296.0,1,-nbitq), 
to_sfixed(143589826.0/4294967296.0,1,-nbitq), 
to_sfixed(618010703.0/4294967296.0,1,-nbitq), 
to_sfixed(225355326.0/4294967296.0,1,-nbitq), 
to_sfixed(-350347943.0/4294967296.0,1,-nbitq), 
to_sfixed(-290566988.0/4294967296.0,1,-nbitq), 
to_sfixed(392799259.0/4294967296.0,1,-nbitq), 
to_sfixed(-185010924.0/4294967296.0,1,-nbitq), 
to_sfixed(142510457.0/4294967296.0,1,-nbitq), 
to_sfixed(-1001922328.0/4294967296.0,1,-nbitq), 
to_sfixed(50814927.0/4294967296.0,1,-nbitq), 
to_sfixed(110442099.0/4294967296.0,1,-nbitq), 
to_sfixed(-63002829.0/4294967296.0,1,-nbitq), 
to_sfixed(-883059568.0/4294967296.0,1,-nbitq), 
to_sfixed(384756746.0/4294967296.0,1,-nbitq), 
to_sfixed(-158301203.0/4294967296.0,1,-nbitq), 
to_sfixed(-98825155.0/4294967296.0,1,-nbitq), 
to_sfixed(126781971.0/4294967296.0,1,-nbitq), 
to_sfixed(262133309.0/4294967296.0,1,-nbitq), 
to_sfixed(-192155871.0/4294967296.0,1,-nbitq), 
to_sfixed(231323837.0/4294967296.0,1,-nbitq), 
to_sfixed(-271437005.0/4294967296.0,1,-nbitq), 
to_sfixed(-311344784.0/4294967296.0,1,-nbitq), 
to_sfixed(964149302.0/4294967296.0,1,-nbitq), 
to_sfixed(-168696210.0/4294967296.0,1,-nbitq), 
to_sfixed(-708775532.0/4294967296.0,1,-nbitq), 
to_sfixed(803725870.0/4294967296.0,1,-nbitq), 
to_sfixed(88652154.0/4294967296.0,1,-nbitq), 
to_sfixed(85131400.0/4294967296.0,1,-nbitq), 
to_sfixed(368040885.0/4294967296.0,1,-nbitq), 
to_sfixed(9566454.0/4294967296.0,1,-nbitq), 
to_sfixed(-605550095.0/4294967296.0,1,-nbitq), 
to_sfixed(-8977090.0/4294967296.0,1,-nbitq), 
to_sfixed(327033273.0/4294967296.0,1,-nbitq), 
to_sfixed(-427875669.0/4294967296.0,1,-nbitq), 
to_sfixed(-589724297.0/4294967296.0,1,-nbitq), 
to_sfixed(-150372507.0/4294967296.0,1,-nbitq), 
to_sfixed(465479058.0/4294967296.0,1,-nbitq), 
to_sfixed(150009982.0/4294967296.0,1,-nbitq), 
to_sfixed(321014055.0/4294967296.0,1,-nbitq), 
to_sfixed(472289308.0/4294967296.0,1,-nbitq), 
to_sfixed(176663822.0/4294967296.0,1,-nbitq), 
to_sfixed(-25159426.0/4294967296.0,1,-nbitq), 
to_sfixed(607831400.0/4294967296.0,1,-nbitq), 
to_sfixed(-9310649.0/4294967296.0,1,-nbitq), 
to_sfixed(-488128839.0/4294967296.0,1,-nbitq), 
to_sfixed(-24583966.0/4294967296.0,1,-nbitq), 
to_sfixed(118193350.0/4294967296.0,1,-nbitq), 
to_sfixed(-552130533.0/4294967296.0,1,-nbitq), 
to_sfixed(-246183085.0/4294967296.0,1,-nbitq), 
to_sfixed(204513847.0/4294967296.0,1,-nbitq), 
to_sfixed(95328086.0/4294967296.0,1,-nbitq), 
to_sfixed(262507778.0/4294967296.0,1,-nbitq), 
to_sfixed(-53384884.0/4294967296.0,1,-nbitq), 
to_sfixed(39247630.0/4294967296.0,1,-nbitq), 
to_sfixed(116409843.0/4294967296.0,1,-nbitq), 
to_sfixed(348986135.0/4294967296.0,1,-nbitq), 
to_sfixed(-344061207.0/4294967296.0,1,-nbitq), 
to_sfixed(-136445860.0/4294967296.0,1,-nbitq), 
to_sfixed(10757883.0/4294967296.0,1,-nbitq), 
to_sfixed(156463792.0/4294967296.0,1,-nbitq), 
to_sfixed(-229429065.0/4294967296.0,1,-nbitq), 
to_sfixed(-64720319.0/4294967296.0,1,-nbitq), 
to_sfixed(-255594322.0/4294967296.0,1,-nbitq), 
to_sfixed(-526922652.0/4294967296.0,1,-nbitq), 
to_sfixed(-169778142.0/4294967296.0,1,-nbitq), 
to_sfixed(-28923908.0/4294967296.0,1,-nbitq), 
to_sfixed(160094297.0/4294967296.0,1,-nbitq), 
to_sfixed(420447545.0/4294967296.0,1,-nbitq), 
to_sfixed(-34456747.0/4294967296.0,1,-nbitq), 
to_sfixed(-725161374.0/4294967296.0,1,-nbitq), 
to_sfixed(-69336045.0/4294967296.0,1,-nbitq), 
to_sfixed(-10487795.0/4294967296.0,1,-nbitq), 
to_sfixed(124013087.0/4294967296.0,1,-nbitq), 
to_sfixed(-248135193.0/4294967296.0,1,-nbitq), 
to_sfixed(35483227.0/4294967296.0,1,-nbitq), 
to_sfixed(-17499593.0/4294967296.0,1,-nbitq), 
to_sfixed(180561209.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(104191723.0/4294967296.0,1,-nbitq), 
to_sfixed(-311340925.0/4294967296.0,1,-nbitq), 
to_sfixed(-242849457.0/4294967296.0,1,-nbitq), 
to_sfixed(604565419.0/4294967296.0,1,-nbitq), 
to_sfixed(652626033.0/4294967296.0,1,-nbitq), 
to_sfixed(230096257.0/4294967296.0,1,-nbitq), 
to_sfixed(24221489.0/4294967296.0,1,-nbitq), 
to_sfixed(34175962.0/4294967296.0,1,-nbitq), 
to_sfixed(744379008.0/4294967296.0,1,-nbitq), 
to_sfixed(202114184.0/4294967296.0,1,-nbitq), 
to_sfixed(-95307605.0/4294967296.0,1,-nbitq), 
to_sfixed(-80742126.0/4294967296.0,1,-nbitq), 
to_sfixed(548755159.0/4294967296.0,1,-nbitq), 
to_sfixed(186989226.0/4294967296.0,1,-nbitq), 
to_sfixed(291577332.0/4294967296.0,1,-nbitq), 
to_sfixed(-920892699.0/4294967296.0,1,-nbitq), 
to_sfixed(-407857730.0/4294967296.0,1,-nbitq), 
to_sfixed(-298886725.0/4294967296.0,1,-nbitq), 
to_sfixed(30287614.0/4294967296.0,1,-nbitq), 
to_sfixed(92712732.0/4294967296.0,1,-nbitq), 
to_sfixed(359603067.0/4294967296.0,1,-nbitq), 
to_sfixed(351604868.0/4294967296.0,1,-nbitq), 
to_sfixed(278900016.0/4294967296.0,1,-nbitq), 
to_sfixed(390762212.0/4294967296.0,1,-nbitq), 
to_sfixed(189522392.0/4294967296.0,1,-nbitq), 
to_sfixed(525593890.0/4294967296.0,1,-nbitq), 
to_sfixed(-403486731.0/4294967296.0,1,-nbitq), 
to_sfixed(174947058.0/4294967296.0,1,-nbitq), 
to_sfixed(430200907.0/4294967296.0,1,-nbitq), 
to_sfixed(82583938.0/4294967296.0,1,-nbitq), 
to_sfixed(-538993275.0/4294967296.0,1,-nbitq), 
to_sfixed(-102599731.0/4294967296.0,1,-nbitq), 
to_sfixed(-32500397.0/4294967296.0,1,-nbitq), 
to_sfixed(-104314998.0/4294967296.0,1,-nbitq), 
to_sfixed(559443438.0/4294967296.0,1,-nbitq), 
to_sfixed(265350703.0/4294967296.0,1,-nbitq), 
to_sfixed(299359121.0/4294967296.0,1,-nbitq), 
to_sfixed(-607922790.0/4294967296.0,1,-nbitq), 
to_sfixed(221589656.0/4294967296.0,1,-nbitq), 
to_sfixed(115883659.0/4294967296.0,1,-nbitq), 
to_sfixed(429114264.0/4294967296.0,1,-nbitq), 
to_sfixed(364619942.0/4294967296.0,1,-nbitq), 
to_sfixed(184974127.0/4294967296.0,1,-nbitq), 
to_sfixed(293873148.0/4294967296.0,1,-nbitq), 
to_sfixed(63181047.0/4294967296.0,1,-nbitq), 
to_sfixed(739191090.0/4294967296.0,1,-nbitq), 
to_sfixed(-346406016.0/4294967296.0,1,-nbitq), 
to_sfixed(-386818476.0/4294967296.0,1,-nbitq), 
to_sfixed(-205548640.0/4294967296.0,1,-nbitq), 
to_sfixed(40655325.0/4294967296.0,1,-nbitq), 
to_sfixed(42255728.0/4294967296.0,1,-nbitq), 
to_sfixed(64234058.0/4294967296.0,1,-nbitq), 
to_sfixed(493631706.0/4294967296.0,1,-nbitq), 
to_sfixed(377136564.0/4294967296.0,1,-nbitq), 
to_sfixed(-275184590.0/4294967296.0,1,-nbitq), 
to_sfixed(-564612914.0/4294967296.0,1,-nbitq), 
to_sfixed(-361017541.0/4294967296.0,1,-nbitq), 
to_sfixed(314297308.0/4294967296.0,1,-nbitq), 
to_sfixed(-246261074.0/4294967296.0,1,-nbitq), 
to_sfixed(137273615.0/4294967296.0,1,-nbitq), 
to_sfixed(-12319211.0/4294967296.0,1,-nbitq), 
to_sfixed(-29414080.0/4294967296.0,1,-nbitq), 
to_sfixed(113292788.0/4294967296.0,1,-nbitq), 
to_sfixed(-174253428.0/4294967296.0,1,-nbitq), 
to_sfixed(112551121.0/4294967296.0,1,-nbitq), 
to_sfixed(120891176.0/4294967296.0,1,-nbitq), 
to_sfixed(-12783822.0/4294967296.0,1,-nbitq), 
to_sfixed(-93109471.0/4294967296.0,1,-nbitq), 
to_sfixed(204412841.0/4294967296.0,1,-nbitq), 
to_sfixed(-5497420.0/4294967296.0,1,-nbitq), 
to_sfixed(941389217.0/4294967296.0,1,-nbitq), 
to_sfixed(434445158.0/4294967296.0,1,-nbitq), 
to_sfixed(-654332223.0/4294967296.0,1,-nbitq), 
to_sfixed(-131724073.0/4294967296.0,1,-nbitq), 
to_sfixed(599728400.0/4294967296.0,1,-nbitq), 
to_sfixed(-418993084.0/4294967296.0,1,-nbitq), 
to_sfixed(156366689.0/4294967296.0,1,-nbitq), 
to_sfixed(18952234.0/4294967296.0,1,-nbitq), 
to_sfixed(44715895.0/4294967296.0,1,-nbitq), 
to_sfixed(-50776072.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-334691786.0/4294967296.0,1,-nbitq), 
to_sfixed(-540039666.0/4294967296.0,1,-nbitq), 
to_sfixed(-209579167.0/4294967296.0,1,-nbitq), 
to_sfixed(273478370.0/4294967296.0,1,-nbitq), 
to_sfixed(-98091801.0/4294967296.0,1,-nbitq), 
to_sfixed(-51678821.0/4294967296.0,1,-nbitq), 
to_sfixed(79606689.0/4294967296.0,1,-nbitq), 
to_sfixed(-51627302.0/4294967296.0,1,-nbitq), 
to_sfixed(-103319574.0/4294967296.0,1,-nbitq), 
to_sfixed(423312222.0/4294967296.0,1,-nbitq), 
to_sfixed(47358819.0/4294967296.0,1,-nbitq), 
to_sfixed(163067828.0/4294967296.0,1,-nbitq), 
to_sfixed(660858500.0/4294967296.0,1,-nbitq), 
to_sfixed(-355185867.0/4294967296.0,1,-nbitq), 
to_sfixed(-149995487.0/4294967296.0,1,-nbitq), 
to_sfixed(-540537686.0/4294967296.0,1,-nbitq), 
to_sfixed(153196185.0/4294967296.0,1,-nbitq), 
to_sfixed(-251474565.0/4294967296.0,1,-nbitq), 
to_sfixed(399195110.0/4294967296.0,1,-nbitq), 
to_sfixed(133073713.0/4294967296.0,1,-nbitq), 
to_sfixed(-31435027.0/4294967296.0,1,-nbitq), 
to_sfixed(482166563.0/4294967296.0,1,-nbitq), 
to_sfixed(595203263.0/4294967296.0,1,-nbitq), 
to_sfixed(-114897432.0/4294967296.0,1,-nbitq), 
to_sfixed(299485853.0/4294967296.0,1,-nbitq), 
to_sfixed(92927673.0/4294967296.0,1,-nbitq), 
to_sfixed(11055594.0/4294967296.0,1,-nbitq), 
to_sfixed(-486686659.0/4294967296.0,1,-nbitq), 
to_sfixed(341760570.0/4294967296.0,1,-nbitq), 
to_sfixed(-136710310.0/4294967296.0,1,-nbitq), 
to_sfixed(342237088.0/4294967296.0,1,-nbitq), 
to_sfixed(-226865757.0/4294967296.0,1,-nbitq), 
to_sfixed(281825398.0/4294967296.0,1,-nbitq), 
to_sfixed(363923055.0/4294967296.0,1,-nbitq), 
to_sfixed(273481848.0/4294967296.0,1,-nbitq), 
to_sfixed(-50489715.0/4294967296.0,1,-nbitq), 
to_sfixed(327355137.0/4294967296.0,1,-nbitq), 
to_sfixed(-761613860.0/4294967296.0,1,-nbitq), 
to_sfixed(156459912.0/4294967296.0,1,-nbitq), 
to_sfixed(517104390.0/4294967296.0,1,-nbitq), 
to_sfixed(265447783.0/4294967296.0,1,-nbitq), 
to_sfixed(400588393.0/4294967296.0,1,-nbitq), 
to_sfixed(-274204611.0/4294967296.0,1,-nbitq), 
to_sfixed(261088190.0/4294967296.0,1,-nbitq), 
to_sfixed(402364004.0/4294967296.0,1,-nbitq), 
to_sfixed(274522472.0/4294967296.0,1,-nbitq), 
to_sfixed(272439363.0/4294967296.0,1,-nbitq), 
to_sfixed(-177013532.0/4294967296.0,1,-nbitq), 
to_sfixed(-5664272.0/4294967296.0,1,-nbitq), 
to_sfixed(38613931.0/4294967296.0,1,-nbitq), 
to_sfixed(41492768.0/4294967296.0,1,-nbitq), 
to_sfixed(-132644381.0/4294967296.0,1,-nbitq), 
to_sfixed(378469867.0/4294967296.0,1,-nbitq), 
to_sfixed(-11740869.0/4294967296.0,1,-nbitq), 
to_sfixed(211164774.0/4294967296.0,1,-nbitq), 
to_sfixed(-189131836.0/4294967296.0,1,-nbitq), 
to_sfixed(-590982038.0/4294967296.0,1,-nbitq), 
to_sfixed(180159205.0/4294967296.0,1,-nbitq), 
to_sfixed(275403553.0/4294967296.0,1,-nbitq), 
to_sfixed(-95430228.0/4294967296.0,1,-nbitq), 
to_sfixed(-37370973.0/4294967296.0,1,-nbitq), 
to_sfixed(-198105491.0/4294967296.0,1,-nbitq), 
to_sfixed(393293806.0/4294967296.0,1,-nbitq), 
to_sfixed(222702705.0/4294967296.0,1,-nbitq), 
to_sfixed(340477702.0/4294967296.0,1,-nbitq), 
to_sfixed(-405217999.0/4294967296.0,1,-nbitq), 
to_sfixed(-377152390.0/4294967296.0,1,-nbitq), 
to_sfixed(-100869101.0/4294967296.0,1,-nbitq), 
to_sfixed(272470734.0/4294967296.0,1,-nbitq), 
to_sfixed(-74532470.0/4294967296.0,1,-nbitq), 
to_sfixed(11238897.0/4294967296.0,1,-nbitq), 
to_sfixed(-134924398.0/4294967296.0,1,-nbitq), 
to_sfixed(91947857.0/4294967296.0,1,-nbitq), 
to_sfixed(-112734175.0/4294967296.0,1,-nbitq), 
to_sfixed(194706841.0/4294967296.0,1,-nbitq), 
to_sfixed(-577720112.0/4294967296.0,1,-nbitq), 
to_sfixed(512623116.0/4294967296.0,1,-nbitq), 
to_sfixed(-24431441.0/4294967296.0,1,-nbitq), 
to_sfixed(-220545038.0/4294967296.0,1,-nbitq), 
to_sfixed(-342976002.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(114901121.0/4294967296.0,1,-nbitq), 
to_sfixed(-473486750.0/4294967296.0,1,-nbitq), 
to_sfixed(348979587.0/4294967296.0,1,-nbitq), 
to_sfixed(-90221522.0/4294967296.0,1,-nbitq), 
to_sfixed(222683771.0/4294967296.0,1,-nbitq), 
to_sfixed(148930842.0/4294967296.0,1,-nbitq), 
to_sfixed(-248642922.0/4294967296.0,1,-nbitq), 
to_sfixed(-529445262.0/4294967296.0,1,-nbitq), 
to_sfixed(80214751.0/4294967296.0,1,-nbitq), 
to_sfixed(-303922949.0/4294967296.0,1,-nbitq), 
to_sfixed(-408979414.0/4294967296.0,1,-nbitq), 
to_sfixed(-184584519.0/4294967296.0,1,-nbitq), 
to_sfixed(-62191998.0/4294967296.0,1,-nbitq), 
to_sfixed(-360955664.0/4294967296.0,1,-nbitq), 
to_sfixed(-321901905.0/4294967296.0,1,-nbitq), 
to_sfixed(-37189554.0/4294967296.0,1,-nbitq), 
to_sfixed(-270829304.0/4294967296.0,1,-nbitq), 
to_sfixed(-53650525.0/4294967296.0,1,-nbitq), 
to_sfixed(595777306.0/4294967296.0,1,-nbitq), 
to_sfixed(-442245793.0/4294967296.0,1,-nbitq), 
to_sfixed(196553019.0/4294967296.0,1,-nbitq), 
to_sfixed(-173243920.0/4294967296.0,1,-nbitq), 
to_sfixed(30507088.0/4294967296.0,1,-nbitq), 
to_sfixed(107925871.0/4294967296.0,1,-nbitq), 
to_sfixed(-25345855.0/4294967296.0,1,-nbitq), 
to_sfixed(657329489.0/4294967296.0,1,-nbitq), 
to_sfixed(109410590.0/4294967296.0,1,-nbitq), 
to_sfixed(-411964525.0/4294967296.0,1,-nbitq), 
to_sfixed(94157663.0/4294967296.0,1,-nbitq), 
to_sfixed(367935163.0/4294967296.0,1,-nbitq), 
to_sfixed(-273482404.0/4294967296.0,1,-nbitq), 
to_sfixed(238304754.0/4294967296.0,1,-nbitq), 
to_sfixed(163326018.0/4294967296.0,1,-nbitq), 
to_sfixed(146775768.0/4294967296.0,1,-nbitq), 
to_sfixed(540254532.0/4294967296.0,1,-nbitq), 
to_sfixed(-319472688.0/4294967296.0,1,-nbitq), 
to_sfixed(-210435125.0/4294967296.0,1,-nbitq), 
to_sfixed(-151982178.0/4294967296.0,1,-nbitq), 
to_sfixed(-194199695.0/4294967296.0,1,-nbitq), 
to_sfixed(172410750.0/4294967296.0,1,-nbitq), 
to_sfixed(268669665.0/4294967296.0,1,-nbitq), 
to_sfixed(315233402.0/4294967296.0,1,-nbitq), 
to_sfixed(466061424.0/4294967296.0,1,-nbitq), 
to_sfixed(-112947924.0/4294967296.0,1,-nbitq), 
to_sfixed(449402946.0/4294967296.0,1,-nbitq), 
to_sfixed(-89713816.0/4294967296.0,1,-nbitq), 
to_sfixed(-146546234.0/4294967296.0,1,-nbitq), 
to_sfixed(21198046.0/4294967296.0,1,-nbitq), 
to_sfixed(-19979882.0/4294967296.0,1,-nbitq), 
to_sfixed(-196053153.0/4294967296.0,1,-nbitq), 
to_sfixed(55073493.0/4294967296.0,1,-nbitq), 
to_sfixed(-75150327.0/4294967296.0,1,-nbitq), 
to_sfixed(-98821287.0/4294967296.0,1,-nbitq), 
to_sfixed(136538021.0/4294967296.0,1,-nbitq), 
to_sfixed(92012481.0/4294967296.0,1,-nbitq), 
to_sfixed(-161067519.0/4294967296.0,1,-nbitq), 
to_sfixed(-166046395.0/4294967296.0,1,-nbitq), 
to_sfixed(158988726.0/4294967296.0,1,-nbitq), 
to_sfixed(190277895.0/4294967296.0,1,-nbitq), 
to_sfixed(-246210804.0/4294967296.0,1,-nbitq), 
to_sfixed(-267908080.0/4294967296.0,1,-nbitq), 
to_sfixed(5235785.0/4294967296.0,1,-nbitq), 
to_sfixed(168080447.0/4294967296.0,1,-nbitq), 
to_sfixed(-275911751.0/4294967296.0,1,-nbitq), 
to_sfixed(-77934733.0/4294967296.0,1,-nbitq), 
to_sfixed(302894212.0/4294967296.0,1,-nbitq), 
to_sfixed(57442554.0/4294967296.0,1,-nbitq), 
to_sfixed(333227013.0/4294967296.0,1,-nbitq), 
to_sfixed(257221532.0/4294967296.0,1,-nbitq), 
to_sfixed(-268336897.0/4294967296.0,1,-nbitq), 
to_sfixed(276576306.0/4294967296.0,1,-nbitq), 
to_sfixed(111810314.0/4294967296.0,1,-nbitq), 
to_sfixed(-136545124.0/4294967296.0,1,-nbitq), 
to_sfixed(278528206.0/4294967296.0,1,-nbitq), 
to_sfixed(-276456977.0/4294967296.0,1,-nbitq), 
to_sfixed(-327874571.0/4294967296.0,1,-nbitq), 
to_sfixed(-190761536.0/4294967296.0,1,-nbitq), 
to_sfixed(-189158289.0/4294967296.0,1,-nbitq), 
to_sfixed(-431410507.0/4294967296.0,1,-nbitq), 
to_sfixed(213954957.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(223562220.0/4294967296.0,1,-nbitq), 
to_sfixed(-8898600.0/4294967296.0,1,-nbitq), 
to_sfixed(-186914009.0/4294967296.0,1,-nbitq), 
to_sfixed(73939796.0/4294967296.0,1,-nbitq), 
to_sfixed(-226118267.0/4294967296.0,1,-nbitq), 
to_sfixed(247126174.0/4294967296.0,1,-nbitq), 
to_sfixed(-392404166.0/4294967296.0,1,-nbitq), 
to_sfixed(47004539.0/4294967296.0,1,-nbitq), 
to_sfixed(112318056.0/4294967296.0,1,-nbitq), 
to_sfixed(184498317.0/4294967296.0,1,-nbitq), 
to_sfixed(-460867826.0/4294967296.0,1,-nbitq), 
to_sfixed(-141012145.0/4294967296.0,1,-nbitq), 
to_sfixed(5224342.0/4294967296.0,1,-nbitq), 
to_sfixed(-263381160.0/4294967296.0,1,-nbitq), 
to_sfixed(122319879.0/4294967296.0,1,-nbitq), 
to_sfixed(-557947160.0/4294967296.0,1,-nbitq), 
to_sfixed(35421028.0/4294967296.0,1,-nbitq), 
to_sfixed(-29271853.0/4294967296.0,1,-nbitq), 
to_sfixed(512726029.0/4294967296.0,1,-nbitq), 
to_sfixed(128758660.0/4294967296.0,1,-nbitq), 
to_sfixed(20400354.0/4294967296.0,1,-nbitq), 
to_sfixed(72417757.0/4294967296.0,1,-nbitq), 
to_sfixed(269056040.0/4294967296.0,1,-nbitq), 
to_sfixed(-81457052.0/4294967296.0,1,-nbitq), 
to_sfixed(-184248950.0/4294967296.0,1,-nbitq), 
to_sfixed(279597675.0/4294967296.0,1,-nbitq), 
to_sfixed(193074668.0/4294967296.0,1,-nbitq), 
to_sfixed(-428225082.0/4294967296.0,1,-nbitq), 
to_sfixed(179520363.0/4294967296.0,1,-nbitq), 
to_sfixed(-313152053.0/4294967296.0,1,-nbitq), 
to_sfixed(-28605220.0/4294967296.0,1,-nbitq), 
to_sfixed(-367461679.0/4294967296.0,1,-nbitq), 
to_sfixed(-26698364.0/4294967296.0,1,-nbitq), 
to_sfixed(3933302.0/4294967296.0,1,-nbitq), 
to_sfixed(377803995.0/4294967296.0,1,-nbitq), 
to_sfixed(-311756779.0/4294967296.0,1,-nbitq), 
to_sfixed(-161258541.0/4294967296.0,1,-nbitq), 
to_sfixed(224388188.0/4294967296.0,1,-nbitq), 
to_sfixed(-151654623.0/4294967296.0,1,-nbitq), 
to_sfixed(-200262325.0/4294967296.0,1,-nbitq), 
to_sfixed(82265951.0/4294967296.0,1,-nbitq), 
to_sfixed(323399657.0/4294967296.0,1,-nbitq), 
to_sfixed(-62787375.0/4294967296.0,1,-nbitq), 
to_sfixed(414577453.0/4294967296.0,1,-nbitq), 
to_sfixed(55867403.0/4294967296.0,1,-nbitq), 
to_sfixed(327993839.0/4294967296.0,1,-nbitq), 
to_sfixed(59834417.0/4294967296.0,1,-nbitq), 
to_sfixed(97504129.0/4294967296.0,1,-nbitq), 
to_sfixed(95637743.0/4294967296.0,1,-nbitq), 
to_sfixed(-2739398.0/4294967296.0,1,-nbitq), 
to_sfixed(236143183.0/4294967296.0,1,-nbitq), 
to_sfixed(385163840.0/4294967296.0,1,-nbitq), 
to_sfixed(-527773493.0/4294967296.0,1,-nbitq), 
to_sfixed(443608450.0/4294967296.0,1,-nbitq), 
to_sfixed(250282074.0/4294967296.0,1,-nbitq), 
to_sfixed(319450144.0/4294967296.0,1,-nbitq), 
to_sfixed(-202358904.0/4294967296.0,1,-nbitq), 
to_sfixed(-517906789.0/4294967296.0,1,-nbitq), 
to_sfixed(-72008495.0/4294967296.0,1,-nbitq), 
to_sfixed(-288187777.0/4294967296.0,1,-nbitq), 
to_sfixed(222915730.0/4294967296.0,1,-nbitq), 
to_sfixed(-225160526.0/4294967296.0,1,-nbitq), 
to_sfixed(145189892.0/4294967296.0,1,-nbitq), 
to_sfixed(-334459609.0/4294967296.0,1,-nbitq), 
to_sfixed(284381655.0/4294967296.0,1,-nbitq), 
to_sfixed(-271217596.0/4294967296.0,1,-nbitq), 
to_sfixed(-171263475.0/4294967296.0,1,-nbitq), 
to_sfixed(-415655306.0/4294967296.0,1,-nbitq), 
to_sfixed(265504828.0/4294967296.0,1,-nbitq), 
to_sfixed(-279598375.0/4294967296.0,1,-nbitq), 
to_sfixed(108786141.0/4294967296.0,1,-nbitq), 
to_sfixed(257444085.0/4294967296.0,1,-nbitq), 
to_sfixed(7883419.0/4294967296.0,1,-nbitq), 
to_sfixed(139436425.0/4294967296.0,1,-nbitq), 
to_sfixed(-55027083.0/4294967296.0,1,-nbitq), 
to_sfixed(-82236562.0/4294967296.0,1,-nbitq), 
to_sfixed(316261107.0/4294967296.0,1,-nbitq), 
to_sfixed(-74286496.0/4294967296.0,1,-nbitq), 
to_sfixed(-608469116.0/4294967296.0,1,-nbitq), 
to_sfixed(96533621.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(106692208.0/4294967296.0,1,-nbitq), 
to_sfixed(-489198069.0/4294967296.0,1,-nbitq), 
to_sfixed(-116964147.0/4294967296.0,1,-nbitq), 
to_sfixed(57913654.0/4294967296.0,1,-nbitq), 
to_sfixed(-73801560.0/4294967296.0,1,-nbitq), 
to_sfixed(194941307.0/4294967296.0,1,-nbitq), 
to_sfixed(291793676.0/4294967296.0,1,-nbitq), 
to_sfixed(-484655186.0/4294967296.0,1,-nbitq), 
to_sfixed(179357348.0/4294967296.0,1,-nbitq), 
to_sfixed(346535603.0/4294967296.0,1,-nbitq), 
to_sfixed(331473371.0/4294967296.0,1,-nbitq), 
to_sfixed(-197019827.0/4294967296.0,1,-nbitq), 
to_sfixed(-89727206.0/4294967296.0,1,-nbitq), 
to_sfixed(173277297.0/4294967296.0,1,-nbitq), 
to_sfixed(-4930189.0/4294967296.0,1,-nbitq), 
to_sfixed(-115505610.0/4294967296.0,1,-nbitq), 
to_sfixed(-288448275.0/4294967296.0,1,-nbitq), 
to_sfixed(371196324.0/4294967296.0,1,-nbitq), 
to_sfixed(269966837.0/4294967296.0,1,-nbitq), 
to_sfixed(-409670295.0/4294967296.0,1,-nbitq), 
to_sfixed(23914655.0/4294967296.0,1,-nbitq), 
to_sfixed(407532432.0/4294967296.0,1,-nbitq), 
to_sfixed(620376439.0/4294967296.0,1,-nbitq), 
to_sfixed(-327403961.0/4294967296.0,1,-nbitq), 
to_sfixed(-28218370.0/4294967296.0,1,-nbitq), 
to_sfixed(128849212.0/4294967296.0,1,-nbitq), 
to_sfixed(-228280037.0/4294967296.0,1,-nbitq), 
to_sfixed(-524202531.0/4294967296.0,1,-nbitq), 
to_sfixed(-275688814.0/4294967296.0,1,-nbitq), 
to_sfixed(362074329.0/4294967296.0,1,-nbitq), 
to_sfixed(-66245546.0/4294967296.0,1,-nbitq), 
to_sfixed(-258271862.0/4294967296.0,1,-nbitq), 
to_sfixed(-150093707.0/4294967296.0,1,-nbitq), 
to_sfixed(107167800.0/4294967296.0,1,-nbitq), 
to_sfixed(140159481.0/4294967296.0,1,-nbitq), 
to_sfixed(37303895.0/4294967296.0,1,-nbitq), 
to_sfixed(-200229306.0/4294967296.0,1,-nbitq), 
to_sfixed(-285693368.0/4294967296.0,1,-nbitq), 
to_sfixed(84311259.0/4294967296.0,1,-nbitq), 
to_sfixed(-239138422.0/4294967296.0,1,-nbitq), 
to_sfixed(-13230288.0/4294967296.0,1,-nbitq), 
to_sfixed(-267264425.0/4294967296.0,1,-nbitq), 
to_sfixed(201090423.0/4294967296.0,1,-nbitq), 
to_sfixed(96418021.0/4294967296.0,1,-nbitq), 
to_sfixed(136519345.0/4294967296.0,1,-nbitq), 
to_sfixed(304074842.0/4294967296.0,1,-nbitq), 
to_sfixed(-305309670.0/4294967296.0,1,-nbitq), 
to_sfixed(-40276708.0/4294967296.0,1,-nbitq), 
to_sfixed(227717038.0/4294967296.0,1,-nbitq), 
to_sfixed(488674697.0/4294967296.0,1,-nbitq), 
to_sfixed(127710999.0/4294967296.0,1,-nbitq), 
to_sfixed(185791919.0/4294967296.0,1,-nbitq), 
to_sfixed(176373549.0/4294967296.0,1,-nbitq), 
to_sfixed(-281803147.0/4294967296.0,1,-nbitq), 
to_sfixed(269791481.0/4294967296.0,1,-nbitq), 
to_sfixed(-135977292.0/4294967296.0,1,-nbitq), 
to_sfixed(381376754.0/4294967296.0,1,-nbitq), 
to_sfixed(-466069094.0/4294967296.0,1,-nbitq), 
to_sfixed(-319435291.0/4294967296.0,1,-nbitq), 
to_sfixed(-245407773.0/4294967296.0,1,-nbitq), 
to_sfixed(363958947.0/4294967296.0,1,-nbitq), 
to_sfixed(-193884943.0/4294967296.0,1,-nbitq), 
to_sfixed(289277123.0/4294967296.0,1,-nbitq), 
to_sfixed(-275226740.0/4294967296.0,1,-nbitq), 
to_sfixed(-134944899.0/4294967296.0,1,-nbitq), 
to_sfixed(-106779013.0/4294967296.0,1,-nbitq), 
to_sfixed(118006894.0/4294967296.0,1,-nbitq), 
to_sfixed(237075053.0/4294967296.0,1,-nbitq), 
to_sfixed(-184164585.0/4294967296.0,1,-nbitq), 
to_sfixed(-212950533.0/4294967296.0,1,-nbitq), 
to_sfixed(1408585.0/4294967296.0,1,-nbitq), 
to_sfixed(-386841564.0/4294967296.0,1,-nbitq), 
to_sfixed(191869754.0/4294967296.0,1,-nbitq), 
to_sfixed(236521255.0/4294967296.0,1,-nbitq), 
to_sfixed(423651750.0/4294967296.0,1,-nbitq), 
to_sfixed(-125645291.0/4294967296.0,1,-nbitq), 
to_sfixed(205978350.0/4294967296.0,1,-nbitq), 
to_sfixed(184745101.0/4294967296.0,1,-nbitq), 
to_sfixed(-415319811.0/4294967296.0,1,-nbitq), 
to_sfixed(6902715.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-125021618.0/4294967296.0,1,-nbitq), 
to_sfixed(-249984615.0/4294967296.0,1,-nbitq), 
to_sfixed(199355390.0/4294967296.0,1,-nbitq), 
to_sfixed(-48058840.0/4294967296.0,1,-nbitq), 
to_sfixed(-14493726.0/4294967296.0,1,-nbitq), 
to_sfixed(207823808.0/4294967296.0,1,-nbitq), 
to_sfixed(3684383.0/4294967296.0,1,-nbitq), 
to_sfixed(-452595956.0/4294967296.0,1,-nbitq), 
to_sfixed(176461116.0/4294967296.0,1,-nbitq), 
to_sfixed(-67306837.0/4294967296.0,1,-nbitq), 
to_sfixed(-148066287.0/4294967296.0,1,-nbitq), 
to_sfixed(-264124274.0/4294967296.0,1,-nbitq), 
to_sfixed(351174834.0/4294967296.0,1,-nbitq), 
to_sfixed(78635850.0/4294967296.0,1,-nbitq), 
to_sfixed(-145856304.0/4294967296.0,1,-nbitq), 
to_sfixed(-124199640.0/4294967296.0,1,-nbitq), 
to_sfixed(-191466068.0/4294967296.0,1,-nbitq), 
to_sfixed(-18686382.0/4294967296.0,1,-nbitq), 
to_sfixed(-200547668.0/4294967296.0,1,-nbitq), 
to_sfixed(-339177464.0/4294967296.0,1,-nbitq), 
to_sfixed(-372082317.0/4294967296.0,1,-nbitq), 
to_sfixed(-44092158.0/4294967296.0,1,-nbitq), 
to_sfixed(610938207.0/4294967296.0,1,-nbitq), 
to_sfixed(421630525.0/4294967296.0,1,-nbitq), 
to_sfixed(30824171.0/4294967296.0,1,-nbitq), 
to_sfixed(-85493418.0/4294967296.0,1,-nbitq), 
to_sfixed(-161439869.0/4294967296.0,1,-nbitq), 
to_sfixed(-4543057.0/4294967296.0,1,-nbitq), 
to_sfixed(384710576.0/4294967296.0,1,-nbitq), 
to_sfixed(-269240425.0/4294967296.0,1,-nbitq), 
to_sfixed(-315566331.0/4294967296.0,1,-nbitq), 
to_sfixed(-145367134.0/4294967296.0,1,-nbitq), 
to_sfixed(-127362615.0/4294967296.0,1,-nbitq), 
to_sfixed(43172913.0/4294967296.0,1,-nbitq), 
to_sfixed(96245113.0/4294967296.0,1,-nbitq), 
to_sfixed(723352.0/4294967296.0,1,-nbitq), 
to_sfixed(178350837.0/4294967296.0,1,-nbitq), 
to_sfixed(-66234861.0/4294967296.0,1,-nbitq), 
to_sfixed(121785800.0/4294967296.0,1,-nbitq), 
to_sfixed(-241762339.0/4294967296.0,1,-nbitq), 
to_sfixed(275493298.0/4294967296.0,1,-nbitq), 
to_sfixed(366592958.0/4294967296.0,1,-nbitq), 
to_sfixed(69584247.0/4294967296.0,1,-nbitq), 
to_sfixed(92650190.0/4294967296.0,1,-nbitq), 
to_sfixed(-9993289.0/4294967296.0,1,-nbitq), 
to_sfixed(-148417691.0/4294967296.0,1,-nbitq), 
to_sfixed(-418546069.0/4294967296.0,1,-nbitq), 
to_sfixed(-114460932.0/4294967296.0,1,-nbitq), 
to_sfixed(104454001.0/4294967296.0,1,-nbitq), 
to_sfixed(234536247.0/4294967296.0,1,-nbitq), 
to_sfixed(220170353.0/4294967296.0,1,-nbitq), 
to_sfixed(-296905279.0/4294967296.0,1,-nbitq), 
to_sfixed(-527039696.0/4294967296.0,1,-nbitq), 
to_sfixed(45442328.0/4294967296.0,1,-nbitq), 
to_sfixed(78762601.0/4294967296.0,1,-nbitq), 
to_sfixed(399578732.0/4294967296.0,1,-nbitq), 
to_sfixed(228651183.0/4294967296.0,1,-nbitq), 
to_sfixed(183941068.0/4294967296.0,1,-nbitq), 
to_sfixed(-111693578.0/4294967296.0,1,-nbitq), 
to_sfixed(293394635.0/4294967296.0,1,-nbitq), 
to_sfixed(-388023593.0/4294967296.0,1,-nbitq), 
to_sfixed(206112945.0/4294967296.0,1,-nbitq), 
to_sfixed(-246604950.0/4294967296.0,1,-nbitq), 
to_sfixed(211981826.0/4294967296.0,1,-nbitq), 
to_sfixed(-25365954.0/4294967296.0,1,-nbitq), 
to_sfixed(265674177.0/4294967296.0,1,-nbitq), 
to_sfixed(775318322.0/4294967296.0,1,-nbitq), 
to_sfixed(-92692243.0/4294967296.0,1,-nbitq), 
to_sfixed(-73673905.0/4294967296.0,1,-nbitq), 
to_sfixed(114273521.0/4294967296.0,1,-nbitq), 
to_sfixed(-321596133.0/4294967296.0,1,-nbitq), 
to_sfixed(-163826227.0/4294967296.0,1,-nbitq), 
to_sfixed(57419494.0/4294967296.0,1,-nbitq), 
to_sfixed(244052448.0/4294967296.0,1,-nbitq), 
to_sfixed(397870451.0/4294967296.0,1,-nbitq), 
to_sfixed(-246423542.0/4294967296.0,1,-nbitq), 
to_sfixed(-58207737.0/4294967296.0,1,-nbitq), 
to_sfixed(-489372618.0/4294967296.0,1,-nbitq), 
to_sfixed(-566079401.0/4294967296.0,1,-nbitq), 
to_sfixed(-287556757.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(26046966.0/4294967296.0,1,-nbitq), 
to_sfixed(-310167104.0/4294967296.0,1,-nbitq), 
to_sfixed(-209122823.0/4294967296.0,1,-nbitq), 
to_sfixed(307129255.0/4294967296.0,1,-nbitq), 
to_sfixed(354450758.0/4294967296.0,1,-nbitq), 
to_sfixed(-287873381.0/4294967296.0,1,-nbitq), 
to_sfixed(-161625364.0/4294967296.0,1,-nbitq), 
to_sfixed(-253521598.0/4294967296.0,1,-nbitq), 
to_sfixed(192761833.0/4294967296.0,1,-nbitq), 
to_sfixed(257940998.0/4294967296.0,1,-nbitq), 
to_sfixed(-414388236.0/4294967296.0,1,-nbitq), 
to_sfixed(14236268.0/4294967296.0,1,-nbitq), 
to_sfixed(135280842.0/4294967296.0,1,-nbitq), 
to_sfixed(398940433.0/4294967296.0,1,-nbitq), 
to_sfixed(239346993.0/4294967296.0,1,-nbitq), 
to_sfixed(-270673761.0/4294967296.0,1,-nbitq), 
to_sfixed(-172404444.0/4294967296.0,1,-nbitq), 
to_sfixed(-63231425.0/4294967296.0,1,-nbitq), 
to_sfixed(426877426.0/4294967296.0,1,-nbitq), 
to_sfixed(-400595694.0/4294967296.0,1,-nbitq), 
to_sfixed(-1727719.0/4294967296.0,1,-nbitq), 
to_sfixed(509330368.0/4294967296.0,1,-nbitq), 
to_sfixed(480402745.0/4294967296.0,1,-nbitq), 
to_sfixed(264679052.0/4294967296.0,1,-nbitq), 
to_sfixed(-65731445.0/4294967296.0,1,-nbitq), 
to_sfixed(55440242.0/4294967296.0,1,-nbitq), 
to_sfixed(-319580108.0/4294967296.0,1,-nbitq), 
to_sfixed(-513309080.0/4294967296.0,1,-nbitq), 
to_sfixed(50416185.0/4294967296.0,1,-nbitq), 
to_sfixed(34371267.0/4294967296.0,1,-nbitq), 
to_sfixed(-573955265.0/4294967296.0,1,-nbitq), 
to_sfixed(-345023995.0/4294967296.0,1,-nbitq), 
to_sfixed(121085936.0/4294967296.0,1,-nbitq), 
to_sfixed(-119552377.0/4294967296.0,1,-nbitq), 
to_sfixed(-131764387.0/4294967296.0,1,-nbitq), 
to_sfixed(-279643908.0/4294967296.0,1,-nbitq), 
to_sfixed(56061368.0/4294967296.0,1,-nbitq), 
to_sfixed(102208482.0/4294967296.0,1,-nbitq), 
to_sfixed(1869743.0/4294967296.0,1,-nbitq), 
to_sfixed(-293237351.0/4294967296.0,1,-nbitq), 
to_sfixed(-370224454.0/4294967296.0,1,-nbitq), 
to_sfixed(50553516.0/4294967296.0,1,-nbitq), 
to_sfixed(-257717914.0/4294967296.0,1,-nbitq), 
to_sfixed(-266348312.0/4294967296.0,1,-nbitq), 
to_sfixed(-276138591.0/4294967296.0,1,-nbitq), 
to_sfixed(-23711536.0/4294967296.0,1,-nbitq), 
to_sfixed(209893299.0/4294967296.0,1,-nbitq), 
to_sfixed(-474020696.0/4294967296.0,1,-nbitq), 
to_sfixed(-198465315.0/4294967296.0,1,-nbitq), 
to_sfixed(-205064048.0/4294967296.0,1,-nbitq), 
to_sfixed(-348192515.0/4294967296.0,1,-nbitq), 
to_sfixed(-163656427.0/4294967296.0,1,-nbitq), 
to_sfixed(-203315433.0/4294967296.0,1,-nbitq), 
to_sfixed(-257386742.0/4294967296.0,1,-nbitq), 
to_sfixed(186286560.0/4294967296.0,1,-nbitq), 
to_sfixed(-102834880.0/4294967296.0,1,-nbitq), 
to_sfixed(133383763.0/4294967296.0,1,-nbitq), 
to_sfixed(-28426117.0/4294967296.0,1,-nbitq), 
to_sfixed(227616365.0/4294967296.0,1,-nbitq), 
to_sfixed(388892621.0/4294967296.0,1,-nbitq), 
to_sfixed(306626804.0/4294967296.0,1,-nbitq), 
to_sfixed(-203997660.0/4294967296.0,1,-nbitq), 
to_sfixed(-459960613.0/4294967296.0,1,-nbitq), 
to_sfixed(-53681106.0/4294967296.0,1,-nbitq), 
to_sfixed(141094475.0/4294967296.0,1,-nbitq), 
to_sfixed(147876111.0/4294967296.0,1,-nbitq), 
to_sfixed(629333630.0/4294967296.0,1,-nbitq), 
to_sfixed(-87881115.0/4294967296.0,1,-nbitq), 
to_sfixed(-78478259.0/4294967296.0,1,-nbitq), 
to_sfixed(-187880258.0/4294967296.0,1,-nbitq), 
to_sfixed(-105706568.0/4294967296.0,1,-nbitq), 
to_sfixed(-243857836.0/4294967296.0,1,-nbitq), 
to_sfixed(-15094409.0/4294967296.0,1,-nbitq), 
to_sfixed(316323785.0/4294967296.0,1,-nbitq), 
to_sfixed(401252532.0/4294967296.0,1,-nbitq), 
to_sfixed(-481260107.0/4294967296.0,1,-nbitq), 
to_sfixed(-117688338.0/4294967296.0,1,-nbitq), 
to_sfixed(-343491971.0/4294967296.0,1,-nbitq), 
to_sfixed(-201958599.0/4294967296.0,1,-nbitq), 
to_sfixed(-326655344.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-141484765.0/4294967296.0,1,-nbitq), 
to_sfixed(137624469.0/4294967296.0,1,-nbitq), 
to_sfixed(-9421901.0/4294967296.0,1,-nbitq), 
to_sfixed(180311347.0/4294967296.0,1,-nbitq), 
to_sfixed(-269402051.0/4294967296.0,1,-nbitq), 
to_sfixed(-66127735.0/4294967296.0,1,-nbitq), 
to_sfixed(151336683.0/4294967296.0,1,-nbitq), 
to_sfixed(16031923.0/4294967296.0,1,-nbitq), 
to_sfixed(-354350197.0/4294967296.0,1,-nbitq), 
to_sfixed(24034162.0/4294967296.0,1,-nbitq), 
to_sfixed(-217752122.0/4294967296.0,1,-nbitq), 
to_sfixed(223924702.0/4294967296.0,1,-nbitq), 
to_sfixed(271382498.0/4294967296.0,1,-nbitq), 
to_sfixed(420500429.0/4294967296.0,1,-nbitq), 
to_sfixed(-316302839.0/4294967296.0,1,-nbitq), 
to_sfixed(-485524448.0/4294967296.0,1,-nbitq), 
to_sfixed(5106052.0/4294967296.0,1,-nbitq), 
to_sfixed(326424922.0/4294967296.0,1,-nbitq), 
to_sfixed(-56100185.0/4294967296.0,1,-nbitq), 
to_sfixed(24871875.0/4294967296.0,1,-nbitq), 
to_sfixed(-98696141.0/4294967296.0,1,-nbitq), 
to_sfixed(14939791.0/4294967296.0,1,-nbitq), 
to_sfixed(149543073.0/4294967296.0,1,-nbitq), 
to_sfixed(133202235.0/4294967296.0,1,-nbitq), 
to_sfixed(-299550097.0/4294967296.0,1,-nbitq), 
to_sfixed(89677489.0/4294967296.0,1,-nbitq), 
to_sfixed(268775747.0/4294967296.0,1,-nbitq), 
to_sfixed(-240832989.0/4294967296.0,1,-nbitq), 
to_sfixed(-180920524.0/4294967296.0,1,-nbitq), 
to_sfixed(-233796902.0/4294967296.0,1,-nbitq), 
to_sfixed(-479984252.0/4294967296.0,1,-nbitq), 
to_sfixed(-434359087.0/4294967296.0,1,-nbitq), 
to_sfixed(367266254.0/4294967296.0,1,-nbitq), 
to_sfixed(-448822759.0/4294967296.0,1,-nbitq), 
to_sfixed(-174911393.0/4294967296.0,1,-nbitq), 
to_sfixed(-231292177.0/4294967296.0,1,-nbitq), 
to_sfixed(393716296.0/4294967296.0,1,-nbitq), 
to_sfixed(227306427.0/4294967296.0,1,-nbitq), 
to_sfixed(63849492.0/4294967296.0,1,-nbitq), 
to_sfixed(193175771.0/4294967296.0,1,-nbitq), 
to_sfixed(-115859751.0/4294967296.0,1,-nbitq), 
to_sfixed(250521588.0/4294967296.0,1,-nbitq), 
to_sfixed(-70336570.0/4294967296.0,1,-nbitq), 
to_sfixed(-270442812.0/4294967296.0,1,-nbitq), 
to_sfixed(-123653991.0/4294967296.0,1,-nbitq), 
to_sfixed(139863655.0/4294967296.0,1,-nbitq), 
to_sfixed(309803437.0/4294967296.0,1,-nbitq), 
to_sfixed(180406344.0/4294967296.0,1,-nbitq), 
to_sfixed(-186928360.0/4294967296.0,1,-nbitq), 
to_sfixed(-92979539.0/4294967296.0,1,-nbitq), 
to_sfixed(9986820.0/4294967296.0,1,-nbitq), 
to_sfixed(141973045.0/4294967296.0,1,-nbitq), 
to_sfixed(152134219.0/4294967296.0,1,-nbitq), 
to_sfixed(-37460559.0/4294967296.0,1,-nbitq), 
to_sfixed(325096233.0/4294967296.0,1,-nbitq), 
to_sfixed(233996250.0/4294967296.0,1,-nbitq), 
to_sfixed(376344115.0/4294967296.0,1,-nbitq), 
to_sfixed(149686539.0/4294967296.0,1,-nbitq), 
to_sfixed(-15332623.0/4294967296.0,1,-nbitq), 
to_sfixed(276159181.0/4294967296.0,1,-nbitq), 
to_sfixed(-401967265.0/4294967296.0,1,-nbitq), 
to_sfixed(-177852870.0/4294967296.0,1,-nbitq), 
to_sfixed(-259765476.0/4294967296.0,1,-nbitq), 
to_sfixed(-18980924.0/4294967296.0,1,-nbitq), 
to_sfixed(244533129.0/4294967296.0,1,-nbitq), 
to_sfixed(-446874279.0/4294967296.0,1,-nbitq), 
to_sfixed(201792843.0/4294967296.0,1,-nbitq), 
to_sfixed(-81078319.0/4294967296.0,1,-nbitq), 
to_sfixed(275750685.0/4294967296.0,1,-nbitq), 
to_sfixed(-48911151.0/4294967296.0,1,-nbitq), 
to_sfixed(-464393391.0/4294967296.0,1,-nbitq), 
to_sfixed(117059447.0/4294967296.0,1,-nbitq), 
to_sfixed(-493006003.0/4294967296.0,1,-nbitq), 
to_sfixed(-145248845.0/4294967296.0,1,-nbitq), 
to_sfixed(287833672.0/4294967296.0,1,-nbitq), 
to_sfixed(-597111317.0/4294967296.0,1,-nbitq), 
to_sfixed(301719947.0/4294967296.0,1,-nbitq), 
to_sfixed(-13757892.0/4294967296.0,1,-nbitq), 
to_sfixed(-507207852.0/4294967296.0,1,-nbitq), 
to_sfixed(348104368.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(9839719.0/4294967296.0,1,-nbitq), 
to_sfixed(-44502707.0/4294967296.0,1,-nbitq), 
to_sfixed(526284078.0/4294967296.0,1,-nbitq), 
to_sfixed(-221084471.0/4294967296.0,1,-nbitq), 
to_sfixed(-260655771.0/4294967296.0,1,-nbitq), 
to_sfixed(304677220.0/4294967296.0,1,-nbitq), 
to_sfixed(-392033810.0/4294967296.0,1,-nbitq), 
to_sfixed(-498945219.0/4294967296.0,1,-nbitq), 
to_sfixed(6988081.0/4294967296.0,1,-nbitq), 
to_sfixed(-38947557.0/4294967296.0,1,-nbitq), 
to_sfixed(-193409292.0/4294967296.0,1,-nbitq), 
to_sfixed(15103177.0/4294967296.0,1,-nbitq), 
to_sfixed(-112551414.0/4294967296.0,1,-nbitq), 
to_sfixed(-324321445.0/4294967296.0,1,-nbitq), 
to_sfixed(197637736.0/4294967296.0,1,-nbitq), 
to_sfixed(-547483070.0/4294967296.0,1,-nbitq), 
to_sfixed(-168116379.0/4294967296.0,1,-nbitq), 
to_sfixed(396362148.0/4294967296.0,1,-nbitq), 
to_sfixed(173804784.0/4294967296.0,1,-nbitq), 
to_sfixed(217314316.0/4294967296.0,1,-nbitq), 
to_sfixed(-231048760.0/4294967296.0,1,-nbitq), 
to_sfixed(117667213.0/4294967296.0,1,-nbitq), 
to_sfixed(531744.0/4294967296.0,1,-nbitq), 
to_sfixed(433081661.0/4294967296.0,1,-nbitq), 
to_sfixed(260885588.0/4294967296.0,1,-nbitq), 
to_sfixed(313786170.0/4294967296.0,1,-nbitq), 
to_sfixed(-193478532.0/4294967296.0,1,-nbitq), 
to_sfixed(-235743516.0/4294967296.0,1,-nbitq), 
to_sfixed(221578962.0/4294967296.0,1,-nbitq), 
to_sfixed(225091499.0/4294967296.0,1,-nbitq), 
to_sfixed(-366781024.0/4294967296.0,1,-nbitq), 
to_sfixed(-782138897.0/4294967296.0,1,-nbitq), 
to_sfixed(-32353412.0/4294967296.0,1,-nbitq), 
to_sfixed(-400783683.0/4294967296.0,1,-nbitq), 
to_sfixed(-311106275.0/4294967296.0,1,-nbitq), 
to_sfixed(-13718095.0/4294967296.0,1,-nbitq), 
to_sfixed(433958930.0/4294967296.0,1,-nbitq), 
to_sfixed(-232296083.0/4294967296.0,1,-nbitq), 
to_sfixed(-3663998.0/4294967296.0,1,-nbitq), 
to_sfixed(105825243.0/4294967296.0,1,-nbitq), 
to_sfixed(-165308244.0/4294967296.0,1,-nbitq), 
to_sfixed(-265500317.0/4294967296.0,1,-nbitq), 
to_sfixed(-15574436.0/4294967296.0,1,-nbitq), 
to_sfixed(-325536507.0/4294967296.0,1,-nbitq), 
to_sfixed(608044898.0/4294967296.0,1,-nbitq), 
to_sfixed(312141403.0/4294967296.0,1,-nbitq), 
to_sfixed(-98928258.0/4294967296.0,1,-nbitq), 
to_sfixed(-337611118.0/4294967296.0,1,-nbitq), 
to_sfixed(-112689331.0/4294967296.0,1,-nbitq), 
to_sfixed(-43304325.0/4294967296.0,1,-nbitq), 
to_sfixed(-8892309.0/4294967296.0,1,-nbitq), 
to_sfixed(-413108658.0/4294967296.0,1,-nbitq), 
to_sfixed(115756901.0/4294967296.0,1,-nbitq), 
to_sfixed(28969639.0/4294967296.0,1,-nbitq), 
to_sfixed(-225451995.0/4294967296.0,1,-nbitq), 
to_sfixed(-57177900.0/4294967296.0,1,-nbitq), 
to_sfixed(420606761.0/4294967296.0,1,-nbitq), 
to_sfixed(-347928970.0/4294967296.0,1,-nbitq), 
to_sfixed(368090853.0/4294967296.0,1,-nbitq), 
to_sfixed(233410229.0/4294967296.0,1,-nbitq), 
to_sfixed(33116325.0/4294967296.0,1,-nbitq), 
to_sfixed(176980096.0/4294967296.0,1,-nbitq), 
to_sfixed(185898288.0/4294967296.0,1,-nbitq), 
to_sfixed(151202199.0/4294967296.0,1,-nbitq), 
to_sfixed(-262041941.0/4294967296.0,1,-nbitq), 
to_sfixed(205421612.0/4294967296.0,1,-nbitq), 
to_sfixed(158580319.0/4294967296.0,1,-nbitq), 
to_sfixed(-151638735.0/4294967296.0,1,-nbitq), 
to_sfixed(420301024.0/4294967296.0,1,-nbitq), 
to_sfixed(99497385.0/4294967296.0,1,-nbitq), 
to_sfixed(-582290566.0/4294967296.0,1,-nbitq), 
to_sfixed(320771101.0/4294967296.0,1,-nbitq), 
to_sfixed(262977704.0/4294967296.0,1,-nbitq), 
to_sfixed(148557640.0/4294967296.0,1,-nbitq), 
to_sfixed(45631298.0/4294967296.0,1,-nbitq), 
to_sfixed(-457680587.0/4294967296.0,1,-nbitq), 
to_sfixed(67003951.0/4294967296.0,1,-nbitq), 
to_sfixed(-423889444.0/4294967296.0,1,-nbitq), 
to_sfixed(-71410754.0/4294967296.0,1,-nbitq), 
to_sfixed(136339130.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-396898628.0/4294967296.0,1,-nbitq), 
to_sfixed(16109032.0/4294967296.0,1,-nbitq), 
to_sfixed(439813395.0/4294967296.0,1,-nbitq), 
to_sfixed(495257811.0/4294967296.0,1,-nbitq), 
to_sfixed(229935440.0/4294967296.0,1,-nbitq), 
to_sfixed(75188974.0/4294967296.0,1,-nbitq), 
to_sfixed(40377940.0/4294967296.0,1,-nbitq), 
to_sfixed(102153602.0/4294967296.0,1,-nbitq), 
to_sfixed(-12033057.0/4294967296.0,1,-nbitq), 
to_sfixed(-156160137.0/4294967296.0,1,-nbitq), 
to_sfixed(-74256364.0/4294967296.0,1,-nbitq), 
to_sfixed(178766522.0/4294967296.0,1,-nbitq), 
to_sfixed(-426901970.0/4294967296.0,1,-nbitq), 
to_sfixed(-490160836.0/4294967296.0,1,-nbitq), 
to_sfixed(-56555723.0/4294967296.0,1,-nbitq), 
to_sfixed(-492848488.0/4294967296.0,1,-nbitq), 
to_sfixed(-280109719.0/4294967296.0,1,-nbitq), 
to_sfixed(-252278298.0/4294967296.0,1,-nbitq), 
to_sfixed(-156948855.0/4294967296.0,1,-nbitq), 
to_sfixed(110303228.0/4294967296.0,1,-nbitq), 
to_sfixed(-286541617.0/4294967296.0,1,-nbitq), 
to_sfixed(411682810.0/4294967296.0,1,-nbitq), 
to_sfixed(209306807.0/4294967296.0,1,-nbitq), 
to_sfixed(202490610.0/4294967296.0,1,-nbitq), 
to_sfixed(83436513.0/4294967296.0,1,-nbitq), 
to_sfixed(356642273.0/4294967296.0,1,-nbitq), 
to_sfixed(-56231470.0/4294967296.0,1,-nbitq), 
to_sfixed(319179956.0/4294967296.0,1,-nbitq), 
to_sfixed(-40543165.0/4294967296.0,1,-nbitq), 
to_sfixed(-377896436.0/4294967296.0,1,-nbitq), 
to_sfixed(397457715.0/4294967296.0,1,-nbitq), 
to_sfixed(-640167135.0/4294967296.0,1,-nbitq), 
to_sfixed(36033319.0/4294967296.0,1,-nbitq), 
to_sfixed(334942571.0/4294967296.0,1,-nbitq), 
to_sfixed(41555418.0/4294967296.0,1,-nbitq), 
to_sfixed(-71014768.0/4294967296.0,1,-nbitq), 
to_sfixed(-152160918.0/4294967296.0,1,-nbitq), 
to_sfixed(-43659315.0/4294967296.0,1,-nbitq), 
to_sfixed(110848872.0/4294967296.0,1,-nbitq), 
to_sfixed(321933139.0/4294967296.0,1,-nbitq), 
to_sfixed(488042726.0/4294967296.0,1,-nbitq), 
to_sfixed(-291521056.0/4294967296.0,1,-nbitq), 
to_sfixed(142613571.0/4294967296.0,1,-nbitq), 
to_sfixed(-689877647.0/4294967296.0,1,-nbitq), 
to_sfixed(7129060.0/4294967296.0,1,-nbitq), 
to_sfixed(678017065.0/4294967296.0,1,-nbitq), 
to_sfixed(-439720678.0/4294967296.0,1,-nbitq), 
to_sfixed(760621304.0/4294967296.0,1,-nbitq), 
to_sfixed(-143460212.0/4294967296.0,1,-nbitq), 
to_sfixed(-32802002.0/4294967296.0,1,-nbitq), 
to_sfixed(-99858015.0/4294967296.0,1,-nbitq), 
to_sfixed(-492153739.0/4294967296.0,1,-nbitq), 
to_sfixed(414718517.0/4294967296.0,1,-nbitq), 
to_sfixed(-302986090.0/4294967296.0,1,-nbitq), 
to_sfixed(231184508.0/4294967296.0,1,-nbitq), 
to_sfixed(442490260.0/4294967296.0,1,-nbitq), 
to_sfixed(387618172.0/4294967296.0,1,-nbitq), 
to_sfixed(97790400.0/4294967296.0,1,-nbitq), 
to_sfixed(127627522.0/4294967296.0,1,-nbitq), 
to_sfixed(-65744478.0/4294967296.0,1,-nbitq), 
to_sfixed(145477131.0/4294967296.0,1,-nbitq), 
to_sfixed(-110399582.0/4294967296.0,1,-nbitq), 
to_sfixed(99026146.0/4294967296.0,1,-nbitq), 
to_sfixed(600660910.0/4294967296.0,1,-nbitq), 
to_sfixed(-351326489.0/4294967296.0,1,-nbitq), 
to_sfixed(222652925.0/4294967296.0,1,-nbitq), 
to_sfixed(-440514993.0/4294967296.0,1,-nbitq), 
to_sfixed(-30140085.0/4294967296.0,1,-nbitq), 
to_sfixed(343415324.0/4294967296.0,1,-nbitq), 
to_sfixed(-226468366.0/4294967296.0,1,-nbitq), 
to_sfixed(-662128140.0/4294967296.0,1,-nbitq), 
to_sfixed(-495293318.0/4294967296.0,1,-nbitq), 
to_sfixed(137878897.0/4294967296.0,1,-nbitq), 
to_sfixed(-54554597.0/4294967296.0,1,-nbitq), 
to_sfixed(265078880.0/4294967296.0,1,-nbitq), 
to_sfixed(-735704772.0/4294967296.0,1,-nbitq), 
to_sfixed(718851002.0/4294967296.0,1,-nbitq), 
to_sfixed(-45634981.0/4294967296.0,1,-nbitq), 
to_sfixed(123737013.0/4294967296.0,1,-nbitq), 
to_sfixed(89660416.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(542523691.0/4294967296.0,1,-nbitq), 
to_sfixed(-426224813.0/4294967296.0,1,-nbitq), 
to_sfixed(553367802.0/4294967296.0,1,-nbitq), 
to_sfixed(549703498.0/4294967296.0,1,-nbitq), 
to_sfixed(-276655894.0/4294967296.0,1,-nbitq), 
to_sfixed(434980790.0/4294967296.0,1,-nbitq), 
to_sfixed(328827380.0/4294967296.0,1,-nbitq), 
to_sfixed(-106438686.0/4294967296.0,1,-nbitq), 
to_sfixed(420793562.0/4294967296.0,1,-nbitq), 
to_sfixed(-254021382.0/4294967296.0,1,-nbitq), 
to_sfixed(537041374.0/4294967296.0,1,-nbitq), 
to_sfixed(-130659301.0/4294967296.0,1,-nbitq), 
to_sfixed(-1273332103.0/4294967296.0,1,-nbitq), 
to_sfixed(-422019778.0/4294967296.0,1,-nbitq), 
to_sfixed(160909991.0/4294967296.0,1,-nbitq), 
to_sfixed(-212618954.0/4294967296.0,1,-nbitq), 
to_sfixed(306910479.0/4294967296.0,1,-nbitq), 
to_sfixed(345256817.0/4294967296.0,1,-nbitq), 
to_sfixed(142829179.0/4294967296.0,1,-nbitq), 
to_sfixed(409876471.0/4294967296.0,1,-nbitq), 
to_sfixed(-167298400.0/4294967296.0,1,-nbitq), 
to_sfixed(-314811230.0/4294967296.0,1,-nbitq), 
to_sfixed(268513740.0/4294967296.0,1,-nbitq), 
to_sfixed(-643832130.0/4294967296.0,1,-nbitq), 
to_sfixed(-4957028.0/4294967296.0,1,-nbitq), 
to_sfixed(4443709.0/4294967296.0,1,-nbitq), 
to_sfixed(220970212.0/4294967296.0,1,-nbitq), 
to_sfixed(-37288724.0/4294967296.0,1,-nbitq), 
to_sfixed(-867421938.0/4294967296.0,1,-nbitq), 
to_sfixed(-262609180.0/4294967296.0,1,-nbitq), 
to_sfixed(269115076.0/4294967296.0,1,-nbitq), 
to_sfixed(-737610112.0/4294967296.0,1,-nbitq), 
to_sfixed(-279522141.0/4294967296.0,1,-nbitq), 
to_sfixed(408709515.0/4294967296.0,1,-nbitq), 
to_sfixed(-6110425.0/4294967296.0,1,-nbitq), 
to_sfixed(-327073959.0/4294967296.0,1,-nbitq), 
to_sfixed(-231106104.0/4294967296.0,1,-nbitq), 
to_sfixed(-44108606.0/4294967296.0,1,-nbitq), 
to_sfixed(-223758749.0/4294967296.0,1,-nbitq), 
to_sfixed(567265319.0/4294967296.0,1,-nbitq), 
to_sfixed(213579804.0/4294967296.0,1,-nbitq), 
to_sfixed(-79663896.0/4294967296.0,1,-nbitq), 
to_sfixed(821473920.0/4294967296.0,1,-nbitq), 
to_sfixed(-893128683.0/4294967296.0,1,-nbitq), 
to_sfixed(151711788.0/4294967296.0,1,-nbitq), 
to_sfixed(39294761.0/4294967296.0,1,-nbitq), 
to_sfixed(269077183.0/4294967296.0,1,-nbitq), 
to_sfixed(821166942.0/4294967296.0,1,-nbitq), 
to_sfixed(140675306.0/4294967296.0,1,-nbitq), 
to_sfixed(-113469267.0/4294967296.0,1,-nbitq), 
to_sfixed(-61417819.0/4294967296.0,1,-nbitq), 
to_sfixed(-31630987.0/4294967296.0,1,-nbitq), 
to_sfixed(208305218.0/4294967296.0,1,-nbitq), 
to_sfixed(-533051482.0/4294967296.0,1,-nbitq), 
to_sfixed(-151460786.0/4294967296.0,1,-nbitq), 
to_sfixed(32312005.0/4294967296.0,1,-nbitq), 
to_sfixed(-225278176.0/4294967296.0,1,-nbitq), 
to_sfixed(-351814277.0/4294967296.0,1,-nbitq), 
to_sfixed(65357251.0/4294967296.0,1,-nbitq), 
to_sfixed(-339765711.0/4294967296.0,1,-nbitq), 
to_sfixed(335019660.0/4294967296.0,1,-nbitq), 
to_sfixed(198633564.0/4294967296.0,1,-nbitq), 
to_sfixed(218753619.0/4294967296.0,1,-nbitq), 
to_sfixed(432000428.0/4294967296.0,1,-nbitq), 
to_sfixed(-85554992.0/4294967296.0,1,-nbitq), 
to_sfixed(-170961458.0/4294967296.0,1,-nbitq), 
to_sfixed(-546767884.0/4294967296.0,1,-nbitq), 
to_sfixed(-201233230.0/4294967296.0,1,-nbitq), 
to_sfixed(-275382247.0/4294967296.0,1,-nbitq), 
to_sfixed(-176291472.0/4294967296.0,1,-nbitq), 
to_sfixed(-657830653.0/4294967296.0,1,-nbitq), 
to_sfixed(-41863384.0/4294967296.0,1,-nbitq), 
to_sfixed(329682611.0/4294967296.0,1,-nbitq), 
to_sfixed(31637612.0/4294967296.0,1,-nbitq), 
to_sfixed(365382645.0/4294967296.0,1,-nbitq), 
to_sfixed(-622166467.0/4294967296.0,1,-nbitq), 
to_sfixed(443030044.0/4294967296.0,1,-nbitq), 
to_sfixed(210037310.0/4294967296.0,1,-nbitq), 
to_sfixed(81367182.0/4294967296.0,1,-nbitq), 
to_sfixed(-176539724.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(559439047.0/4294967296.0,1,-nbitq), 
to_sfixed(-98267406.0/4294967296.0,1,-nbitq), 
to_sfixed(337191092.0/4294967296.0,1,-nbitq), 
to_sfixed(814098895.0/4294967296.0,1,-nbitq), 
to_sfixed(312389129.0/4294967296.0,1,-nbitq), 
to_sfixed(-101890053.0/4294967296.0,1,-nbitq), 
to_sfixed(336270117.0/4294967296.0,1,-nbitq), 
to_sfixed(154779906.0/4294967296.0,1,-nbitq), 
to_sfixed(-190077512.0/4294967296.0,1,-nbitq), 
to_sfixed(379135351.0/4294967296.0,1,-nbitq), 
to_sfixed(515294296.0/4294967296.0,1,-nbitq), 
to_sfixed(-246768507.0/4294967296.0,1,-nbitq), 
to_sfixed(-1309092005.0/4294967296.0,1,-nbitq), 
to_sfixed(-960997670.0/4294967296.0,1,-nbitq), 
to_sfixed(51909784.0/4294967296.0,1,-nbitq), 
to_sfixed(-667220707.0/4294967296.0,1,-nbitq), 
to_sfixed(-172392928.0/4294967296.0,1,-nbitq), 
to_sfixed(373083369.0/4294967296.0,1,-nbitq), 
to_sfixed(470102672.0/4294967296.0,1,-nbitq), 
to_sfixed(283128239.0/4294967296.0,1,-nbitq), 
to_sfixed(-417832384.0/4294967296.0,1,-nbitq), 
to_sfixed(240778105.0/4294967296.0,1,-nbitq), 
to_sfixed(138670672.0/4294967296.0,1,-nbitq), 
to_sfixed(-973017154.0/4294967296.0,1,-nbitq), 
to_sfixed(393837504.0/4294967296.0,1,-nbitq), 
to_sfixed(-149814251.0/4294967296.0,1,-nbitq), 
to_sfixed(-81628765.0/4294967296.0,1,-nbitq), 
to_sfixed(304716903.0/4294967296.0,1,-nbitq), 
to_sfixed(-693103140.0/4294967296.0,1,-nbitq), 
to_sfixed(-1529236766.0/4294967296.0,1,-nbitq), 
to_sfixed(77054482.0/4294967296.0,1,-nbitq), 
to_sfixed(17135776.0/4294967296.0,1,-nbitq), 
to_sfixed(219923196.0/4294967296.0,1,-nbitq), 
to_sfixed(436300720.0/4294967296.0,1,-nbitq), 
to_sfixed(-419301072.0/4294967296.0,1,-nbitq), 
to_sfixed(-518273316.0/4294967296.0,1,-nbitq), 
to_sfixed(421378073.0/4294967296.0,1,-nbitq), 
to_sfixed(47008055.0/4294967296.0,1,-nbitq), 
to_sfixed(-304119452.0/4294967296.0,1,-nbitq), 
to_sfixed(-11019314.0/4294967296.0,1,-nbitq), 
to_sfixed(368219891.0/4294967296.0,1,-nbitq), 
to_sfixed(-165654314.0/4294967296.0,1,-nbitq), 
to_sfixed(578059497.0/4294967296.0,1,-nbitq), 
to_sfixed(-927934563.0/4294967296.0,1,-nbitq), 
to_sfixed(508923339.0/4294967296.0,1,-nbitq), 
to_sfixed(-41560012.0/4294967296.0,1,-nbitq), 
to_sfixed(-140750899.0/4294967296.0,1,-nbitq), 
to_sfixed(1185593063.0/4294967296.0,1,-nbitq), 
to_sfixed(339911322.0/4294967296.0,1,-nbitq), 
to_sfixed(221836523.0/4294967296.0,1,-nbitq), 
to_sfixed(-19688871.0/4294967296.0,1,-nbitq), 
to_sfixed(699044927.0/4294967296.0,1,-nbitq), 
to_sfixed(501571951.0/4294967296.0,1,-nbitq), 
to_sfixed(-206436351.0/4294967296.0,1,-nbitq), 
to_sfixed(-408665701.0/4294967296.0,1,-nbitq), 
to_sfixed(666144620.0/4294967296.0,1,-nbitq), 
to_sfixed(66918040.0/4294967296.0,1,-nbitq), 
to_sfixed(87124924.0/4294967296.0,1,-nbitq), 
to_sfixed(211356830.0/4294967296.0,1,-nbitq), 
to_sfixed(32378974.0/4294967296.0,1,-nbitq), 
to_sfixed(436110088.0/4294967296.0,1,-nbitq), 
to_sfixed(83783223.0/4294967296.0,1,-nbitq), 
to_sfixed(114562759.0/4294967296.0,1,-nbitq), 
to_sfixed(1108572941.0/4294967296.0,1,-nbitq), 
to_sfixed(120083663.0/4294967296.0,1,-nbitq), 
to_sfixed(-114154199.0/4294967296.0,1,-nbitq), 
to_sfixed(-533501350.0/4294967296.0,1,-nbitq), 
to_sfixed(-881423764.0/4294967296.0,1,-nbitq), 
to_sfixed(-68878589.0/4294967296.0,1,-nbitq), 
to_sfixed(-392404624.0/4294967296.0,1,-nbitq), 
to_sfixed(-1552284927.0/4294967296.0,1,-nbitq), 
to_sfixed(130826561.0/4294967296.0,1,-nbitq), 
to_sfixed(196193104.0/4294967296.0,1,-nbitq), 
to_sfixed(172036964.0/4294967296.0,1,-nbitq), 
to_sfixed(414949429.0/4294967296.0,1,-nbitq), 
to_sfixed(-538251791.0/4294967296.0,1,-nbitq), 
to_sfixed(-65955799.0/4294967296.0,1,-nbitq), 
to_sfixed(63956309.0/4294967296.0,1,-nbitq), 
to_sfixed(136670249.0/4294967296.0,1,-nbitq), 
to_sfixed(328876964.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(160060726.0/4294967296.0,1,-nbitq), 
to_sfixed(235067267.0/4294967296.0,1,-nbitq), 
to_sfixed(-83062305.0/4294967296.0,1,-nbitq), 
to_sfixed(933281227.0/4294967296.0,1,-nbitq), 
to_sfixed(230937146.0/4294967296.0,1,-nbitq), 
to_sfixed(367185526.0/4294967296.0,1,-nbitq), 
to_sfixed(219793994.0/4294967296.0,1,-nbitq), 
to_sfixed(-310200102.0/4294967296.0,1,-nbitq), 
to_sfixed(252314209.0/4294967296.0,1,-nbitq), 
to_sfixed(381729262.0/4294967296.0,1,-nbitq), 
to_sfixed(810071921.0/4294967296.0,1,-nbitq), 
to_sfixed(169777241.0/4294967296.0,1,-nbitq), 
to_sfixed(-693086524.0/4294967296.0,1,-nbitq), 
to_sfixed(-857918336.0/4294967296.0,1,-nbitq), 
to_sfixed(194106591.0/4294967296.0,1,-nbitq), 
to_sfixed(-188672674.0/4294967296.0,1,-nbitq), 
to_sfixed(54697737.0/4294967296.0,1,-nbitq), 
to_sfixed(-297279797.0/4294967296.0,1,-nbitq), 
to_sfixed(497811467.0/4294967296.0,1,-nbitq), 
to_sfixed(242269644.0/4294967296.0,1,-nbitq), 
to_sfixed(-287733741.0/4294967296.0,1,-nbitq), 
to_sfixed(-36920247.0/4294967296.0,1,-nbitq), 
to_sfixed(97784753.0/4294967296.0,1,-nbitq), 
to_sfixed(-1179896955.0/4294967296.0,1,-nbitq), 
to_sfixed(332632233.0/4294967296.0,1,-nbitq), 
to_sfixed(-135783060.0/4294967296.0,1,-nbitq), 
to_sfixed(-33548254.0/4294967296.0,1,-nbitq), 
to_sfixed(568672001.0/4294967296.0,1,-nbitq), 
to_sfixed(-711699278.0/4294967296.0,1,-nbitq), 
to_sfixed(-1126911858.0/4294967296.0,1,-nbitq), 
to_sfixed(357123735.0/4294967296.0,1,-nbitq), 
to_sfixed(-155422794.0/4294967296.0,1,-nbitq), 
to_sfixed(-531058232.0/4294967296.0,1,-nbitq), 
to_sfixed(64210372.0/4294967296.0,1,-nbitq), 
to_sfixed(-544207908.0/4294967296.0,1,-nbitq), 
to_sfixed(-415515162.0/4294967296.0,1,-nbitq), 
to_sfixed(108199444.0/4294967296.0,1,-nbitq), 
to_sfixed(-593918168.0/4294967296.0,1,-nbitq), 
to_sfixed(-284529515.0/4294967296.0,1,-nbitq), 
to_sfixed(481218569.0/4294967296.0,1,-nbitq), 
to_sfixed(536741803.0/4294967296.0,1,-nbitq), 
to_sfixed(137525983.0/4294967296.0,1,-nbitq), 
to_sfixed(44136371.0/4294967296.0,1,-nbitq), 
to_sfixed(-1589954889.0/4294967296.0,1,-nbitq), 
to_sfixed(951682114.0/4294967296.0,1,-nbitq), 
to_sfixed(-155767063.0/4294967296.0,1,-nbitq), 
to_sfixed(-12781701.0/4294967296.0,1,-nbitq), 
to_sfixed(1026135991.0/4294967296.0,1,-nbitq), 
to_sfixed(-173109141.0/4294967296.0,1,-nbitq), 
to_sfixed(12571780.0/4294967296.0,1,-nbitq), 
to_sfixed(83842469.0/4294967296.0,1,-nbitq), 
to_sfixed(85040706.0/4294967296.0,1,-nbitq), 
to_sfixed(-54087065.0/4294967296.0,1,-nbitq), 
to_sfixed(-1488018908.0/4294967296.0,1,-nbitq), 
to_sfixed(171180176.0/4294967296.0,1,-nbitq), 
to_sfixed(394213518.0/4294967296.0,1,-nbitq), 
to_sfixed(-110852677.0/4294967296.0,1,-nbitq), 
to_sfixed(-36194038.0/4294967296.0,1,-nbitq), 
to_sfixed(-210282345.0/4294967296.0,1,-nbitq), 
to_sfixed(329696457.0/4294967296.0,1,-nbitq), 
to_sfixed(285575473.0/4294967296.0,1,-nbitq), 
to_sfixed(-319899171.0/4294967296.0,1,-nbitq), 
to_sfixed(994455886.0/4294967296.0,1,-nbitq), 
to_sfixed(296178537.0/4294967296.0,1,-nbitq), 
to_sfixed(15569993.0/4294967296.0,1,-nbitq), 
to_sfixed(158417600.0/4294967296.0,1,-nbitq), 
to_sfixed(-571463543.0/4294967296.0,1,-nbitq), 
to_sfixed(-808406518.0/4294967296.0,1,-nbitq), 
to_sfixed(258706719.0/4294967296.0,1,-nbitq), 
to_sfixed(-395214304.0/4294967296.0,1,-nbitq), 
to_sfixed(-1170460052.0/4294967296.0,1,-nbitq), 
to_sfixed(-236105338.0/4294967296.0,1,-nbitq), 
to_sfixed(483231127.0/4294967296.0,1,-nbitq), 
to_sfixed(-288847222.0/4294967296.0,1,-nbitq), 
to_sfixed(169347012.0/4294967296.0,1,-nbitq), 
to_sfixed(-630025285.0/4294967296.0,1,-nbitq), 
to_sfixed(540347805.0/4294967296.0,1,-nbitq), 
to_sfixed(-30380800.0/4294967296.0,1,-nbitq), 
to_sfixed(149489787.0/4294967296.0,1,-nbitq), 
to_sfixed(135512806.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-138207290.0/4294967296.0,1,-nbitq), 
to_sfixed(-471500312.0/4294967296.0,1,-nbitq), 
to_sfixed(1004118186.0/4294967296.0,1,-nbitq), 
to_sfixed(660969227.0/4294967296.0,1,-nbitq), 
to_sfixed(761488834.0/4294967296.0,1,-nbitq), 
to_sfixed(110011723.0/4294967296.0,1,-nbitq), 
to_sfixed(2639902.0/4294967296.0,1,-nbitq), 
to_sfixed(-574274988.0/4294967296.0,1,-nbitq), 
to_sfixed(739088053.0/4294967296.0,1,-nbitq), 
to_sfixed(-304882755.0/4294967296.0,1,-nbitq), 
to_sfixed(1387307396.0/4294967296.0,1,-nbitq), 
to_sfixed(347829113.0/4294967296.0,1,-nbitq), 
to_sfixed(-789814222.0/4294967296.0,1,-nbitq), 
to_sfixed(-1040547225.0/4294967296.0,1,-nbitq), 
to_sfixed(24703934.0/4294967296.0,1,-nbitq), 
to_sfixed(-647212403.0/4294967296.0,1,-nbitq), 
to_sfixed(-106156155.0/4294967296.0,1,-nbitq), 
to_sfixed(140687365.0/4294967296.0,1,-nbitq), 
to_sfixed(432329845.0/4294967296.0,1,-nbitq), 
to_sfixed(671279343.0/4294967296.0,1,-nbitq), 
to_sfixed(-362267553.0/4294967296.0,1,-nbitq), 
to_sfixed(551999349.0/4294967296.0,1,-nbitq), 
to_sfixed(110625121.0/4294967296.0,1,-nbitq), 
to_sfixed(-930568509.0/4294967296.0,1,-nbitq), 
to_sfixed(-284487253.0/4294967296.0,1,-nbitq), 
to_sfixed(-192952924.0/4294967296.0,1,-nbitq), 
to_sfixed(-172594644.0/4294967296.0,1,-nbitq), 
to_sfixed(38562147.0/4294967296.0,1,-nbitq), 
to_sfixed(-709729845.0/4294967296.0,1,-nbitq), 
to_sfixed(-718280366.0/4294967296.0,1,-nbitq), 
to_sfixed(642303839.0/4294967296.0,1,-nbitq), 
to_sfixed(-166628699.0/4294967296.0,1,-nbitq), 
to_sfixed(-582317302.0/4294967296.0,1,-nbitq), 
to_sfixed(341104997.0/4294967296.0,1,-nbitq), 
to_sfixed(-359545966.0/4294967296.0,1,-nbitq), 
to_sfixed(98580795.0/4294967296.0,1,-nbitq), 
to_sfixed(-412763994.0/4294967296.0,1,-nbitq), 
to_sfixed(-246383403.0/4294967296.0,1,-nbitq), 
to_sfixed(-359075128.0/4294967296.0,1,-nbitq), 
to_sfixed(757145912.0/4294967296.0,1,-nbitq), 
to_sfixed(-84719624.0/4294967296.0,1,-nbitq), 
to_sfixed(-91502054.0/4294967296.0,1,-nbitq), 
to_sfixed(119738739.0/4294967296.0,1,-nbitq), 
to_sfixed(-1975226834.0/4294967296.0,1,-nbitq), 
to_sfixed(-74716021.0/4294967296.0,1,-nbitq), 
to_sfixed(430694424.0/4294967296.0,1,-nbitq), 
to_sfixed(-119270621.0/4294967296.0,1,-nbitq), 
to_sfixed(1006042374.0/4294967296.0,1,-nbitq), 
to_sfixed(-143439871.0/4294967296.0,1,-nbitq), 
to_sfixed(256553537.0/4294967296.0,1,-nbitq), 
to_sfixed(308621004.0/4294967296.0,1,-nbitq), 
to_sfixed(918311036.0/4294967296.0,1,-nbitq), 
to_sfixed(-2912413.0/4294967296.0,1,-nbitq), 
to_sfixed(-1421933993.0/4294967296.0,1,-nbitq), 
to_sfixed(-150486029.0/4294967296.0,1,-nbitq), 
to_sfixed(34964632.0/4294967296.0,1,-nbitq), 
to_sfixed(-383807600.0/4294967296.0,1,-nbitq), 
to_sfixed(592906844.0/4294967296.0,1,-nbitq), 
to_sfixed(-328850320.0/4294967296.0,1,-nbitq), 
to_sfixed(213141324.0/4294967296.0,1,-nbitq), 
to_sfixed(-161673023.0/4294967296.0,1,-nbitq), 
to_sfixed(-565349415.0/4294967296.0,1,-nbitq), 
to_sfixed(1021863013.0/4294967296.0,1,-nbitq), 
to_sfixed(433784337.0/4294967296.0,1,-nbitq), 
to_sfixed(-506083902.0/4294967296.0,1,-nbitq), 
to_sfixed(77587133.0/4294967296.0,1,-nbitq), 
to_sfixed(-748934582.0/4294967296.0,1,-nbitq), 
to_sfixed(-1550485946.0/4294967296.0,1,-nbitq), 
to_sfixed(131688351.0/4294967296.0,1,-nbitq), 
to_sfixed(-560759028.0/4294967296.0,1,-nbitq), 
to_sfixed(-981244445.0/4294967296.0,1,-nbitq), 
to_sfixed(-274237453.0/4294967296.0,1,-nbitq), 
to_sfixed(-29694541.0/4294967296.0,1,-nbitq), 
to_sfixed(-43145013.0/4294967296.0,1,-nbitq), 
to_sfixed(-37038457.0/4294967296.0,1,-nbitq), 
to_sfixed(-765224580.0/4294967296.0,1,-nbitq), 
to_sfixed(848993138.0/4294967296.0,1,-nbitq), 
to_sfixed(22268448.0/4294967296.0,1,-nbitq), 
to_sfixed(226445020.0/4294967296.0,1,-nbitq), 
to_sfixed(-165316336.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(78947520.0/4294967296.0,1,-nbitq), 
to_sfixed(-482192540.0/4294967296.0,1,-nbitq), 
to_sfixed(1326403885.0/4294967296.0,1,-nbitq), 
to_sfixed(363092304.0/4294967296.0,1,-nbitq), 
to_sfixed(140730813.0/4294967296.0,1,-nbitq), 
to_sfixed(52259842.0/4294967296.0,1,-nbitq), 
to_sfixed(-384640809.0/4294967296.0,1,-nbitq), 
to_sfixed(-786825297.0/4294967296.0,1,-nbitq), 
to_sfixed(928150130.0/4294967296.0,1,-nbitq), 
to_sfixed(-39770704.0/4294967296.0,1,-nbitq), 
to_sfixed(1021027900.0/4294967296.0,1,-nbitq), 
to_sfixed(-339110614.0/4294967296.0,1,-nbitq), 
to_sfixed(-552407173.0/4294967296.0,1,-nbitq), 
to_sfixed(-501196025.0/4294967296.0,1,-nbitq), 
to_sfixed(-99069353.0/4294967296.0,1,-nbitq), 
to_sfixed(-613459731.0/4294967296.0,1,-nbitq), 
to_sfixed(-566381.0/4294967296.0,1,-nbitq), 
to_sfixed(-185588764.0/4294967296.0,1,-nbitq), 
to_sfixed(457976453.0/4294967296.0,1,-nbitq), 
to_sfixed(325537603.0/4294967296.0,1,-nbitq), 
to_sfixed(189804410.0/4294967296.0,1,-nbitq), 
to_sfixed(204582141.0/4294967296.0,1,-nbitq), 
to_sfixed(86031104.0/4294967296.0,1,-nbitq), 
to_sfixed(-612137763.0/4294967296.0,1,-nbitq), 
to_sfixed(242433406.0/4294967296.0,1,-nbitq), 
to_sfixed(-688892148.0/4294967296.0,1,-nbitq), 
to_sfixed(-434809175.0/4294967296.0,1,-nbitq), 
to_sfixed(512069408.0/4294967296.0,1,-nbitq), 
to_sfixed(-948776687.0/4294967296.0,1,-nbitq), 
to_sfixed(-1081023650.0/4294967296.0,1,-nbitq), 
to_sfixed(217948836.0/4294967296.0,1,-nbitq), 
to_sfixed(449833247.0/4294967296.0,1,-nbitq), 
to_sfixed(104376991.0/4294967296.0,1,-nbitq), 
to_sfixed(173470469.0/4294967296.0,1,-nbitq), 
to_sfixed(-230745771.0/4294967296.0,1,-nbitq), 
to_sfixed(-62235680.0/4294967296.0,1,-nbitq), 
to_sfixed(-338366820.0/4294967296.0,1,-nbitq), 
to_sfixed(-235121344.0/4294967296.0,1,-nbitq), 
to_sfixed(-642205251.0/4294967296.0,1,-nbitq), 
to_sfixed(654455528.0/4294967296.0,1,-nbitq), 
to_sfixed(75397123.0/4294967296.0,1,-nbitq), 
to_sfixed(302767815.0/4294967296.0,1,-nbitq), 
to_sfixed(193037547.0/4294967296.0,1,-nbitq), 
to_sfixed(-1792523875.0/4294967296.0,1,-nbitq), 
to_sfixed(58230701.0/4294967296.0,1,-nbitq), 
to_sfixed(703716360.0/4294967296.0,1,-nbitq), 
to_sfixed(-235858498.0/4294967296.0,1,-nbitq), 
to_sfixed(662600288.0/4294967296.0,1,-nbitq), 
to_sfixed(-537004715.0/4294967296.0,1,-nbitq), 
to_sfixed(202643107.0/4294967296.0,1,-nbitq), 
to_sfixed(482896165.0/4294967296.0,1,-nbitq), 
to_sfixed(828082501.0/4294967296.0,1,-nbitq), 
to_sfixed(318673945.0/4294967296.0,1,-nbitq), 
to_sfixed(-1293375428.0/4294967296.0,1,-nbitq), 
to_sfixed(-141157149.0/4294967296.0,1,-nbitq), 
to_sfixed(86357289.0/4294967296.0,1,-nbitq), 
to_sfixed(-144601386.0/4294967296.0,1,-nbitq), 
to_sfixed(446100786.0/4294967296.0,1,-nbitq), 
to_sfixed(308946058.0/4294967296.0,1,-nbitq), 
to_sfixed(-276677276.0/4294967296.0,1,-nbitq), 
to_sfixed(117032752.0/4294967296.0,1,-nbitq), 
to_sfixed(-705681929.0/4294967296.0,1,-nbitq), 
to_sfixed(1028706119.0/4294967296.0,1,-nbitq), 
to_sfixed(111783197.0/4294967296.0,1,-nbitq), 
to_sfixed(-113460436.0/4294967296.0,1,-nbitq), 
to_sfixed(136171409.0/4294967296.0,1,-nbitq), 
to_sfixed(-555742112.0/4294967296.0,1,-nbitq), 
to_sfixed(-1989876256.0/4294967296.0,1,-nbitq), 
to_sfixed(-295209701.0/4294967296.0,1,-nbitq), 
to_sfixed(-847909044.0/4294967296.0,1,-nbitq), 
to_sfixed(-1337125498.0/4294967296.0,1,-nbitq), 
to_sfixed(175282750.0/4294967296.0,1,-nbitq), 
to_sfixed(462009509.0/4294967296.0,1,-nbitq), 
to_sfixed(-347360761.0/4294967296.0,1,-nbitq), 
to_sfixed(226839261.0/4294967296.0,1,-nbitq), 
to_sfixed(-410133940.0/4294967296.0,1,-nbitq), 
to_sfixed(1518075713.0/4294967296.0,1,-nbitq), 
to_sfixed(331144791.0/4294967296.0,1,-nbitq), 
to_sfixed(107340435.0/4294967296.0,1,-nbitq), 
to_sfixed(-331224303.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-151284700.0/4294967296.0,1,-nbitq), 
to_sfixed(-100297437.0/4294967296.0,1,-nbitq), 
to_sfixed(388173568.0/4294967296.0,1,-nbitq), 
to_sfixed(533603594.0/4294967296.0,1,-nbitq), 
to_sfixed(735067597.0/4294967296.0,1,-nbitq), 
to_sfixed(-308842123.0/4294967296.0,1,-nbitq), 
to_sfixed(-100884558.0/4294967296.0,1,-nbitq), 
to_sfixed(-430364225.0/4294967296.0,1,-nbitq), 
to_sfixed(961833145.0/4294967296.0,1,-nbitq), 
to_sfixed(331077891.0/4294967296.0,1,-nbitq), 
to_sfixed(1125723984.0/4294967296.0,1,-nbitq), 
to_sfixed(-96711337.0/4294967296.0,1,-nbitq), 
to_sfixed(-666786165.0/4294967296.0,1,-nbitq), 
to_sfixed(-217741576.0/4294967296.0,1,-nbitq), 
to_sfixed(-366359618.0/4294967296.0,1,-nbitq), 
to_sfixed(-76171600.0/4294967296.0,1,-nbitq), 
to_sfixed(111426498.0/4294967296.0,1,-nbitq), 
to_sfixed(51778385.0/4294967296.0,1,-nbitq), 
to_sfixed(640588464.0/4294967296.0,1,-nbitq), 
to_sfixed(284829938.0/4294967296.0,1,-nbitq), 
to_sfixed(270049940.0/4294967296.0,1,-nbitq), 
to_sfixed(103040167.0/4294967296.0,1,-nbitq), 
to_sfixed(547895330.0/4294967296.0,1,-nbitq), 
to_sfixed(-861859981.0/4294967296.0,1,-nbitq), 
to_sfixed(408110129.0/4294967296.0,1,-nbitq), 
to_sfixed(-528548721.0/4294967296.0,1,-nbitq), 
to_sfixed(-137070581.0/4294967296.0,1,-nbitq), 
to_sfixed(-244878703.0/4294967296.0,1,-nbitq), 
to_sfixed(-704963211.0/4294967296.0,1,-nbitq), 
to_sfixed(-1056276913.0/4294967296.0,1,-nbitq), 
to_sfixed(323686339.0/4294967296.0,1,-nbitq), 
to_sfixed(754478536.0/4294967296.0,1,-nbitq), 
to_sfixed(198920466.0/4294967296.0,1,-nbitq), 
to_sfixed(346627497.0/4294967296.0,1,-nbitq), 
to_sfixed(-284489654.0/4294967296.0,1,-nbitq), 
to_sfixed(228945755.0/4294967296.0,1,-nbitq), 
to_sfixed(-109715919.0/4294967296.0,1,-nbitq), 
to_sfixed(-691710831.0/4294967296.0,1,-nbitq), 
to_sfixed(-97955903.0/4294967296.0,1,-nbitq), 
to_sfixed(18259494.0/4294967296.0,1,-nbitq), 
to_sfixed(415304479.0/4294967296.0,1,-nbitq), 
to_sfixed(279559373.0/4294967296.0,1,-nbitq), 
to_sfixed(148509205.0/4294967296.0,1,-nbitq), 
to_sfixed(-602473357.0/4294967296.0,1,-nbitq), 
to_sfixed(-34228517.0/4294967296.0,1,-nbitq), 
to_sfixed(557299465.0/4294967296.0,1,-nbitq), 
to_sfixed(-201831324.0/4294967296.0,1,-nbitq), 
to_sfixed(478788435.0/4294967296.0,1,-nbitq), 
to_sfixed(-60607379.0/4294967296.0,1,-nbitq), 
to_sfixed(115910192.0/4294967296.0,1,-nbitq), 
to_sfixed(-299405915.0/4294967296.0,1,-nbitq), 
to_sfixed(230072870.0/4294967296.0,1,-nbitq), 
to_sfixed(-32029171.0/4294967296.0,1,-nbitq), 
to_sfixed(-752234621.0/4294967296.0,1,-nbitq), 
to_sfixed(-680115594.0/4294967296.0,1,-nbitq), 
to_sfixed(-152776848.0/4294967296.0,1,-nbitq), 
to_sfixed(261135080.0/4294967296.0,1,-nbitq), 
to_sfixed(-167940355.0/4294967296.0,1,-nbitq), 
to_sfixed(-195138816.0/4294967296.0,1,-nbitq), 
to_sfixed(329568759.0/4294967296.0,1,-nbitq), 
to_sfixed(-456812691.0/4294967296.0,1,-nbitq), 
to_sfixed(163722934.0/4294967296.0,1,-nbitq), 
to_sfixed(962885077.0/4294967296.0,1,-nbitq), 
to_sfixed(-23005086.0/4294967296.0,1,-nbitq), 
to_sfixed(-47551662.0/4294967296.0,1,-nbitq), 
to_sfixed(-409808904.0/4294967296.0,1,-nbitq), 
to_sfixed(4143015.0/4294967296.0,1,-nbitq), 
to_sfixed(-1153030705.0/4294967296.0,1,-nbitq), 
to_sfixed(57466295.0/4294967296.0,1,-nbitq), 
to_sfixed(-373132680.0/4294967296.0,1,-nbitq), 
to_sfixed(-454195713.0/4294967296.0,1,-nbitq), 
to_sfixed(-509963.0/4294967296.0,1,-nbitq), 
to_sfixed(660967893.0/4294967296.0,1,-nbitq), 
to_sfixed(16507769.0/4294967296.0,1,-nbitq), 
to_sfixed(50834104.0/4294967296.0,1,-nbitq), 
to_sfixed(432351859.0/4294967296.0,1,-nbitq), 
to_sfixed(1652602389.0/4294967296.0,1,-nbitq), 
to_sfixed(-101940880.0/4294967296.0,1,-nbitq), 
to_sfixed(317658106.0/4294967296.0,1,-nbitq), 
to_sfixed(355792113.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-8960609.0/4294967296.0,1,-nbitq), 
to_sfixed(334606743.0/4294967296.0,1,-nbitq), 
to_sfixed(744530538.0/4294967296.0,1,-nbitq), 
to_sfixed(93824404.0/4294967296.0,1,-nbitq), 
to_sfixed(1142931525.0/4294967296.0,1,-nbitq), 
to_sfixed(-982609874.0/4294967296.0,1,-nbitq), 
to_sfixed(-281713984.0/4294967296.0,1,-nbitq), 
to_sfixed(-825380286.0/4294967296.0,1,-nbitq), 
to_sfixed(1189855864.0/4294967296.0,1,-nbitq), 
to_sfixed(-277834501.0/4294967296.0,1,-nbitq), 
to_sfixed(-87253095.0/4294967296.0,1,-nbitq), 
to_sfixed(-206277114.0/4294967296.0,1,-nbitq), 
to_sfixed(-500135466.0/4294967296.0,1,-nbitq), 
to_sfixed(-303644435.0/4294967296.0,1,-nbitq), 
to_sfixed(173913226.0/4294967296.0,1,-nbitq), 
to_sfixed(-56970382.0/4294967296.0,1,-nbitq), 
to_sfixed(-69113656.0/4294967296.0,1,-nbitq), 
to_sfixed(81879187.0/4294967296.0,1,-nbitq), 
to_sfixed(353446338.0/4294967296.0,1,-nbitq), 
to_sfixed(114195921.0/4294967296.0,1,-nbitq), 
to_sfixed(260099552.0/4294967296.0,1,-nbitq), 
to_sfixed(741115390.0/4294967296.0,1,-nbitq), 
to_sfixed(384433160.0/4294967296.0,1,-nbitq), 
to_sfixed(-989188318.0/4294967296.0,1,-nbitq), 
to_sfixed(285615873.0/4294967296.0,1,-nbitq), 
to_sfixed(-371013361.0/4294967296.0,1,-nbitq), 
to_sfixed(-7515777.0/4294967296.0,1,-nbitq), 
to_sfixed(-145172658.0/4294967296.0,1,-nbitq), 
to_sfixed(-442432336.0/4294967296.0,1,-nbitq), 
to_sfixed(-512171902.0/4294967296.0,1,-nbitq), 
to_sfixed(564366956.0/4294967296.0,1,-nbitq), 
to_sfixed(671325703.0/4294967296.0,1,-nbitq), 
to_sfixed(-143185746.0/4294967296.0,1,-nbitq), 
to_sfixed(504546254.0/4294967296.0,1,-nbitq), 
to_sfixed(74737284.0/4294967296.0,1,-nbitq), 
to_sfixed(554500168.0/4294967296.0,1,-nbitq), 
to_sfixed(170984267.0/4294967296.0,1,-nbitq), 
to_sfixed(-7280089.0/4294967296.0,1,-nbitq), 
to_sfixed(-168354390.0/4294967296.0,1,-nbitq), 
to_sfixed(582419764.0/4294967296.0,1,-nbitq), 
to_sfixed(-271545230.0/4294967296.0,1,-nbitq), 
to_sfixed(356845035.0/4294967296.0,1,-nbitq), 
to_sfixed(304928729.0/4294967296.0,1,-nbitq), 
to_sfixed(50036365.0/4294967296.0,1,-nbitq), 
to_sfixed(200802517.0/4294967296.0,1,-nbitq), 
to_sfixed(892847190.0/4294967296.0,1,-nbitq), 
to_sfixed(-362268389.0/4294967296.0,1,-nbitq), 
to_sfixed(339908482.0/4294967296.0,1,-nbitq), 
to_sfixed(-76532865.0/4294967296.0,1,-nbitq), 
to_sfixed(-54789926.0/4294967296.0,1,-nbitq), 
to_sfixed(294336561.0/4294967296.0,1,-nbitq), 
to_sfixed(-157445630.0/4294967296.0,1,-nbitq), 
to_sfixed(421849530.0/4294967296.0,1,-nbitq), 
to_sfixed(270644234.0/4294967296.0,1,-nbitq), 
to_sfixed(-506254958.0/4294967296.0,1,-nbitq), 
to_sfixed(-536923618.0/4294967296.0,1,-nbitq), 
to_sfixed(219071065.0/4294967296.0,1,-nbitq), 
to_sfixed(-289786669.0/4294967296.0,1,-nbitq), 
to_sfixed(-119294929.0/4294967296.0,1,-nbitq), 
to_sfixed(108176249.0/4294967296.0,1,-nbitq), 
to_sfixed(168209092.0/4294967296.0,1,-nbitq), 
to_sfixed(154303191.0/4294967296.0,1,-nbitq), 
to_sfixed(774647249.0/4294967296.0,1,-nbitq), 
to_sfixed(-547254809.0/4294967296.0,1,-nbitq), 
to_sfixed(-257596202.0/4294967296.0,1,-nbitq), 
to_sfixed(164677668.0/4294967296.0,1,-nbitq), 
to_sfixed(172386847.0/4294967296.0,1,-nbitq), 
to_sfixed(-820068623.0/4294967296.0,1,-nbitq), 
to_sfixed(226031011.0/4294967296.0,1,-nbitq), 
to_sfixed(-391642603.0/4294967296.0,1,-nbitq), 
to_sfixed(-159055051.0/4294967296.0,1,-nbitq), 
to_sfixed(5617289.0/4294967296.0,1,-nbitq), 
to_sfixed(478487114.0/4294967296.0,1,-nbitq), 
to_sfixed(-29106418.0/4294967296.0,1,-nbitq), 
to_sfixed(223761602.0/4294967296.0,1,-nbitq), 
to_sfixed(72404155.0/4294967296.0,1,-nbitq), 
to_sfixed(930381933.0/4294967296.0,1,-nbitq), 
to_sfixed(-4923823.0/4294967296.0,1,-nbitq), 
to_sfixed(-292263230.0/4294967296.0,1,-nbitq), 
to_sfixed(-190552232.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(10754251.0/4294967296.0,1,-nbitq), 
to_sfixed(70531751.0/4294967296.0,1,-nbitq), 
to_sfixed(1011659721.0/4294967296.0,1,-nbitq), 
to_sfixed(-215894920.0/4294967296.0,1,-nbitq), 
to_sfixed(383884315.0/4294967296.0,1,-nbitq), 
to_sfixed(-1563007621.0/4294967296.0,1,-nbitq), 
to_sfixed(-337386089.0/4294967296.0,1,-nbitq), 
to_sfixed(-1078689610.0/4294967296.0,1,-nbitq), 
to_sfixed(597072093.0/4294967296.0,1,-nbitq), 
to_sfixed(307817570.0/4294967296.0,1,-nbitq), 
to_sfixed(-714201759.0/4294967296.0,1,-nbitq), 
to_sfixed(-679868160.0/4294967296.0,1,-nbitq), 
to_sfixed(256461324.0/4294967296.0,1,-nbitq), 
to_sfixed(-539799751.0/4294967296.0,1,-nbitq), 
to_sfixed(-263497571.0/4294967296.0,1,-nbitq), 
to_sfixed(361384547.0/4294967296.0,1,-nbitq), 
to_sfixed(120530102.0/4294967296.0,1,-nbitq), 
to_sfixed(16325284.0/4294967296.0,1,-nbitq), 
to_sfixed(392842389.0/4294967296.0,1,-nbitq), 
to_sfixed(-21227366.0/4294967296.0,1,-nbitq), 
to_sfixed(352337716.0/4294967296.0,1,-nbitq), 
to_sfixed(287353828.0/4294967296.0,1,-nbitq), 
to_sfixed(39397693.0/4294967296.0,1,-nbitq), 
to_sfixed(-753205901.0/4294967296.0,1,-nbitq), 
to_sfixed(394178200.0/4294967296.0,1,-nbitq), 
to_sfixed(-285318286.0/4294967296.0,1,-nbitq), 
to_sfixed(-197055105.0/4294967296.0,1,-nbitq), 
to_sfixed(408680455.0/4294967296.0,1,-nbitq), 
to_sfixed(-159494372.0/4294967296.0,1,-nbitq), 
to_sfixed(-241950896.0/4294967296.0,1,-nbitq), 
to_sfixed(64607284.0/4294967296.0,1,-nbitq), 
to_sfixed(458630258.0/4294967296.0,1,-nbitq), 
to_sfixed(411764468.0/4294967296.0,1,-nbitq), 
to_sfixed(132012825.0/4294967296.0,1,-nbitq), 
to_sfixed(-214746774.0/4294967296.0,1,-nbitq), 
to_sfixed(-384081013.0/4294967296.0,1,-nbitq), 
to_sfixed(474652278.0/4294967296.0,1,-nbitq), 
to_sfixed(-268186743.0/4294967296.0,1,-nbitq), 
to_sfixed(-18898036.0/4294967296.0,1,-nbitq), 
to_sfixed(16617275.0/4294967296.0,1,-nbitq), 
to_sfixed(-300369683.0/4294967296.0,1,-nbitq), 
to_sfixed(-396920555.0/4294967296.0,1,-nbitq), 
to_sfixed(415524442.0/4294967296.0,1,-nbitq), 
to_sfixed(-411944779.0/4294967296.0,1,-nbitq), 
to_sfixed(303318158.0/4294967296.0,1,-nbitq), 
to_sfixed(430421049.0/4294967296.0,1,-nbitq), 
to_sfixed(-225962318.0/4294967296.0,1,-nbitq), 
to_sfixed(152310612.0/4294967296.0,1,-nbitq), 
to_sfixed(118974044.0/4294967296.0,1,-nbitq), 
to_sfixed(-51821876.0/4294967296.0,1,-nbitq), 
to_sfixed(-81982318.0/4294967296.0,1,-nbitq), 
to_sfixed(185790070.0/4294967296.0,1,-nbitq), 
to_sfixed(237385913.0/4294967296.0,1,-nbitq), 
to_sfixed(-661376457.0/4294967296.0,1,-nbitq), 
to_sfixed(-248247474.0/4294967296.0,1,-nbitq), 
to_sfixed(-534129770.0/4294967296.0,1,-nbitq), 
to_sfixed(255231265.0/4294967296.0,1,-nbitq), 
to_sfixed(86238302.0/4294967296.0,1,-nbitq), 
to_sfixed(-128873566.0/4294967296.0,1,-nbitq), 
to_sfixed(47498117.0/4294967296.0,1,-nbitq), 
to_sfixed(-262726182.0/4294967296.0,1,-nbitq), 
to_sfixed(412087385.0/4294967296.0,1,-nbitq), 
to_sfixed(952170974.0/4294967296.0,1,-nbitq), 
to_sfixed(-76269450.0/4294967296.0,1,-nbitq), 
to_sfixed(59519245.0/4294967296.0,1,-nbitq), 
to_sfixed(-84759940.0/4294967296.0,1,-nbitq), 
to_sfixed(-290395697.0/4294967296.0,1,-nbitq), 
to_sfixed(-30002584.0/4294967296.0,1,-nbitq), 
to_sfixed(82976471.0/4294967296.0,1,-nbitq), 
to_sfixed(982574.0/4294967296.0,1,-nbitq), 
to_sfixed(116634565.0/4294967296.0,1,-nbitq), 
to_sfixed(66067376.0/4294967296.0,1,-nbitq), 
to_sfixed(889353127.0/4294967296.0,1,-nbitq), 
to_sfixed(57169803.0/4294967296.0,1,-nbitq), 
to_sfixed(-194072085.0/4294967296.0,1,-nbitq), 
to_sfixed(-117484824.0/4294967296.0,1,-nbitq), 
to_sfixed(1014667929.0/4294967296.0,1,-nbitq), 
to_sfixed(164194019.0/4294967296.0,1,-nbitq), 
to_sfixed(-489931035.0/4294967296.0,1,-nbitq), 
to_sfixed(-125067014.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(299968620.0/4294967296.0,1,-nbitq), 
to_sfixed(-307965122.0/4294967296.0,1,-nbitq), 
to_sfixed(494449924.0/4294967296.0,1,-nbitq), 
to_sfixed(-79095124.0/4294967296.0,1,-nbitq), 
to_sfixed(176595766.0/4294967296.0,1,-nbitq), 
to_sfixed(-1390431114.0/4294967296.0,1,-nbitq), 
to_sfixed(-441461184.0/4294967296.0,1,-nbitq), 
to_sfixed(-504580630.0/4294967296.0,1,-nbitq), 
to_sfixed(688089349.0/4294967296.0,1,-nbitq), 
to_sfixed(65158006.0/4294967296.0,1,-nbitq), 
to_sfixed(-274239811.0/4294967296.0,1,-nbitq), 
to_sfixed(212634798.0/4294967296.0,1,-nbitq), 
to_sfixed(-89677147.0/4294967296.0,1,-nbitq), 
to_sfixed(-68274478.0/4294967296.0,1,-nbitq), 
to_sfixed(-94334023.0/4294967296.0,1,-nbitq), 
to_sfixed(530615.0/4294967296.0,1,-nbitq), 
to_sfixed(-136348281.0/4294967296.0,1,-nbitq), 
to_sfixed(-223420863.0/4294967296.0,1,-nbitq), 
to_sfixed(570108783.0/4294967296.0,1,-nbitq), 
to_sfixed(312877161.0/4294967296.0,1,-nbitq), 
to_sfixed(315463750.0/4294967296.0,1,-nbitq), 
to_sfixed(221302181.0/4294967296.0,1,-nbitq), 
to_sfixed(800130067.0/4294967296.0,1,-nbitq), 
to_sfixed(-225092635.0/4294967296.0,1,-nbitq), 
to_sfixed(-242332463.0/4294967296.0,1,-nbitq), 
to_sfixed(395918271.0/4294967296.0,1,-nbitq), 
to_sfixed(-388160425.0/4294967296.0,1,-nbitq), 
to_sfixed(-298397164.0/4294967296.0,1,-nbitq), 
to_sfixed(-167204268.0/4294967296.0,1,-nbitq), 
to_sfixed(-331752819.0/4294967296.0,1,-nbitq), 
to_sfixed(-218401382.0/4294967296.0,1,-nbitq), 
to_sfixed(132789659.0/4294967296.0,1,-nbitq), 
to_sfixed(-335185415.0/4294967296.0,1,-nbitq), 
to_sfixed(61958797.0/4294967296.0,1,-nbitq), 
to_sfixed(-12579700.0/4294967296.0,1,-nbitq), 
to_sfixed(-159378589.0/4294967296.0,1,-nbitq), 
to_sfixed(171249337.0/4294967296.0,1,-nbitq), 
to_sfixed(-998946666.0/4294967296.0,1,-nbitq), 
to_sfixed(-228192731.0/4294967296.0,1,-nbitq), 
to_sfixed(691010600.0/4294967296.0,1,-nbitq), 
to_sfixed(-452584693.0/4294967296.0,1,-nbitq), 
to_sfixed(90674567.0/4294967296.0,1,-nbitq), 
to_sfixed(798379603.0/4294967296.0,1,-nbitq), 
to_sfixed(-12957815.0/4294967296.0,1,-nbitq), 
to_sfixed(240534238.0/4294967296.0,1,-nbitq), 
to_sfixed(6119774.0/4294967296.0,1,-nbitq), 
to_sfixed(17142594.0/4294967296.0,1,-nbitq), 
to_sfixed(106134029.0/4294967296.0,1,-nbitq), 
to_sfixed(-16324961.0/4294967296.0,1,-nbitq), 
to_sfixed(-287542719.0/4294967296.0,1,-nbitq), 
to_sfixed(-167542256.0/4294967296.0,1,-nbitq), 
to_sfixed(621956323.0/4294967296.0,1,-nbitq), 
to_sfixed(88939526.0/4294967296.0,1,-nbitq), 
to_sfixed(-134655227.0/4294967296.0,1,-nbitq), 
to_sfixed(-132938468.0/4294967296.0,1,-nbitq), 
to_sfixed(-461859272.0/4294967296.0,1,-nbitq), 
to_sfixed(-268252793.0/4294967296.0,1,-nbitq), 
to_sfixed(392336720.0/4294967296.0,1,-nbitq), 
to_sfixed(183281254.0/4294967296.0,1,-nbitq), 
to_sfixed(-18963270.0/4294967296.0,1,-nbitq), 
to_sfixed(-27731754.0/4294967296.0,1,-nbitq), 
to_sfixed(-10280195.0/4294967296.0,1,-nbitq), 
to_sfixed(722330593.0/4294967296.0,1,-nbitq), 
to_sfixed(-160457610.0/4294967296.0,1,-nbitq), 
to_sfixed(-371217033.0/4294967296.0,1,-nbitq), 
to_sfixed(-220104184.0/4294967296.0,1,-nbitq), 
to_sfixed(-522050855.0/4294967296.0,1,-nbitq), 
to_sfixed(-240346193.0/4294967296.0,1,-nbitq), 
to_sfixed(18482347.0/4294967296.0,1,-nbitq), 
to_sfixed(-182769798.0/4294967296.0,1,-nbitq), 
to_sfixed(212882238.0/4294967296.0,1,-nbitq), 
to_sfixed(142973832.0/4294967296.0,1,-nbitq), 
to_sfixed(92044530.0/4294967296.0,1,-nbitq), 
to_sfixed(-170412196.0/4294967296.0,1,-nbitq), 
to_sfixed(396207512.0/4294967296.0,1,-nbitq), 
to_sfixed(263234318.0/4294967296.0,1,-nbitq), 
to_sfixed(981610808.0/4294967296.0,1,-nbitq), 
to_sfixed(114041888.0/4294967296.0,1,-nbitq), 
to_sfixed(-321753189.0/4294967296.0,1,-nbitq), 
to_sfixed(218262327.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-124193036.0/4294967296.0,1,-nbitq), 
to_sfixed(-175595319.0/4294967296.0,1,-nbitq), 
to_sfixed(728919215.0/4294967296.0,1,-nbitq), 
to_sfixed(-72013966.0/4294967296.0,1,-nbitq), 
to_sfixed(-49740256.0/4294967296.0,1,-nbitq), 
to_sfixed(-1425375122.0/4294967296.0,1,-nbitq), 
to_sfixed(-14556744.0/4294967296.0,1,-nbitq), 
to_sfixed(-7156308.0/4294967296.0,1,-nbitq), 
to_sfixed(1123663143.0/4294967296.0,1,-nbitq), 
to_sfixed(215111881.0/4294967296.0,1,-nbitq), 
to_sfixed(-145086218.0/4294967296.0,1,-nbitq), 
to_sfixed(282318965.0/4294967296.0,1,-nbitq), 
to_sfixed(-899856310.0/4294967296.0,1,-nbitq), 
to_sfixed(236440463.0/4294967296.0,1,-nbitq), 
to_sfixed(250681120.0/4294967296.0,1,-nbitq), 
to_sfixed(628562081.0/4294967296.0,1,-nbitq), 
to_sfixed(341915225.0/4294967296.0,1,-nbitq), 
to_sfixed(-141891518.0/4294967296.0,1,-nbitq), 
to_sfixed(244467484.0/4294967296.0,1,-nbitq), 
to_sfixed(293147596.0/4294967296.0,1,-nbitq), 
to_sfixed(-365886558.0/4294967296.0,1,-nbitq), 
to_sfixed(12103187.0/4294967296.0,1,-nbitq), 
to_sfixed(333084935.0/4294967296.0,1,-nbitq), 
to_sfixed(-507981931.0/4294967296.0,1,-nbitq), 
to_sfixed(397112233.0/4294967296.0,1,-nbitq), 
to_sfixed(-52025051.0/4294967296.0,1,-nbitq), 
to_sfixed(67245468.0/4294967296.0,1,-nbitq), 
to_sfixed(83696417.0/4294967296.0,1,-nbitq), 
to_sfixed(-246307109.0/4294967296.0,1,-nbitq), 
to_sfixed(-1141931081.0/4294967296.0,1,-nbitq), 
to_sfixed(-93965778.0/4294967296.0,1,-nbitq), 
to_sfixed(258431693.0/4294967296.0,1,-nbitq), 
to_sfixed(-332099661.0/4294967296.0,1,-nbitq), 
to_sfixed(444264089.0/4294967296.0,1,-nbitq), 
to_sfixed(-33489795.0/4294967296.0,1,-nbitq), 
to_sfixed(-322367315.0/4294967296.0,1,-nbitq), 
to_sfixed(-23333469.0/4294967296.0,1,-nbitq), 
to_sfixed(-871642768.0/4294967296.0,1,-nbitq), 
to_sfixed(68628493.0/4294967296.0,1,-nbitq), 
to_sfixed(531180439.0/4294967296.0,1,-nbitq), 
to_sfixed(234423351.0/4294967296.0,1,-nbitq), 
to_sfixed(255676674.0/4294967296.0,1,-nbitq), 
to_sfixed(346772444.0/4294967296.0,1,-nbitq), 
to_sfixed(253745049.0/4294967296.0,1,-nbitq), 
to_sfixed(96551530.0/4294967296.0,1,-nbitq), 
to_sfixed(678886557.0/4294967296.0,1,-nbitq), 
to_sfixed(-322587293.0/4294967296.0,1,-nbitq), 
to_sfixed(448802499.0/4294967296.0,1,-nbitq), 
to_sfixed(157748741.0/4294967296.0,1,-nbitq), 
to_sfixed(-671833001.0/4294967296.0,1,-nbitq), 
to_sfixed(-313405998.0/4294967296.0,1,-nbitq), 
to_sfixed(549994341.0/4294967296.0,1,-nbitq), 
to_sfixed(-379876049.0/4294967296.0,1,-nbitq), 
to_sfixed(356677068.0/4294967296.0,1,-nbitq), 
to_sfixed(13668140.0/4294967296.0,1,-nbitq), 
to_sfixed(-12920124.0/4294967296.0,1,-nbitq), 
to_sfixed(-358140005.0/4294967296.0,1,-nbitq), 
to_sfixed(233876417.0/4294967296.0,1,-nbitq), 
to_sfixed(325837771.0/4294967296.0,1,-nbitq), 
to_sfixed(109597951.0/4294967296.0,1,-nbitq), 
to_sfixed(41057535.0/4294967296.0,1,-nbitq), 
to_sfixed(224744798.0/4294967296.0,1,-nbitq), 
to_sfixed(603495448.0/4294967296.0,1,-nbitq), 
to_sfixed(322856553.0/4294967296.0,1,-nbitq), 
to_sfixed(168673800.0/4294967296.0,1,-nbitq), 
to_sfixed(-168153110.0/4294967296.0,1,-nbitq), 
to_sfixed(-775162524.0/4294967296.0,1,-nbitq), 
to_sfixed(-124401622.0/4294967296.0,1,-nbitq), 
to_sfixed(174647007.0/4294967296.0,1,-nbitq), 
to_sfixed(-434726638.0/4294967296.0,1,-nbitq), 
to_sfixed(264687524.0/4294967296.0,1,-nbitq), 
to_sfixed(503652032.0/4294967296.0,1,-nbitq), 
to_sfixed(-30493074.0/4294967296.0,1,-nbitq), 
to_sfixed(86561596.0/4294967296.0,1,-nbitq), 
to_sfixed(328912417.0/4294967296.0,1,-nbitq), 
to_sfixed(202678563.0/4294967296.0,1,-nbitq), 
to_sfixed(1248023213.0/4294967296.0,1,-nbitq), 
to_sfixed(-97877050.0/4294967296.0,1,-nbitq), 
to_sfixed(-160115521.0/4294967296.0,1,-nbitq), 
to_sfixed(152777391.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(654879957.0/4294967296.0,1,-nbitq), 
to_sfixed(-301158420.0/4294967296.0,1,-nbitq), 
to_sfixed(417238932.0/4294967296.0,1,-nbitq), 
to_sfixed(678816538.0/4294967296.0,1,-nbitq), 
to_sfixed(313861161.0/4294967296.0,1,-nbitq), 
to_sfixed(-956214480.0/4294967296.0,1,-nbitq), 
to_sfixed(-53259545.0/4294967296.0,1,-nbitq), 
to_sfixed(-111541337.0/4294967296.0,1,-nbitq), 
to_sfixed(403185950.0/4294967296.0,1,-nbitq), 
to_sfixed(407793541.0/4294967296.0,1,-nbitq), 
to_sfixed(-425837832.0/4294967296.0,1,-nbitq), 
to_sfixed(-516203089.0/4294967296.0,1,-nbitq), 
to_sfixed(-701652993.0/4294967296.0,1,-nbitq), 
to_sfixed(240284527.0/4294967296.0,1,-nbitq), 
to_sfixed(-336458189.0/4294967296.0,1,-nbitq), 
to_sfixed(371186263.0/4294967296.0,1,-nbitq), 
to_sfixed(-343855547.0/4294967296.0,1,-nbitq), 
to_sfixed(-291488783.0/4294967296.0,1,-nbitq), 
to_sfixed(-634644535.0/4294967296.0,1,-nbitq), 
to_sfixed(201549860.0/4294967296.0,1,-nbitq), 
to_sfixed(-178421299.0/4294967296.0,1,-nbitq), 
to_sfixed(68833143.0/4294967296.0,1,-nbitq), 
to_sfixed(-42253951.0/4294967296.0,1,-nbitq), 
to_sfixed(-134048930.0/4294967296.0,1,-nbitq), 
to_sfixed(82519156.0/4294967296.0,1,-nbitq), 
to_sfixed(146147839.0/4294967296.0,1,-nbitq), 
to_sfixed(433442818.0/4294967296.0,1,-nbitq), 
to_sfixed(-492009724.0/4294967296.0,1,-nbitq), 
to_sfixed(290852665.0/4294967296.0,1,-nbitq), 
to_sfixed(-530643400.0/4294967296.0,1,-nbitq), 
to_sfixed(-16898839.0/4294967296.0,1,-nbitq), 
to_sfixed(324956905.0/4294967296.0,1,-nbitq), 
to_sfixed(107904634.0/4294967296.0,1,-nbitq), 
to_sfixed(399203821.0/4294967296.0,1,-nbitq), 
to_sfixed(319871512.0/4294967296.0,1,-nbitq), 
to_sfixed(310141778.0/4294967296.0,1,-nbitq), 
to_sfixed(528899657.0/4294967296.0,1,-nbitq), 
to_sfixed(-243819930.0/4294967296.0,1,-nbitq), 
to_sfixed(-299945743.0/4294967296.0,1,-nbitq), 
to_sfixed(531643124.0/4294967296.0,1,-nbitq), 
to_sfixed(-126650433.0/4294967296.0,1,-nbitq), 
to_sfixed(865642021.0/4294967296.0,1,-nbitq), 
to_sfixed(1025855513.0/4294967296.0,1,-nbitq), 
to_sfixed(1007301815.0/4294967296.0,1,-nbitq), 
to_sfixed(-313299998.0/4294967296.0,1,-nbitq), 
to_sfixed(780603645.0/4294967296.0,1,-nbitq), 
to_sfixed(94818646.0/4294967296.0,1,-nbitq), 
to_sfixed(-455325660.0/4294967296.0,1,-nbitq), 
to_sfixed(83389832.0/4294967296.0,1,-nbitq), 
to_sfixed(-788044927.0/4294967296.0,1,-nbitq), 
to_sfixed(-257762352.0/4294967296.0,1,-nbitq), 
to_sfixed(484443640.0/4294967296.0,1,-nbitq), 
to_sfixed(-294543922.0/4294967296.0,1,-nbitq), 
to_sfixed(103571726.0/4294967296.0,1,-nbitq), 
to_sfixed(-433571210.0/4294967296.0,1,-nbitq), 
to_sfixed(-413562461.0/4294967296.0,1,-nbitq), 
to_sfixed(-500291907.0/4294967296.0,1,-nbitq), 
to_sfixed(704205131.0/4294967296.0,1,-nbitq), 
to_sfixed(65698218.0/4294967296.0,1,-nbitq), 
to_sfixed(15316661.0/4294967296.0,1,-nbitq), 
to_sfixed(-79149981.0/4294967296.0,1,-nbitq), 
to_sfixed(402876142.0/4294967296.0,1,-nbitq), 
to_sfixed(259127296.0/4294967296.0,1,-nbitq), 
to_sfixed(779328065.0/4294967296.0,1,-nbitq), 
to_sfixed(-168332375.0/4294967296.0,1,-nbitq), 
to_sfixed(409231906.0/4294967296.0,1,-nbitq), 
to_sfixed(-601915413.0/4294967296.0,1,-nbitq), 
to_sfixed(-257545785.0/4294967296.0,1,-nbitq), 
to_sfixed(149079304.0/4294967296.0,1,-nbitq), 
to_sfixed(-845963423.0/4294967296.0,1,-nbitq), 
to_sfixed(461745497.0/4294967296.0,1,-nbitq), 
to_sfixed(227358794.0/4294967296.0,1,-nbitq), 
to_sfixed(-570485046.0/4294967296.0,1,-nbitq), 
to_sfixed(-239091783.0/4294967296.0,1,-nbitq), 
to_sfixed(17515296.0/4294967296.0,1,-nbitq), 
to_sfixed(168431888.0/4294967296.0,1,-nbitq), 
to_sfixed(1299215416.0/4294967296.0,1,-nbitq), 
to_sfixed(488034037.0/4294967296.0,1,-nbitq), 
to_sfixed(441478377.0/4294967296.0,1,-nbitq), 
to_sfixed(-67607458.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-220682609.0/4294967296.0,1,-nbitq), 
to_sfixed(-558841008.0/4294967296.0,1,-nbitq), 
to_sfixed(66419374.0/4294967296.0,1,-nbitq), 
to_sfixed(-38261089.0/4294967296.0,1,-nbitq), 
to_sfixed(82341290.0/4294967296.0,1,-nbitq), 
to_sfixed(-628591789.0/4294967296.0,1,-nbitq), 
to_sfixed(11110706.0/4294967296.0,1,-nbitq), 
to_sfixed(-519078101.0/4294967296.0,1,-nbitq), 
to_sfixed(138216768.0/4294967296.0,1,-nbitq), 
to_sfixed(-303390108.0/4294967296.0,1,-nbitq), 
to_sfixed(-523418209.0/4294967296.0,1,-nbitq), 
to_sfixed(-756503771.0/4294967296.0,1,-nbitq), 
to_sfixed(-578091691.0/4294967296.0,1,-nbitq), 
to_sfixed(254168938.0/4294967296.0,1,-nbitq), 
to_sfixed(100938796.0/4294967296.0,1,-nbitq), 
to_sfixed(161623395.0/4294967296.0,1,-nbitq), 
to_sfixed(390807043.0/4294967296.0,1,-nbitq), 
to_sfixed(-285035507.0/4294967296.0,1,-nbitq), 
to_sfixed(-304211630.0/4294967296.0,1,-nbitq), 
to_sfixed(-375791312.0/4294967296.0,1,-nbitq), 
to_sfixed(185853496.0/4294967296.0,1,-nbitq), 
to_sfixed(-168151042.0/4294967296.0,1,-nbitq), 
to_sfixed(287789366.0/4294967296.0,1,-nbitq), 
to_sfixed(-358035721.0/4294967296.0,1,-nbitq), 
to_sfixed(-229203744.0/4294967296.0,1,-nbitq), 
to_sfixed(23269549.0/4294967296.0,1,-nbitq), 
to_sfixed(86074854.0/4294967296.0,1,-nbitq), 
to_sfixed(-641352321.0/4294967296.0,1,-nbitq), 
to_sfixed(-27297054.0/4294967296.0,1,-nbitq), 
to_sfixed(-536907589.0/4294967296.0,1,-nbitq), 
to_sfixed(-822567941.0/4294967296.0,1,-nbitq), 
to_sfixed(-91273124.0/4294967296.0,1,-nbitq), 
to_sfixed(-185528799.0/4294967296.0,1,-nbitq), 
to_sfixed(-160547558.0/4294967296.0,1,-nbitq), 
to_sfixed(705859980.0/4294967296.0,1,-nbitq), 
to_sfixed(314471675.0/4294967296.0,1,-nbitq), 
to_sfixed(189090175.0/4294967296.0,1,-nbitq), 
to_sfixed(221499734.0/4294967296.0,1,-nbitq), 
to_sfixed(72419576.0/4294967296.0,1,-nbitq), 
to_sfixed(685956369.0/4294967296.0,1,-nbitq), 
to_sfixed(-527619121.0/4294967296.0,1,-nbitq), 
to_sfixed(791896753.0/4294967296.0,1,-nbitq), 
to_sfixed(408017844.0/4294967296.0,1,-nbitq), 
to_sfixed(1176964747.0/4294967296.0,1,-nbitq), 
to_sfixed(-60857549.0/4294967296.0,1,-nbitq), 
to_sfixed(195111845.0/4294967296.0,1,-nbitq), 
to_sfixed(-109030075.0/4294967296.0,1,-nbitq), 
to_sfixed(-680543515.0/4294967296.0,1,-nbitq), 
to_sfixed(668058.0/4294967296.0,1,-nbitq), 
to_sfixed(-55236196.0/4294967296.0,1,-nbitq), 
to_sfixed(210517332.0/4294967296.0,1,-nbitq), 
to_sfixed(271099010.0/4294967296.0,1,-nbitq), 
to_sfixed(-264891432.0/4294967296.0,1,-nbitq), 
to_sfixed(61236560.0/4294967296.0,1,-nbitq), 
to_sfixed(283680758.0/4294967296.0,1,-nbitq), 
to_sfixed(255845715.0/4294967296.0,1,-nbitq), 
to_sfixed(-753450954.0/4294967296.0,1,-nbitq), 
to_sfixed(352766676.0/4294967296.0,1,-nbitq), 
to_sfixed(369291109.0/4294967296.0,1,-nbitq), 
to_sfixed(325268286.0/4294967296.0,1,-nbitq), 
to_sfixed(-390578812.0/4294967296.0,1,-nbitq), 
to_sfixed(322672422.0/4294967296.0,1,-nbitq), 
to_sfixed(388938030.0/4294967296.0,1,-nbitq), 
to_sfixed(787034755.0/4294967296.0,1,-nbitq), 
to_sfixed(309021665.0/4294967296.0,1,-nbitq), 
to_sfixed(-364128379.0/4294967296.0,1,-nbitq), 
to_sfixed(-115420359.0/4294967296.0,1,-nbitq), 
to_sfixed(-193586329.0/4294967296.0,1,-nbitq), 
to_sfixed(51737054.0/4294967296.0,1,-nbitq), 
to_sfixed(12881153.0/4294967296.0,1,-nbitq), 
to_sfixed(970304169.0/4294967296.0,1,-nbitq), 
to_sfixed(214721924.0/4294967296.0,1,-nbitq), 
to_sfixed(-582213392.0/4294967296.0,1,-nbitq), 
to_sfixed(81291383.0/4294967296.0,1,-nbitq), 
to_sfixed(172097023.0/4294967296.0,1,-nbitq), 
to_sfixed(355646921.0/4294967296.0,1,-nbitq), 
to_sfixed(547150360.0/4294967296.0,1,-nbitq), 
to_sfixed(65327959.0/4294967296.0,1,-nbitq), 
to_sfixed(56483892.0/4294967296.0,1,-nbitq), 
to_sfixed(400241787.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-327778949.0/4294967296.0,1,-nbitq), 
to_sfixed(-312481496.0/4294967296.0,1,-nbitq), 
to_sfixed(427550928.0/4294967296.0,1,-nbitq), 
to_sfixed(-132471031.0/4294967296.0,1,-nbitq), 
to_sfixed(692720843.0/4294967296.0,1,-nbitq), 
to_sfixed(231041968.0/4294967296.0,1,-nbitq), 
to_sfixed(264579858.0/4294967296.0,1,-nbitq), 
to_sfixed(-530762488.0/4294967296.0,1,-nbitq), 
to_sfixed(176508211.0/4294967296.0,1,-nbitq), 
to_sfixed(-377600143.0/4294967296.0,1,-nbitq), 
to_sfixed(147879169.0/4294967296.0,1,-nbitq), 
to_sfixed(-749294344.0/4294967296.0,1,-nbitq), 
to_sfixed(-387224648.0/4294967296.0,1,-nbitq), 
to_sfixed(753016572.0/4294967296.0,1,-nbitq), 
to_sfixed(54839214.0/4294967296.0,1,-nbitq), 
to_sfixed(-482482718.0/4294967296.0,1,-nbitq), 
to_sfixed(-242468393.0/4294967296.0,1,-nbitq), 
to_sfixed(229788099.0/4294967296.0,1,-nbitq), 
to_sfixed(227167006.0/4294967296.0,1,-nbitq), 
to_sfixed(222327977.0/4294967296.0,1,-nbitq), 
to_sfixed(-189012788.0/4294967296.0,1,-nbitq), 
to_sfixed(556272424.0/4294967296.0,1,-nbitq), 
to_sfixed(-15993244.0/4294967296.0,1,-nbitq), 
to_sfixed(239248892.0/4294967296.0,1,-nbitq), 
to_sfixed(39211258.0/4294967296.0,1,-nbitq), 
to_sfixed(723542521.0/4294967296.0,1,-nbitq), 
to_sfixed(-119553078.0/4294967296.0,1,-nbitq), 
to_sfixed(-41440210.0/4294967296.0,1,-nbitq), 
to_sfixed(532202776.0/4294967296.0,1,-nbitq), 
to_sfixed(209705322.0/4294967296.0,1,-nbitq), 
to_sfixed(-1026031268.0/4294967296.0,1,-nbitq), 
to_sfixed(363246630.0/4294967296.0,1,-nbitq), 
to_sfixed(192827401.0/4294967296.0,1,-nbitq), 
to_sfixed(-54339191.0/4294967296.0,1,-nbitq), 
to_sfixed(905542506.0/4294967296.0,1,-nbitq), 
to_sfixed(-94629871.0/4294967296.0,1,-nbitq), 
to_sfixed(810891.0/4294967296.0,1,-nbitq), 
to_sfixed(533803681.0/4294967296.0,1,-nbitq), 
to_sfixed(-54705929.0/4294967296.0,1,-nbitq), 
to_sfixed(581701669.0/4294967296.0,1,-nbitq), 
to_sfixed(-381531188.0/4294967296.0,1,-nbitq), 
to_sfixed(538623693.0/4294967296.0,1,-nbitq), 
to_sfixed(423821212.0/4294967296.0,1,-nbitq), 
to_sfixed(326970935.0/4294967296.0,1,-nbitq), 
to_sfixed(331231132.0/4294967296.0,1,-nbitq), 
to_sfixed(-112318137.0/4294967296.0,1,-nbitq), 
to_sfixed(42569317.0/4294967296.0,1,-nbitq), 
to_sfixed(-59323880.0/4294967296.0,1,-nbitq), 
to_sfixed(-182474797.0/4294967296.0,1,-nbitq), 
to_sfixed(-186142496.0/4294967296.0,1,-nbitq), 
to_sfixed(-88933176.0/4294967296.0,1,-nbitq), 
to_sfixed(-652027681.0/4294967296.0,1,-nbitq), 
to_sfixed(-663457228.0/4294967296.0,1,-nbitq), 
to_sfixed(372390246.0/4294967296.0,1,-nbitq), 
to_sfixed(427827664.0/4294967296.0,1,-nbitq), 
to_sfixed(169676800.0/4294967296.0,1,-nbitq), 
to_sfixed(68840786.0/4294967296.0,1,-nbitq), 
to_sfixed(-174592989.0/4294967296.0,1,-nbitq), 
to_sfixed(-51201558.0/4294967296.0,1,-nbitq), 
to_sfixed(28832604.0/4294967296.0,1,-nbitq), 
to_sfixed(225277512.0/4294967296.0,1,-nbitq), 
to_sfixed(-189030198.0/4294967296.0,1,-nbitq), 
to_sfixed(-165487491.0/4294967296.0,1,-nbitq), 
to_sfixed(54929254.0/4294967296.0,1,-nbitq), 
to_sfixed(86275003.0/4294967296.0,1,-nbitq), 
to_sfixed(-417425993.0/4294967296.0,1,-nbitq), 
to_sfixed(-414376481.0/4294967296.0,1,-nbitq), 
to_sfixed(-264405282.0/4294967296.0,1,-nbitq), 
to_sfixed(226647172.0/4294967296.0,1,-nbitq), 
to_sfixed(87239672.0/4294967296.0,1,-nbitq), 
to_sfixed(738199492.0/4294967296.0,1,-nbitq), 
to_sfixed(346703603.0/4294967296.0,1,-nbitq), 
to_sfixed(-884365453.0/4294967296.0,1,-nbitq), 
to_sfixed(-109219646.0/4294967296.0,1,-nbitq), 
to_sfixed(372255124.0/4294967296.0,1,-nbitq), 
to_sfixed(-93698261.0/4294967296.0,1,-nbitq), 
to_sfixed(123762783.0/4294967296.0,1,-nbitq), 
to_sfixed(257044594.0/4294967296.0,1,-nbitq), 
to_sfixed(-368904335.0/4294967296.0,1,-nbitq), 
to_sfixed(345543555.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(370336220.0/4294967296.0,1,-nbitq), 
to_sfixed(-541481381.0/4294967296.0,1,-nbitq), 
to_sfixed(-174454169.0/4294967296.0,1,-nbitq), 
to_sfixed(72751166.0/4294967296.0,1,-nbitq), 
to_sfixed(388409960.0/4294967296.0,1,-nbitq), 
to_sfixed(382611754.0/4294967296.0,1,-nbitq), 
to_sfixed(17001197.0/4294967296.0,1,-nbitq), 
to_sfixed(-598156927.0/4294967296.0,1,-nbitq), 
to_sfixed(-54223197.0/4294967296.0,1,-nbitq), 
to_sfixed(-256848669.0/4294967296.0,1,-nbitq), 
to_sfixed(131092414.0/4294967296.0,1,-nbitq), 
to_sfixed(-649332085.0/4294967296.0,1,-nbitq), 
to_sfixed(466621881.0/4294967296.0,1,-nbitq), 
to_sfixed(178861948.0/4294967296.0,1,-nbitq), 
to_sfixed(165406395.0/4294967296.0,1,-nbitq), 
to_sfixed(-553100119.0/4294967296.0,1,-nbitq), 
to_sfixed(293159842.0/4294967296.0,1,-nbitq), 
to_sfixed(-302035770.0/4294967296.0,1,-nbitq), 
to_sfixed(163893438.0/4294967296.0,1,-nbitq), 
to_sfixed(-92857623.0/4294967296.0,1,-nbitq), 
to_sfixed(69264020.0/4294967296.0,1,-nbitq), 
to_sfixed(595836384.0/4294967296.0,1,-nbitq), 
to_sfixed(-88148618.0/4294967296.0,1,-nbitq), 
to_sfixed(-30899095.0/4294967296.0,1,-nbitq), 
to_sfixed(-316337544.0/4294967296.0,1,-nbitq), 
to_sfixed(562251829.0/4294967296.0,1,-nbitq), 
to_sfixed(43835742.0/4294967296.0,1,-nbitq), 
to_sfixed(-409253469.0/4294967296.0,1,-nbitq), 
to_sfixed(-102014318.0/4294967296.0,1,-nbitq), 
to_sfixed(-275640400.0/4294967296.0,1,-nbitq), 
to_sfixed(-83342605.0/4294967296.0,1,-nbitq), 
to_sfixed(-283940418.0/4294967296.0,1,-nbitq), 
to_sfixed(4800280.0/4294967296.0,1,-nbitq), 
to_sfixed(-434042801.0/4294967296.0,1,-nbitq), 
to_sfixed(508099509.0/4294967296.0,1,-nbitq), 
to_sfixed(40198523.0/4294967296.0,1,-nbitq), 
to_sfixed(-208575743.0/4294967296.0,1,-nbitq), 
to_sfixed(-343287652.0/4294967296.0,1,-nbitq), 
to_sfixed(-10167379.0/4294967296.0,1,-nbitq), 
to_sfixed(447846087.0/4294967296.0,1,-nbitq), 
to_sfixed(63176731.0/4294967296.0,1,-nbitq), 
to_sfixed(552458519.0/4294967296.0,1,-nbitq), 
to_sfixed(43377949.0/4294967296.0,1,-nbitq), 
to_sfixed(370260062.0/4294967296.0,1,-nbitq), 
to_sfixed(453547707.0/4294967296.0,1,-nbitq), 
to_sfixed(831348635.0/4294967296.0,1,-nbitq), 
to_sfixed(70192198.0/4294967296.0,1,-nbitq), 
to_sfixed(37634360.0/4294967296.0,1,-nbitq), 
to_sfixed(407792614.0/4294967296.0,1,-nbitq), 
to_sfixed(258830423.0/4294967296.0,1,-nbitq), 
to_sfixed(-400875041.0/4294967296.0,1,-nbitq), 
to_sfixed(-606687113.0/4294967296.0,1,-nbitq), 
to_sfixed(24724691.0/4294967296.0,1,-nbitq), 
to_sfixed(-367205415.0/4294967296.0,1,-nbitq), 
to_sfixed(-97757844.0/4294967296.0,1,-nbitq), 
to_sfixed(-120438193.0/4294967296.0,1,-nbitq), 
to_sfixed(-360899607.0/4294967296.0,1,-nbitq), 
to_sfixed(-123331558.0/4294967296.0,1,-nbitq), 
to_sfixed(222907167.0/4294967296.0,1,-nbitq), 
to_sfixed(-307196728.0/4294967296.0,1,-nbitq), 
to_sfixed(104598831.0/4294967296.0,1,-nbitq), 
to_sfixed(38627047.0/4294967296.0,1,-nbitq), 
to_sfixed(75808255.0/4294967296.0,1,-nbitq), 
to_sfixed(-11563393.0/4294967296.0,1,-nbitq), 
to_sfixed(379512806.0/4294967296.0,1,-nbitq), 
to_sfixed(111722361.0/4294967296.0,1,-nbitq), 
to_sfixed(-87981854.0/4294967296.0,1,-nbitq), 
to_sfixed(-399922883.0/4294967296.0,1,-nbitq), 
to_sfixed(418531707.0/4294967296.0,1,-nbitq), 
to_sfixed(74510935.0/4294967296.0,1,-nbitq), 
to_sfixed(391046647.0/4294967296.0,1,-nbitq), 
to_sfixed(443181655.0/4294967296.0,1,-nbitq), 
to_sfixed(-146438867.0/4294967296.0,1,-nbitq), 
to_sfixed(-307582514.0/4294967296.0,1,-nbitq), 
to_sfixed(-128441690.0/4294967296.0,1,-nbitq), 
to_sfixed(-130927643.0/4294967296.0,1,-nbitq), 
to_sfixed(-44957148.0/4294967296.0,1,-nbitq), 
to_sfixed(151295560.0/4294967296.0,1,-nbitq), 
to_sfixed(86181453.0/4294967296.0,1,-nbitq), 
to_sfixed(-80899774.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-96728059.0/4294967296.0,1,-nbitq), 
to_sfixed(-629385474.0/4294967296.0,1,-nbitq), 
to_sfixed(396370290.0/4294967296.0,1,-nbitq), 
to_sfixed(-38934640.0/4294967296.0,1,-nbitq), 
to_sfixed(332066666.0/4294967296.0,1,-nbitq), 
to_sfixed(-403237559.0/4294967296.0,1,-nbitq), 
to_sfixed(169588208.0/4294967296.0,1,-nbitq), 
to_sfixed(-444669955.0/4294967296.0,1,-nbitq), 
to_sfixed(275349149.0/4294967296.0,1,-nbitq), 
to_sfixed(-265715446.0/4294967296.0,1,-nbitq), 
to_sfixed(-124300356.0/4294967296.0,1,-nbitq), 
to_sfixed(48244997.0/4294967296.0,1,-nbitq), 
to_sfixed(-191471377.0/4294967296.0,1,-nbitq), 
to_sfixed(180220450.0/4294967296.0,1,-nbitq), 
to_sfixed(-67302345.0/4294967296.0,1,-nbitq), 
to_sfixed(-808399198.0/4294967296.0,1,-nbitq), 
to_sfixed(-10502830.0/4294967296.0,1,-nbitq), 
to_sfixed(132067078.0/4294967296.0,1,-nbitq), 
to_sfixed(84037672.0/4294967296.0,1,-nbitq), 
to_sfixed(-275585796.0/4294967296.0,1,-nbitq), 
to_sfixed(-338523252.0/4294967296.0,1,-nbitq), 
to_sfixed(185135459.0/4294967296.0,1,-nbitq), 
to_sfixed(-93541900.0/4294967296.0,1,-nbitq), 
to_sfixed(378136051.0/4294967296.0,1,-nbitq), 
to_sfixed(-228539331.0/4294967296.0,1,-nbitq), 
to_sfixed(68898518.0/4294967296.0,1,-nbitq), 
to_sfixed(287007379.0/4294967296.0,1,-nbitq), 
to_sfixed(63496148.0/4294967296.0,1,-nbitq), 
to_sfixed(213592104.0/4294967296.0,1,-nbitq), 
to_sfixed(129484723.0/4294967296.0,1,-nbitq), 
to_sfixed(-250451176.0/4294967296.0,1,-nbitq), 
to_sfixed(41921865.0/4294967296.0,1,-nbitq), 
to_sfixed(600966470.0/4294967296.0,1,-nbitq), 
to_sfixed(268488560.0/4294967296.0,1,-nbitq), 
to_sfixed(560827458.0/4294967296.0,1,-nbitq), 
to_sfixed(-169046436.0/4294967296.0,1,-nbitq), 
to_sfixed(20724422.0/4294967296.0,1,-nbitq), 
to_sfixed(-323211917.0/4294967296.0,1,-nbitq), 
to_sfixed(216774184.0/4294967296.0,1,-nbitq), 
to_sfixed(-135098001.0/4294967296.0,1,-nbitq), 
to_sfixed(502000847.0/4294967296.0,1,-nbitq), 
to_sfixed(-257073341.0/4294967296.0,1,-nbitq), 
to_sfixed(317048869.0/4294967296.0,1,-nbitq), 
to_sfixed(268625114.0/4294967296.0,1,-nbitq), 
to_sfixed(280307099.0/4294967296.0,1,-nbitq), 
to_sfixed(464634205.0/4294967296.0,1,-nbitq), 
to_sfixed(-424974974.0/4294967296.0,1,-nbitq), 
to_sfixed(-267845804.0/4294967296.0,1,-nbitq), 
to_sfixed(-372259169.0/4294967296.0,1,-nbitq), 
to_sfixed(-20646588.0/4294967296.0,1,-nbitq), 
to_sfixed(-420411625.0/4294967296.0,1,-nbitq), 
to_sfixed(-9778578.0/4294967296.0,1,-nbitq), 
to_sfixed(214404905.0/4294967296.0,1,-nbitq), 
to_sfixed(198233392.0/4294967296.0,1,-nbitq), 
to_sfixed(-131659719.0/4294967296.0,1,-nbitq), 
to_sfixed(-626863560.0/4294967296.0,1,-nbitq), 
to_sfixed(-236652890.0/4294967296.0,1,-nbitq), 
to_sfixed(-144882073.0/4294967296.0,1,-nbitq), 
to_sfixed(1111051.0/4294967296.0,1,-nbitq), 
to_sfixed(-8673044.0/4294967296.0,1,-nbitq), 
to_sfixed(-320405501.0/4294967296.0,1,-nbitq), 
to_sfixed(-339069268.0/4294967296.0,1,-nbitq), 
to_sfixed(63440339.0/4294967296.0,1,-nbitq), 
to_sfixed(119430632.0/4294967296.0,1,-nbitq), 
to_sfixed(-25575955.0/4294967296.0,1,-nbitq), 
to_sfixed(-374884133.0/4294967296.0,1,-nbitq), 
to_sfixed(-221393601.0/4294967296.0,1,-nbitq), 
to_sfixed(-371462149.0/4294967296.0,1,-nbitq), 
to_sfixed(373040869.0/4294967296.0,1,-nbitq), 
to_sfixed(327306978.0/4294967296.0,1,-nbitq), 
to_sfixed(86434069.0/4294967296.0,1,-nbitq), 
to_sfixed(904813.0/4294967296.0,1,-nbitq), 
to_sfixed(65693381.0/4294967296.0,1,-nbitq), 
to_sfixed(-101146580.0/4294967296.0,1,-nbitq), 
to_sfixed(173186688.0/4294967296.0,1,-nbitq), 
to_sfixed(-458535226.0/4294967296.0,1,-nbitq), 
to_sfixed(258987247.0/4294967296.0,1,-nbitq), 
to_sfixed(305307941.0/4294967296.0,1,-nbitq), 
to_sfixed(332069653.0/4294967296.0,1,-nbitq), 
to_sfixed(-21246893.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(91365154.0/4294967296.0,1,-nbitq), 
to_sfixed(38086349.0/4294967296.0,1,-nbitq), 
to_sfixed(596077355.0/4294967296.0,1,-nbitq), 
to_sfixed(-412409743.0/4294967296.0,1,-nbitq), 
to_sfixed(41875.0/4294967296.0,1,-nbitq), 
to_sfixed(-55072818.0/4294967296.0,1,-nbitq), 
to_sfixed(35515374.0/4294967296.0,1,-nbitq), 
to_sfixed(-30394407.0/4294967296.0,1,-nbitq), 
to_sfixed(100017807.0/4294967296.0,1,-nbitq), 
to_sfixed(-81898501.0/4294967296.0,1,-nbitq), 
to_sfixed(-413351774.0/4294967296.0,1,-nbitq), 
to_sfixed(438232875.0/4294967296.0,1,-nbitq), 
to_sfixed(-56085304.0/4294967296.0,1,-nbitq), 
to_sfixed(-314218731.0/4294967296.0,1,-nbitq), 
to_sfixed(260937132.0/4294967296.0,1,-nbitq), 
to_sfixed(-610106000.0/4294967296.0,1,-nbitq), 
to_sfixed(383861819.0/4294967296.0,1,-nbitq), 
to_sfixed(311844918.0/4294967296.0,1,-nbitq), 
to_sfixed(286591061.0/4294967296.0,1,-nbitq), 
to_sfixed(-209685986.0/4294967296.0,1,-nbitq), 
to_sfixed(75546254.0/4294967296.0,1,-nbitq), 
to_sfixed(76819375.0/4294967296.0,1,-nbitq), 
to_sfixed(260837738.0/4294967296.0,1,-nbitq), 
to_sfixed(278744305.0/4294967296.0,1,-nbitq), 
to_sfixed(384560969.0/4294967296.0,1,-nbitq), 
to_sfixed(283423656.0/4294967296.0,1,-nbitq), 
to_sfixed(-78085345.0/4294967296.0,1,-nbitq), 
to_sfixed(-595002783.0/4294967296.0,1,-nbitq), 
to_sfixed(73418414.0/4294967296.0,1,-nbitq), 
to_sfixed(-280165246.0/4294967296.0,1,-nbitq), 
to_sfixed(-463484616.0/4294967296.0,1,-nbitq), 
to_sfixed(-30142304.0/4294967296.0,1,-nbitq), 
to_sfixed(499607037.0/4294967296.0,1,-nbitq), 
to_sfixed(482045617.0/4294967296.0,1,-nbitq), 
to_sfixed(186343015.0/4294967296.0,1,-nbitq), 
to_sfixed(178923876.0/4294967296.0,1,-nbitq), 
to_sfixed(347423672.0/4294967296.0,1,-nbitq), 
to_sfixed(-462610022.0/4294967296.0,1,-nbitq), 
to_sfixed(254437240.0/4294967296.0,1,-nbitq), 
to_sfixed(76959618.0/4294967296.0,1,-nbitq), 
to_sfixed(-231485738.0/4294967296.0,1,-nbitq), 
to_sfixed(353777215.0/4294967296.0,1,-nbitq), 
to_sfixed(-177330509.0/4294967296.0,1,-nbitq), 
to_sfixed(194686207.0/4294967296.0,1,-nbitq), 
to_sfixed(152757746.0/4294967296.0,1,-nbitq), 
to_sfixed(529231358.0/4294967296.0,1,-nbitq), 
to_sfixed(272045629.0/4294967296.0,1,-nbitq), 
to_sfixed(-398386754.0/4294967296.0,1,-nbitq), 
to_sfixed(149517507.0/4294967296.0,1,-nbitq), 
to_sfixed(67434656.0/4294967296.0,1,-nbitq), 
to_sfixed(-311543941.0/4294967296.0,1,-nbitq), 
to_sfixed(131729902.0/4294967296.0,1,-nbitq), 
to_sfixed(241115828.0/4294967296.0,1,-nbitq), 
to_sfixed(92737431.0/4294967296.0,1,-nbitq), 
to_sfixed(411065623.0/4294967296.0,1,-nbitq), 
to_sfixed(-369319113.0/4294967296.0,1,-nbitq), 
to_sfixed(283523709.0/4294967296.0,1,-nbitq), 
to_sfixed(241207755.0/4294967296.0,1,-nbitq), 
to_sfixed(-10115672.0/4294967296.0,1,-nbitq), 
to_sfixed(-217536264.0/4294967296.0,1,-nbitq), 
to_sfixed(-119369420.0/4294967296.0,1,-nbitq), 
to_sfixed(-317672785.0/4294967296.0,1,-nbitq), 
to_sfixed(-328901890.0/4294967296.0,1,-nbitq), 
to_sfixed(-42814688.0/4294967296.0,1,-nbitq), 
to_sfixed(-353952841.0/4294967296.0,1,-nbitq), 
to_sfixed(-388118160.0/4294967296.0,1,-nbitq), 
to_sfixed(467813259.0/4294967296.0,1,-nbitq), 
to_sfixed(-35188597.0/4294967296.0,1,-nbitq), 
to_sfixed(-303839732.0/4294967296.0,1,-nbitq), 
to_sfixed(218727857.0/4294967296.0,1,-nbitq), 
to_sfixed(-160277594.0/4294967296.0,1,-nbitq), 
to_sfixed(-107144478.0/4294967296.0,1,-nbitq), 
to_sfixed(160753178.0/4294967296.0,1,-nbitq), 
to_sfixed(-236575494.0/4294967296.0,1,-nbitq), 
to_sfixed(438494484.0/4294967296.0,1,-nbitq), 
to_sfixed(108356306.0/4294967296.0,1,-nbitq), 
to_sfixed(550660213.0/4294967296.0,1,-nbitq), 
to_sfixed(-280707429.0/4294967296.0,1,-nbitq), 
to_sfixed(-113030989.0/4294967296.0,1,-nbitq), 
to_sfixed(357162382.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(181535832.0/4294967296.0,1,-nbitq), 
to_sfixed(-569535253.0/4294967296.0,1,-nbitq), 
to_sfixed(375259343.0/4294967296.0,1,-nbitq), 
to_sfixed(-252746376.0/4294967296.0,1,-nbitq), 
to_sfixed(418789857.0/4294967296.0,1,-nbitq), 
to_sfixed(-451574131.0/4294967296.0,1,-nbitq), 
to_sfixed(-24190774.0/4294967296.0,1,-nbitq), 
to_sfixed(19822027.0/4294967296.0,1,-nbitq), 
to_sfixed(-396605614.0/4294967296.0,1,-nbitq), 
to_sfixed(-361640659.0/4294967296.0,1,-nbitq), 
to_sfixed(81153018.0/4294967296.0,1,-nbitq), 
to_sfixed(-7506616.0/4294967296.0,1,-nbitq), 
to_sfixed(40552523.0/4294967296.0,1,-nbitq), 
to_sfixed(-90653546.0/4294967296.0,1,-nbitq), 
to_sfixed(389796896.0/4294967296.0,1,-nbitq), 
to_sfixed(-210114863.0/4294967296.0,1,-nbitq), 
to_sfixed(-254398378.0/4294967296.0,1,-nbitq), 
to_sfixed(-29736380.0/4294967296.0,1,-nbitq), 
to_sfixed(222629277.0/4294967296.0,1,-nbitq), 
to_sfixed(-268187990.0/4294967296.0,1,-nbitq), 
to_sfixed(-73919619.0/4294967296.0,1,-nbitq), 
to_sfixed(-52947878.0/4294967296.0,1,-nbitq), 
to_sfixed(-16299187.0/4294967296.0,1,-nbitq), 
to_sfixed(291810734.0/4294967296.0,1,-nbitq), 
to_sfixed(383707814.0/4294967296.0,1,-nbitq), 
to_sfixed(412695670.0/4294967296.0,1,-nbitq), 
to_sfixed(186669429.0/4294967296.0,1,-nbitq), 
to_sfixed(-460611570.0/4294967296.0,1,-nbitq), 
to_sfixed(-3712098.0/4294967296.0,1,-nbitq), 
to_sfixed(-311185262.0/4294967296.0,1,-nbitq), 
to_sfixed(-472066509.0/4294967296.0,1,-nbitq), 
to_sfixed(-485143584.0/4294967296.0,1,-nbitq), 
to_sfixed(-39735468.0/4294967296.0,1,-nbitq), 
to_sfixed(-335168948.0/4294967296.0,1,-nbitq), 
to_sfixed(445882589.0/4294967296.0,1,-nbitq), 
to_sfixed(46248717.0/4294967296.0,1,-nbitq), 
to_sfixed(197585315.0/4294967296.0,1,-nbitq), 
to_sfixed(-482090226.0/4294967296.0,1,-nbitq), 
to_sfixed(241776479.0/4294967296.0,1,-nbitq), 
to_sfixed(54058365.0/4294967296.0,1,-nbitq), 
to_sfixed(-177754982.0/4294967296.0,1,-nbitq), 
to_sfixed(469746850.0/4294967296.0,1,-nbitq), 
to_sfixed(40649911.0/4294967296.0,1,-nbitq), 
to_sfixed(548164633.0/4294967296.0,1,-nbitq), 
to_sfixed(328817999.0/4294967296.0,1,-nbitq), 
to_sfixed(785845790.0/4294967296.0,1,-nbitq), 
to_sfixed(-192214852.0/4294967296.0,1,-nbitq), 
to_sfixed(-617048478.0/4294967296.0,1,-nbitq), 
to_sfixed(-383177698.0/4294967296.0,1,-nbitq), 
to_sfixed(60144998.0/4294967296.0,1,-nbitq), 
to_sfixed(-106280142.0/4294967296.0,1,-nbitq), 
to_sfixed(-190551238.0/4294967296.0,1,-nbitq), 
to_sfixed(-111378012.0/4294967296.0,1,-nbitq), 
to_sfixed(156806696.0/4294967296.0,1,-nbitq), 
to_sfixed(178613489.0/4294967296.0,1,-nbitq), 
to_sfixed(-490023980.0/4294967296.0,1,-nbitq), 
to_sfixed(186485787.0/4294967296.0,1,-nbitq), 
to_sfixed(-331895139.0/4294967296.0,1,-nbitq), 
to_sfixed(-85931402.0/4294967296.0,1,-nbitq), 
to_sfixed(113939161.0/4294967296.0,1,-nbitq), 
to_sfixed(282166155.0/4294967296.0,1,-nbitq), 
to_sfixed(340684566.0/4294967296.0,1,-nbitq), 
to_sfixed(38144596.0/4294967296.0,1,-nbitq), 
to_sfixed(26019157.0/4294967296.0,1,-nbitq), 
to_sfixed(-338706755.0/4294967296.0,1,-nbitq), 
to_sfixed(-444575257.0/4294967296.0,1,-nbitq), 
to_sfixed(-57640061.0/4294967296.0,1,-nbitq), 
to_sfixed(268358921.0/4294967296.0,1,-nbitq), 
to_sfixed(-319190741.0/4294967296.0,1,-nbitq), 
to_sfixed(-59872382.0/4294967296.0,1,-nbitq), 
to_sfixed(-134285595.0/4294967296.0,1,-nbitq), 
to_sfixed(157048961.0/4294967296.0,1,-nbitq), 
to_sfixed(167824135.0/4294967296.0,1,-nbitq), 
to_sfixed(-40301202.0/4294967296.0,1,-nbitq), 
to_sfixed(-278895582.0/4294967296.0,1,-nbitq), 
to_sfixed(-463632680.0/4294967296.0,1,-nbitq), 
to_sfixed(247740854.0/4294967296.0,1,-nbitq), 
to_sfixed(202949458.0/4294967296.0,1,-nbitq), 
to_sfixed(140939798.0/4294967296.0,1,-nbitq), 
to_sfixed(237700219.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-218933102.0/4294967296.0,1,-nbitq), 
to_sfixed(-23958015.0/4294967296.0,1,-nbitq), 
to_sfixed(-129408463.0/4294967296.0,1,-nbitq), 
to_sfixed(-82523214.0/4294967296.0,1,-nbitq), 
to_sfixed(276445058.0/4294967296.0,1,-nbitq), 
to_sfixed(-293921307.0/4294967296.0,1,-nbitq), 
to_sfixed(115456246.0/4294967296.0,1,-nbitq), 
to_sfixed(73138156.0/4294967296.0,1,-nbitq), 
to_sfixed(262969522.0/4294967296.0,1,-nbitq), 
to_sfixed(-21202708.0/4294967296.0,1,-nbitq), 
to_sfixed(-520386642.0/4294967296.0,1,-nbitq), 
to_sfixed(165004347.0/4294967296.0,1,-nbitq), 
to_sfixed(135556384.0/4294967296.0,1,-nbitq), 
to_sfixed(67292387.0/4294967296.0,1,-nbitq), 
to_sfixed(-180156258.0/4294967296.0,1,-nbitq), 
to_sfixed(66160688.0/4294967296.0,1,-nbitq), 
to_sfixed(-344450736.0/4294967296.0,1,-nbitq), 
to_sfixed(260715640.0/4294967296.0,1,-nbitq), 
to_sfixed(543017650.0/4294967296.0,1,-nbitq), 
to_sfixed(-389145873.0/4294967296.0,1,-nbitq), 
to_sfixed(366325080.0/4294967296.0,1,-nbitq), 
to_sfixed(79497996.0/4294967296.0,1,-nbitq), 
to_sfixed(491067572.0/4294967296.0,1,-nbitq), 
to_sfixed(337382179.0/4294967296.0,1,-nbitq), 
to_sfixed(-224668489.0/4294967296.0,1,-nbitq), 
to_sfixed(479873736.0/4294967296.0,1,-nbitq), 
to_sfixed(173433679.0/4294967296.0,1,-nbitq), 
to_sfixed(-475114534.0/4294967296.0,1,-nbitq), 
to_sfixed(199911552.0/4294967296.0,1,-nbitq), 
to_sfixed(115856761.0/4294967296.0,1,-nbitq), 
to_sfixed(-288475947.0/4294967296.0,1,-nbitq), 
to_sfixed(151310742.0/4294967296.0,1,-nbitq), 
to_sfixed(-212149482.0/4294967296.0,1,-nbitq), 
to_sfixed(136466963.0/4294967296.0,1,-nbitq), 
to_sfixed(131420980.0/4294967296.0,1,-nbitq), 
to_sfixed(-99513918.0/4294967296.0,1,-nbitq), 
to_sfixed(300951744.0/4294967296.0,1,-nbitq), 
to_sfixed(-7328389.0/4294967296.0,1,-nbitq), 
to_sfixed(-293625328.0/4294967296.0,1,-nbitq), 
to_sfixed(-243933732.0/4294967296.0,1,-nbitq), 
to_sfixed(-317240581.0/4294967296.0,1,-nbitq), 
to_sfixed(431766765.0/4294967296.0,1,-nbitq), 
to_sfixed(396261652.0/4294967296.0,1,-nbitq), 
to_sfixed(-302801862.0/4294967296.0,1,-nbitq), 
to_sfixed(103428652.0/4294967296.0,1,-nbitq), 
to_sfixed(627628998.0/4294967296.0,1,-nbitq), 
to_sfixed(-357407088.0/4294967296.0,1,-nbitq), 
to_sfixed(-12027096.0/4294967296.0,1,-nbitq), 
to_sfixed(-395848433.0/4294967296.0,1,-nbitq), 
to_sfixed(444272618.0/4294967296.0,1,-nbitq), 
to_sfixed(-302360411.0/4294967296.0,1,-nbitq), 
to_sfixed(417600901.0/4294967296.0,1,-nbitq), 
to_sfixed(-301888239.0/4294967296.0,1,-nbitq), 
to_sfixed(-88896334.0/4294967296.0,1,-nbitq), 
to_sfixed(449095726.0/4294967296.0,1,-nbitq), 
to_sfixed(-240633810.0/4294967296.0,1,-nbitq), 
to_sfixed(-160371322.0/4294967296.0,1,-nbitq), 
to_sfixed(-231977501.0/4294967296.0,1,-nbitq), 
to_sfixed(-79506362.0/4294967296.0,1,-nbitq), 
to_sfixed(21047739.0/4294967296.0,1,-nbitq), 
to_sfixed(-299326189.0/4294967296.0,1,-nbitq), 
to_sfixed(263455319.0/4294967296.0,1,-nbitq), 
to_sfixed(-481077321.0/4294967296.0,1,-nbitq), 
to_sfixed(-92821119.0/4294967296.0,1,-nbitq), 
to_sfixed(384939914.0/4294967296.0,1,-nbitq), 
to_sfixed(154196172.0/4294967296.0,1,-nbitq), 
to_sfixed(429627235.0/4294967296.0,1,-nbitq), 
to_sfixed(-171089157.0/4294967296.0,1,-nbitq), 
to_sfixed(275129229.0/4294967296.0,1,-nbitq), 
to_sfixed(396470685.0/4294967296.0,1,-nbitq), 
to_sfixed(-344364503.0/4294967296.0,1,-nbitq), 
to_sfixed(150044848.0/4294967296.0,1,-nbitq), 
to_sfixed(123309237.0/4294967296.0,1,-nbitq), 
to_sfixed(396552431.0/4294967296.0,1,-nbitq), 
to_sfixed(-267473730.0/4294967296.0,1,-nbitq), 
to_sfixed(-480880255.0/4294967296.0,1,-nbitq), 
to_sfixed(-230356527.0/4294967296.0,1,-nbitq), 
to_sfixed(-363732487.0/4294967296.0,1,-nbitq), 
to_sfixed(-161385593.0/4294967296.0,1,-nbitq), 
to_sfixed(-344359776.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-94922869.0/4294967296.0,1,-nbitq), 
to_sfixed(-168466183.0/4294967296.0,1,-nbitq), 
to_sfixed(238044213.0/4294967296.0,1,-nbitq), 
to_sfixed(-50134220.0/4294967296.0,1,-nbitq), 
to_sfixed(333288157.0/4294967296.0,1,-nbitq), 
to_sfixed(-179543240.0/4294967296.0,1,-nbitq), 
to_sfixed(129290288.0/4294967296.0,1,-nbitq), 
to_sfixed(56525505.0/4294967296.0,1,-nbitq), 
to_sfixed(-350371368.0/4294967296.0,1,-nbitq), 
to_sfixed(-342375554.0/4294967296.0,1,-nbitq), 
to_sfixed(10387569.0/4294967296.0,1,-nbitq), 
to_sfixed(-186924727.0/4294967296.0,1,-nbitq), 
to_sfixed(-72090018.0/4294967296.0,1,-nbitq), 
to_sfixed(-126342647.0/4294967296.0,1,-nbitq), 
to_sfixed(-2763568.0/4294967296.0,1,-nbitq), 
to_sfixed(121162524.0/4294967296.0,1,-nbitq), 
to_sfixed(-360368753.0/4294967296.0,1,-nbitq), 
to_sfixed(-246372514.0/4294967296.0,1,-nbitq), 
to_sfixed(235079185.0/4294967296.0,1,-nbitq), 
to_sfixed(-72815042.0/4294967296.0,1,-nbitq), 
to_sfixed(-32388557.0/4294967296.0,1,-nbitq), 
to_sfixed(97473318.0/4294967296.0,1,-nbitq), 
to_sfixed(317823921.0/4294967296.0,1,-nbitq), 
to_sfixed(-71028023.0/4294967296.0,1,-nbitq), 
to_sfixed(-257201947.0/4294967296.0,1,-nbitq), 
to_sfixed(-43734251.0/4294967296.0,1,-nbitq), 
to_sfixed(-349859524.0/4294967296.0,1,-nbitq), 
to_sfixed(-6100855.0/4294967296.0,1,-nbitq), 
to_sfixed(238805993.0/4294967296.0,1,-nbitq), 
to_sfixed(314094616.0/4294967296.0,1,-nbitq), 
to_sfixed(-206488633.0/4294967296.0,1,-nbitq), 
to_sfixed(-285930319.0/4294967296.0,1,-nbitq), 
to_sfixed(320331953.0/4294967296.0,1,-nbitq), 
to_sfixed(23807500.0/4294967296.0,1,-nbitq), 
to_sfixed(426019082.0/4294967296.0,1,-nbitq), 
to_sfixed(-244993871.0/4294967296.0,1,-nbitq), 
to_sfixed(-135884833.0/4294967296.0,1,-nbitq), 
to_sfixed(-39074565.0/4294967296.0,1,-nbitq), 
to_sfixed(260977663.0/4294967296.0,1,-nbitq), 
to_sfixed(310226347.0/4294967296.0,1,-nbitq), 
to_sfixed(-148386622.0/4294967296.0,1,-nbitq), 
to_sfixed(-51946810.0/4294967296.0,1,-nbitq), 
to_sfixed(243775244.0/4294967296.0,1,-nbitq), 
to_sfixed(258873041.0/4294967296.0,1,-nbitq), 
to_sfixed(186431386.0/4294967296.0,1,-nbitq), 
to_sfixed(77562192.0/4294967296.0,1,-nbitq), 
to_sfixed(-71101123.0/4294967296.0,1,-nbitq), 
to_sfixed(-501127784.0/4294967296.0,1,-nbitq), 
to_sfixed(142299052.0/4294967296.0,1,-nbitq), 
to_sfixed(-66652212.0/4294967296.0,1,-nbitq), 
to_sfixed(-89823144.0/4294967296.0,1,-nbitq), 
to_sfixed(291813792.0/4294967296.0,1,-nbitq), 
to_sfixed(-297219518.0/4294967296.0,1,-nbitq), 
to_sfixed(94039729.0/4294967296.0,1,-nbitq), 
to_sfixed(349067458.0/4294967296.0,1,-nbitq), 
to_sfixed(-426668339.0/4294967296.0,1,-nbitq), 
to_sfixed(-328143970.0/4294967296.0,1,-nbitq), 
to_sfixed(186854438.0/4294967296.0,1,-nbitq), 
to_sfixed(235637287.0/4294967296.0,1,-nbitq), 
to_sfixed(49768517.0/4294967296.0,1,-nbitq), 
to_sfixed(387559836.0/4294967296.0,1,-nbitq), 
to_sfixed(375650257.0/4294967296.0,1,-nbitq), 
to_sfixed(-158295755.0/4294967296.0,1,-nbitq), 
to_sfixed(414641058.0/4294967296.0,1,-nbitq), 
to_sfixed(-242212107.0/4294967296.0,1,-nbitq), 
to_sfixed(-475289450.0/4294967296.0,1,-nbitq), 
to_sfixed(609108658.0/4294967296.0,1,-nbitq), 
to_sfixed(139302380.0/4294967296.0,1,-nbitq), 
to_sfixed(146682288.0/4294967296.0,1,-nbitq), 
to_sfixed(342323966.0/4294967296.0,1,-nbitq), 
to_sfixed(-488781004.0/4294967296.0,1,-nbitq), 
to_sfixed(-349796847.0/4294967296.0,1,-nbitq), 
to_sfixed(44185115.0/4294967296.0,1,-nbitq), 
to_sfixed(-28989216.0/4294967296.0,1,-nbitq), 
to_sfixed(-145665072.0/4294967296.0,1,-nbitq), 
to_sfixed(-254775695.0/4294967296.0,1,-nbitq), 
to_sfixed(-67281858.0/4294967296.0,1,-nbitq), 
to_sfixed(280862521.0/4294967296.0,1,-nbitq), 
to_sfixed(170941645.0/4294967296.0,1,-nbitq), 
to_sfixed(-169648550.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-343480273.0/4294967296.0,1,-nbitq), 
to_sfixed(-395439191.0/4294967296.0,1,-nbitq), 
to_sfixed(399335385.0/4294967296.0,1,-nbitq), 
to_sfixed(-103856302.0/4294967296.0,1,-nbitq), 
to_sfixed(40665048.0/4294967296.0,1,-nbitq), 
to_sfixed(-169093119.0/4294967296.0,1,-nbitq), 
to_sfixed(-220819065.0/4294967296.0,1,-nbitq), 
to_sfixed(-71951716.0/4294967296.0,1,-nbitq), 
to_sfixed(71554624.0/4294967296.0,1,-nbitq), 
to_sfixed(-50513849.0/4294967296.0,1,-nbitq), 
to_sfixed(247458140.0/4294967296.0,1,-nbitq), 
to_sfixed(-40199868.0/4294967296.0,1,-nbitq), 
to_sfixed(139731820.0/4294967296.0,1,-nbitq), 
to_sfixed(304209721.0/4294967296.0,1,-nbitq), 
to_sfixed(-283150883.0/4294967296.0,1,-nbitq), 
to_sfixed(-233176868.0/4294967296.0,1,-nbitq), 
to_sfixed(-181426428.0/4294967296.0,1,-nbitq), 
to_sfixed(-12938267.0/4294967296.0,1,-nbitq), 
to_sfixed(-174819967.0/4294967296.0,1,-nbitq), 
to_sfixed(-31793092.0/4294967296.0,1,-nbitq), 
to_sfixed(-116666536.0/4294967296.0,1,-nbitq), 
to_sfixed(-45430378.0/4294967296.0,1,-nbitq), 
to_sfixed(524955659.0/4294967296.0,1,-nbitq), 
to_sfixed(-125714587.0/4294967296.0,1,-nbitq), 
to_sfixed(268906116.0/4294967296.0,1,-nbitq), 
to_sfixed(463108904.0/4294967296.0,1,-nbitq), 
to_sfixed(119724035.0/4294967296.0,1,-nbitq), 
to_sfixed(-605948345.0/4294967296.0,1,-nbitq), 
to_sfixed(2603963.0/4294967296.0,1,-nbitq), 
to_sfixed(306170573.0/4294967296.0,1,-nbitq), 
to_sfixed(-426103594.0/4294967296.0,1,-nbitq), 
to_sfixed(-541271650.0/4294967296.0,1,-nbitq), 
to_sfixed(-251282898.0/4294967296.0,1,-nbitq), 
to_sfixed(-514075962.0/4294967296.0,1,-nbitq), 
to_sfixed(541521637.0/4294967296.0,1,-nbitq), 
to_sfixed(33421783.0/4294967296.0,1,-nbitq), 
to_sfixed(358883200.0/4294967296.0,1,-nbitq), 
to_sfixed(-796424.0/4294967296.0,1,-nbitq), 
to_sfixed(-295103797.0/4294967296.0,1,-nbitq), 
to_sfixed(-56827054.0/4294967296.0,1,-nbitq), 
to_sfixed(-482221688.0/4294967296.0,1,-nbitq), 
to_sfixed(435935825.0/4294967296.0,1,-nbitq), 
to_sfixed(102516630.0/4294967296.0,1,-nbitq), 
to_sfixed(-363147410.0/4294967296.0,1,-nbitq), 
to_sfixed(102669361.0/4294967296.0,1,-nbitq), 
to_sfixed(161694769.0/4294967296.0,1,-nbitq), 
to_sfixed(-377991737.0/4294967296.0,1,-nbitq), 
to_sfixed(54887975.0/4294967296.0,1,-nbitq), 
to_sfixed(85293531.0/4294967296.0,1,-nbitq), 
to_sfixed(132864175.0/4294967296.0,1,-nbitq), 
to_sfixed(-165049063.0/4294967296.0,1,-nbitq), 
to_sfixed(-44696675.0/4294967296.0,1,-nbitq), 
to_sfixed(-325149358.0/4294967296.0,1,-nbitq), 
to_sfixed(433594974.0/4294967296.0,1,-nbitq), 
to_sfixed(85442462.0/4294967296.0,1,-nbitq), 
to_sfixed(-68406546.0/4294967296.0,1,-nbitq), 
to_sfixed(109415970.0/4294967296.0,1,-nbitq), 
to_sfixed(-101583386.0/4294967296.0,1,-nbitq), 
to_sfixed(-272661721.0/4294967296.0,1,-nbitq), 
to_sfixed(118811078.0/4294967296.0,1,-nbitq), 
to_sfixed(-130448723.0/4294967296.0,1,-nbitq), 
to_sfixed(-223250200.0/4294967296.0,1,-nbitq), 
to_sfixed(164353187.0/4294967296.0,1,-nbitq), 
to_sfixed(90108426.0/4294967296.0,1,-nbitq), 
to_sfixed(-298589222.0/4294967296.0,1,-nbitq), 
to_sfixed(-444344670.0/4294967296.0,1,-nbitq), 
to_sfixed(863014894.0/4294967296.0,1,-nbitq), 
to_sfixed(-205366102.0/4294967296.0,1,-nbitq), 
to_sfixed(-71977975.0/4294967296.0,1,-nbitq), 
to_sfixed(12647024.0/4294967296.0,1,-nbitq), 
to_sfixed(5989016.0/4294967296.0,1,-nbitq), 
to_sfixed(318711089.0/4294967296.0,1,-nbitq), 
to_sfixed(-317113061.0/4294967296.0,1,-nbitq), 
to_sfixed(-189536693.0/4294967296.0,1,-nbitq), 
to_sfixed(-152084395.0/4294967296.0,1,-nbitq), 
to_sfixed(-516568413.0/4294967296.0,1,-nbitq), 
to_sfixed(-225899967.0/4294967296.0,1,-nbitq), 
to_sfixed(109125569.0/4294967296.0,1,-nbitq), 
to_sfixed(-281050167.0/4294967296.0,1,-nbitq), 
to_sfixed(-89208374.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-400665890.0/4294967296.0,1,-nbitq), 
to_sfixed(-359009756.0/4294967296.0,1,-nbitq), 
to_sfixed(-5774487.0/4294967296.0,1,-nbitq), 
to_sfixed(-292955463.0/4294967296.0,1,-nbitq), 
to_sfixed(513527288.0/4294967296.0,1,-nbitq), 
to_sfixed(-108587499.0/4294967296.0,1,-nbitq), 
to_sfixed(361682749.0/4294967296.0,1,-nbitq), 
to_sfixed(-85302930.0/4294967296.0,1,-nbitq), 
to_sfixed(88128843.0/4294967296.0,1,-nbitq), 
to_sfixed(-40620566.0/4294967296.0,1,-nbitq), 
to_sfixed(-286936105.0/4294967296.0,1,-nbitq), 
to_sfixed(-122590857.0/4294967296.0,1,-nbitq), 
to_sfixed(-83311689.0/4294967296.0,1,-nbitq), 
to_sfixed(137343657.0/4294967296.0,1,-nbitq), 
to_sfixed(81660774.0/4294967296.0,1,-nbitq), 
to_sfixed(318072610.0/4294967296.0,1,-nbitq), 
to_sfixed(-156844809.0/4294967296.0,1,-nbitq), 
to_sfixed(-169172602.0/4294967296.0,1,-nbitq), 
to_sfixed(329456922.0/4294967296.0,1,-nbitq), 
to_sfixed(-153870226.0/4294967296.0,1,-nbitq), 
to_sfixed(-402737025.0/4294967296.0,1,-nbitq), 
to_sfixed(226442535.0/4294967296.0,1,-nbitq), 
to_sfixed(139584179.0/4294967296.0,1,-nbitq), 
to_sfixed(-281514675.0/4294967296.0,1,-nbitq), 
to_sfixed(22792710.0/4294967296.0,1,-nbitq), 
to_sfixed(-120117145.0/4294967296.0,1,-nbitq), 
to_sfixed(91465388.0/4294967296.0,1,-nbitq), 
to_sfixed(-496487267.0/4294967296.0,1,-nbitq), 
to_sfixed(-177956038.0/4294967296.0,1,-nbitq), 
to_sfixed(-45079117.0/4294967296.0,1,-nbitq), 
to_sfixed(110736895.0/4294967296.0,1,-nbitq), 
to_sfixed(-207855022.0/4294967296.0,1,-nbitq), 
to_sfixed(-12142669.0/4294967296.0,1,-nbitq), 
to_sfixed(-256011070.0/4294967296.0,1,-nbitq), 
to_sfixed(-134374524.0/4294967296.0,1,-nbitq), 
to_sfixed(-313901892.0/4294967296.0,1,-nbitq), 
to_sfixed(171830089.0/4294967296.0,1,-nbitq), 
to_sfixed(77955327.0/4294967296.0,1,-nbitq), 
to_sfixed(-275471399.0/4294967296.0,1,-nbitq), 
to_sfixed(182017337.0/4294967296.0,1,-nbitq), 
to_sfixed(-360584658.0/4294967296.0,1,-nbitq), 
to_sfixed(147094506.0/4294967296.0,1,-nbitq), 
to_sfixed(-54510417.0/4294967296.0,1,-nbitq), 
to_sfixed(-72956883.0/4294967296.0,1,-nbitq), 
to_sfixed(19308713.0/4294967296.0,1,-nbitq), 
to_sfixed(138579376.0/4294967296.0,1,-nbitq), 
to_sfixed(102621676.0/4294967296.0,1,-nbitq), 
to_sfixed(-33420868.0/4294967296.0,1,-nbitq), 
to_sfixed(-384263144.0/4294967296.0,1,-nbitq), 
to_sfixed(426766578.0/4294967296.0,1,-nbitq), 
to_sfixed(328386263.0/4294967296.0,1,-nbitq), 
to_sfixed(344361393.0/4294967296.0,1,-nbitq), 
to_sfixed(-309099813.0/4294967296.0,1,-nbitq), 
to_sfixed(221508894.0/4294967296.0,1,-nbitq), 
to_sfixed(-4361721.0/4294967296.0,1,-nbitq), 
to_sfixed(-38252163.0/4294967296.0,1,-nbitq), 
to_sfixed(-9700427.0/4294967296.0,1,-nbitq), 
to_sfixed(-73563655.0/4294967296.0,1,-nbitq), 
to_sfixed(-244820690.0/4294967296.0,1,-nbitq), 
to_sfixed(124462851.0/4294967296.0,1,-nbitq), 
to_sfixed(-76693717.0/4294967296.0,1,-nbitq), 
to_sfixed(280306108.0/4294967296.0,1,-nbitq), 
to_sfixed(-120708698.0/4294967296.0,1,-nbitq), 
to_sfixed(329149776.0/4294967296.0,1,-nbitq), 
to_sfixed(-195934613.0/4294967296.0,1,-nbitq), 
to_sfixed(-280714377.0/4294967296.0,1,-nbitq), 
to_sfixed(462737350.0/4294967296.0,1,-nbitq), 
to_sfixed(53621609.0/4294967296.0,1,-nbitq), 
to_sfixed(79131606.0/4294967296.0,1,-nbitq), 
to_sfixed(205524708.0/4294967296.0,1,-nbitq), 
to_sfixed(-473278234.0/4294967296.0,1,-nbitq), 
to_sfixed(-309795254.0/4294967296.0,1,-nbitq), 
to_sfixed(136114994.0/4294967296.0,1,-nbitq), 
to_sfixed(17195994.0/4294967296.0,1,-nbitq), 
to_sfixed(-109292302.0/4294967296.0,1,-nbitq), 
to_sfixed(-548762272.0/4294967296.0,1,-nbitq), 
to_sfixed(-296731481.0/4294967296.0,1,-nbitq), 
to_sfixed(-78633152.0/4294967296.0,1,-nbitq), 
to_sfixed(-327876519.0/4294967296.0,1,-nbitq), 
to_sfixed(-258944241.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-102294817.0/4294967296.0,1,-nbitq), 
to_sfixed(239736633.0/4294967296.0,1,-nbitq), 
to_sfixed(-67528621.0/4294967296.0,1,-nbitq), 
to_sfixed(-233053513.0/4294967296.0,1,-nbitq), 
to_sfixed(440938182.0/4294967296.0,1,-nbitq), 
to_sfixed(-85001474.0/4294967296.0,1,-nbitq), 
to_sfixed(-33161863.0/4294967296.0,1,-nbitq), 
to_sfixed(227529170.0/4294967296.0,1,-nbitq), 
to_sfixed(-424396424.0/4294967296.0,1,-nbitq), 
to_sfixed(-12140751.0/4294967296.0,1,-nbitq), 
to_sfixed(-463662393.0/4294967296.0,1,-nbitq), 
to_sfixed(5748246.0/4294967296.0,1,-nbitq), 
to_sfixed(333926953.0/4294967296.0,1,-nbitq), 
to_sfixed(-144012665.0/4294967296.0,1,-nbitq), 
to_sfixed(96140884.0/4294967296.0,1,-nbitq), 
to_sfixed(71306392.0/4294967296.0,1,-nbitq), 
to_sfixed(350217949.0/4294967296.0,1,-nbitq), 
to_sfixed(8478453.0/4294967296.0,1,-nbitq), 
to_sfixed(467096164.0/4294967296.0,1,-nbitq), 
to_sfixed(322547698.0/4294967296.0,1,-nbitq), 
to_sfixed(-400967137.0/4294967296.0,1,-nbitq), 
to_sfixed(-2880126.0/4294967296.0,1,-nbitq), 
to_sfixed(148743116.0/4294967296.0,1,-nbitq), 
to_sfixed(155642694.0/4294967296.0,1,-nbitq), 
to_sfixed(5346381.0/4294967296.0,1,-nbitq), 
to_sfixed(591581872.0/4294967296.0,1,-nbitq), 
to_sfixed(-157786976.0/4294967296.0,1,-nbitq), 
to_sfixed(-444758985.0/4294967296.0,1,-nbitq), 
to_sfixed(200843743.0/4294967296.0,1,-nbitq), 
to_sfixed(-43109762.0/4294967296.0,1,-nbitq), 
to_sfixed(-141879980.0/4294967296.0,1,-nbitq), 
to_sfixed(-399390376.0/4294967296.0,1,-nbitq), 
to_sfixed(453675613.0/4294967296.0,1,-nbitq), 
to_sfixed(-50542178.0/4294967296.0,1,-nbitq), 
to_sfixed(308951811.0/4294967296.0,1,-nbitq), 
to_sfixed(240312793.0/4294967296.0,1,-nbitq), 
to_sfixed(-242876421.0/4294967296.0,1,-nbitq), 
to_sfixed(202013153.0/4294967296.0,1,-nbitq), 
to_sfixed(-167928835.0/4294967296.0,1,-nbitq), 
to_sfixed(-34697020.0/4294967296.0,1,-nbitq), 
to_sfixed(-465041409.0/4294967296.0,1,-nbitq), 
to_sfixed(122995877.0/4294967296.0,1,-nbitq), 
to_sfixed(238427021.0/4294967296.0,1,-nbitq), 
to_sfixed(-82238837.0/4294967296.0,1,-nbitq), 
to_sfixed(-49569930.0/4294967296.0,1,-nbitq), 
to_sfixed(475220846.0/4294967296.0,1,-nbitq), 
to_sfixed(102080053.0/4294967296.0,1,-nbitq), 
to_sfixed(-157351314.0/4294967296.0,1,-nbitq), 
to_sfixed(205960695.0/4294967296.0,1,-nbitq), 
to_sfixed(154867963.0/4294967296.0,1,-nbitq), 
to_sfixed(348548727.0/4294967296.0,1,-nbitq), 
to_sfixed(128082979.0/4294967296.0,1,-nbitq), 
to_sfixed(-451393199.0/4294967296.0,1,-nbitq), 
to_sfixed(222894188.0/4294967296.0,1,-nbitq), 
to_sfixed(-19877411.0/4294967296.0,1,-nbitq), 
to_sfixed(209911987.0/4294967296.0,1,-nbitq), 
to_sfixed(-221347777.0/4294967296.0,1,-nbitq), 
to_sfixed(-217645342.0/4294967296.0,1,-nbitq), 
to_sfixed(388355056.0/4294967296.0,1,-nbitq), 
to_sfixed(-273959285.0/4294967296.0,1,-nbitq), 
to_sfixed(-97048010.0/4294967296.0,1,-nbitq), 
to_sfixed(457505300.0/4294967296.0,1,-nbitq), 
to_sfixed(-194911654.0/4294967296.0,1,-nbitq), 
to_sfixed(389775028.0/4294967296.0,1,-nbitq), 
to_sfixed(-272627257.0/4294967296.0,1,-nbitq), 
to_sfixed(-300524507.0/4294967296.0,1,-nbitq), 
to_sfixed(198964851.0/4294967296.0,1,-nbitq), 
to_sfixed(-397503825.0/4294967296.0,1,-nbitq), 
to_sfixed(-226636681.0/4294967296.0,1,-nbitq), 
to_sfixed(257780517.0/4294967296.0,1,-nbitq), 
to_sfixed(-414221009.0/4294967296.0,1,-nbitq), 
to_sfixed(173862960.0/4294967296.0,1,-nbitq), 
to_sfixed(37612924.0/4294967296.0,1,-nbitq), 
to_sfixed(-231855064.0/4294967296.0,1,-nbitq), 
to_sfixed(-217823522.0/4294967296.0,1,-nbitq), 
to_sfixed(-642258226.0/4294967296.0,1,-nbitq), 
to_sfixed(-52347419.0/4294967296.0,1,-nbitq), 
to_sfixed(-86959797.0/4294967296.0,1,-nbitq), 
to_sfixed(-530014931.0/4294967296.0,1,-nbitq), 
to_sfixed(378725430.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-297836672.0/4294967296.0,1,-nbitq), 
to_sfixed(-244246953.0/4294967296.0,1,-nbitq), 
to_sfixed(-317467727.0/4294967296.0,1,-nbitq), 
to_sfixed(-112284485.0/4294967296.0,1,-nbitq), 
to_sfixed(447788429.0/4294967296.0,1,-nbitq), 
to_sfixed(-13826618.0/4294967296.0,1,-nbitq), 
to_sfixed(357853812.0/4294967296.0,1,-nbitq), 
to_sfixed(201860901.0/4294967296.0,1,-nbitq), 
to_sfixed(-10045586.0/4294967296.0,1,-nbitq), 
to_sfixed(-5003083.0/4294967296.0,1,-nbitq), 
to_sfixed(5295251.0/4294967296.0,1,-nbitq), 
to_sfixed(99810698.0/4294967296.0,1,-nbitq), 
to_sfixed(-157863843.0/4294967296.0,1,-nbitq), 
to_sfixed(59027306.0/4294967296.0,1,-nbitq), 
to_sfixed(466603523.0/4294967296.0,1,-nbitq), 
to_sfixed(-62179525.0/4294967296.0,1,-nbitq), 
to_sfixed(-107529335.0/4294967296.0,1,-nbitq), 
to_sfixed(-11927662.0/4294967296.0,1,-nbitq), 
to_sfixed(690605768.0/4294967296.0,1,-nbitq), 
to_sfixed(-226436830.0/4294967296.0,1,-nbitq), 
to_sfixed(-196418051.0/4294967296.0,1,-nbitq), 
to_sfixed(464323695.0/4294967296.0,1,-nbitq), 
to_sfixed(565585362.0/4294967296.0,1,-nbitq), 
to_sfixed(-194563107.0/4294967296.0,1,-nbitq), 
to_sfixed(-9104968.0/4294967296.0,1,-nbitq), 
to_sfixed(543319329.0/4294967296.0,1,-nbitq), 
to_sfixed(320647443.0/4294967296.0,1,-nbitq), 
to_sfixed(187396933.0/4294967296.0,1,-nbitq), 
to_sfixed(-245122142.0/4294967296.0,1,-nbitq), 
to_sfixed(280116918.0/4294967296.0,1,-nbitq), 
to_sfixed(192361969.0/4294967296.0,1,-nbitq), 
to_sfixed(80433754.0/4294967296.0,1,-nbitq), 
to_sfixed(118392568.0/4294967296.0,1,-nbitq), 
to_sfixed(-353994456.0/4294967296.0,1,-nbitq), 
to_sfixed(420826453.0/4294967296.0,1,-nbitq), 
to_sfixed(-20429042.0/4294967296.0,1,-nbitq), 
to_sfixed(-264046210.0/4294967296.0,1,-nbitq), 
to_sfixed(-458939401.0/4294967296.0,1,-nbitq), 
to_sfixed(245007680.0/4294967296.0,1,-nbitq), 
to_sfixed(-104550262.0/4294967296.0,1,-nbitq), 
to_sfixed(-183440296.0/4294967296.0,1,-nbitq), 
to_sfixed(418404109.0/4294967296.0,1,-nbitq), 
to_sfixed(304954617.0/4294967296.0,1,-nbitq), 
to_sfixed(-253005134.0/4294967296.0,1,-nbitq), 
to_sfixed(17789859.0/4294967296.0,1,-nbitq), 
to_sfixed(231566848.0/4294967296.0,1,-nbitq), 
to_sfixed(277925848.0/4294967296.0,1,-nbitq), 
to_sfixed(296687673.0/4294967296.0,1,-nbitq), 
to_sfixed(-137457862.0/4294967296.0,1,-nbitq), 
to_sfixed(177829114.0/4294967296.0,1,-nbitq), 
to_sfixed(302670888.0/4294967296.0,1,-nbitq), 
to_sfixed(-207437480.0/4294967296.0,1,-nbitq), 
to_sfixed(154217356.0/4294967296.0,1,-nbitq), 
to_sfixed(-180537440.0/4294967296.0,1,-nbitq), 
to_sfixed(393540965.0/4294967296.0,1,-nbitq), 
to_sfixed(88933255.0/4294967296.0,1,-nbitq), 
to_sfixed(521136974.0/4294967296.0,1,-nbitq), 
to_sfixed(-519398403.0/4294967296.0,1,-nbitq), 
to_sfixed(-355188585.0/4294967296.0,1,-nbitq), 
to_sfixed(305813175.0/4294967296.0,1,-nbitq), 
to_sfixed(92116391.0/4294967296.0,1,-nbitq), 
to_sfixed(-307025102.0/4294967296.0,1,-nbitq), 
to_sfixed(-175636904.0/4294967296.0,1,-nbitq), 
to_sfixed(-91594460.0/4294967296.0,1,-nbitq), 
to_sfixed(-20743062.0/4294967296.0,1,-nbitq), 
to_sfixed(-44436515.0/4294967296.0,1,-nbitq), 
to_sfixed(564662996.0/4294967296.0,1,-nbitq), 
to_sfixed(-20242218.0/4294967296.0,1,-nbitq), 
to_sfixed(144658453.0/4294967296.0,1,-nbitq), 
to_sfixed(146793391.0/4294967296.0,1,-nbitq), 
to_sfixed(-394297097.0/4294967296.0,1,-nbitq), 
to_sfixed(-330129746.0/4294967296.0,1,-nbitq), 
to_sfixed(-44397945.0/4294967296.0,1,-nbitq), 
to_sfixed(-135575583.0/4294967296.0,1,-nbitq), 
to_sfixed(366399549.0/4294967296.0,1,-nbitq), 
to_sfixed(-233852126.0/4294967296.0,1,-nbitq), 
to_sfixed(96751882.0/4294967296.0,1,-nbitq), 
to_sfixed(249766045.0/4294967296.0,1,-nbitq), 
to_sfixed(274519095.0/4294967296.0,1,-nbitq), 
to_sfixed(290730670.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(150828770.0/4294967296.0,1,-nbitq), 
to_sfixed(-189578411.0/4294967296.0,1,-nbitq), 
to_sfixed(-205035681.0/4294967296.0,1,-nbitq), 
to_sfixed(18305786.0/4294967296.0,1,-nbitq), 
to_sfixed(40788.0/4294967296.0,1,-nbitq), 
to_sfixed(-190240212.0/4294967296.0,1,-nbitq), 
to_sfixed(-263948036.0/4294967296.0,1,-nbitq), 
to_sfixed(246983377.0/4294967296.0,1,-nbitq), 
to_sfixed(-8649301.0/4294967296.0,1,-nbitq), 
to_sfixed(-34589821.0/4294967296.0,1,-nbitq), 
to_sfixed(-56941557.0/4294967296.0,1,-nbitq), 
to_sfixed(188713243.0/4294967296.0,1,-nbitq), 
to_sfixed(-140562158.0/4294967296.0,1,-nbitq), 
to_sfixed(-75987842.0/4294967296.0,1,-nbitq), 
to_sfixed(-185205573.0/4294967296.0,1,-nbitq), 
to_sfixed(-515286777.0/4294967296.0,1,-nbitq), 
to_sfixed(-298791807.0/4294967296.0,1,-nbitq), 
to_sfixed(-244038296.0/4294967296.0,1,-nbitq), 
to_sfixed(53846645.0/4294967296.0,1,-nbitq), 
to_sfixed(-42768415.0/4294967296.0,1,-nbitq), 
to_sfixed(-187869264.0/4294967296.0,1,-nbitq), 
to_sfixed(364221530.0/4294967296.0,1,-nbitq), 
to_sfixed(150124507.0/4294967296.0,1,-nbitq), 
to_sfixed(-23010944.0/4294967296.0,1,-nbitq), 
to_sfixed(291732523.0/4294967296.0,1,-nbitq), 
to_sfixed(265034301.0/4294967296.0,1,-nbitq), 
to_sfixed(-180652491.0/4294967296.0,1,-nbitq), 
to_sfixed(265053277.0/4294967296.0,1,-nbitq), 
to_sfixed(60494485.0/4294967296.0,1,-nbitq), 
to_sfixed(38803294.0/4294967296.0,1,-nbitq), 
to_sfixed(-366731231.0/4294967296.0,1,-nbitq), 
to_sfixed(-197724015.0/4294967296.0,1,-nbitq), 
to_sfixed(-230861607.0/4294967296.0,1,-nbitq), 
to_sfixed(127509873.0/4294967296.0,1,-nbitq), 
to_sfixed(-14654443.0/4294967296.0,1,-nbitq), 
to_sfixed(21212421.0/4294967296.0,1,-nbitq), 
to_sfixed(42304830.0/4294967296.0,1,-nbitq), 
to_sfixed(-441086327.0/4294967296.0,1,-nbitq), 
to_sfixed(-131288714.0/4294967296.0,1,-nbitq), 
to_sfixed(43355736.0/4294967296.0,1,-nbitq), 
to_sfixed(481146426.0/4294967296.0,1,-nbitq), 
to_sfixed(233152349.0/4294967296.0,1,-nbitq), 
to_sfixed(246807102.0/4294967296.0,1,-nbitq), 
to_sfixed(-493413489.0/4294967296.0,1,-nbitq), 
to_sfixed(366911331.0/4294967296.0,1,-nbitq), 
to_sfixed(447211554.0/4294967296.0,1,-nbitq), 
to_sfixed(159973435.0/4294967296.0,1,-nbitq), 
to_sfixed(-30004739.0/4294967296.0,1,-nbitq), 
to_sfixed(61360638.0/4294967296.0,1,-nbitq), 
to_sfixed(426001901.0/4294967296.0,1,-nbitq), 
to_sfixed(128965381.0/4294967296.0,1,-nbitq), 
to_sfixed(-163947029.0/4294967296.0,1,-nbitq), 
to_sfixed(-185143593.0/4294967296.0,1,-nbitq), 
to_sfixed(-73490680.0/4294967296.0,1,-nbitq), 
to_sfixed(168332676.0/4294967296.0,1,-nbitq), 
to_sfixed(424332556.0/4294967296.0,1,-nbitq), 
to_sfixed(461280351.0/4294967296.0,1,-nbitq), 
to_sfixed(-662909461.0/4294967296.0,1,-nbitq), 
to_sfixed(-338979725.0/4294967296.0,1,-nbitq), 
to_sfixed(197145432.0/4294967296.0,1,-nbitq), 
to_sfixed(151266744.0/4294967296.0,1,-nbitq), 
to_sfixed(18780965.0/4294967296.0,1,-nbitq), 
to_sfixed(-285663390.0/4294967296.0,1,-nbitq), 
to_sfixed(-272776254.0/4294967296.0,1,-nbitq), 
to_sfixed(138780160.0/4294967296.0,1,-nbitq), 
to_sfixed(-156811750.0/4294967296.0,1,-nbitq), 
to_sfixed(567583798.0/4294967296.0,1,-nbitq), 
to_sfixed(231749844.0/4294967296.0,1,-nbitq), 
to_sfixed(253287571.0/4294967296.0,1,-nbitq), 
to_sfixed(237255108.0/4294967296.0,1,-nbitq), 
to_sfixed(-506939349.0/4294967296.0,1,-nbitq), 
to_sfixed(277836508.0/4294967296.0,1,-nbitq), 
to_sfixed(-90525258.0/4294967296.0,1,-nbitq), 
to_sfixed(-40973707.0/4294967296.0,1,-nbitq), 
to_sfixed(492430378.0/4294967296.0,1,-nbitq), 
to_sfixed(-652838319.0/4294967296.0,1,-nbitq), 
to_sfixed(316502877.0/4294967296.0,1,-nbitq), 
to_sfixed(-347761788.0/4294967296.0,1,-nbitq), 
to_sfixed(54451316.0/4294967296.0,1,-nbitq), 
to_sfixed(-92435262.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-325957654.0/4294967296.0,1,-nbitq), 
to_sfixed(86475874.0/4294967296.0,1,-nbitq), 
to_sfixed(-428494506.0/4294967296.0,1,-nbitq), 
to_sfixed(169370199.0/4294967296.0,1,-nbitq), 
to_sfixed(-98856127.0/4294967296.0,1,-nbitq), 
to_sfixed(355085121.0/4294967296.0,1,-nbitq), 
to_sfixed(-183079298.0/4294967296.0,1,-nbitq), 
to_sfixed(-198237167.0/4294967296.0,1,-nbitq), 
to_sfixed(-381463891.0/4294967296.0,1,-nbitq), 
to_sfixed(371322563.0/4294967296.0,1,-nbitq), 
to_sfixed(200478982.0/4294967296.0,1,-nbitq), 
to_sfixed(-236124949.0/4294967296.0,1,-nbitq), 
to_sfixed(215132196.0/4294967296.0,1,-nbitq), 
to_sfixed(-186491656.0/4294967296.0,1,-nbitq), 
to_sfixed(283233473.0/4294967296.0,1,-nbitq), 
to_sfixed(-319478183.0/4294967296.0,1,-nbitq), 
to_sfixed(-129695678.0/4294967296.0,1,-nbitq), 
to_sfixed(355111898.0/4294967296.0,1,-nbitq), 
to_sfixed(386533358.0/4294967296.0,1,-nbitq), 
to_sfixed(66144469.0/4294967296.0,1,-nbitq), 
to_sfixed(-176152597.0/4294967296.0,1,-nbitq), 
to_sfixed(529704885.0/4294967296.0,1,-nbitq), 
to_sfixed(565732469.0/4294967296.0,1,-nbitq), 
to_sfixed(-145382215.0/4294967296.0,1,-nbitq), 
to_sfixed(-289639750.0/4294967296.0,1,-nbitq), 
to_sfixed(371470923.0/4294967296.0,1,-nbitq), 
to_sfixed(-63539442.0/4294967296.0,1,-nbitq), 
to_sfixed(-124518478.0/4294967296.0,1,-nbitq), 
to_sfixed(18215017.0/4294967296.0,1,-nbitq), 
to_sfixed(-554880644.0/4294967296.0,1,-nbitq), 
to_sfixed(-165277593.0/4294967296.0,1,-nbitq), 
to_sfixed(-398725311.0/4294967296.0,1,-nbitq), 
to_sfixed(-116178736.0/4294967296.0,1,-nbitq), 
to_sfixed(-419099451.0/4294967296.0,1,-nbitq), 
to_sfixed(-373969545.0/4294967296.0,1,-nbitq), 
to_sfixed(206351831.0/4294967296.0,1,-nbitq), 
to_sfixed(516740186.0/4294967296.0,1,-nbitq), 
to_sfixed(171771959.0/4294967296.0,1,-nbitq), 
to_sfixed(130071270.0/4294967296.0,1,-nbitq), 
to_sfixed(155311637.0/4294967296.0,1,-nbitq), 
to_sfixed(-107954987.0/4294967296.0,1,-nbitq), 
to_sfixed(-82866387.0/4294967296.0,1,-nbitq), 
to_sfixed(-44731943.0/4294967296.0,1,-nbitq), 
to_sfixed(-679359642.0/4294967296.0,1,-nbitq), 
to_sfixed(386144616.0/4294967296.0,1,-nbitq), 
to_sfixed(324575996.0/4294967296.0,1,-nbitq), 
to_sfixed(225653271.0/4294967296.0,1,-nbitq), 
to_sfixed(-97098109.0/4294967296.0,1,-nbitq), 
to_sfixed(88910767.0/4294967296.0,1,-nbitq), 
to_sfixed(173903587.0/4294967296.0,1,-nbitq), 
to_sfixed(122587753.0/4294967296.0,1,-nbitq), 
to_sfixed(-292009361.0/4294967296.0,1,-nbitq), 
to_sfixed(55839384.0/4294967296.0,1,-nbitq), 
to_sfixed(-263864610.0/4294967296.0,1,-nbitq), 
to_sfixed(369481038.0/4294967296.0,1,-nbitq), 
to_sfixed(266907561.0/4294967296.0,1,-nbitq), 
to_sfixed(375941385.0/4294967296.0,1,-nbitq), 
to_sfixed(-329413517.0/4294967296.0,1,-nbitq), 
to_sfixed(252748391.0/4294967296.0,1,-nbitq), 
to_sfixed(388227215.0/4294967296.0,1,-nbitq), 
to_sfixed(223686373.0/4294967296.0,1,-nbitq), 
to_sfixed(34074263.0/4294967296.0,1,-nbitq), 
to_sfixed(-289021432.0/4294967296.0,1,-nbitq), 
to_sfixed(-147775270.0/4294967296.0,1,-nbitq), 
to_sfixed(-243746329.0/4294967296.0,1,-nbitq), 
to_sfixed(-238886692.0/4294967296.0,1,-nbitq), 
to_sfixed(306252157.0/4294967296.0,1,-nbitq), 
to_sfixed(118271821.0/4294967296.0,1,-nbitq), 
to_sfixed(-347406434.0/4294967296.0,1,-nbitq), 
to_sfixed(-107351855.0/4294967296.0,1,-nbitq), 
to_sfixed(-646024808.0/4294967296.0,1,-nbitq), 
to_sfixed(-306228566.0/4294967296.0,1,-nbitq), 
to_sfixed(209180799.0/4294967296.0,1,-nbitq), 
to_sfixed(100987823.0/4294967296.0,1,-nbitq), 
to_sfixed(82943615.0/4294967296.0,1,-nbitq), 
to_sfixed(-56729135.0/4294967296.0,1,-nbitq), 
to_sfixed(-109295926.0/4294967296.0,1,-nbitq), 
to_sfixed(-322958727.0/4294967296.0,1,-nbitq), 
to_sfixed(287537480.0/4294967296.0,1,-nbitq), 
to_sfixed(-154813415.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(79778737.0/4294967296.0,1,-nbitq), 
to_sfixed(-294777635.0/4294967296.0,1,-nbitq), 
to_sfixed(465876186.0/4294967296.0,1,-nbitq), 
to_sfixed(-368022546.0/4294967296.0,1,-nbitq), 
to_sfixed(167309966.0/4294967296.0,1,-nbitq), 
to_sfixed(94592637.0/4294967296.0,1,-nbitq), 
to_sfixed(339120015.0/4294967296.0,1,-nbitq), 
to_sfixed(-351301856.0/4294967296.0,1,-nbitq), 
to_sfixed(26803561.0/4294967296.0,1,-nbitq), 
to_sfixed(268252975.0/4294967296.0,1,-nbitq), 
to_sfixed(939176638.0/4294967296.0,1,-nbitq), 
to_sfixed(-152213246.0/4294967296.0,1,-nbitq), 
to_sfixed(-1061531901.0/4294967296.0,1,-nbitq), 
to_sfixed(-596177050.0/4294967296.0,1,-nbitq), 
to_sfixed(-151727640.0/4294967296.0,1,-nbitq), 
to_sfixed(-341456531.0/4294967296.0,1,-nbitq), 
to_sfixed(16158.0/4294967296.0,1,-nbitq), 
to_sfixed(366088851.0/4294967296.0,1,-nbitq), 
to_sfixed(695447041.0/4294967296.0,1,-nbitq), 
to_sfixed(-28548121.0/4294967296.0,1,-nbitq), 
to_sfixed(223518843.0/4294967296.0,1,-nbitq), 
to_sfixed(267306524.0/4294967296.0,1,-nbitq), 
to_sfixed(721520084.0/4294967296.0,1,-nbitq), 
to_sfixed(-125700315.0/4294967296.0,1,-nbitq), 
to_sfixed(-302752379.0/4294967296.0,1,-nbitq), 
to_sfixed(571597081.0/4294967296.0,1,-nbitq), 
to_sfixed(437226914.0/4294967296.0,1,-nbitq), 
to_sfixed(527440459.0/4294967296.0,1,-nbitq), 
to_sfixed(-287106118.0/4294967296.0,1,-nbitq), 
to_sfixed(-659750192.0/4294967296.0,1,-nbitq), 
to_sfixed(-163533888.0/4294967296.0,1,-nbitq), 
to_sfixed(-216796917.0/4294967296.0,1,-nbitq), 
to_sfixed(-203130351.0/4294967296.0,1,-nbitq), 
to_sfixed(435112855.0/4294967296.0,1,-nbitq), 
to_sfixed(222679161.0/4294967296.0,1,-nbitq), 
to_sfixed(-610163118.0/4294967296.0,1,-nbitq), 
to_sfixed(274679841.0/4294967296.0,1,-nbitq), 
to_sfixed(-587780543.0/4294967296.0,1,-nbitq), 
to_sfixed(171358385.0/4294967296.0,1,-nbitq), 
to_sfixed(122811779.0/4294967296.0,1,-nbitq), 
to_sfixed(-57039923.0/4294967296.0,1,-nbitq), 
to_sfixed(-261039979.0/4294967296.0,1,-nbitq), 
to_sfixed(209025470.0/4294967296.0,1,-nbitq), 
to_sfixed(-821471102.0/4294967296.0,1,-nbitq), 
to_sfixed(543413936.0/4294967296.0,1,-nbitq), 
to_sfixed(516860343.0/4294967296.0,1,-nbitq), 
to_sfixed(199004206.0/4294967296.0,1,-nbitq), 
to_sfixed(717784775.0/4294967296.0,1,-nbitq), 
to_sfixed(-237537638.0/4294967296.0,1,-nbitq), 
to_sfixed(-93951265.0/4294967296.0,1,-nbitq), 
to_sfixed(244361.0/4294967296.0,1,-nbitq), 
to_sfixed(582361488.0/4294967296.0,1,-nbitq), 
to_sfixed(-43030274.0/4294967296.0,1,-nbitq), 
to_sfixed(-823554184.0/4294967296.0,1,-nbitq), 
to_sfixed(-561941098.0/4294967296.0,1,-nbitq), 
to_sfixed(-878068.0/4294967296.0,1,-nbitq), 
to_sfixed(267369914.0/4294967296.0,1,-nbitq), 
to_sfixed(-737038756.0/4294967296.0,1,-nbitq), 
to_sfixed(232449783.0/4294967296.0,1,-nbitq), 
to_sfixed(-117609730.0/4294967296.0,1,-nbitq), 
to_sfixed(113769726.0/4294967296.0,1,-nbitq), 
to_sfixed(-535676061.0/4294967296.0,1,-nbitq), 
to_sfixed(342743717.0/4294967296.0,1,-nbitq), 
to_sfixed(-153961136.0/4294967296.0,1,-nbitq), 
to_sfixed(-321738466.0/4294967296.0,1,-nbitq), 
to_sfixed(145699495.0/4294967296.0,1,-nbitq), 
to_sfixed(-209269979.0/4294967296.0,1,-nbitq), 
to_sfixed(-76679305.0/4294967296.0,1,-nbitq), 
to_sfixed(29348711.0/4294967296.0,1,-nbitq), 
to_sfixed(-564525923.0/4294967296.0,1,-nbitq), 
to_sfixed(-478429732.0/4294967296.0,1,-nbitq), 
to_sfixed(-345042879.0/4294967296.0,1,-nbitq), 
to_sfixed(-19176807.0/4294967296.0,1,-nbitq), 
to_sfixed(270253994.0/4294967296.0,1,-nbitq), 
to_sfixed(73133532.0/4294967296.0,1,-nbitq), 
to_sfixed(-218027390.0/4294967296.0,1,-nbitq), 
to_sfixed(-3779695.0/4294967296.0,1,-nbitq), 
to_sfixed(-270860730.0/4294967296.0,1,-nbitq), 
to_sfixed(288052386.0/4294967296.0,1,-nbitq), 
to_sfixed(353577362.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-75031191.0/4294967296.0,1,-nbitq), 
to_sfixed(397058192.0/4294967296.0,1,-nbitq), 
to_sfixed(101360006.0/4294967296.0,1,-nbitq), 
to_sfixed(-370335689.0/4294967296.0,1,-nbitq), 
to_sfixed(-94570390.0/4294967296.0,1,-nbitq), 
to_sfixed(381806988.0/4294967296.0,1,-nbitq), 
to_sfixed(-293710299.0/4294967296.0,1,-nbitq), 
to_sfixed(-534340523.0/4294967296.0,1,-nbitq), 
to_sfixed(79985652.0/4294967296.0,1,-nbitq), 
to_sfixed(-265743610.0/4294967296.0,1,-nbitq), 
to_sfixed(1052015187.0/4294967296.0,1,-nbitq), 
to_sfixed(-22273052.0/4294967296.0,1,-nbitq), 
to_sfixed(-872362436.0/4294967296.0,1,-nbitq), 
to_sfixed(-490361363.0/4294967296.0,1,-nbitq), 
to_sfixed(-172961268.0/4294967296.0,1,-nbitq), 
to_sfixed(-1034777875.0/4294967296.0,1,-nbitq), 
to_sfixed(-378718043.0/4294967296.0,1,-nbitq), 
to_sfixed(96890408.0/4294967296.0,1,-nbitq), 
to_sfixed(638904378.0/4294967296.0,1,-nbitq), 
to_sfixed(-99994010.0/4294967296.0,1,-nbitq), 
to_sfixed(-214440996.0/4294967296.0,1,-nbitq), 
to_sfixed(472967032.0/4294967296.0,1,-nbitq), 
to_sfixed(240685888.0/4294967296.0,1,-nbitq), 
to_sfixed(-388261819.0/4294967296.0,1,-nbitq), 
to_sfixed(175499626.0/4294967296.0,1,-nbitq), 
to_sfixed(-152269478.0/4294967296.0,1,-nbitq), 
to_sfixed(259793025.0/4294967296.0,1,-nbitq), 
to_sfixed(367297259.0/4294967296.0,1,-nbitq), 
to_sfixed(-961375434.0/4294967296.0,1,-nbitq), 
to_sfixed(-608102697.0/4294967296.0,1,-nbitq), 
to_sfixed(372115704.0/4294967296.0,1,-nbitq), 
to_sfixed(-291205093.0/4294967296.0,1,-nbitq), 
to_sfixed(-407614554.0/4294967296.0,1,-nbitq), 
to_sfixed(65809394.0/4294967296.0,1,-nbitq), 
to_sfixed(-260653334.0/4294967296.0,1,-nbitq), 
to_sfixed(-899776426.0/4294967296.0,1,-nbitq), 
to_sfixed(-234702568.0/4294967296.0,1,-nbitq), 
to_sfixed(-156858745.0/4294967296.0,1,-nbitq), 
to_sfixed(351399415.0/4294967296.0,1,-nbitq), 
to_sfixed(-10225041.0/4294967296.0,1,-nbitq), 
to_sfixed(-141567488.0/4294967296.0,1,-nbitq), 
to_sfixed(543044539.0/4294967296.0,1,-nbitq), 
to_sfixed(21087559.0/4294967296.0,1,-nbitq), 
to_sfixed(-924339305.0/4294967296.0,1,-nbitq), 
to_sfixed(392614204.0/4294967296.0,1,-nbitq), 
to_sfixed(510332340.0/4294967296.0,1,-nbitq), 
to_sfixed(-290954579.0/4294967296.0,1,-nbitq), 
to_sfixed(919481239.0/4294967296.0,1,-nbitq), 
to_sfixed(-291207046.0/4294967296.0,1,-nbitq), 
to_sfixed(-114230731.0/4294967296.0,1,-nbitq), 
to_sfixed(250868889.0/4294967296.0,1,-nbitq), 
to_sfixed(314770299.0/4294967296.0,1,-nbitq), 
to_sfixed(205145039.0/4294967296.0,1,-nbitq), 
to_sfixed(-1093812516.0/4294967296.0,1,-nbitq), 
to_sfixed(-423374236.0/4294967296.0,1,-nbitq), 
to_sfixed(129726786.0/4294967296.0,1,-nbitq), 
to_sfixed(108331646.0/4294967296.0,1,-nbitq), 
to_sfixed(-330852936.0/4294967296.0,1,-nbitq), 
to_sfixed(212646447.0/4294967296.0,1,-nbitq), 
to_sfixed(399216133.0/4294967296.0,1,-nbitq), 
to_sfixed(263265075.0/4294967296.0,1,-nbitq), 
to_sfixed(-637194614.0/4294967296.0,1,-nbitq), 
to_sfixed(556335822.0/4294967296.0,1,-nbitq), 
to_sfixed(-149642027.0/4294967296.0,1,-nbitq), 
to_sfixed(110337521.0/4294967296.0,1,-nbitq), 
to_sfixed(-372443131.0/4294967296.0,1,-nbitq), 
to_sfixed(-524381553.0/4294967296.0,1,-nbitq), 
to_sfixed(-392375496.0/4294967296.0,1,-nbitq), 
to_sfixed(-299673973.0/4294967296.0,1,-nbitq), 
to_sfixed(-569966496.0/4294967296.0,1,-nbitq), 
to_sfixed(-694603587.0/4294967296.0,1,-nbitq), 
to_sfixed(-534805477.0/4294967296.0,1,-nbitq), 
to_sfixed(23112506.0/4294967296.0,1,-nbitq), 
to_sfixed(-301849722.0/4294967296.0,1,-nbitq), 
to_sfixed(262273645.0/4294967296.0,1,-nbitq), 
to_sfixed(-384466690.0/4294967296.0,1,-nbitq), 
to_sfixed(653836177.0/4294967296.0,1,-nbitq), 
to_sfixed(-341121215.0/4294967296.0,1,-nbitq), 
to_sfixed(531010888.0/4294967296.0,1,-nbitq), 
to_sfixed(191366730.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(367591997.0/4294967296.0,1,-nbitq), 
to_sfixed(-44369436.0/4294967296.0,1,-nbitq), 
to_sfixed(102440163.0/4294967296.0,1,-nbitq), 
to_sfixed(342902131.0/4294967296.0,1,-nbitq), 
to_sfixed(462774709.0/4294967296.0,1,-nbitq), 
to_sfixed(-244552365.0/4294967296.0,1,-nbitq), 
to_sfixed(319084009.0/4294967296.0,1,-nbitq), 
to_sfixed(-538057008.0/4294967296.0,1,-nbitq), 
to_sfixed(-27640047.0/4294967296.0,1,-nbitq), 
to_sfixed(-251765821.0/4294967296.0,1,-nbitq), 
to_sfixed(636756080.0/4294967296.0,1,-nbitq), 
to_sfixed(278244469.0/4294967296.0,1,-nbitq), 
to_sfixed(-903232616.0/4294967296.0,1,-nbitq), 
to_sfixed(-1405942680.0/4294967296.0,1,-nbitq), 
to_sfixed(-102924333.0/4294967296.0,1,-nbitq), 
to_sfixed(-765745335.0/4294967296.0,1,-nbitq), 
to_sfixed(-81586325.0/4294967296.0,1,-nbitq), 
to_sfixed(-239242648.0/4294967296.0,1,-nbitq), 
to_sfixed(1194138.0/4294967296.0,1,-nbitq), 
to_sfixed(9659730.0/4294967296.0,1,-nbitq), 
to_sfixed(-1600584.0/4294967296.0,1,-nbitq), 
to_sfixed(120361651.0/4294967296.0,1,-nbitq), 
to_sfixed(534438034.0/4294967296.0,1,-nbitq), 
to_sfixed(-1023348392.0/4294967296.0,1,-nbitq), 
to_sfixed(-167162032.0/4294967296.0,1,-nbitq), 
to_sfixed(-568555258.0/4294967296.0,1,-nbitq), 
to_sfixed(86799652.0/4294967296.0,1,-nbitq), 
to_sfixed(637334714.0/4294967296.0,1,-nbitq), 
to_sfixed(-501348197.0/4294967296.0,1,-nbitq), 
to_sfixed(-985559710.0/4294967296.0,1,-nbitq), 
to_sfixed(61817029.0/4294967296.0,1,-nbitq), 
to_sfixed(-210731134.0/4294967296.0,1,-nbitq), 
to_sfixed(134026797.0/4294967296.0,1,-nbitq), 
to_sfixed(429045847.0/4294967296.0,1,-nbitq), 
to_sfixed(-129509646.0/4294967296.0,1,-nbitq), 
to_sfixed(-452706819.0/4294967296.0,1,-nbitq), 
to_sfixed(123029003.0/4294967296.0,1,-nbitq), 
to_sfixed(-571932335.0/4294967296.0,1,-nbitq), 
to_sfixed(-438054814.0/4294967296.0,1,-nbitq), 
to_sfixed(451289165.0/4294967296.0,1,-nbitq), 
to_sfixed(327108135.0/4294967296.0,1,-nbitq), 
to_sfixed(401012792.0/4294967296.0,1,-nbitq), 
to_sfixed(-67213936.0/4294967296.0,1,-nbitq), 
to_sfixed(-1263725006.0/4294967296.0,1,-nbitq), 
to_sfixed(594772915.0/4294967296.0,1,-nbitq), 
to_sfixed(28914752.0/4294967296.0,1,-nbitq), 
to_sfixed(-323179371.0/4294967296.0,1,-nbitq), 
to_sfixed(965053140.0/4294967296.0,1,-nbitq), 
to_sfixed(-231647614.0/4294967296.0,1,-nbitq), 
to_sfixed(340417782.0/4294967296.0,1,-nbitq), 
to_sfixed(159786538.0/4294967296.0,1,-nbitq), 
to_sfixed(325900622.0/4294967296.0,1,-nbitq), 
to_sfixed(307042373.0/4294967296.0,1,-nbitq), 
to_sfixed(-566551967.0/4294967296.0,1,-nbitq), 
to_sfixed(-471891396.0/4294967296.0,1,-nbitq), 
to_sfixed(85856891.0/4294967296.0,1,-nbitq), 
to_sfixed(-108569691.0/4294967296.0,1,-nbitq), 
to_sfixed(206278635.0/4294967296.0,1,-nbitq), 
to_sfixed(333070263.0/4294967296.0,1,-nbitq), 
to_sfixed(200488078.0/4294967296.0,1,-nbitq), 
to_sfixed(-242679312.0/4294967296.0,1,-nbitq), 
to_sfixed(-266890721.0/4294967296.0,1,-nbitq), 
to_sfixed(299743414.0/4294967296.0,1,-nbitq), 
to_sfixed(437306481.0/4294967296.0,1,-nbitq), 
to_sfixed(56436140.0/4294967296.0,1,-nbitq), 
to_sfixed(-158355171.0/4294967296.0,1,-nbitq), 
to_sfixed(-1019685509.0/4294967296.0,1,-nbitq), 
to_sfixed(-875724489.0/4294967296.0,1,-nbitq), 
to_sfixed(129866207.0/4294967296.0,1,-nbitq), 
to_sfixed(-687559485.0/4294967296.0,1,-nbitq), 
to_sfixed(-888652511.0/4294967296.0,1,-nbitq), 
to_sfixed(-470119238.0/4294967296.0,1,-nbitq), 
to_sfixed(412569438.0/4294967296.0,1,-nbitq), 
to_sfixed(392140143.0/4294967296.0,1,-nbitq), 
to_sfixed(387762299.0/4294967296.0,1,-nbitq), 
to_sfixed(182438243.0/4294967296.0,1,-nbitq), 
to_sfixed(725562436.0/4294967296.0,1,-nbitq), 
to_sfixed(-65716474.0/4294967296.0,1,-nbitq), 
to_sfixed(219767089.0/4294967296.0,1,-nbitq), 
to_sfixed(117156929.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(19239205.0/4294967296.0,1,-nbitq), 
to_sfixed(-42864804.0/4294967296.0,1,-nbitq), 
to_sfixed(140649146.0/4294967296.0,1,-nbitq), 
to_sfixed(-324830517.0/4294967296.0,1,-nbitq), 
to_sfixed(344845519.0/4294967296.0,1,-nbitq), 
to_sfixed(306529496.0/4294967296.0,1,-nbitq), 
to_sfixed(-109465248.0/4294967296.0,1,-nbitq), 
to_sfixed(-364583333.0/4294967296.0,1,-nbitq), 
to_sfixed(189824496.0/4294967296.0,1,-nbitq), 
to_sfixed(209034397.0/4294967296.0,1,-nbitq), 
to_sfixed(862105208.0/4294967296.0,1,-nbitq), 
to_sfixed(569157751.0/4294967296.0,1,-nbitq), 
to_sfixed(-969278869.0/4294967296.0,1,-nbitq), 
to_sfixed(-1113056427.0/4294967296.0,1,-nbitq), 
to_sfixed(-93192823.0/4294967296.0,1,-nbitq), 
to_sfixed(-910287567.0/4294967296.0,1,-nbitq), 
to_sfixed(-272381989.0/4294967296.0,1,-nbitq), 
to_sfixed(-328071524.0/4294967296.0,1,-nbitq), 
to_sfixed(263200024.0/4294967296.0,1,-nbitq), 
to_sfixed(-111550818.0/4294967296.0,1,-nbitq), 
to_sfixed(-169897913.0/4294967296.0,1,-nbitq), 
to_sfixed(614234183.0/4294967296.0,1,-nbitq), 
to_sfixed(862628163.0/4294967296.0,1,-nbitq), 
to_sfixed(-425305246.0/4294967296.0,1,-nbitq), 
to_sfixed(-37584814.0/4294967296.0,1,-nbitq), 
to_sfixed(-855238657.0/4294967296.0,1,-nbitq), 
to_sfixed(-10378809.0/4294967296.0,1,-nbitq), 
to_sfixed(460429278.0/4294967296.0,1,-nbitq), 
to_sfixed(-637125066.0/4294967296.0,1,-nbitq), 
to_sfixed(-693350079.0/4294967296.0,1,-nbitq), 
to_sfixed(13510372.0/4294967296.0,1,-nbitq), 
to_sfixed(-584918614.0/4294967296.0,1,-nbitq), 
to_sfixed(-145846223.0/4294967296.0,1,-nbitq), 
to_sfixed(69234241.0/4294967296.0,1,-nbitq), 
to_sfixed(-394623082.0/4294967296.0,1,-nbitq), 
to_sfixed(-367709472.0/4294967296.0,1,-nbitq), 
to_sfixed(287049721.0/4294967296.0,1,-nbitq), 
to_sfixed(-578888628.0/4294967296.0,1,-nbitq), 
to_sfixed(-7102824.0/4294967296.0,1,-nbitq), 
to_sfixed(239726455.0/4294967296.0,1,-nbitq), 
to_sfixed(16743693.0/4294967296.0,1,-nbitq), 
to_sfixed(581163568.0/4294967296.0,1,-nbitq), 
to_sfixed(584691979.0/4294967296.0,1,-nbitq), 
to_sfixed(-1119343936.0/4294967296.0,1,-nbitq), 
to_sfixed(233319665.0/4294967296.0,1,-nbitq), 
to_sfixed(695456713.0/4294967296.0,1,-nbitq), 
to_sfixed(-241717185.0/4294967296.0,1,-nbitq), 
to_sfixed(828443023.0/4294967296.0,1,-nbitq), 
to_sfixed(-414759385.0/4294967296.0,1,-nbitq), 
to_sfixed(201588638.0/4294967296.0,1,-nbitq), 
to_sfixed(-245751874.0/4294967296.0,1,-nbitq), 
to_sfixed(225187553.0/4294967296.0,1,-nbitq), 
to_sfixed(-52491091.0/4294967296.0,1,-nbitq), 
to_sfixed(-1138139326.0/4294967296.0,1,-nbitq), 
to_sfixed(113891536.0/4294967296.0,1,-nbitq), 
to_sfixed(-112771282.0/4294967296.0,1,-nbitq), 
to_sfixed(-307935447.0/4294967296.0,1,-nbitq), 
to_sfixed(207576346.0/4294967296.0,1,-nbitq), 
to_sfixed(402016323.0/4294967296.0,1,-nbitq), 
to_sfixed(-256336483.0/4294967296.0,1,-nbitq), 
to_sfixed(67712494.0/4294967296.0,1,-nbitq), 
to_sfixed(-520172783.0/4294967296.0,1,-nbitq), 
to_sfixed(535324963.0/4294967296.0,1,-nbitq), 
to_sfixed(-186275446.0/4294967296.0,1,-nbitq), 
to_sfixed(-118762677.0/4294967296.0,1,-nbitq), 
to_sfixed(8846789.0/4294967296.0,1,-nbitq), 
to_sfixed(-503850773.0/4294967296.0,1,-nbitq), 
to_sfixed(-763398980.0/4294967296.0,1,-nbitq), 
to_sfixed(-305044009.0/4294967296.0,1,-nbitq), 
to_sfixed(-543680075.0/4294967296.0,1,-nbitq), 
to_sfixed(-345112812.0/4294967296.0,1,-nbitq), 
to_sfixed(-325101032.0/4294967296.0,1,-nbitq), 
to_sfixed(-10172243.0/4294967296.0,1,-nbitq), 
to_sfixed(213791995.0/4294967296.0,1,-nbitq), 
to_sfixed(182796985.0/4294967296.0,1,-nbitq), 
to_sfixed(-234055234.0/4294967296.0,1,-nbitq), 
to_sfixed(454576504.0/4294967296.0,1,-nbitq), 
to_sfixed(-20196679.0/4294967296.0,1,-nbitq), 
to_sfixed(72423745.0/4294967296.0,1,-nbitq), 
to_sfixed(248856678.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(242282527.0/4294967296.0,1,-nbitq), 
to_sfixed(-667175149.0/4294967296.0,1,-nbitq), 
to_sfixed(491797224.0/4294967296.0,1,-nbitq), 
to_sfixed(-747643881.0/4294967296.0,1,-nbitq), 
to_sfixed(265967857.0/4294967296.0,1,-nbitq), 
to_sfixed(-75062170.0/4294967296.0,1,-nbitq), 
to_sfixed(-84934023.0/4294967296.0,1,-nbitq), 
to_sfixed(110652465.0/4294967296.0,1,-nbitq), 
to_sfixed(879310673.0/4294967296.0,1,-nbitq), 
to_sfixed(-1915265.0/4294967296.0,1,-nbitq), 
to_sfixed(-129417573.0/4294967296.0,1,-nbitq), 
to_sfixed(158518724.0/4294967296.0,1,-nbitq), 
to_sfixed(-958244584.0/4294967296.0,1,-nbitq), 
to_sfixed(-779854149.0/4294967296.0,1,-nbitq), 
to_sfixed(-99281513.0/4294967296.0,1,-nbitq), 
to_sfixed(-549643739.0/4294967296.0,1,-nbitq), 
to_sfixed(340798445.0/4294967296.0,1,-nbitq), 
to_sfixed(-176135778.0/4294967296.0,1,-nbitq), 
to_sfixed(37699717.0/4294967296.0,1,-nbitq), 
to_sfixed(-127401023.0/4294967296.0,1,-nbitq), 
to_sfixed(-103512041.0/4294967296.0,1,-nbitq), 
to_sfixed(867848149.0/4294967296.0,1,-nbitq), 
to_sfixed(503361902.0/4294967296.0,1,-nbitq), 
to_sfixed(-384076307.0/4294967296.0,1,-nbitq), 
to_sfixed(-201536987.0/4294967296.0,1,-nbitq), 
to_sfixed(-859457229.0/4294967296.0,1,-nbitq), 
to_sfixed(304072101.0/4294967296.0,1,-nbitq), 
to_sfixed(384132855.0/4294967296.0,1,-nbitq), 
to_sfixed(-676495423.0/4294967296.0,1,-nbitq), 
to_sfixed(-840299473.0/4294967296.0,1,-nbitq), 
to_sfixed(251885828.0/4294967296.0,1,-nbitq), 
to_sfixed(113255377.0/4294967296.0,1,-nbitq), 
to_sfixed(290326661.0/4294967296.0,1,-nbitq), 
to_sfixed(416584619.0/4294967296.0,1,-nbitq), 
to_sfixed(-142499325.0/4294967296.0,1,-nbitq), 
to_sfixed(168696626.0/4294967296.0,1,-nbitq), 
to_sfixed(195456742.0/4294967296.0,1,-nbitq), 
to_sfixed(-914507859.0/4294967296.0,1,-nbitq), 
to_sfixed(-362462890.0/4294967296.0,1,-nbitq), 
to_sfixed(625220316.0/4294967296.0,1,-nbitq), 
to_sfixed(59790077.0/4294967296.0,1,-nbitq), 
to_sfixed(87247137.0/4294967296.0,1,-nbitq), 
to_sfixed(112286149.0/4294967296.0,1,-nbitq), 
to_sfixed(-547711821.0/4294967296.0,1,-nbitq), 
to_sfixed(406329226.0/4294967296.0,1,-nbitq), 
to_sfixed(1135046618.0/4294967296.0,1,-nbitq), 
to_sfixed(-387227917.0/4294967296.0,1,-nbitq), 
to_sfixed(13472921.0/4294967296.0,1,-nbitq), 
to_sfixed(-339257129.0/4294967296.0,1,-nbitq), 
to_sfixed(-223356660.0/4294967296.0,1,-nbitq), 
to_sfixed(-209233918.0/4294967296.0,1,-nbitq), 
to_sfixed(229660712.0/4294967296.0,1,-nbitq), 
to_sfixed(-283823889.0/4294967296.0,1,-nbitq), 
to_sfixed(-869328369.0/4294967296.0,1,-nbitq), 
to_sfixed(-80363076.0/4294967296.0,1,-nbitq), 
to_sfixed(-12488467.0/4294967296.0,1,-nbitq), 
to_sfixed(109880283.0/4294967296.0,1,-nbitq), 
to_sfixed(167515734.0/4294967296.0,1,-nbitq), 
to_sfixed(-250991030.0/4294967296.0,1,-nbitq), 
to_sfixed(-45407721.0/4294967296.0,1,-nbitq), 
to_sfixed(-345093119.0/4294967296.0,1,-nbitq), 
to_sfixed(-395721024.0/4294967296.0,1,-nbitq), 
to_sfixed(873751847.0/4294967296.0,1,-nbitq), 
to_sfixed(-503439942.0/4294967296.0,1,-nbitq), 
to_sfixed(-108694432.0/4294967296.0,1,-nbitq), 
to_sfixed(167116645.0/4294967296.0,1,-nbitq), 
to_sfixed(-216252496.0/4294967296.0,1,-nbitq), 
to_sfixed(-798775925.0/4294967296.0,1,-nbitq), 
to_sfixed(256168005.0/4294967296.0,1,-nbitq), 
to_sfixed(-372046917.0/4294967296.0,1,-nbitq), 
to_sfixed(-775496819.0/4294967296.0,1,-nbitq), 
to_sfixed(-107146270.0/4294967296.0,1,-nbitq), 
to_sfixed(512477172.0/4294967296.0,1,-nbitq), 
to_sfixed(366726989.0/4294967296.0,1,-nbitq), 
to_sfixed(580816192.0/4294967296.0,1,-nbitq), 
to_sfixed(15880422.0/4294967296.0,1,-nbitq), 
to_sfixed(531686049.0/4294967296.0,1,-nbitq), 
to_sfixed(440754028.0/4294967296.0,1,-nbitq), 
to_sfixed(482686684.0/4294967296.0,1,-nbitq), 
to_sfixed(274534343.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-168945717.0/4294967296.0,1,-nbitq), 
to_sfixed(-287769509.0/4294967296.0,1,-nbitq), 
to_sfixed(932005914.0/4294967296.0,1,-nbitq), 
to_sfixed(-690778500.0/4294967296.0,1,-nbitq), 
to_sfixed(763836991.0/4294967296.0,1,-nbitq), 
to_sfixed(-360088691.0/4294967296.0,1,-nbitq), 
to_sfixed(-341385252.0/4294967296.0,1,-nbitq), 
to_sfixed(182899916.0/4294967296.0,1,-nbitq), 
to_sfixed(666569821.0/4294967296.0,1,-nbitq), 
to_sfixed(-157530530.0/4294967296.0,1,-nbitq), 
to_sfixed(-258233650.0/4294967296.0,1,-nbitq), 
to_sfixed(-369263581.0/4294967296.0,1,-nbitq), 
to_sfixed(-337165309.0/4294967296.0,1,-nbitq), 
to_sfixed(163019417.0/4294967296.0,1,-nbitq), 
to_sfixed(196473143.0/4294967296.0,1,-nbitq), 
to_sfixed(-304158287.0/4294967296.0,1,-nbitq), 
to_sfixed(-106567588.0/4294967296.0,1,-nbitq), 
to_sfixed(-349252608.0/4294967296.0,1,-nbitq), 
to_sfixed(832618381.0/4294967296.0,1,-nbitq), 
to_sfixed(129555323.0/4294967296.0,1,-nbitq), 
to_sfixed(-81395561.0/4294967296.0,1,-nbitq), 
to_sfixed(731107165.0/4294967296.0,1,-nbitq), 
to_sfixed(672747805.0/4294967296.0,1,-nbitq), 
to_sfixed(-513679725.0/4294967296.0,1,-nbitq), 
to_sfixed(-321299375.0/4294967296.0,1,-nbitq), 
to_sfixed(-487650960.0/4294967296.0,1,-nbitq), 
to_sfixed(-287411244.0/4294967296.0,1,-nbitq), 
to_sfixed(343220309.0/4294967296.0,1,-nbitq), 
to_sfixed(-199071741.0/4294967296.0,1,-nbitq), 
to_sfixed(-738877127.0/4294967296.0,1,-nbitq), 
to_sfixed(-57841762.0/4294967296.0,1,-nbitq), 
to_sfixed(273010033.0/4294967296.0,1,-nbitq), 
to_sfixed(421769543.0/4294967296.0,1,-nbitq), 
to_sfixed(419296094.0/4294967296.0,1,-nbitq), 
to_sfixed(-125346802.0/4294967296.0,1,-nbitq), 
to_sfixed(-198352463.0/4294967296.0,1,-nbitq), 
to_sfixed(85286263.0/4294967296.0,1,-nbitq), 
to_sfixed(-157715687.0/4294967296.0,1,-nbitq), 
to_sfixed(-26812404.0/4294967296.0,1,-nbitq), 
to_sfixed(505076151.0/4294967296.0,1,-nbitq), 
to_sfixed(-152434462.0/4294967296.0,1,-nbitq), 
to_sfixed(182856357.0/4294967296.0,1,-nbitq), 
to_sfixed(-92188807.0/4294967296.0,1,-nbitq), 
to_sfixed(-83776886.0/4294967296.0,1,-nbitq), 
to_sfixed(683313009.0/4294967296.0,1,-nbitq), 
to_sfixed(302463726.0/4294967296.0,1,-nbitq), 
to_sfixed(43044902.0/4294967296.0,1,-nbitq), 
to_sfixed(-402898136.0/4294967296.0,1,-nbitq), 
to_sfixed(-193775142.0/4294967296.0,1,-nbitq), 
to_sfixed(-156536679.0/4294967296.0,1,-nbitq), 
to_sfixed(-261632361.0/4294967296.0,1,-nbitq), 
to_sfixed(110237946.0/4294967296.0,1,-nbitq), 
to_sfixed(-219341730.0/4294967296.0,1,-nbitq), 
to_sfixed(-71644148.0/4294967296.0,1,-nbitq), 
to_sfixed(16704591.0/4294967296.0,1,-nbitq), 
to_sfixed(-350716883.0/4294967296.0,1,-nbitq), 
to_sfixed(-122177956.0/4294967296.0,1,-nbitq), 
to_sfixed(401953303.0/4294967296.0,1,-nbitq), 
to_sfixed(-344872894.0/4294967296.0,1,-nbitq), 
to_sfixed(-274231482.0/4294967296.0,1,-nbitq), 
to_sfixed(-351036994.0/4294967296.0,1,-nbitq), 
to_sfixed(254385603.0/4294967296.0,1,-nbitq), 
to_sfixed(307536130.0/4294967296.0,1,-nbitq), 
to_sfixed(-42390565.0/4294967296.0,1,-nbitq), 
to_sfixed(-185711528.0/4294967296.0,1,-nbitq), 
to_sfixed(-14122674.0/4294967296.0,1,-nbitq), 
to_sfixed(-26557566.0/4294967296.0,1,-nbitq), 
to_sfixed(-939187883.0/4294967296.0,1,-nbitq), 
to_sfixed(-133176530.0/4294967296.0,1,-nbitq), 
to_sfixed(-468609428.0/4294967296.0,1,-nbitq), 
to_sfixed(-434464062.0/4294967296.0,1,-nbitq), 
to_sfixed(-193032173.0/4294967296.0,1,-nbitq), 
to_sfixed(690243939.0/4294967296.0,1,-nbitq), 
to_sfixed(118097179.0/4294967296.0,1,-nbitq), 
to_sfixed(480165133.0/4294967296.0,1,-nbitq), 
to_sfixed(110750242.0/4294967296.0,1,-nbitq), 
to_sfixed(773686511.0/4294967296.0,1,-nbitq), 
to_sfixed(61021448.0/4294967296.0,1,-nbitq), 
to_sfixed(101740590.0/4294967296.0,1,-nbitq), 
to_sfixed(-276069360.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(87836380.0/4294967296.0,1,-nbitq), 
to_sfixed(-386325792.0/4294967296.0,1,-nbitq), 
to_sfixed(474689053.0/4294967296.0,1,-nbitq), 
to_sfixed(-224650244.0/4294967296.0,1,-nbitq), 
to_sfixed(454768835.0/4294967296.0,1,-nbitq), 
to_sfixed(-510369692.0/4294967296.0,1,-nbitq), 
to_sfixed(-21996126.0/4294967296.0,1,-nbitq), 
to_sfixed(-414482310.0/4294967296.0,1,-nbitq), 
to_sfixed(498557560.0/4294967296.0,1,-nbitq), 
to_sfixed(2091091.0/4294967296.0,1,-nbitq), 
to_sfixed(-344450612.0/4294967296.0,1,-nbitq), 
to_sfixed(-241470278.0/4294967296.0,1,-nbitq), 
to_sfixed(-691882509.0/4294967296.0,1,-nbitq), 
to_sfixed(-239520054.0/4294967296.0,1,-nbitq), 
to_sfixed(122812347.0/4294967296.0,1,-nbitq), 
to_sfixed(-537048675.0/4294967296.0,1,-nbitq), 
to_sfixed(-174154427.0/4294967296.0,1,-nbitq), 
to_sfixed(209076351.0/4294967296.0,1,-nbitq), 
to_sfixed(250583661.0/4294967296.0,1,-nbitq), 
to_sfixed(18834871.0/4294967296.0,1,-nbitq), 
to_sfixed(-72199467.0/4294967296.0,1,-nbitq), 
to_sfixed(513722888.0/4294967296.0,1,-nbitq), 
to_sfixed(106535153.0/4294967296.0,1,-nbitq), 
to_sfixed(-436032037.0/4294967296.0,1,-nbitq), 
to_sfixed(285749429.0/4294967296.0,1,-nbitq), 
to_sfixed(-311489368.0/4294967296.0,1,-nbitq), 
to_sfixed(-53961323.0/4294967296.0,1,-nbitq), 
to_sfixed(-169345956.0/4294967296.0,1,-nbitq), 
to_sfixed(-515937607.0/4294967296.0,1,-nbitq), 
to_sfixed(-266642536.0/4294967296.0,1,-nbitq), 
to_sfixed(-212435320.0/4294967296.0,1,-nbitq), 
to_sfixed(339604363.0/4294967296.0,1,-nbitq), 
to_sfixed(-57064972.0/4294967296.0,1,-nbitq), 
to_sfixed(299677119.0/4294967296.0,1,-nbitq), 
to_sfixed(-332758941.0/4294967296.0,1,-nbitq), 
to_sfixed(-551730166.0/4294967296.0,1,-nbitq), 
to_sfixed(325484310.0/4294967296.0,1,-nbitq), 
to_sfixed(-244422696.0/4294967296.0,1,-nbitq), 
to_sfixed(163660614.0/4294967296.0,1,-nbitq), 
to_sfixed(303489677.0/4294967296.0,1,-nbitq), 
to_sfixed(370671393.0/4294967296.0,1,-nbitq), 
to_sfixed(-126451872.0/4294967296.0,1,-nbitq), 
to_sfixed(398167387.0/4294967296.0,1,-nbitq), 
to_sfixed(226319920.0/4294967296.0,1,-nbitq), 
to_sfixed(73432562.0/4294967296.0,1,-nbitq), 
to_sfixed(356156845.0/4294967296.0,1,-nbitq), 
to_sfixed(-435430333.0/4294967296.0,1,-nbitq), 
to_sfixed(144609153.0/4294967296.0,1,-nbitq), 
to_sfixed(362819463.0/4294967296.0,1,-nbitq), 
to_sfixed(-663129827.0/4294967296.0,1,-nbitq), 
to_sfixed(229464117.0/4294967296.0,1,-nbitq), 
to_sfixed(-475700415.0/4294967296.0,1,-nbitq), 
to_sfixed(-432733701.0/4294967296.0,1,-nbitq), 
to_sfixed(-356840841.0/4294967296.0,1,-nbitq), 
to_sfixed(-34072143.0/4294967296.0,1,-nbitq), 
to_sfixed(-667417785.0/4294967296.0,1,-nbitq), 
to_sfixed(-232948933.0/4294967296.0,1,-nbitq), 
to_sfixed(73524687.0/4294967296.0,1,-nbitq), 
to_sfixed(75079799.0/4294967296.0,1,-nbitq), 
to_sfixed(-320308541.0/4294967296.0,1,-nbitq), 
to_sfixed(-57438115.0/4294967296.0,1,-nbitq), 
to_sfixed(-321500291.0/4294967296.0,1,-nbitq), 
to_sfixed(503262045.0/4294967296.0,1,-nbitq), 
to_sfixed(-154717198.0/4294967296.0,1,-nbitq), 
to_sfixed(152816515.0/4294967296.0,1,-nbitq), 
to_sfixed(-415671184.0/4294967296.0,1,-nbitq), 
to_sfixed(75455543.0/4294967296.0,1,-nbitq), 
to_sfixed(-678009102.0/4294967296.0,1,-nbitq), 
to_sfixed(-222404451.0/4294967296.0,1,-nbitq), 
to_sfixed(-171915103.0/4294967296.0,1,-nbitq), 
to_sfixed(79375206.0/4294967296.0,1,-nbitq), 
to_sfixed(408271509.0/4294967296.0,1,-nbitq), 
to_sfixed(-61303445.0/4294967296.0,1,-nbitq), 
to_sfixed(351351802.0/4294967296.0,1,-nbitq), 
to_sfixed(149959.0/4294967296.0,1,-nbitq), 
to_sfixed(-515476803.0/4294967296.0,1,-nbitq), 
to_sfixed(725936839.0/4294967296.0,1,-nbitq), 
to_sfixed(351685654.0/4294967296.0,1,-nbitq), 
to_sfixed(23926528.0/4294967296.0,1,-nbitq), 
to_sfixed(41368037.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(26344721.0/4294967296.0,1,-nbitq), 
to_sfixed(-508767357.0/4294967296.0,1,-nbitq), 
to_sfixed(-292556279.0/4294967296.0,1,-nbitq), 
to_sfixed(-31513768.0/4294967296.0,1,-nbitq), 
to_sfixed(491888420.0/4294967296.0,1,-nbitq), 
to_sfixed(-523861854.0/4294967296.0,1,-nbitq), 
to_sfixed(-297324375.0/4294967296.0,1,-nbitq), 
to_sfixed(-423713031.0/4294967296.0,1,-nbitq), 
to_sfixed(597452453.0/4294967296.0,1,-nbitq), 
to_sfixed(-91400877.0/4294967296.0,1,-nbitq), 
to_sfixed(-169451617.0/4294967296.0,1,-nbitq), 
to_sfixed(-305636696.0/4294967296.0,1,-nbitq), 
to_sfixed(-261108691.0/4294967296.0,1,-nbitq), 
to_sfixed(-87197168.0/4294967296.0,1,-nbitq), 
to_sfixed(35748583.0/4294967296.0,1,-nbitq), 
to_sfixed(-316619420.0/4294967296.0,1,-nbitq), 
to_sfixed(-386894001.0/4294967296.0,1,-nbitq), 
to_sfixed(-310915471.0/4294967296.0,1,-nbitq), 
to_sfixed(501077166.0/4294967296.0,1,-nbitq), 
to_sfixed(203065612.0/4294967296.0,1,-nbitq), 
to_sfixed(125381231.0/4294967296.0,1,-nbitq), 
to_sfixed(-118500666.0/4294967296.0,1,-nbitq), 
to_sfixed(398948850.0/4294967296.0,1,-nbitq), 
to_sfixed(-173403867.0/4294967296.0,1,-nbitq), 
to_sfixed(268814832.0/4294967296.0,1,-nbitq), 
to_sfixed(-176109502.0/4294967296.0,1,-nbitq), 
to_sfixed(134618484.0/4294967296.0,1,-nbitq), 
to_sfixed(150422523.0/4294967296.0,1,-nbitq), 
to_sfixed(-318799024.0/4294967296.0,1,-nbitq), 
to_sfixed(-312099248.0/4294967296.0,1,-nbitq), 
to_sfixed(-161737373.0/4294967296.0,1,-nbitq), 
to_sfixed(76405741.0/4294967296.0,1,-nbitq), 
to_sfixed(38877246.0/4294967296.0,1,-nbitq), 
to_sfixed(105945560.0/4294967296.0,1,-nbitq), 
to_sfixed(110775459.0/4294967296.0,1,-nbitq), 
to_sfixed(-319531612.0/4294967296.0,1,-nbitq), 
to_sfixed(-90780126.0/4294967296.0,1,-nbitq), 
to_sfixed(-306577518.0/4294967296.0,1,-nbitq), 
to_sfixed(76170157.0/4294967296.0,1,-nbitq), 
to_sfixed(302912624.0/4294967296.0,1,-nbitq), 
to_sfixed(-46231057.0/4294967296.0,1,-nbitq), 
to_sfixed(258028547.0/4294967296.0,1,-nbitq), 
to_sfixed(485085247.0/4294967296.0,1,-nbitq), 
to_sfixed(267505315.0/4294967296.0,1,-nbitq), 
to_sfixed(426133326.0/4294967296.0,1,-nbitq), 
to_sfixed(321816171.0/4294967296.0,1,-nbitq), 
to_sfixed(-64330786.0/4294967296.0,1,-nbitq), 
to_sfixed(234153216.0/4294967296.0,1,-nbitq), 
to_sfixed(-424668389.0/4294967296.0,1,-nbitq), 
to_sfixed(-746881600.0/4294967296.0,1,-nbitq), 
to_sfixed(-230787441.0/4294967296.0,1,-nbitq), 
to_sfixed(-287503253.0/4294967296.0,1,-nbitq), 
to_sfixed(-615393968.0/4294967296.0,1,-nbitq), 
to_sfixed(-65453150.0/4294967296.0,1,-nbitq), 
to_sfixed(118467282.0/4294967296.0,1,-nbitq), 
to_sfixed(25378246.0/4294967296.0,1,-nbitq), 
to_sfixed(-580563152.0/4294967296.0,1,-nbitq), 
to_sfixed(477853101.0/4294967296.0,1,-nbitq), 
to_sfixed(-153210649.0/4294967296.0,1,-nbitq), 
to_sfixed(260912210.0/4294967296.0,1,-nbitq), 
to_sfixed(168148604.0/4294967296.0,1,-nbitq), 
to_sfixed(104318376.0/4294967296.0,1,-nbitq), 
to_sfixed(798999506.0/4294967296.0,1,-nbitq), 
to_sfixed(-257546266.0/4294967296.0,1,-nbitq), 
to_sfixed(-54353700.0/4294967296.0,1,-nbitq), 
to_sfixed(-168865378.0/4294967296.0,1,-nbitq), 
to_sfixed(-336437468.0/4294967296.0,1,-nbitq), 
to_sfixed(-126362585.0/4294967296.0,1,-nbitq), 
to_sfixed(-224164417.0/4294967296.0,1,-nbitq), 
to_sfixed(-179017562.0/4294967296.0,1,-nbitq), 
to_sfixed(180672901.0/4294967296.0,1,-nbitq), 
to_sfixed(43656518.0/4294967296.0,1,-nbitq), 
to_sfixed(13417230.0/4294967296.0,1,-nbitq), 
to_sfixed(-192006156.0/4294967296.0,1,-nbitq), 
to_sfixed(455574442.0/4294967296.0,1,-nbitq), 
to_sfixed(106517287.0/4294967296.0,1,-nbitq), 
to_sfixed(825378505.0/4294967296.0,1,-nbitq), 
to_sfixed(-35762856.0/4294967296.0,1,-nbitq), 
to_sfixed(-522772015.0/4294967296.0,1,-nbitq), 
to_sfixed(-260525102.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-282282137.0/4294967296.0,1,-nbitq), 
to_sfixed(-85486806.0/4294967296.0,1,-nbitq), 
to_sfixed(512885632.0/4294967296.0,1,-nbitq), 
to_sfixed(399634042.0/4294967296.0,1,-nbitq), 
to_sfixed(187668823.0/4294967296.0,1,-nbitq), 
to_sfixed(-1191340620.0/4294967296.0,1,-nbitq), 
to_sfixed(-281074786.0/4294967296.0,1,-nbitq), 
to_sfixed(-144105219.0/4294967296.0,1,-nbitq), 
to_sfixed(1036178362.0/4294967296.0,1,-nbitq), 
to_sfixed(-92657185.0/4294967296.0,1,-nbitq), 
to_sfixed(-324677765.0/4294967296.0,1,-nbitq), 
to_sfixed(-22655333.0/4294967296.0,1,-nbitq), 
to_sfixed(-293369146.0/4294967296.0,1,-nbitq), 
to_sfixed(454788479.0/4294967296.0,1,-nbitq), 
to_sfixed(331541479.0/4294967296.0,1,-nbitq), 
to_sfixed(-573037463.0/4294967296.0,1,-nbitq), 
to_sfixed(-382836637.0/4294967296.0,1,-nbitq), 
to_sfixed(-355749605.0/4294967296.0,1,-nbitq), 
to_sfixed(-149771200.0/4294967296.0,1,-nbitq), 
to_sfixed(99089658.0/4294967296.0,1,-nbitq), 
to_sfixed(68157157.0/4294967296.0,1,-nbitq), 
to_sfixed(-23538489.0/4294967296.0,1,-nbitq), 
to_sfixed(125073131.0/4294967296.0,1,-nbitq), 
to_sfixed(-460112082.0/4294967296.0,1,-nbitq), 
to_sfixed(98612531.0/4294967296.0,1,-nbitq), 
to_sfixed(-51105733.0/4294967296.0,1,-nbitq), 
to_sfixed(-186641145.0/4294967296.0,1,-nbitq), 
to_sfixed(-479252086.0/4294967296.0,1,-nbitq), 
to_sfixed(-84916631.0/4294967296.0,1,-nbitq), 
to_sfixed(-1004360142.0/4294967296.0,1,-nbitq), 
to_sfixed(-484788759.0/4294967296.0,1,-nbitq), 
to_sfixed(61819648.0/4294967296.0,1,-nbitq), 
to_sfixed(-103864546.0/4294967296.0,1,-nbitq), 
to_sfixed(-282510952.0/4294967296.0,1,-nbitq), 
to_sfixed(-46613928.0/4294967296.0,1,-nbitq), 
to_sfixed(-233356780.0/4294967296.0,1,-nbitq), 
to_sfixed(386380644.0/4294967296.0,1,-nbitq), 
to_sfixed(-276492762.0/4294967296.0,1,-nbitq), 
to_sfixed(-39104071.0/4294967296.0,1,-nbitq), 
to_sfixed(440931177.0/4294967296.0,1,-nbitq), 
to_sfixed(402631965.0/4294967296.0,1,-nbitq), 
to_sfixed(285253283.0/4294967296.0,1,-nbitq), 
to_sfixed(474166406.0/4294967296.0,1,-nbitq), 
to_sfixed(-146097103.0/4294967296.0,1,-nbitq), 
to_sfixed(368662859.0/4294967296.0,1,-nbitq), 
to_sfixed(716739040.0/4294967296.0,1,-nbitq), 
to_sfixed(126408850.0/4294967296.0,1,-nbitq), 
to_sfixed(-158474982.0/4294967296.0,1,-nbitq), 
to_sfixed(-125768289.0/4294967296.0,1,-nbitq), 
to_sfixed(-78667834.0/4294967296.0,1,-nbitq), 
to_sfixed(171597565.0/4294967296.0,1,-nbitq), 
to_sfixed(-73988620.0/4294967296.0,1,-nbitq), 
to_sfixed(-428062342.0/4294967296.0,1,-nbitq), 
to_sfixed(-125400206.0/4294967296.0,1,-nbitq), 
to_sfixed(-332891052.0/4294967296.0,1,-nbitq), 
to_sfixed(-337255542.0/4294967296.0,1,-nbitq), 
to_sfixed(-726093240.0/4294967296.0,1,-nbitq), 
to_sfixed(6318569.0/4294967296.0,1,-nbitq), 
to_sfixed(-53072630.0/4294967296.0,1,-nbitq), 
to_sfixed(360814674.0/4294967296.0,1,-nbitq), 
to_sfixed(344077206.0/4294967296.0,1,-nbitq), 
to_sfixed(264244435.0/4294967296.0,1,-nbitq), 
to_sfixed(-84045864.0/4294967296.0,1,-nbitq), 
to_sfixed(-118809.0/4294967296.0,1,-nbitq), 
to_sfixed(-346615847.0/4294967296.0,1,-nbitq), 
to_sfixed(-435063704.0/4294967296.0,1,-nbitq), 
to_sfixed(-101992725.0/4294967296.0,1,-nbitq), 
to_sfixed(-303776453.0/4294967296.0,1,-nbitq), 
to_sfixed(-319454101.0/4294967296.0,1,-nbitq), 
to_sfixed(-17986571.0/4294967296.0,1,-nbitq), 
to_sfixed(-79157004.0/4294967296.0,1,-nbitq), 
to_sfixed(-119096679.0/4294967296.0,1,-nbitq), 
to_sfixed(-69705311.0/4294967296.0,1,-nbitq), 
to_sfixed(123839200.0/4294967296.0,1,-nbitq), 
to_sfixed(-8559996.0/4294967296.0,1,-nbitq), 
to_sfixed(375266378.0/4294967296.0,1,-nbitq), 
to_sfixed(967297107.0/4294967296.0,1,-nbitq), 
to_sfixed(-236065036.0/4294967296.0,1,-nbitq), 
to_sfixed(-192261223.0/4294967296.0,1,-nbitq), 
to_sfixed(128840897.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(434081214.0/4294967296.0,1,-nbitq), 
to_sfixed(-603736741.0/4294967296.0,1,-nbitq), 
to_sfixed(622679494.0/4294967296.0,1,-nbitq), 
to_sfixed(308721420.0/4294967296.0,1,-nbitq), 
to_sfixed(519431446.0/4294967296.0,1,-nbitq), 
to_sfixed(-393330785.0/4294967296.0,1,-nbitq), 
to_sfixed(33786632.0/4294967296.0,1,-nbitq), 
to_sfixed(-240804238.0/4294967296.0,1,-nbitq), 
to_sfixed(741227283.0/4294967296.0,1,-nbitq), 
to_sfixed(256853409.0/4294967296.0,1,-nbitq), 
to_sfixed(243741855.0/4294967296.0,1,-nbitq), 
to_sfixed(-184740510.0/4294967296.0,1,-nbitq), 
to_sfixed(-894846551.0/4294967296.0,1,-nbitq), 
to_sfixed(-206082069.0/4294967296.0,1,-nbitq), 
to_sfixed(322716379.0/4294967296.0,1,-nbitq), 
to_sfixed(93311481.0/4294967296.0,1,-nbitq), 
to_sfixed(200849454.0/4294967296.0,1,-nbitq), 
to_sfixed(112034078.0/4294967296.0,1,-nbitq), 
to_sfixed(-332198960.0/4294967296.0,1,-nbitq), 
to_sfixed(-63380825.0/4294967296.0,1,-nbitq), 
to_sfixed(39031189.0/4294967296.0,1,-nbitq), 
to_sfixed(560671648.0/4294967296.0,1,-nbitq), 
to_sfixed(334890812.0/4294967296.0,1,-nbitq), 
to_sfixed(239013243.0/4294967296.0,1,-nbitq), 
to_sfixed(62059628.0/4294967296.0,1,-nbitq), 
to_sfixed(-614187038.0/4294967296.0,1,-nbitq), 
to_sfixed(223578369.0/4294967296.0,1,-nbitq), 
to_sfixed(-491722546.0/4294967296.0,1,-nbitq), 
to_sfixed(291158335.0/4294967296.0,1,-nbitq), 
to_sfixed(-430845399.0/4294967296.0,1,-nbitq), 
to_sfixed(-612080553.0/4294967296.0,1,-nbitq), 
to_sfixed(235863896.0/4294967296.0,1,-nbitq), 
to_sfixed(-140839379.0/4294967296.0,1,-nbitq), 
to_sfixed(292426943.0/4294967296.0,1,-nbitq), 
to_sfixed(252810378.0/4294967296.0,1,-nbitq), 
to_sfixed(155661093.0/4294967296.0,1,-nbitq), 
to_sfixed(58901416.0/4294967296.0,1,-nbitq), 
to_sfixed(231266521.0/4294967296.0,1,-nbitq), 
to_sfixed(25051262.0/4294967296.0,1,-nbitq), 
to_sfixed(-39774829.0/4294967296.0,1,-nbitq), 
to_sfixed(189470787.0/4294967296.0,1,-nbitq), 
to_sfixed(561720053.0/4294967296.0,1,-nbitq), 
to_sfixed(62497220.0/4294967296.0,1,-nbitq), 
to_sfixed(587733214.0/4294967296.0,1,-nbitq), 
to_sfixed(47699917.0/4294967296.0,1,-nbitq), 
to_sfixed(223488224.0/4294967296.0,1,-nbitq), 
to_sfixed(100719294.0/4294967296.0,1,-nbitq), 
to_sfixed(-419281822.0/4294967296.0,1,-nbitq), 
to_sfixed(-251915439.0/4294967296.0,1,-nbitq), 
to_sfixed(-163078554.0/4294967296.0,1,-nbitq), 
to_sfixed(-470433737.0/4294967296.0,1,-nbitq), 
to_sfixed(307597618.0/4294967296.0,1,-nbitq), 
to_sfixed(-337053521.0/4294967296.0,1,-nbitq), 
to_sfixed(263978822.0/4294967296.0,1,-nbitq), 
to_sfixed(311432759.0/4294967296.0,1,-nbitq), 
to_sfixed(437374197.0/4294967296.0,1,-nbitq), 
to_sfixed(-260519769.0/4294967296.0,1,-nbitq), 
to_sfixed(1132658.0/4294967296.0,1,-nbitq), 
to_sfixed(-316185224.0/4294967296.0,1,-nbitq), 
to_sfixed(-125064466.0/4294967296.0,1,-nbitq), 
to_sfixed(364287058.0/4294967296.0,1,-nbitq), 
to_sfixed(-227510598.0/4294967296.0,1,-nbitq), 
to_sfixed(297305841.0/4294967296.0,1,-nbitq), 
to_sfixed(282841748.0/4294967296.0,1,-nbitq), 
to_sfixed(345168233.0/4294967296.0,1,-nbitq), 
to_sfixed(338884337.0/4294967296.0,1,-nbitq), 
to_sfixed(453442989.0/4294967296.0,1,-nbitq), 
to_sfixed(-474650004.0/4294967296.0,1,-nbitq), 
to_sfixed(34191430.0/4294967296.0,1,-nbitq), 
to_sfixed(-637914494.0/4294967296.0,1,-nbitq), 
to_sfixed(429894045.0/4294967296.0,1,-nbitq), 
to_sfixed(486672354.0/4294967296.0,1,-nbitq), 
to_sfixed(-211145634.0/4294967296.0,1,-nbitq), 
to_sfixed(349757528.0/4294967296.0,1,-nbitq), 
to_sfixed(-219711933.0/4294967296.0,1,-nbitq), 
to_sfixed(124403875.0/4294967296.0,1,-nbitq), 
to_sfixed(150147052.0/4294967296.0,1,-nbitq), 
to_sfixed(199169074.0/4294967296.0,1,-nbitq), 
to_sfixed(682275960.0/4294967296.0,1,-nbitq), 
to_sfixed(307384955.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(237163679.0/4294967296.0,1,-nbitq), 
to_sfixed(-11765452.0/4294967296.0,1,-nbitq), 
to_sfixed(9603025.0/4294967296.0,1,-nbitq), 
to_sfixed(120836290.0/4294967296.0,1,-nbitq), 
to_sfixed(208849698.0/4294967296.0,1,-nbitq), 
to_sfixed(-73982470.0/4294967296.0,1,-nbitq), 
to_sfixed(252985898.0/4294967296.0,1,-nbitq), 
to_sfixed(-324068054.0/4294967296.0,1,-nbitq), 
to_sfixed(-203839746.0/4294967296.0,1,-nbitq), 
to_sfixed(18975932.0/4294967296.0,1,-nbitq), 
to_sfixed(86250330.0/4294967296.0,1,-nbitq), 
to_sfixed(-64717166.0/4294967296.0,1,-nbitq), 
to_sfixed(-956155982.0/4294967296.0,1,-nbitq), 
to_sfixed(-31103104.0/4294967296.0,1,-nbitq), 
to_sfixed(-282408389.0/4294967296.0,1,-nbitq), 
to_sfixed(-105183225.0/4294967296.0,1,-nbitq), 
to_sfixed(-227466900.0/4294967296.0,1,-nbitq), 
to_sfixed(-290129407.0/4294967296.0,1,-nbitq), 
to_sfixed(-173228633.0/4294967296.0,1,-nbitq), 
to_sfixed(-156997046.0/4294967296.0,1,-nbitq), 
to_sfixed(-80777892.0/4294967296.0,1,-nbitq), 
to_sfixed(554152191.0/4294967296.0,1,-nbitq), 
to_sfixed(314840424.0/4294967296.0,1,-nbitq), 
to_sfixed(-99832777.0/4294967296.0,1,-nbitq), 
to_sfixed(-113993640.0/4294967296.0,1,-nbitq), 
to_sfixed(222482978.0/4294967296.0,1,-nbitq), 
to_sfixed(190699475.0/4294967296.0,1,-nbitq), 
to_sfixed(-358825370.0/4294967296.0,1,-nbitq), 
to_sfixed(-108509220.0/4294967296.0,1,-nbitq), 
to_sfixed(-705302090.0/4294967296.0,1,-nbitq), 
to_sfixed(-533783780.0/4294967296.0,1,-nbitq), 
to_sfixed(235933400.0/4294967296.0,1,-nbitq), 
to_sfixed(435127541.0/4294967296.0,1,-nbitq), 
to_sfixed(-45912209.0/4294967296.0,1,-nbitq), 
to_sfixed(562405924.0/4294967296.0,1,-nbitq), 
to_sfixed(74531102.0/4294967296.0,1,-nbitq), 
to_sfixed(17094445.0/4294967296.0,1,-nbitq), 
to_sfixed(646938527.0/4294967296.0,1,-nbitq), 
to_sfixed(-59513640.0/4294967296.0,1,-nbitq), 
to_sfixed(-92896056.0/4294967296.0,1,-nbitq), 
to_sfixed(-729462599.0/4294967296.0,1,-nbitq), 
to_sfixed(307914935.0/4294967296.0,1,-nbitq), 
to_sfixed(407983539.0/4294967296.0,1,-nbitq), 
to_sfixed(799384796.0/4294967296.0,1,-nbitq), 
to_sfixed(263771891.0/4294967296.0,1,-nbitq), 
to_sfixed(404706458.0/4294967296.0,1,-nbitq), 
to_sfixed(-225216298.0/4294967296.0,1,-nbitq), 
to_sfixed(-917442550.0/4294967296.0,1,-nbitq), 
to_sfixed(150156097.0/4294967296.0,1,-nbitq), 
to_sfixed(-272416475.0/4294967296.0,1,-nbitq), 
to_sfixed(-144208922.0/4294967296.0,1,-nbitq), 
to_sfixed(-636698907.0/4294967296.0,1,-nbitq), 
to_sfixed(-520531747.0/4294967296.0,1,-nbitq), 
to_sfixed(110361194.0/4294967296.0,1,-nbitq), 
to_sfixed(-189296507.0/4294967296.0,1,-nbitq), 
to_sfixed(-384311829.0/4294967296.0,1,-nbitq), 
to_sfixed(-886313685.0/4294967296.0,1,-nbitq), 
to_sfixed(390494159.0/4294967296.0,1,-nbitq), 
to_sfixed(-113764221.0/4294967296.0,1,-nbitq), 
to_sfixed(-30442818.0/4294967296.0,1,-nbitq), 
to_sfixed(-79090398.0/4294967296.0,1,-nbitq), 
to_sfixed(569048256.0/4294967296.0,1,-nbitq), 
to_sfixed(233267926.0/4294967296.0,1,-nbitq), 
to_sfixed(227178462.0/4294967296.0,1,-nbitq), 
to_sfixed(420990072.0/4294967296.0,1,-nbitq), 
to_sfixed(237564569.0/4294967296.0,1,-nbitq), 
to_sfixed(268278107.0/4294967296.0,1,-nbitq), 
to_sfixed(-244052590.0/4294967296.0,1,-nbitq), 
to_sfixed(-26503510.0/4294967296.0,1,-nbitq), 
to_sfixed(-314311966.0/4294967296.0,1,-nbitq), 
to_sfixed(868604039.0/4294967296.0,1,-nbitq), 
to_sfixed(364200060.0/4294967296.0,1,-nbitq), 
to_sfixed(-595399272.0/4294967296.0,1,-nbitq), 
to_sfixed(-208989514.0/4294967296.0,1,-nbitq), 
to_sfixed(210419720.0/4294967296.0,1,-nbitq), 
to_sfixed(-334373527.0/4294967296.0,1,-nbitq), 
to_sfixed(704176327.0/4294967296.0,1,-nbitq), 
to_sfixed(243354033.0/4294967296.0,1,-nbitq), 
to_sfixed(231095459.0/4294967296.0,1,-nbitq), 
to_sfixed(248850087.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-176311069.0/4294967296.0,1,-nbitq), 
to_sfixed(-259267686.0/4294967296.0,1,-nbitq), 
to_sfixed(362840582.0/4294967296.0,1,-nbitq), 
to_sfixed(-835555560.0/4294967296.0,1,-nbitq), 
to_sfixed(417810926.0/4294967296.0,1,-nbitq), 
to_sfixed(398456713.0/4294967296.0,1,-nbitq), 
to_sfixed(-207792186.0/4294967296.0,1,-nbitq), 
to_sfixed(-399363687.0/4294967296.0,1,-nbitq), 
to_sfixed(-148300581.0/4294967296.0,1,-nbitq), 
to_sfixed(235952948.0/4294967296.0,1,-nbitq), 
to_sfixed(-202716248.0/4294967296.0,1,-nbitq), 
to_sfixed(64622357.0/4294967296.0,1,-nbitq), 
to_sfixed(-370176092.0/4294967296.0,1,-nbitq), 
to_sfixed(275679172.0/4294967296.0,1,-nbitq), 
to_sfixed(-20479773.0/4294967296.0,1,-nbitq), 
to_sfixed(-581908117.0/4294967296.0,1,-nbitq), 
to_sfixed(47335603.0/4294967296.0,1,-nbitq), 
to_sfixed(124751476.0/4294967296.0,1,-nbitq), 
to_sfixed(-259742083.0/4294967296.0,1,-nbitq), 
to_sfixed(147528161.0/4294967296.0,1,-nbitq), 
to_sfixed(-325931558.0/4294967296.0,1,-nbitq), 
to_sfixed(198547123.0/4294967296.0,1,-nbitq), 
to_sfixed(408666793.0/4294967296.0,1,-nbitq), 
to_sfixed(299326362.0/4294967296.0,1,-nbitq), 
to_sfixed(-199775705.0/4294967296.0,1,-nbitq), 
to_sfixed(224710859.0/4294967296.0,1,-nbitq), 
to_sfixed(377842559.0/4294967296.0,1,-nbitq), 
to_sfixed(-73574601.0/4294967296.0,1,-nbitq), 
to_sfixed(486523334.0/4294967296.0,1,-nbitq), 
to_sfixed(-309099311.0/4294967296.0,1,-nbitq), 
to_sfixed(-961471031.0/4294967296.0,1,-nbitq), 
to_sfixed(-299568705.0/4294967296.0,1,-nbitq), 
to_sfixed(95006859.0/4294967296.0,1,-nbitq), 
to_sfixed(22194999.0/4294967296.0,1,-nbitq), 
to_sfixed(457790459.0/4294967296.0,1,-nbitq), 
to_sfixed(280861469.0/4294967296.0,1,-nbitq), 
to_sfixed(-162345583.0/4294967296.0,1,-nbitq), 
to_sfixed(119456487.0/4294967296.0,1,-nbitq), 
to_sfixed(69660666.0/4294967296.0,1,-nbitq), 
to_sfixed(15572370.0/4294967296.0,1,-nbitq), 
to_sfixed(-387384566.0/4294967296.0,1,-nbitq), 
to_sfixed(268739001.0/4294967296.0,1,-nbitq), 
to_sfixed(-47289184.0/4294967296.0,1,-nbitq), 
to_sfixed(393642741.0/4294967296.0,1,-nbitq), 
to_sfixed(264584191.0/4294967296.0,1,-nbitq), 
to_sfixed(-77223275.0/4294967296.0,1,-nbitq), 
to_sfixed(-177042331.0/4294967296.0,1,-nbitq), 
to_sfixed(-671501798.0/4294967296.0,1,-nbitq), 
to_sfixed(12622355.0/4294967296.0,1,-nbitq), 
to_sfixed(-285458024.0/4294967296.0,1,-nbitq), 
to_sfixed(-217539707.0/4294967296.0,1,-nbitq), 
to_sfixed(-763979323.0/4294967296.0,1,-nbitq), 
to_sfixed(280548724.0/4294967296.0,1,-nbitq), 
to_sfixed(-155713775.0/4294967296.0,1,-nbitq), 
to_sfixed(-306580022.0/4294967296.0,1,-nbitq), 
to_sfixed(67031589.0/4294967296.0,1,-nbitq), 
to_sfixed(27917130.0/4294967296.0,1,-nbitq), 
to_sfixed(-83465730.0/4294967296.0,1,-nbitq), 
to_sfixed(33556792.0/4294967296.0,1,-nbitq), 
to_sfixed(258816012.0/4294967296.0,1,-nbitq), 
to_sfixed(336864406.0/4294967296.0,1,-nbitq), 
to_sfixed(386760818.0/4294967296.0,1,-nbitq), 
to_sfixed(-179407956.0/4294967296.0,1,-nbitq), 
to_sfixed(-55170806.0/4294967296.0,1,-nbitq), 
to_sfixed(-299514382.0/4294967296.0,1,-nbitq), 
to_sfixed(115513780.0/4294967296.0,1,-nbitq), 
to_sfixed(-71314816.0/4294967296.0,1,-nbitq), 
to_sfixed(-191119763.0/4294967296.0,1,-nbitq), 
to_sfixed(199797734.0/4294967296.0,1,-nbitq), 
to_sfixed(326086253.0/4294967296.0,1,-nbitq), 
to_sfixed(600848786.0/4294967296.0,1,-nbitq), 
to_sfixed(9980196.0/4294967296.0,1,-nbitq), 
to_sfixed(-515458813.0/4294967296.0,1,-nbitq), 
to_sfixed(-270471113.0/4294967296.0,1,-nbitq), 
to_sfixed(595739016.0/4294967296.0,1,-nbitq), 
to_sfixed(-538569771.0/4294967296.0,1,-nbitq), 
to_sfixed(-84273835.0/4294967296.0,1,-nbitq), 
to_sfixed(-284933849.0/4294967296.0,1,-nbitq), 
to_sfixed(347761543.0/4294967296.0,1,-nbitq), 
to_sfixed(138177209.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-354342931.0/4294967296.0,1,-nbitq), 
to_sfixed(-202211454.0/4294967296.0,1,-nbitq), 
to_sfixed(-139087133.0/4294967296.0,1,-nbitq), 
to_sfixed(-100709119.0/4294967296.0,1,-nbitq), 
to_sfixed(-26200688.0/4294967296.0,1,-nbitq), 
to_sfixed(82358897.0/4294967296.0,1,-nbitq), 
to_sfixed(-234118527.0/4294967296.0,1,-nbitq), 
to_sfixed(-649269337.0/4294967296.0,1,-nbitq), 
to_sfixed(-352672464.0/4294967296.0,1,-nbitq), 
to_sfixed(-287406935.0/4294967296.0,1,-nbitq), 
to_sfixed(-227137235.0/4294967296.0,1,-nbitq), 
to_sfixed(-148817765.0/4294967296.0,1,-nbitq), 
to_sfixed(97491704.0/4294967296.0,1,-nbitq), 
to_sfixed(165967703.0/4294967296.0,1,-nbitq), 
to_sfixed(-217296393.0/4294967296.0,1,-nbitq), 
to_sfixed(81674456.0/4294967296.0,1,-nbitq), 
to_sfixed(-220235806.0/4294967296.0,1,-nbitq), 
to_sfixed(-105602868.0/4294967296.0,1,-nbitq), 
to_sfixed(515942415.0/4294967296.0,1,-nbitq), 
to_sfixed(153004547.0/4294967296.0,1,-nbitq), 
to_sfixed(-360310569.0/4294967296.0,1,-nbitq), 
to_sfixed(-97680809.0/4294967296.0,1,-nbitq), 
to_sfixed(43445532.0/4294967296.0,1,-nbitq), 
to_sfixed(-253188331.0/4294967296.0,1,-nbitq), 
to_sfixed(-36572973.0/4294967296.0,1,-nbitq), 
to_sfixed(-5499394.0/4294967296.0,1,-nbitq), 
to_sfixed(344058371.0/4294967296.0,1,-nbitq), 
to_sfixed(-353289585.0/4294967296.0,1,-nbitq), 
to_sfixed(503527928.0/4294967296.0,1,-nbitq), 
to_sfixed(154876433.0/4294967296.0,1,-nbitq), 
to_sfixed(-722230361.0/4294967296.0,1,-nbitq), 
to_sfixed(330633734.0/4294967296.0,1,-nbitq), 
to_sfixed(-71190692.0/4294967296.0,1,-nbitq), 
to_sfixed(237445506.0/4294967296.0,1,-nbitq), 
to_sfixed(431107992.0/4294967296.0,1,-nbitq), 
to_sfixed(487313220.0/4294967296.0,1,-nbitq), 
to_sfixed(100863610.0/4294967296.0,1,-nbitq), 
to_sfixed(62526779.0/4294967296.0,1,-nbitq), 
to_sfixed(3415152.0/4294967296.0,1,-nbitq), 
to_sfixed(436536052.0/4294967296.0,1,-nbitq), 
to_sfixed(343194883.0/4294967296.0,1,-nbitq), 
to_sfixed(184492185.0/4294967296.0,1,-nbitq), 
to_sfixed(373126465.0/4294967296.0,1,-nbitq), 
to_sfixed(198963968.0/4294967296.0,1,-nbitq), 
to_sfixed(-270930890.0/4294967296.0,1,-nbitq), 
to_sfixed(896455142.0/4294967296.0,1,-nbitq), 
to_sfixed(-415402362.0/4294967296.0,1,-nbitq), 
to_sfixed(-319213199.0/4294967296.0,1,-nbitq), 
to_sfixed(18299311.0/4294967296.0,1,-nbitq), 
to_sfixed(321122443.0/4294967296.0,1,-nbitq), 
to_sfixed(-230408791.0/4294967296.0,1,-nbitq), 
to_sfixed(-291482337.0/4294967296.0,1,-nbitq), 
to_sfixed(83742620.0/4294967296.0,1,-nbitq), 
to_sfixed(-151349821.0/4294967296.0,1,-nbitq), 
to_sfixed(-296145079.0/4294967296.0,1,-nbitq), 
to_sfixed(-411961093.0/4294967296.0,1,-nbitq), 
to_sfixed(-245767741.0/4294967296.0,1,-nbitq), 
to_sfixed(-392718673.0/4294967296.0,1,-nbitq), 
to_sfixed(-72626895.0/4294967296.0,1,-nbitq), 
to_sfixed(185912058.0/4294967296.0,1,-nbitq), 
to_sfixed(121572891.0/4294967296.0,1,-nbitq), 
to_sfixed(120635742.0/4294967296.0,1,-nbitq), 
to_sfixed(351868968.0/4294967296.0,1,-nbitq), 
to_sfixed(225704967.0/4294967296.0,1,-nbitq), 
to_sfixed(281846684.0/4294967296.0,1,-nbitq), 
to_sfixed(-303440155.0/4294967296.0,1,-nbitq), 
to_sfixed(237192835.0/4294967296.0,1,-nbitq), 
to_sfixed(-584869475.0/4294967296.0,1,-nbitq), 
to_sfixed(310574401.0/4294967296.0,1,-nbitq), 
to_sfixed(-33876427.0/4294967296.0,1,-nbitq), 
to_sfixed(-148761407.0/4294967296.0,1,-nbitq), 
to_sfixed(459083093.0/4294967296.0,1,-nbitq), 
to_sfixed(-11427439.0/4294967296.0,1,-nbitq), 
to_sfixed(-76483735.0/4294967296.0,1,-nbitq), 
to_sfixed(9589377.0/4294967296.0,1,-nbitq), 
to_sfixed(-113276135.0/4294967296.0,1,-nbitq), 
to_sfixed(37243742.0/4294967296.0,1,-nbitq), 
to_sfixed(353830675.0/4294967296.0,1,-nbitq), 
to_sfixed(143197983.0/4294967296.0,1,-nbitq), 
to_sfixed(123779270.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-349397422.0/4294967296.0,1,-nbitq), 
to_sfixed(-607114421.0/4294967296.0,1,-nbitq), 
to_sfixed(-188488539.0/4294967296.0,1,-nbitq), 
to_sfixed(-520122125.0/4294967296.0,1,-nbitq), 
to_sfixed(-248745153.0/4294967296.0,1,-nbitq), 
to_sfixed(-130548869.0/4294967296.0,1,-nbitq), 
to_sfixed(296161776.0/4294967296.0,1,-nbitq), 
to_sfixed(-128212990.0/4294967296.0,1,-nbitq), 
to_sfixed(-450218994.0/4294967296.0,1,-nbitq), 
to_sfixed(160374680.0/4294967296.0,1,-nbitq), 
to_sfixed(-234323134.0/4294967296.0,1,-nbitq), 
to_sfixed(415458542.0/4294967296.0,1,-nbitq), 
to_sfixed(-103482141.0/4294967296.0,1,-nbitq), 
to_sfixed(-382712258.0/4294967296.0,1,-nbitq), 
to_sfixed(268009867.0/4294967296.0,1,-nbitq), 
to_sfixed(30121501.0/4294967296.0,1,-nbitq), 
to_sfixed(-313034128.0/4294967296.0,1,-nbitq), 
to_sfixed(82403275.0/4294967296.0,1,-nbitq), 
to_sfixed(21601717.0/4294967296.0,1,-nbitq), 
to_sfixed(255152396.0/4294967296.0,1,-nbitq), 
to_sfixed(57820670.0/4294967296.0,1,-nbitq), 
to_sfixed(512479672.0/4294967296.0,1,-nbitq), 
to_sfixed(-67788073.0/4294967296.0,1,-nbitq), 
to_sfixed(258724096.0/4294967296.0,1,-nbitq), 
to_sfixed(424424122.0/4294967296.0,1,-nbitq), 
to_sfixed(-347249359.0/4294967296.0,1,-nbitq), 
to_sfixed(280801277.0/4294967296.0,1,-nbitq), 
to_sfixed(-361483081.0/4294967296.0,1,-nbitq), 
to_sfixed(-248744068.0/4294967296.0,1,-nbitq), 
to_sfixed(240974839.0/4294967296.0,1,-nbitq), 
to_sfixed(-143990196.0/4294967296.0,1,-nbitq), 
to_sfixed(-511171989.0/4294967296.0,1,-nbitq), 
to_sfixed(374582441.0/4294967296.0,1,-nbitq), 
to_sfixed(508640511.0/4294967296.0,1,-nbitq), 
to_sfixed(349713761.0/4294967296.0,1,-nbitq), 
to_sfixed(313940614.0/4294967296.0,1,-nbitq), 
to_sfixed(-152425423.0/4294967296.0,1,-nbitq), 
to_sfixed(-41374021.0/4294967296.0,1,-nbitq), 
to_sfixed(224394152.0/4294967296.0,1,-nbitq), 
to_sfixed(-14154932.0/4294967296.0,1,-nbitq), 
to_sfixed(291475414.0/4294967296.0,1,-nbitq), 
to_sfixed(-50163556.0/4294967296.0,1,-nbitq), 
to_sfixed(162441810.0/4294967296.0,1,-nbitq), 
to_sfixed(15960012.0/4294967296.0,1,-nbitq), 
to_sfixed(262754021.0/4294967296.0,1,-nbitq), 
to_sfixed(545316963.0/4294967296.0,1,-nbitq), 
to_sfixed(-448011587.0/4294967296.0,1,-nbitq), 
to_sfixed(-377994646.0/4294967296.0,1,-nbitq), 
to_sfixed(282832003.0/4294967296.0,1,-nbitq), 
to_sfixed(434091345.0/4294967296.0,1,-nbitq), 
to_sfixed(292930378.0/4294967296.0,1,-nbitq), 
to_sfixed(-182282840.0/4294967296.0,1,-nbitq), 
to_sfixed(-423311933.0/4294967296.0,1,-nbitq), 
to_sfixed(-288733349.0/4294967296.0,1,-nbitq), 
to_sfixed(-348839717.0/4294967296.0,1,-nbitq), 
to_sfixed(-7236935.0/4294967296.0,1,-nbitq), 
to_sfixed(303823078.0/4294967296.0,1,-nbitq), 
to_sfixed(-74203195.0/4294967296.0,1,-nbitq), 
to_sfixed(-332904664.0/4294967296.0,1,-nbitq), 
to_sfixed(409957955.0/4294967296.0,1,-nbitq), 
to_sfixed(45991634.0/4294967296.0,1,-nbitq), 
to_sfixed(387414769.0/4294967296.0,1,-nbitq), 
to_sfixed(36056961.0/4294967296.0,1,-nbitq), 
to_sfixed(261525534.0/4294967296.0,1,-nbitq), 
to_sfixed(-254398152.0/4294967296.0,1,-nbitq), 
to_sfixed(6496635.0/4294967296.0,1,-nbitq), 
to_sfixed(389929490.0/4294967296.0,1,-nbitq), 
to_sfixed(-515409115.0/4294967296.0,1,-nbitq), 
to_sfixed(-153370572.0/4294967296.0,1,-nbitq), 
to_sfixed(-219258557.0/4294967296.0,1,-nbitq), 
to_sfixed(-144383297.0/4294967296.0,1,-nbitq), 
to_sfixed(-270263356.0/4294967296.0,1,-nbitq), 
to_sfixed(-420251462.0/4294967296.0,1,-nbitq), 
to_sfixed(-77602457.0/4294967296.0,1,-nbitq), 
to_sfixed(470662159.0/4294967296.0,1,-nbitq), 
to_sfixed(-429818225.0/4294967296.0,1,-nbitq), 
to_sfixed(151485555.0/4294967296.0,1,-nbitq), 
to_sfixed(-77774403.0/4294967296.0,1,-nbitq), 
to_sfixed(-247829322.0/4294967296.0,1,-nbitq), 
to_sfixed(-294729293.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(39774448.0/4294967296.0,1,-nbitq), 
to_sfixed(-359075995.0/4294967296.0,1,-nbitq), 
to_sfixed(458858702.0/4294967296.0,1,-nbitq), 
to_sfixed(142891745.0/4294967296.0,1,-nbitq), 
to_sfixed(297147568.0/4294967296.0,1,-nbitq), 
to_sfixed(140984587.0/4294967296.0,1,-nbitq), 
to_sfixed(312580013.0/4294967296.0,1,-nbitq), 
to_sfixed(-211022154.0/4294967296.0,1,-nbitq), 
to_sfixed(-115149933.0/4294967296.0,1,-nbitq), 
to_sfixed(-176466938.0/4294967296.0,1,-nbitq), 
to_sfixed(287388878.0/4294967296.0,1,-nbitq), 
to_sfixed(70459554.0/4294967296.0,1,-nbitq), 
to_sfixed(1345973.0/4294967296.0,1,-nbitq), 
to_sfixed(39480639.0/4294967296.0,1,-nbitq), 
to_sfixed(284994492.0/4294967296.0,1,-nbitq), 
to_sfixed(187751176.0/4294967296.0,1,-nbitq), 
to_sfixed(276014684.0/4294967296.0,1,-nbitq), 
to_sfixed(-315757671.0/4294967296.0,1,-nbitq), 
to_sfixed(261543568.0/4294967296.0,1,-nbitq), 
to_sfixed(271709628.0/4294967296.0,1,-nbitq), 
to_sfixed(210233513.0/4294967296.0,1,-nbitq), 
to_sfixed(475323666.0/4294967296.0,1,-nbitq), 
to_sfixed(-102924638.0/4294967296.0,1,-nbitq), 
to_sfixed(-222529739.0/4294967296.0,1,-nbitq), 
to_sfixed(199781610.0/4294967296.0,1,-nbitq), 
to_sfixed(409737149.0/4294967296.0,1,-nbitq), 
to_sfixed(-15097119.0/4294967296.0,1,-nbitq), 
to_sfixed(-596481343.0/4294967296.0,1,-nbitq), 
to_sfixed(-292202050.0/4294967296.0,1,-nbitq), 
to_sfixed(51665430.0/4294967296.0,1,-nbitq), 
to_sfixed(-208987920.0/4294967296.0,1,-nbitq), 
to_sfixed(-288228503.0/4294967296.0,1,-nbitq), 
to_sfixed(-290740840.0/4294967296.0,1,-nbitq), 
to_sfixed(155667418.0/4294967296.0,1,-nbitq), 
to_sfixed(387287255.0/4294967296.0,1,-nbitq), 
to_sfixed(289319072.0/4294967296.0,1,-nbitq), 
to_sfixed(210121637.0/4294967296.0,1,-nbitq), 
to_sfixed(-184320307.0/4294967296.0,1,-nbitq), 
to_sfixed(-63127362.0/4294967296.0,1,-nbitq), 
to_sfixed(468500162.0/4294967296.0,1,-nbitq), 
to_sfixed(-194587030.0/4294967296.0,1,-nbitq), 
to_sfixed(300775428.0/4294967296.0,1,-nbitq), 
to_sfixed(-141163375.0/4294967296.0,1,-nbitq), 
to_sfixed(80652115.0/4294967296.0,1,-nbitq), 
to_sfixed(175669808.0/4294967296.0,1,-nbitq), 
to_sfixed(-47985975.0/4294967296.0,1,-nbitq), 
to_sfixed(-150812224.0/4294967296.0,1,-nbitq), 
to_sfixed(-145053827.0/4294967296.0,1,-nbitq), 
to_sfixed(-34929623.0/4294967296.0,1,-nbitq), 
to_sfixed(407051642.0/4294967296.0,1,-nbitq), 
to_sfixed(-306583564.0/4294967296.0,1,-nbitq), 
to_sfixed(265030285.0/4294967296.0,1,-nbitq), 
to_sfixed(-12564193.0/4294967296.0,1,-nbitq), 
to_sfixed(-414769964.0/4294967296.0,1,-nbitq), 
to_sfixed(102371410.0/4294967296.0,1,-nbitq), 
to_sfixed(230262124.0/4294967296.0,1,-nbitq), 
to_sfixed(-111749499.0/4294967296.0,1,-nbitq), 
to_sfixed(-233199010.0/4294967296.0,1,-nbitq), 
to_sfixed(16349794.0/4294967296.0,1,-nbitq), 
to_sfixed(-15964495.0/4294967296.0,1,-nbitq), 
to_sfixed(-128854182.0/4294967296.0,1,-nbitq), 
to_sfixed(164686672.0/4294967296.0,1,-nbitq), 
to_sfixed(95265526.0/4294967296.0,1,-nbitq), 
to_sfixed(421821911.0/4294967296.0,1,-nbitq), 
to_sfixed(266788019.0/4294967296.0,1,-nbitq), 
to_sfixed(-116331761.0/4294967296.0,1,-nbitq), 
to_sfixed(377592238.0/4294967296.0,1,-nbitq), 
to_sfixed(177191372.0/4294967296.0,1,-nbitq), 
to_sfixed(38046897.0/4294967296.0,1,-nbitq), 
to_sfixed(114025506.0/4294967296.0,1,-nbitq), 
to_sfixed(-284542619.0/4294967296.0,1,-nbitq), 
to_sfixed(-299168011.0/4294967296.0,1,-nbitq), 
to_sfixed(192736384.0/4294967296.0,1,-nbitq), 
to_sfixed(167971650.0/4294967296.0,1,-nbitq), 
to_sfixed(283056690.0/4294967296.0,1,-nbitq), 
to_sfixed(-605433257.0/4294967296.0,1,-nbitq), 
to_sfixed(-57732300.0/4294967296.0,1,-nbitq), 
to_sfixed(-88809426.0/4294967296.0,1,-nbitq), 
to_sfixed(48621674.0/4294967296.0,1,-nbitq), 
to_sfixed(273250361.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-299062798.0/4294967296.0,1,-nbitq), 
to_sfixed(-125896222.0/4294967296.0,1,-nbitq), 
to_sfixed(261185484.0/4294967296.0,1,-nbitq), 
to_sfixed(-57620646.0/4294967296.0,1,-nbitq), 
to_sfixed(-268656941.0/4294967296.0,1,-nbitq), 
to_sfixed(-80214189.0/4294967296.0,1,-nbitq), 
to_sfixed(-395038725.0/4294967296.0,1,-nbitq), 
to_sfixed(18913818.0/4294967296.0,1,-nbitq), 
to_sfixed(75232473.0/4294967296.0,1,-nbitq), 
to_sfixed(373559449.0/4294967296.0,1,-nbitq), 
to_sfixed(-210053886.0/4294967296.0,1,-nbitq), 
to_sfixed(322101218.0/4294967296.0,1,-nbitq), 
to_sfixed(-170539609.0/4294967296.0,1,-nbitq), 
to_sfixed(358114088.0/4294967296.0,1,-nbitq), 
to_sfixed(-156246273.0/4294967296.0,1,-nbitq), 
to_sfixed(-209990860.0/4294967296.0,1,-nbitq), 
to_sfixed(-117569023.0/4294967296.0,1,-nbitq), 
to_sfixed(379281041.0/4294967296.0,1,-nbitq), 
to_sfixed(-74957525.0/4294967296.0,1,-nbitq), 
to_sfixed(45591836.0/4294967296.0,1,-nbitq), 
to_sfixed(-367789567.0/4294967296.0,1,-nbitq), 
to_sfixed(241480494.0/4294967296.0,1,-nbitq), 
to_sfixed(-44455584.0/4294967296.0,1,-nbitq), 
to_sfixed(41615674.0/4294967296.0,1,-nbitq), 
to_sfixed(363066819.0/4294967296.0,1,-nbitq), 
to_sfixed(106289940.0/4294967296.0,1,-nbitq), 
to_sfixed(-191239218.0/4294967296.0,1,-nbitq), 
to_sfixed(-227768315.0/4294967296.0,1,-nbitq), 
to_sfixed(91208260.0/4294967296.0,1,-nbitq), 
to_sfixed(-216685815.0/4294967296.0,1,-nbitq), 
to_sfixed(-498446025.0/4294967296.0,1,-nbitq), 
to_sfixed(-59839701.0/4294967296.0,1,-nbitq), 
to_sfixed(160348313.0/4294967296.0,1,-nbitq), 
to_sfixed(-29649817.0/4294967296.0,1,-nbitq), 
to_sfixed(-94536690.0/4294967296.0,1,-nbitq), 
to_sfixed(-330535426.0/4294967296.0,1,-nbitq), 
to_sfixed(89198358.0/4294967296.0,1,-nbitq), 
to_sfixed(32386731.0/4294967296.0,1,-nbitq), 
to_sfixed(114890714.0/4294967296.0,1,-nbitq), 
to_sfixed(-293598353.0/4294967296.0,1,-nbitq), 
to_sfixed(-344144978.0/4294967296.0,1,-nbitq), 
to_sfixed(187734774.0/4294967296.0,1,-nbitq), 
to_sfixed(-316695721.0/4294967296.0,1,-nbitq), 
to_sfixed(512155479.0/4294967296.0,1,-nbitq), 
to_sfixed(361995082.0/4294967296.0,1,-nbitq), 
to_sfixed(638377641.0/4294967296.0,1,-nbitq), 
to_sfixed(303816794.0/4294967296.0,1,-nbitq), 
to_sfixed(-22553811.0/4294967296.0,1,-nbitq), 
to_sfixed(160966534.0/4294967296.0,1,-nbitq), 
to_sfixed(535726403.0/4294967296.0,1,-nbitq), 
to_sfixed(336016122.0/4294967296.0,1,-nbitq), 
to_sfixed(192077988.0/4294967296.0,1,-nbitq), 
to_sfixed(45194296.0/4294967296.0,1,-nbitq), 
to_sfixed(-329274052.0/4294967296.0,1,-nbitq), 
to_sfixed(118127748.0/4294967296.0,1,-nbitq), 
to_sfixed(-378749177.0/4294967296.0,1,-nbitq), 
to_sfixed(-63539406.0/4294967296.0,1,-nbitq), 
to_sfixed(-104074301.0/4294967296.0,1,-nbitq), 
to_sfixed(118131376.0/4294967296.0,1,-nbitq), 
to_sfixed(310589172.0/4294967296.0,1,-nbitq), 
to_sfixed(122598909.0/4294967296.0,1,-nbitq), 
to_sfixed(-171163062.0/4294967296.0,1,-nbitq), 
to_sfixed(-492776363.0/4294967296.0,1,-nbitq), 
to_sfixed(-101584713.0/4294967296.0,1,-nbitq), 
to_sfixed(-312188121.0/4294967296.0,1,-nbitq), 
to_sfixed(54761432.0/4294967296.0,1,-nbitq), 
to_sfixed(303939959.0/4294967296.0,1,-nbitq), 
to_sfixed(-335729304.0/4294967296.0,1,-nbitq), 
to_sfixed(245415824.0/4294967296.0,1,-nbitq), 
to_sfixed(192164314.0/4294967296.0,1,-nbitq), 
to_sfixed(-447141377.0/4294967296.0,1,-nbitq), 
to_sfixed(985363.0/4294967296.0,1,-nbitq), 
to_sfixed(-166968908.0/4294967296.0,1,-nbitq), 
to_sfixed(8754031.0/4294967296.0,1,-nbitq), 
to_sfixed(132905634.0/4294967296.0,1,-nbitq), 
to_sfixed(-238187933.0/4294967296.0,1,-nbitq), 
to_sfixed(-260912278.0/4294967296.0,1,-nbitq), 
to_sfixed(-290947606.0/4294967296.0,1,-nbitq), 
to_sfixed(165821317.0/4294967296.0,1,-nbitq), 
to_sfixed(-179522359.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-107625576.0/4294967296.0,1,-nbitq), 
to_sfixed(-308485045.0/4294967296.0,1,-nbitq), 
to_sfixed(200127037.0/4294967296.0,1,-nbitq), 
to_sfixed(-462646868.0/4294967296.0,1,-nbitq), 
to_sfixed(45918141.0/4294967296.0,1,-nbitq), 
to_sfixed(293348158.0/4294967296.0,1,-nbitq), 
to_sfixed(-276134431.0/4294967296.0,1,-nbitq), 
to_sfixed(-110304011.0/4294967296.0,1,-nbitq), 
to_sfixed(120941698.0/4294967296.0,1,-nbitq), 
to_sfixed(-149332078.0/4294967296.0,1,-nbitq), 
to_sfixed(161027140.0/4294967296.0,1,-nbitq), 
to_sfixed(-46841642.0/4294967296.0,1,-nbitq), 
to_sfixed(-226436090.0/4294967296.0,1,-nbitq), 
to_sfixed(462038916.0/4294967296.0,1,-nbitq), 
to_sfixed(-101438862.0/4294967296.0,1,-nbitq), 
to_sfixed(-15090556.0/4294967296.0,1,-nbitq), 
to_sfixed(193599466.0/4294967296.0,1,-nbitq), 
to_sfixed(-252387012.0/4294967296.0,1,-nbitq), 
to_sfixed(-153845927.0/4294967296.0,1,-nbitq), 
to_sfixed(-300797616.0/4294967296.0,1,-nbitq), 
to_sfixed(225057695.0/4294967296.0,1,-nbitq), 
to_sfixed(248008972.0/4294967296.0,1,-nbitq), 
to_sfixed(524568762.0/4294967296.0,1,-nbitq), 
to_sfixed(-278741485.0/4294967296.0,1,-nbitq), 
to_sfixed(-161296280.0/4294967296.0,1,-nbitq), 
to_sfixed(-199529401.0/4294967296.0,1,-nbitq), 
to_sfixed(-119320214.0/4294967296.0,1,-nbitq), 
to_sfixed(-464381186.0/4294967296.0,1,-nbitq), 
to_sfixed(117885861.0/4294967296.0,1,-nbitq), 
to_sfixed(386748844.0/4294967296.0,1,-nbitq), 
to_sfixed(144806035.0/4294967296.0,1,-nbitq), 
to_sfixed(-152684158.0/4294967296.0,1,-nbitq), 
to_sfixed(475853050.0/4294967296.0,1,-nbitq), 
to_sfixed(-236451799.0/4294967296.0,1,-nbitq), 
to_sfixed(48739489.0/4294967296.0,1,-nbitq), 
to_sfixed(34409313.0/4294967296.0,1,-nbitq), 
to_sfixed(304519792.0/4294967296.0,1,-nbitq), 
to_sfixed(-269756328.0/4294967296.0,1,-nbitq), 
to_sfixed(166576565.0/4294967296.0,1,-nbitq), 
to_sfixed(206191974.0/4294967296.0,1,-nbitq), 
to_sfixed(20559541.0/4294967296.0,1,-nbitq), 
to_sfixed(14515936.0/4294967296.0,1,-nbitq), 
to_sfixed(364481888.0/4294967296.0,1,-nbitq), 
to_sfixed(226830841.0/4294967296.0,1,-nbitq), 
to_sfixed(42851853.0/4294967296.0,1,-nbitq), 
to_sfixed(517970378.0/4294967296.0,1,-nbitq), 
to_sfixed(-238654506.0/4294967296.0,1,-nbitq), 
to_sfixed(-232144478.0/4294967296.0,1,-nbitq), 
to_sfixed(104198677.0/4294967296.0,1,-nbitq), 
to_sfixed(-89805664.0/4294967296.0,1,-nbitq), 
to_sfixed(431372987.0/4294967296.0,1,-nbitq), 
to_sfixed(-87526111.0/4294967296.0,1,-nbitq), 
to_sfixed(-164737577.0/4294967296.0,1,-nbitq), 
to_sfixed(171833589.0/4294967296.0,1,-nbitq), 
to_sfixed(-90603780.0/4294967296.0,1,-nbitq), 
to_sfixed(-215891947.0/4294967296.0,1,-nbitq), 
to_sfixed(-262330298.0/4294967296.0,1,-nbitq), 
to_sfixed(-453550533.0/4294967296.0,1,-nbitq), 
to_sfixed(257211576.0/4294967296.0,1,-nbitq), 
to_sfixed(194830734.0/4294967296.0,1,-nbitq), 
to_sfixed(196248290.0/4294967296.0,1,-nbitq), 
to_sfixed(60296478.0/4294967296.0,1,-nbitq), 
to_sfixed(-226904713.0/4294967296.0,1,-nbitq), 
to_sfixed(353690184.0/4294967296.0,1,-nbitq), 
to_sfixed(118395189.0/4294967296.0,1,-nbitq), 
to_sfixed(-395643583.0/4294967296.0,1,-nbitq), 
to_sfixed(391280752.0/4294967296.0,1,-nbitq), 
to_sfixed(-36457534.0/4294967296.0,1,-nbitq), 
to_sfixed(415881732.0/4294967296.0,1,-nbitq), 
to_sfixed(115474979.0/4294967296.0,1,-nbitq), 
to_sfixed(-377106280.0/4294967296.0,1,-nbitq), 
to_sfixed(368598906.0/4294967296.0,1,-nbitq), 
to_sfixed(-421453962.0/4294967296.0,1,-nbitq), 
to_sfixed(286732566.0/4294967296.0,1,-nbitq), 
to_sfixed(316789704.0/4294967296.0,1,-nbitq), 
to_sfixed(64389344.0/4294967296.0,1,-nbitq), 
to_sfixed(320281026.0/4294967296.0,1,-nbitq), 
to_sfixed(245416333.0/4294967296.0,1,-nbitq), 
to_sfixed(129973424.0/4294967296.0,1,-nbitq), 
to_sfixed(-140573903.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(248649110.0/4294967296.0,1,-nbitq), 
to_sfixed(-184585405.0/4294967296.0,1,-nbitq), 
to_sfixed(346835406.0/4294967296.0,1,-nbitq), 
to_sfixed(-158618673.0/4294967296.0,1,-nbitq), 
to_sfixed(-104195732.0/4294967296.0,1,-nbitq), 
to_sfixed(125312408.0/4294967296.0,1,-nbitq), 
to_sfixed(393560588.0/4294967296.0,1,-nbitq), 
to_sfixed(-359465010.0/4294967296.0,1,-nbitq), 
to_sfixed(177678334.0/4294967296.0,1,-nbitq), 
to_sfixed(-69981555.0/4294967296.0,1,-nbitq), 
to_sfixed(272171982.0/4294967296.0,1,-nbitq), 
to_sfixed(514064567.0/4294967296.0,1,-nbitq), 
to_sfixed(309006818.0/4294967296.0,1,-nbitq), 
to_sfixed(-332905843.0/4294967296.0,1,-nbitq), 
to_sfixed(-308942009.0/4294967296.0,1,-nbitq), 
to_sfixed(-281867984.0/4294967296.0,1,-nbitq), 
to_sfixed(-358276079.0/4294967296.0,1,-nbitq), 
to_sfixed(-339695640.0/4294967296.0,1,-nbitq), 
to_sfixed(439418344.0/4294967296.0,1,-nbitq), 
to_sfixed(122077590.0/4294967296.0,1,-nbitq), 
to_sfixed(63847428.0/4294967296.0,1,-nbitq), 
to_sfixed(389149511.0/4294967296.0,1,-nbitq), 
to_sfixed(499328328.0/4294967296.0,1,-nbitq), 
to_sfixed(-62881066.0/4294967296.0,1,-nbitq), 
to_sfixed(-93905295.0/4294967296.0,1,-nbitq), 
to_sfixed(389244661.0/4294967296.0,1,-nbitq), 
to_sfixed(389533290.0/4294967296.0,1,-nbitq), 
to_sfixed(-639881165.0/4294967296.0,1,-nbitq), 
to_sfixed(446551726.0/4294967296.0,1,-nbitq), 
to_sfixed(441921459.0/4294967296.0,1,-nbitq), 
to_sfixed(3896817.0/4294967296.0,1,-nbitq), 
to_sfixed(-24045498.0/4294967296.0,1,-nbitq), 
to_sfixed(292897745.0/4294967296.0,1,-nbitq), 
to_sfixed(217620121.0/4294967296.0,1,-nbitq), 
to_sfixed(495108759.0/4294967296.0,1,-nbitq), 
to_sfixed(5682734.0/4294967296.0,1,-nbitq), 
to_sfixed(154429546.0/4294967296.0,1,-nbitq), 
to_sfixed(263839579.0/4294967296.0,1,-nbitq), 
to_sfixed(-159230911.0/4294967296.0,1,-nbitq), 
to_sfixed(494140541.0/4294967296.0,1,-nbitq), 
to_sfixed(287000072.0/4294967296.0,1,-nbitq), 
to_sfixed(306382367.0/4294967296.0,1,-nbitq), 
to_sfixed(99431495.0/4294967296.0,1,-nbitq), 
to_sfixed(65332789.0/4294967296.0,1,-nbitq), 
to_sfixed(228725434.0/4294967296.0,1,-nbitq), 
to_sfixed(-62216090.0/4294967296.0,1,-nbitq), 
to_sfixed(-271966017.0/4294967296.0,1,-nbitq), 
to_sfixed(-271689196.0/4294967296.0,1,-nbitq), 
to_sfixed(-302953556.0/4294967296.0,1,-nbitq), 
to_sfixed(-163401397.0/4294967296.0,1,-nbitq), 
to_sfixed(-184593647.0/4294967296.0,1,-nbitq), 
to_sfixed(-36521008.0/4294967296.0,1,-nbitq), 
to_sfixed(-75914963.0/4294967296.0,1,-nbitq), 
to_sfixed(-123526980.0/4294967296.0,1,-nbitq), 
to_sfixed(-71622067.0/4294967296.0,1,-nbitq), 
to_sfixed(-422211487.0/4294967296.0,1,-nbitq), 
to_sfixed(200861758.0/4294967296.0,1,-nbitq), 
to_sfixed(-456806597.0/4294967296.0,1,-nbitq), 
to_sfixed(158941747.0/4294967296.0,1,-nbitq), 
to_sfixed(-78404806.0/4294967296.0,1,-nbitq), 
to_sfixed(21871599.0/4294967296.0,1,-nbitq), 
to_sfixed(393412818.0/4294967296.0,1,-nbitq), 
to_sfixed(139461138.0/4294967296.0,1,-nbitq), 
to_sfixed(-61562248.0/4294967296.0,1,-nbitq), 
to_sfixed(-267749582.0/4294967296.0,1,-nbitq), 
to_sfixed(-344451027.0/4294967296.0,1,-nbitq), 
to_sfixed(301630497.0/4294967296.0,1,-nbitq), 
to_sfixed(-370684996.0/4294967296.0,1,-nbitq), 
to_sfixed(72564980.0/4294967296.0,1,-nbitq), 
to_sfixed(166598051.0/4294967296.0,1,-nbitq), 
to_sfixed(-77665661.0/4294967296.0,1,-nbitq), 
to_sfixed(320044708.0/4294967296.0,1,-nbitq), 
to_sfixed(-117594854.0/4294967296.0,1,-nbitq), 
to_sfixed(173895702.0/4294967296.0,1,-nbitq), 
to_sfixed(-113865519.0/4294967296.0,1,-nbitq), 
to_sfixed(-340790914.0/4294967296.0,1,-nbitq), 
to_sfixed(-42508032.0/4294967296.0,1,-nbitq), 
to_sfixed(231336206.0/4294967296.0,1,-nbitq), 
to_sfixed(-430893912.0/4294967296.0,1,-nbitq), 
to_sfixed(242284752.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-336213688.0/4294967296.0,1,-nbitq), 
to_sfixed(-241843880.0/4294967296.0,1,-nbitq), 
to_sfixed(75113316.0/4294967296.0,1,-nbitq), 
to_sfixed(-311267543.0/4294967296.0,1,-nbitq), 
to_sfixed(-230800223.0/4294967296.0,1,-nbitq), 
to_sfixed(-196294183.0/4294967296.0,1,-nbitq), 
to_sfixed(206644934.0/4294967296.0,1,-nbitq), 
to_sfixed(-446227695.0/4294967296.0,1,-nbitq), 
to_sfixed(-241628010.0/4294967296.0,1,-nbitq), 
to_sfixed(48779221.0/4294967296.0,1,-nbitq), 
to_sfixed(190905345.0/4294967296.0,1,-nbitq), 
to_sfixed(-146162598.0/4294967296.0,1,-nbitq), 
to_sfixed(-123589048.0/4294967296.0,1,-nbitq), 
to_sfixed(-245113604.0/4294967296.0,1,-nbitq), 
to_sfixed(-128635444.0/4294967296.0,1,-nbitq), 
to_sfixed(-277227438.0/4294967296.0,1,-nbitq), 
to_sfixed(-357770606.0/4294967296.0,1,-nbitq), 
to_sfixed(386363204.0/4294967296.0,1,-nbitq), 
to_sfixed(301787612.0/4294967296.0,1,-nbitq), 
to_sfixed(75183685.0/4294967296.0,1,-nbitq), 
to_sfixed(-40489329.0/4294967296.0,1,-nbitq), 
to_sfixed(-184471748.0/4294967296.0,1,-nbitq), 
to_sfixed(316503444.0/4294967296.0,1,-nbitq), 
to_sfixed(-101546464.0/4294967296.0,1,-nbitq), 
to_sfixed(249331685.0/4294967296.0,1,-nbitq), 
to_sfixed(265751740.0/4294967296.0,1,-nbitq), 
to_sfixed(-202169535.0/4294967296.0,1,-nbitq), 
to_sfixed(137207494.0/4294967296.0,1,-nbitq), 
to_sfixed(71786326.0/4294967296.0,1,-nbitq), 
to_sfixed(-20472393.0/4294967296.0,1,-nbitq), 
to_sfixed(-407698882.0/4294967296.0,1,-nbitq), 
to_sfixed(-240342154.0/4294967296.0,1,-nbitq), 
to_sfixed(173551518.0/4294967296.0,1,-nbitq), 
to_sfixed(-153749470.0/4294967296.0,1,-nbitq), 
to_sfixed(238866459.0/4294967296.0,1,-nbitq), 
to_sfixed(356551713.0/4294967296.0,1,-nbitq), 
to_sfixed(387003644.0/4294967296.0,1,-nbitq), 
to_sfixed(263806458.0/4294967296.0,1,-nbitq), 
to_sfixed(303894904.0/4294967296.0,1,-nbitq), 
to_sfixed(-118492391.0/4294967296.0,1,-nbitq), 
to_sfixed(-49947141.0/4294967296.0,1,-nbitq), 
to_sfixed(-66863101.0/4294967296.0,1,-nbitq), 
to_sfixed(314846776.0/4294967296.0,1,-nbitq), 
to_sfixed(-166418834.0/4294967296.0,1,-nbitq), 
to_sfixed(1243866.0/4294967296.0,1,-nbitq), 
to_sfixed(-1928375.0/4294967296.0,1,-nbitq), 
to_sfixed(-26638163.0/4294967296.0,1,-nbitq), 
to_sfixed(-390914386.0/4294967296.0,1,-nbitq), 
to_sfixed(315008927.0/4294967296.0,1,-nbitq), 
to_sfixed(-66502384.0/4294967296.0,1,-nbitq), 
to_sfixed(392189480.0/4294967296.0,1,-nbitq), 
to_sfixed(302397174.0/4294967296.0,1,-nbitq), 
to_sfixed(-89571927.0/4294967296.0,1,-nbitq), 
to_sfixed(-127538496.0/4294967296.0,1,-nbitq), 
to_sfixed(462729650.0/4294967296.0,1,-nbitq), 
to_sfixed(251251313.0/4294967296.0,1,-nbitq), 
to_sfixed(405605347.0/4294967296.0,1,-nbitq), 
to_sfixed(8896220.0/4294967296.0,1,-nbitq), 
to_sfixed(167785079.0/4294967296.0,1,-nbitq), 
to_sfixed(161036462.0/4294967296.0,1,-nbitq), 
to_sfixed(67808832.0/4294967296.0,1,-nbitq), 
to_sfixed(-127082857.0/4294967296.0,1,-nbitq), 
to_sfixed(-285344450.0/4294967296.0,1,-nbitq), 
to_sfixed(253115683.0/4294967296.0,1,-nbitq), 
to_sfixed(-8666063.0/4294967296.0,1,-nbitq), 
to_sfixed(-168698576.0/4294967296.0,1,-nbitq), 
to_sfixed(695395832.0/4294967296.0,1,-nbitq), 
to_sfixed(161689112.0/4294967296.0,1,-nbitq), 
to_sfixed(-239265595.0/4294967296.0,1,-nbitq), 
to_sfixed(-200175364.0/4294967296.0,1,-nbitq), 
to_sfixed(-291251130.0/4294967296.0,1,-nbitq), 
to_sfixed(268226623.0/4294967296.0,1,-nbitq), 
to_sfixed(-375467470.0/4294967296.0,1,-nbitq), 
to_sfixed(244067053.0/4294967296.0,1,-nbitq), 
to_sfixed(-152834458.0/4294967296.0,1,-nbitq), 
to_sfixed(-185029252.0/4294967296.0,1,-nbitq), 
to_sfixed(-392661646.0/4294967296.0,1,-nbitq), 
to_sfixed(-255857859.0/4294967296.0,1,-nbitq), 
to_sfixed(-40574704.0/4294967296.0,1,-nbitq), 
to_sfixed(195957055.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(267681357.0/4294967296.0,1,-nbitq), 
to_sfixed(-447262289.0/4294967296.0,1,-nbitq), 
to_sfixed(-180667318.0/4294967296.0,1,-nbitq), 
to_sfixed(-68030366.0/4294967296.0,1,-nbitq), 
to_sfixed(-202059476.0/4294967296.0,1,-nbitq), 
to_sfixed(21597410.0/4294967296.0,1,-nbitq), 
to_sfixed(395117113.0/4294967296.0,1,-nbitq), 
to_sfixed(255719132.0/4294967296.0,1,-nbitq), 
to_sfixed(-412520441.0/4294967296.0,1,-nbitq), 
to_sfixed(-216158493.0/4294967296.0,1,-nbitq), 
to_sfixed(294552778.0/4294967296.0,1,-nbitq), 
to_sfixed(385060985.0/4294967296.0,1,-nbitq), 
to_sfixed(135440274.0/4294967296.0,1,-nbitq), 
to_sfixed(-170334155.0/4294967296.0,1,-nbitq), 
to_sfixed(125712545.0/4294967296.0,1,-nbitq), 
to_sfixed(881868.0/4294967296.0,1,-nbitq), 
to_sfixed(-116360673.0/4294967296.0,1,-nbitq), 
to_sfixed(-370830294.0/4294967296.0,1,-nbitq), 
to_sfixed(148167005.0/4294967296.0,1,-nbitq), 
to_sfixed(319388015.0/4294967296.0,1,-nbitq), 
to_sfixed(-340336842.0/4294967296.0,1,-nbitq), 
to_sfixed(439541128.0/4294967296.0,1,-nbitq), 
to_sfixed(-29072006.0/4294967296.0,1,-nbitq), 
to_sfixed(81423507.0/4294967296.0,1,-nbitq), 
to_sfixed(11879028.0/4294967296.0,1,-nbitq), 
to_sfixed(388800299.0/4294967296.0,1,-nbitq), 
to_sfixed(-149172281.0/4294967296.0,1,-nbitq), 
to_sfixed(125245910.0/4294967296.0,1,-nbitq), 
to_sfixed(468608405.0/4294967296.0,1,-nbitq), 
to_sfixed(31214399.0/4294967296.0,1,-nbitq), 
to_sfixed(-69010049.0/4294967296.0,1,-nbitq), 
to_sfixed(-457073252.0/4294967296.0,1,-nbitq), 
to_sfixed(-318370814.0/4294967296.0,1,-nbitq), 
to_sfixed(59992536.0/4294967296.0,1,-nbitq), 
to_sfixed(353476706.0/4294967296.0,1,-nbitq), 
to_sfixed(-252604499.0/4294967296.0,1,-nbitq), 
to_sfixed(35393653.0/4294967296.0,1,-nbitq), 
to_sfixed(-165521004.0/4294967296.0,1,-nbitq), 
to_sfixed(234907567.0/4294967296.0,1,-nbitq), 
to_sfixed(490073577.0/4294967296.0,1,-nbitq), 
to_sfixed(305636559.0/4294967296.0,1,-nbitq), 
to_sfixed(-115158680.0/4294967296.0,1,-nbitq), 
to_sfixed(283672030.0/4294967296.0,1,-nbitq), 
to_sfixed(-358798605.0/4294967296.0,1,-nbitq), 
to_sfixed(393976620.0/4294967296.0,1,-nbitq), 
to_sfixed(88251613.0/4294967296.0,1,-nbitq), 
to_sfixed(-423113589.0/4294967296.0,1,-nbitq), 
to_sfixed(-154524644.0/4294967296.0,1,-nbitq), 
to_sfixed(-45786233.0/4294967296.0,1,-nbitq), 
to_sfixed(-217791837.0/4294967296.0,1,-nbitq), 
to_sfixed(382547965.0/4294967296.0,1,-nbitq), 
to_sfixed(193210153.0/4294967296.0,1,-nbitq), 
to_sfixed(-105713152.0/4294967296.0,1,-nbitq), 
to_sfixed(-784788.0/4294967296.0,1,-nbitq), 
to_sfixed(535378651.0/4294967296.0,1,-nbitq), 
to_sfixed(55241726.0/4294967296.0,1,-nbitq), 
to_sfixed(386689481.0/4294967296.0,1,-nbitq), 
to_sfixed(-392858948.0/4294967296.0,1,-nbitq), 
to_sfixed(-360326504.0/4294967296.0,1,-nbitq), 
to_sfixed(119888361.0/4294967296.0,1,-nbitq), 
to_sfixed(-28065099.0/4294967296.0,1,-nbitq), 
to_sfixed(-56470721.0/4294967296.0,1,-nbitq), 
to_sfixed(-173107810.0/4294967296.0,1,-nbitq), 
to_sfixed(-12934821.0/4294967296.0,1,-nbitq), 
to_sfixed(-28722167.0/4294967296.0,1,-nbitq), 
to_sfixed(-428189789.0/4294967296.0,1,-nbitq), 
to_sfixed(23878683.0/4294967296.0,1,-nbitq), 
to_sfixed(-440949032.0/4294967296.0,1,-nbitq), 
to_sfixed(14959481.0/4294967296.0,1,-nbitq), 
to_sfixed(-126119155.0/4294967296.0,1,-nbitq), 
to_sfixed(-62226174.0/4294967296.0,1,-nbitq), 
to_sfixed(-103250260.0/4294967296.0,1,-nbitq), 
to_sfixed(-428696515.0/4294967296.0,1,-nbitq), 
to_sfixed(23595957.0/4294967296.0,1,-nbitq), 
to_sfixed(-107783508.0/4294967296.0,1,-nbitq), 
to_sfixed(-439438016.0/4294967296.0,1,-nbitq), 
to_sfixed(-294605431.0/4294967296.0,1,-nbitq), 
to_sfixed(15666148.0/4294967296.0,1,-nbitq), 
to_sfixed(-46178179.0/4294967296.0,1,-nbitq), 
to_sfixed(153953092.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(57658960.0/4294967296.0,1,-nbitq), 
to_sfixed(-138210733.0/4294967296.0,1,-nbitq), 
to_sfixed(233665754.0/4294967296.0,1,-nbitq), 
to_sfixed(-391387434.0/4294967296.0,1,-nbitq), 
to_sfixed(515400932.0/4294967296.0,1,-nbitq), 
to_sfixed(-284416127.0/4294967296.0,1,-nbitq), 
to_sfixed(129915132.0/4294967296.0,1,-nbitq), 
to_sfixed(-341257190.0/4294967296.0,1,-nbitq), 
to_sfixed(-413075994.0/4294967296.0,1,-nbitq), 
to_sfixed(123751781.0/4294967296.0,1,-nbitq), 
to_sfixed(206974357.0/4294967296.0,1,-nbitq), 
to_sfixed(162850325.0/4294967296.0,1,-nbitq), 
to_sfixed(98431631.0/4294967296.0,1,-nbitq), 
to_sfixed(-73890751.0/4294967296.0,1,-nbitq), 
to_sfixed(415588128.0/4294967296.0,1,-nbitq), 
to_sfixed(-166598676.0/4294967296.0,1,-nbitq), 
to_sfixed(-29794299.0/4294967296.0,1,-nbitq), 
to_sfixed(8661959.0/4294967296.0,1,-nbitq), 
to_sfixed(343532960.0/4294967296.0,1,-nbitq), 
to_sfixed(335927754.0/4294967296.0,1,-nbitq), 
to_sfixed(-363348352.0/4294967296.0,1,-nbitq), 
to_sfixed(35730490.0/4294967296.0,1,-nbitq), 
to_sfixed(632872908.0/4294967296.0,1,-nbitq), 
to_sfixed(166549761.0/4294967296.0,1,-nbitq), 
to_sfixed(-115157729.0/4294967296.0,1,-nbitq), 
to_sfixed(329399677.0/4294967296.0,1,-nbitq), 
to_sfixed(293543969.0/4294967296.0,1,-nbitq), 
to_sfixed(53487383.0/4294967296.0,1,-nbitq), 
to_sfixed(-280212970.0/4294967296.0,1,-nbitq), 
to_sfixed(-419059348.0/4294967296.0,1,-nbitq), 
to_sfixed(-459889419.0/4294967296.0,1,-nbitq), 
to_sfixed(-367897337.0/4294967296.0,1,-nbitq), 
to_sfixed(75055020.0/4294967296.0,1,-nbitq), 
to_sfixed(2410050.0/4294967296.0,1,-nbitq), 
to_sfixed(60783390.0/4294967296.0,1,-nbitq), 
to_sfixed(251705150.0/4294967296.0,1,-nbitq), 
to_sfixed(-29864495.0/4294967296.0,1,-nbitq), 
to_sfixed(92941760.0/4294967296.0,1,-nbitq), 
to_sfixed(-341072191.0/4294967296.0,1,-nbitq), 
to_sfixed(415810038.0/4294967296.0,1,-nbitq), 
to_sfixed(49764850.0/4294967296.0,1,-nbitq), 
to_sfixed(28934061.0/4294967296.0,1,-nbitq), 
to_sfixed(-326822877.0/4294967296.0,1,-nbitq), 
to_sfixed(-207594239.0/4294967296.0,1,-nbitq), 
to_sfixed(-122564406.0/4294967296.0,1,-nbitq), 
to_sfixed(539503523.0/4294967296.0,1,-nbitq), 
to_sfixed(312449325.0/4294967296.0,1,-nbitq), 
to_sfixed(18600293.0/4294967296.0,1,-nbitq), 
to_sfixed(356953055.0/4294967296.0,1,-nbitq), 
to_sfixed(336246205.0/4294967296.0,1,-nbitq), 
to_sfixed(249904517.0/4294967296.0,1,-nbitq), 
to_sfixed(-209391457.0/4294967296.0,1,-nbitq), 
to_sfixed(-335784559.0/4294967296.0,1,-nbitq), 
to_sfixed(431407573.0/4294967296.0,1,-nbitq), 
to_sfixed(483479383.0/4294967296.0,1,-nbitq), 
to_sfixed(37444147.0/4294967296.0,1,-nbitq), 
to_sfixed(-50288270.0/4294967296.0,1,-nbitq), 
to_sfixed(-586062172.0/4294967296.0,1,-nbitq), 
to_sfixed(22726968.0/4294967296.0,1,-nbitq), 
to_sfixed(166438462.0/4294967296.0,1,-nbitq), 
to_sfixed(-15174998.0/4294967296.0,1,-nbitq), 
to_sfixed(370168216.0/4294967296.0,1,-nbitq), 
to_sfixed(-222072865.0/4294967296.0,1,-nbitq), 
to_sfixed(-54378699.0/4294967296.0,1,-nbitq), 
to_sfixed(168484131.0/4294967296.0,1,-nbitq), 
to_sfixed(37144053.0/4294967296.0,1,-nbitq), 
to_sfixed(-34473028.0/4294967296.0,1,-nbitq), 
to_sfixed(118959764.0/4294967296.0,1,-nbitq), 
to_sfixed(280725490.0/4294967296.0,1,-nbitq), 
to_sfixed(468309230.0/4294967296.0,1,-nbitq), 
to_sfixed(-424178147.0/4294967296.0,1,-nbitq), 
to_sfixed(193079372.0/4294967296.0,1,-nbitq), 
to_sfixed(-131899244.0/4294967296.0,1,-nbitq), 
to_sfixed(-49180955.0/4294967296.0,1,-nbitq), 
to_sfixed(426021582.0/4294967296.0,1,-nbitq), 
to_sfixed(-526382182.0/4294967296.0,1,-nbitq), 
to_sfixed(-272782814.0/4294967296.0,1,-nbitq), 
to_sfixed(-219779370.0/4294967296.0,1,-nbitq), 
to_sfixed(6155680.0/4294967296.0,1,-nbitq), 
to_sfixed(-134520191.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(263521967.0/4294967296.0,1,-nbitq), 
to_sfixed(-497018989.0/4294967296.0,1,-nbitq), 
to_sfixed(-422792051.0/4294967296.0,1,-nbitq), 
to_sfixed(-404838927.0/4294967296.0,1,-nbitq), 
to_sfixed(103630170.0/4294967296.0,1,-nbitq), 
to_sfixed(219106640.0/4294967296.0,1,-nbitq), 
to_sfixed(341986649.0/4294967296.0,1,-nbitq), 
to_sfixed(-72176099.0/4294967296.0,1,-nbitq), 
to_sfixed(-390616369.0/4294967296.0,1,-nbitq), 
to_sfixed(-158298655.0/4294967296.0,1,-nbitq), 
to_sfixed(-111717046.0/4294967296.0,1,-nbitq), 
to_sfixed(355860333.0/4294967296.0,1,-nbitq), 
to_sfixed(13604564.0/4294967296.0,1,-nbitq), 
to_sfixed(286037679.0/4294967296.0,1,-nbitq), 
to_sfixed(-263120199.0/4294967296.0,1,-nbitq), 
to_sfixed(32098731.0/4294967296.0,1,-nbitq), 
to_sfixed(-280176537.0/4294967296.0,1,-nbitq), 
to_sfixed(-271426060.0/4294967296.0,1,-nbitq), 
to_sfixed(242177036.0/4294967296.0,1,-nbitq), 
to_sfixed(33033537.0/4294967296.0,1,-nbitq), 
to_sfixed(-91202558.0/4294967296.0,1,-nbitq), 
to_sfixed(139523361.0/4294967296.0,1,-nbitq), 
to_sfixed(735676333.0/4294967296.0,1,-nbitq), 
to_sfixed(-189345142.0/4294967296.0,1,-nbitq), 
to_sfixed(-80373548.0/4294967296.0,1,-nbitq), 
to_sfixed(91881491.0/4294967296.0,1,-nbitq), 
to_sfixed(422489493.0/4294967296.0,1,-nbitq), 
to_sfixed(-211751014.0/4294967296.0,1,-nbitq), 
to_sfixed(-195418187.0/4294967296.0,1,-nbitq), 
to_sfixed(197782059.0/4294967296.0,1,-nbitq), 
to_sfixed(-263281085.0/4294967296.0,1,-nbitq), 
to_sfixed(-404347538.0/4294967296.0,1,-nbitq), 
to_sfixed(227171768.0/4294967296.0,1,-nbitq), 
to_sfixed(-415180417.0/4294967296.0,1,-nbitq), 
to_sfixed(473928430.0/4294967296.0,1,-nbitq), 
to_sfixed(-392206990.0/4294967296.0,1,-nbitq), 
to_sfixed(2432674.0/4294967296.0,1,-nbitq), 
to_sfixed(73689342.0/4294967296.0,1,-nbitq), 
to_sfixed(92917689.0/4294967296.0,1,-nbitq), 
to_sfixed(-47300982.0/4294967296.0,1,-nbitq), 
to_sfixed(224939305.0/4294967296.0,1,-nbitq), 
to_sfixed(-88968799.0/4294967296.0,1,-nbitq), 
to_sfixed(355441405.0/4294967296.0,1,-nbitq), 
to_sfixed(-66229699.0/4294967296.0,1,-nbitq), 
to_sfixed(639885570.0/4294967296.0,1,-nbitq), 
to_sfixed(76436913.0/4294967296.0,1,-nbitq), 
to_sfixed(240325924.0/4294967296.0,1,-nbitq), 
to_sfixed(186336825.0/4294967296.0,1,-nbitq), 
to_sfixed(80599948.0/4294967296.0,1,-nbitq), 
to_sfixed(95430149.0/4294967296.0,1,-nbitq), 
to_sfixed(-140426792.0/4294967296.0,1,-nbitq), 
to_sfixed(230217457.0/4294967296.0,1,-nbitq), 
to_sfixed(146888798.0/4294967296.0,1,-nbitq), 
to_sfixed(-421625334.0/4294967296.0,1,-nbitq), 
to_sfixed(118526790.0/4294967296.0,1,-nbitq), 
to_sfixed(-245411450.0/4294967296.0,1,-nbitq), 
to_sfixed(116543326.0/4294967296.0,1,-nbitq), 
to_sfixed(-55244720.0/4294967296.0,1,-nbitq), 
to_sfixed(168555809.0/4294967296.0,1,-nbitq), 
to_sfixed(-364705535.0/4294967296.0,1,-nbitq), 
to_sfixed(-251449342.0/4294967296.0,1,-nbitq), 
to_sfixed(-216565304.0/4294967296.0,1,-nbitq), 
to_sfixed(6903535.0/4294967296.0,1,-nbitq), 
to_sfixed(101858506.0/4294967296.0,1,-nbitq), 
to_sfixed(86208079.0/4294967296.0,1,-nbitq), 
to_sfixed(-190184792.0/4294967296.0,1,-nbitq), 
to_sfixed(492879371.0/4294967296.0,1,-nbitq), 
to_sfixed(316021439.0/4294967296.0,1,-nbitq), 
to_sfixed(-309238382.0/4294967296.0,1,-nbitq), 
to_sfixed(148665389.0/4294967296.0,1,-nbitq), 
to_sfixed(-168300594.0/4294967296.0,1,-nbitq), 
to_sfixed(-143782782.0/4294967296.0,1,-nbitq), 
to_sfixed(-149674920.0/4294967296.0,1,-nbitq), 
to_sfixed(328938570.0/4294967296.0,1,-nbitq), 
to_sfixed(371226931.0/4294967296.0,1,-nbitq), 
to_sfixed(-412419547.0/4294967296.0,1,-nbitq), 
to_sfixed(291719751.0/4294967296.0,1,-nbitq), 
to_sfixed(-231190442.0/4294967296.0,1,-nbitq), 
to_sfixed(-562576732.0/4294967296.0,1,-nbitq), 
to_sfixed(4141864.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(39760710.0/4294967296.0,1,-nbitq), 
to_sfixed(-204018525.0/4294967296.0,1,-nbitq), 
to_sfixed(-329752726.0/4294967296.0,1,-nbitq), 
to_sfixed(71127678.0/4294967296.0,1,-nbitq), 
to_sfixed(-231013521.0/4294967296.0,1,-nbitq), 
to_sfixed(242934030.0/4294967296.0,1,-nbitq), 
to_sfixed(155372294.0/4294967296.0,1,-nbitq), 
to_sfixed(-349944885.0/4294967296.0,1,-nbitq), 
to_sfixed(-62440447.0/4294967296.0,1,-nbitq), 
to_sfixed(201570308.0/4294967296.0,1,-nbitq), 
to_sfixed(-187322447.0/4294967296.0,1,-nbitq), 
to_sfixed(-178181560.0/4294967296.0,1,-nbitq), 
to_sfixed(-316275292.0/4294967296.0,1,-nbitq), 
to_sfixed(-317129603.0/4294967296.0,1,-nbitq), 
to_sfixed(129060868.0/4294967296.0,1,-nbitq), 
to_sfixed(203075566.0/4294967296.0,1,-nbitq), 
to_sfixed(-47073055.0/4294967296.0,1,-nbitq), 
to_sfixed(-7871814.0/4294967296.0,1,-nbitq), 
to_sfixed(737652380.0/4294967296.0,1,-nbitq), 
to_sfixed(174991909.0/4294967296.0,1,-nbitq), 
to_sfixed(-22842645.0/4294967296.0,1,-nbitq), 
to_sfixed(88739384.0/4294967296.0,1,-nbitq), 
to_sfixed(261914401.0/4294967296.0,1,-nbitq), 
to_sfixed(328387720.0/4294967296.0,1,-nbitq), 
to_sfixed(-263307340.0/4294967296.0,1,-nbitq), 
to_sfixed(366889284.0/4294967296.0,1,-nbitq), 
to_sfixed(303430629.0/4294967296.0,1,-nbitq), 
to_sfixed(-395933201.0/4294967296.0,1,-nbitq), 
to_sfixed(-254884225.0/4294967296.0,1,-nbitq), 
to_sfixed(-578673583.0/4294967296.0,1,-nbitq), 
to_sfixed(-58551185.0/4294967296.0,1,-nbitq), 
to_sfixed(270148943.0/4294967296.0,1,-nbitq), 
to_sfixed(157339076.0/4294967296.0,1,-nbitq), 
to_sfixed(176172400.0/4294967296.0,1,-nbitq), 
to_sfixed(-150152631.0/4294967296.0,1,-nbitq), 
to_sfixed(-90881798.0/4294967296.0,1,-nbitq), 
to_sfixed(317369324.0/4294967296.0,1,-nbitq), 
to_sfixed(-201635093.0/4294967296.0,1,-nbitq), 
to_sfixed(-233221921.0/4294967296.0,1,-nbitq), 
to_sfixed(-42820837.0/4294967296.0,1,-nbitq), 
to_sfixed(1284259.0/4294967296.0,1,-nbitq), 
to_sfixed(-259266029.0/4294967296.0,1,-nbitq), 
to_sfixed(180284854.0/4294967296.0,1,-nbitq), 
to_sfixed(69723143.0/4294967296.0,1,-nbitq), 
to_sfixed(43772979.0/4294967296.0,1,-nbitq), 
to_sfixed(478434904.0/4294967296.0,1,-nbitq), 
to_sfixed(70920051.0/4294967296.0,1,-nbitq), 
to_sfixed(321213082.0/4294967296.0,1,-nbitq), 
to_sfixed(-143363113.0/4294967296.0,1,-nbitq), 
to_sfixed(-132589227.0/4294967296.0,1,-nbitq), 
to_sfixed(79184888.0/4294967296.0,1,-nbitq), 
to_sfixed(239216056.0/4294967296.0,1,-nbitq), 
to_sfixed(-350939626.0/4294967296.0,1,-nbitq), 
to_sfixed(-372847835.0/4294967296.0,1,-nbitq), 
to_sfixed(93910978.0/4294967296.0,1,-nbitq), 
to_sfixed(375214683.0/4294967296.0,1,-nbitq), 
to_sfixed(-264523296.0/4294967296.0,1,-nbitq), 
to_sfixed(182180295.0/4294967296.0,1,-nbitq), 
to_sfixed(-299094794.0/4294967296.0,1,-nbitq), 
to_sfixed(-68436213.0/4294967296.0,1,-nbitq), 
to_sfixed(-365222834.0/4294967296.0,1,-nbitq), 
to_sfixed(251793916.0/4294967296.0,1,-nbitq), 
to_sfixed(-367874943.0/4294967296.0,1,-nbitq), 
to_sfixed(142614549.0/4294967296.0,1,-nbitq), 
to_sfixed(-240526383.0/4294967296.0,1,-nbitq), 
to_sfixed(298980715.0/4294967296.0,1,-nbitq), 
to_sfixed(191383527.0/4294967296.0,1,-nbitq), 
to_sfixed(-7652329.0/4294967296.0,1,-nbitq), 
to_sfixed(9109127.0/4294967296.0,1,-nbitq), 
to_sfixed(-255190685.0/4294967296.0,1,-nbitq), 
to_sfixed(-350051747.0/4294967296.0,1,-nbitq), 
to_sfixed(192587004.0/4294967296.0,1,-nbitq), 
to_sfixed(-332008071.0/4294967296.0,1,-nbitq), 
to_sfixed(-202235221.0/4294967296.0,1,-nbitq), 
to_sfixed(103814100.0/4294967296.0,1,-nbitq), 
to_sfixed(-119862106.0/4294967296.0,1,-nbitq), 
to_sfixed(315779536.0/4294967296.0,1,-nbitq), 
to_sfixed(-316724032.0/4294967296.0,1,-nbitq), 
to_sfixed(-154483038.0/4294967296.0,1,-nbitq), 
to_sfixed(-80777867.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(44289346.0/4294967296.0,1,-nbitq), 
to_sfixed(-429760336.0/4294967296.0,1,-nbitq), 
to_sfixed(-52475257.0/4294967296.0,1,-nbitq), 
to_sfixed(414115241.0/4294967296.0,1,-nbitq), 
to_sfixed(454034875.0/4294967296.0,1,-nbitq), 
to_sfixed(-397853077.0/4294967296.0,1,-nbitq), 
to_sfixed(-377732200.0/4294967296.0,1,-nbitq), 
to_sfixed(186310555.0/4294967296.0,1,-nbitq), 
to_sfixed(-201761073.0/4294967296.0,1,-nbitq), 
to_sfixed(118104604.0/4294967296.0,1,-nbitq), 
to_sfixed(178933323.0/4294967296.0,1,-nbitq), 
to_sfixed(-281432005.0/4294967296.0,1,-nbitq), 
to_sfixed(-177329204.0/4294967296.0,1,-nbitq), 
to_sfixed(238905946.0/4294967296.0,1,-nbitq), 
to_sfixed(-97761847.0/4294967296.0,1,-nbitq), 
to_sfixed(-558919353.0/4294967296.0,1,-nbitq), 
to_sfixed(288013509.0/4294967296.0,1,-nbitq), 
to_sfixed(322220041.0/4294967296.0,1,-nbitq), 
to_sfixed(200437160.0/4294967296.0,1,-nbitq), 
to_sfixed(-76531982.0/4294967296.0,1,-nbitq), 
to_sfixed(298920109.0/4294967296.0,1,-nbitq), 
to_sfixed(17786626.0/4294967296.0,1,-nbitq), 
to_sfixed(434677999.0/4294967296.0,1,-nbitq), 
to_sfixed(145318203.0/4294967296.0,1,-nbitq), 
to_sfixed(-328731346.0/4294967296.0,1,-nbitq), 
to_sfixed(519738287.0/4294967296.0,1,-nbitq), 
to_sfixed(-255119794.0/4294967296.0,1,-nbitq), 
to_sfixed(-227783841.0/4294967296.0,1,-nbitq), 
to_sfixed(171462410.0/4294967296.0,1,-nbitq), 
to_sfixed(-117643340.0/4294967296.0,1,-nbitq), 
to_sfixed(-88777037.0/4294967296.0,1,-nbitq), 
to_sfixed(308001359.0/4294967296.0,1,-nbitq), 
to_sfixed(65270619.0/4294967296.0,1,-nbitq), 
to_sfixed(-152001923.0/4294967296.0,1,-nbitq), 
to_sfixed(-133291174.0/4294967296.0,1,-nbitq), 
to_sfixed(-309522955.0/4294967296.0,1,-nbitq), 
to_sfixed(233628373.0/4294967296.0,1,-nbitq), 
to_sfixed(105824992.0/4294967296.0,1,-nbitq), 
to_sfixed(221593947.0/4294967296.0,1,-nbitq), 
to_sfixed(14066746.0/4294967296.0,1,-nbitq), 
to_sfixed(117426837.0/4294967296.0,1,-nbitq), 
to_sfixed(-119522195.0/4294967296.0,1,-nbitq), 
to_sfixed(368170639.0/4294967296.0,1,-nbitq), 
to_sfixed(-499451600.0/4294967296.0,1,-nbitq), 
to_sfixed(511042091.0/4294967296.0,1,-nbitq), 
to_sfixed(23237434.0/4294967296.0,1,-nbitq), 
to_sfixed(-370841288.0/4294967296.0,1,-nbitq), 
to_sfixed(340100301.0/4294967296.0,1,-nbitq), 
to_sfixed(327195106.0/4294967296.0,1,-nbitq), 
to_sfixed(482508937.0/4294967296.0,1,-nbitq), 
to_sfixed(-105028342.0/4294967296.0,1,-nbitq), 
to_sfixed(-163959278.0/4294967296.0,1,-nbitq), 
to_sfixed(-186149189.0/4294967296.0,1,-nbitq), 
to_sfixed(-200014707.0/4294967296.0,1,-nbitq), 
to_sfixed(-290253947.0/4294967296.0,1,-nbitq), 
to_sfixed(-205992443.0/4294967296.0,1,-nbitq), 
to_sfixed(-417961059.0/4294967296.0,1,-nbitq), 
to_sfixed(-36506911.0/4294967296.0,1,-nbitq), 
to_sfixed(-264542353.0/4294967296.0,1,-nbitq), 
to_sfixed(-112533176.0/4294967296.0,1,-nbitq), 
to_sfixed(38785824.0/4294967296.0,1,-nbitq), 
to_sfixed(-254016987.0/4294967296.0,1,-nbitq), 
to_sfixed(34139810.0/4294967296.0,1,-nbitq), 
to_sfixed(-5994720.0/4294967296.0,1,-nbitq), 
to_sfixed(-360336898.0/4294967296.0,1,-nbitq), 
to_sfixed(-326241661.0/4294967296.0,1,-nbitq), 
to_sfixed(530700081.0/4294967296.0,1,-nbitq), 
to_sfixed(-215983873.0/4294967296.0,1,-nbitq), 
to_sfixed(185548623.0/4294967296.0,1,-nbitq), 
to_sfixed(-49763757.0/4294967296.0,1,-nbitq), 
to_sfixed(-537057444.0/4294967296.0,1,-nbitq), 
to_sfixed(-183372063.0/4294967296.0,1,-nbitq), 
to_sfixed(313204302.0/4294967296.0,1,-nbitq), 
to_sfixed(372446316.0/4294967296.0,1,-nbitq), 
to_sfixed(-162246567.0/4294967296.0,1,-nbitq), 
to_sfixed(75115454.0/4294967296.0,1,-nbitq), 
to_sfixed(268547857.0/4294967296.0,1,-nbitq), 
to_sfixed(-91674790.0/4294967296.0,1,-nbitq), 
to_sfixed(-206097325.0/4294967296.0,1,-nbitq), 
to_sfixed(167123096.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(215815622.0/4294967296.0,1,-nbitq), 
to_sfixed(-113242754.0/4294967296.0,1,-nbitq), 
to_sfixed(-50357136.0/4294967296.0,1,-nbitq), 
to_sfixed(120558867.0/4294967296.0,1,-nbitq), 
to_sfixed(-160082068.0/4294967296.0,1,-nbitq), 
to_sfixed(-63590358.0/4294967296.0,1,-nbitq), 
to_sfixed(-195608037.0/4294967296.0,1,-nbitq), 
to_sfixed(130576294.0/4294967296.0,1,-nbitq), 
to_sfixed(-46598614.0/4294967296.0,1,-nbitq), 
to_sfixed(-296725110.0/4294967296.0,1,-nbitq), 
to_sfixed(102981425.0/4294967296.0,1,-nbitq), 
to_sfixed(168575164.0/4294967296.0,1,-nbitq), 
to_sfixed(-547720724.0/4294967296.0,1,-nbitq), 
to_sfixed(-194542078.0/4294967296.0,1,-nbitq), 
to_sfixed(246672843.0/4294967296.0,1,-nbitq), 
to_sfixed(-678438157.0/4294967296.0,1,-nbitq), 
to_sfixed(-90051990.0/4294967296.0,1,-nbitq), 
to_sfixed(-4569093.0/4294967296.0,1,-nbitq), 
to_sfixed(481225909.0/4294967296.0,1,-nbitq), 
to_sfixed(341845248.0/4294967296.0,1,-nbitq), 
to_sfixed(280952545.0/4294967296.0,1,-nbitq), 
to_sfixed(431266505.0/4294967296.0,1,-nbitq), 
to_sfixed(801558944.0/4294967296.0,1,-nbitq), 
to_sfixed(-636909320.0/4294967296.0,1,-nbitq), 
to_sfixed(-272708204.0/4294967296.0,1,-nbitq), 
to_sfixed(10036930.0/4294967296.0,1,-nbitq), 
to_sfixed(-200115859.0/4294967296.0,1,-nbitq), 
to_sfixed(-71029401.0/4294967296.0,1,-nbitq), 
to_sfixed(52519284.0/4294967296.0,1,-nbitq), 
to_sfixed(-639203503.0/4294967296.0,1,-nbitq), 
to_sfixed(173621450.0/4294967296.0,1,-nbitq), 
to_sfixed(43069185.0/4294967296.0,1,-nbitq), 
to_sfixed(-464240722.0/4294967296.0,1,-nbitq), 
to_sfixed(301016285.0/4294967296.0,1,-nbitq), 
to_sfixed(283906157.0/4294967296.0,1,-nbitq), 
to_sfixed(-394688626.0/4294967296.0,1,-nbitq), 
to_sfixed(349740700.0/4294967296.0,1,-nbitq), 
to_sfixed(-496191675.0/4294967296.0,1,-nbitq), 
to_sfixed(27624368.0/4294967296.0,1,-nbitq), 
to_sfixed(152710353.0/4294967296.0,1,-nbitq), 
to_sfixed(398613789.0/4294967296.0,1,-nbitq), 
to_sfixed(-271275347.0/4294967296.0,1,-nbitq), 
to_sfixed(423424667.0/4294967296.0,1,-nbitq), 
to_sfixed(42641233.0/4294967296.0,1,-nbitq), 
to_sfixed(660207794.0/4294967296.0,1,-nbitq), 
to_sfixed(427819521.0/4294967296.0,1,-nbitq), 
to_sfixed(329588293.0/4294967296.0,1,-nbitq), 
to_sfixed(396417614.0/4294967296.0,1,-nbitq), 
to_sfixed(-41820641.0/4294967296.0,1,-nbitq), 
to_sfixed(-28225840.0/4294967296.0,1,-nbitq), 
to_sfixed(-8240804.0/4294967296.0,1,-nbitq), 
to_sfixed(227178489.0/4294967296.0,1,-nbitq), 
to_sfixed(-31682463.0/4294967296.0,1,-nbitq), 
to_sfixed(-646156386.0/4294967296.0,1,-nbitq), 
to_sfixed(341265056.0/4294967296.0,1,-nbitq), 
to_sfixed(186439491.0/4294967296.0,1,-nbitq), 
to_sfixed(-105628480.0/4294967296.0,1,-nbitq), 
to_sfixed(-43566196.0/4294967296.0,1,-nbitq), 
to_sfixed(215880745.0/4294967296.0,1,-nbitq), 
to_sfixed(-107570585.0/4294967296.0,1,-nbitq), 
to_sfixed(-74651756.0/4294967296.0,1,-nbitq), 
to_sfixed(-273756844.0/4294967296.0,1,-nbitq), 
to_sfixed(411930530.0/4294967296.0,1,-nbitq), 
to_sfixed(-215725330.0/4294967296.0,1,-nbitq), 
to_sfixed(311675494.0/4294967296.0,1,-nbitq), 
to_sfixed(16890533.0/4294967296.0,1,-nbitq), 
to_sfixed(218050681.0/4294967296.0,1,-nbitq), 
to_sfixed(-588050871.0/4294967296.0,1,-nbitq), 
to_sfixed(-333260131.0/4294967296.0,1,-nbitq), 
to_sfixed(90316180.0/4294967296.0,1,-nbitq), 
to_sfixed(-393182961.0/4294967296.0,1,-nbitq), 
to_sfixed(-297309173.0/4294967296.0,1,-nbitq), 
to_sfixed(-198234236.0/4294967296.0,1,-nbitq), 
to_sfixed(448282333.0/4294967296.0,1,-nbitq), 
to_sfixed(-112529510.0/4294967296.0,1,-nbitq), 
to_sfixed(-97417945.0/4294967296.0,1,-nbitq), 
to_sfixed(226757793.0/4294967296.0,1,-nbitq), 
to_sfixed(85794321.0/4294967296.0,1,-nbitq), 
to_sfixed(206134146.0/4294967296.0,1,-nbitq), 
to_sfixed(-99244295.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-353328330.0/4294967296.0,1,-nbitq), 
to_sfixed(50336004.0/4294967296.0,1,-nbitq), 
to_sfixed(33861613.0/4294967296.0,1,-nbitq), 
to_sfixed(-10118308.0/4294967296.0,1,-nbitq), 
to_sfixed(-74520898.0/4294967296.0,1,-nbitq), 
to_sfixed(-288781425.0/4294967296.0,1,-nbitq), 
to_sfixed(-285761829.0/4294967296.0,1,-nbitq), 
to_sfixed(-274104919.0/4294967296.0,1,-nbitq), 
to_sfixed(284834593.0/4294967296.0,1,-nbitq), 
to_sfixed(-349547068.0/4294967296.0,1,-nbitq), 
to_sfixed(-86021983.0/4294967296.0,1,-nbitq), 
to_sfixed(401296088.0/4294967296.0,1,-nbitq), 
to_sfixed(-530748678.0/4294967296.0,1,-nbitq), 
to_sfixed(-426976321.0/4294967296.0,1,-nbitq), 
to_sfixed(-188742511.0/4294967296.0,1,-nbitq), 
to_sfixed(-221873590.0/4294967296.0,1,-nbitq), 
to_sfixed(193449414.0/4294967296.0,1,-nbitq), 
to_sfixed(397499526.0/4294967296.0,1,-nbitq), 
to_sfixed(600340405.0/4294967296.0,1,-nbitq), 
to_sfixed(244767992.0/4294967296.0,1,-nbitq), 
to_sfixed(-335390973.0/4294967296.0,1,-nbitq), 
to_sfixed(451588678.0/4294967296.0,1,-nbitq), 
to_sfixed(98086485.0/4294967296.0,1,-nbitq), 
to_sfixed(-224419148.0/4294967296.0,1,-nbitq), 
to_sfixed(319921446.0/4294967296.0,1,-nbitq), 
to_sfixed(-616427526.0/4294967296.0,1,-nbitq), 
to_sfixed(-101112305.0/4294967296.0,1,-nbitq), 
to_sfixed(62624046.0/4294967296.0,1,-nbitq), 
to_sfixed(12443399.0/4294967296.0,1,-nbitq), 
to_sfixed(-120656400.0/4294967296.0,1,-nbitq), 
to_sfixed(-629543176.0/4294967296.0,1,-nbitq), 
to_sfixed(-437906491.0/4294967296.0,1,-nbitq), 
to_sfixed(4157014.0/4294967296.0,1,-nbitq), 
to_sfixed(538798079.0/4294967296.0,1,-nbitq), 
to_sfixed(202746058.0/4294967296.0,1,-nbitq), 
to_sfixed(-694157934.0/4294967296.0,1,-nbitq), 
to_sfixed(19095101.0/4294967296.0,1,-nbitq), 
to_sfixed(-99338058.0/4294967296.0,1,-nbitq), 
to_sfixed(226527453.0/4294967296.0,1,-nbitq), 
to_sfixed(379391613.0/4294967296.0,1,-nbitq), 
to_sfixed(469101267.0/4294967296.0,1,-nbitq), 
to_sfixed(-156439893.0/4294967296.0,1,-nbitq), 
to_sfixed(85741699.0/4294967296.0,1,-nbitq), 
to_sfixed(-224971538.0/4294967296.0,1,-nbitq), 
to_sfixed(-35536899.0/4294967296.0,1,-nbitq), 
to_sfixed(614888756.0/4294967296.0,1,-nbitq), 
to_sfixed(305823976.0/4294967296.0,1,-nbitq), 
to_sfixed(303495805.0/4294967296.0,1,-nbitq), 
to_sfixed(-212110827.0/4294967296.0,1,-nbitq), 
to_sfixed(-17355723.0/4294967296.0,1,-nbitq), 
to_sfixed(189125517.0/4294967296.0,1,-nbitq), 
to_sfixed(-193830947.0/4294967296.0,1,-nbitq), 
to_sfixed(-208128054.0/4294967296.0,1,-nbitq), 
to_sfixed(-630171445.0/4294967296.0,1,-nbitq), 
to_sfixed(-330752031.0/4294967296.0,1,-nbitq), 
to_sfixed(-229968442.0/4294967296.0,1,-nbitq), 
to_sfixed(155604287.0/4294967296.0,1,-nbitq), 
to_sfixed(93301733.0/4294967296.0,1,-nbitq), 
to_sfixed(46650246.0/4294967296.0,1,-nbitq), 
to_sfixed(-194576109.0/4294967296.0,1,-nbitq), 
to_sfixed(198639591.0/4294967296.0,1,-nbitq), 
to_sfixed(-19083444.0/4294967296.0,1,-nbitq), 
to_sfixed(-69227698.0/4294967296.0,1,-nbitq), 
to_sfixed(-19084271.0/4294967296.0,1,-nbitq), 
to_sfixed(326554999.0/4294967296.0,1,-nbitq), 
to_sfixed(16534715.0/4294967296.0,1,-nbitq), 
to_sfixed(627000221.0/4294967296.0,1,-nbitq), 
to_sfixed(-639702080.0/4294967296.0,1,-nbitq), 
to_sfixed(-16110325.0/4294967296.0,1,-nbitq), 
to_sfixed(-365754754.0/4294967296.0,1,-nbitq), 
to_sfixed(-352824581.0/4294967296.0,1,-nbitq), 
to_sfixed(-339496806.0/4294967296.0,1,-nbitq), 
to_sfixed(491413013.0/4294967296.0,1,-nbitq), 
to_sfixed(287001921.0/4294967296.0,1,-nbitq), 
to_sfixed(137171871.0/4294967296.0,1,-nbitq), 
to_sfixed(-253830761.0/4294967296.0,1,-nbitq), 
to_sfixed(258508349.0/4294967296.0,1,-nbitq), 
to_sfixed(-551091460.0/4294967296.0,1,-nbitq), 
to_sfixed(-59628715.0/4294967296.0,1,-nbitq), 
to_sfixed(-353906075.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-373859562.0/4294967296.0,1,-nbitq), 
to_sfixed(28215157.0/4294967296.0,1,-nbitq), 
to_sfixed(-332899684.0/4294967296.0,1,-nbitq), 
to_sfixed(-161467146.0/4294967296.0,1,-nbitq), 
to_sfixed(542629077.0/4294967296.0,1,-nbitq), 
to_sfixed(-364795030.0/4294967296.0,1,-nbitq), 
to_sfixed(93015575.0/4294967296.0,1,-nbitq), 
to_sfixed(6051203.0/4294967296.0,1,-nbitq), 
to_sfixed(189298620.0/4294967296.0,1,-nbitq), 
to_sfixed(273520322.0/4294967296.0,1,-nbitq), 
to_sfixed(-257754281.0/4294967296.0,1,-nbitq), 
to_sfixed(351441723.0/4294967296.0,1,-nbitq), 
to_sfixed(-757421774.0/4294967296.0,1,-nbitq), 
to_sfixed(-601712222.0/4294967296.0,1,-nbitq), 
to_sfixed(24137680.0/4294967296.0,1,-nbitq), 
to_sfixed(-672894823.0/4294967296.0,1,-nbitq), 
to_sfixed(-27263153.0/4294967296.0,1,-nbitq), 
to_sfixed(-27354231.0/4294967296.0,1,-nbitq), 
to_sfixed(710623039.0/4294967296.0,1,-nbitq), 
to_sfixed(-47656410.0/4294967296.0,1,-nbitq), 
to_sfixed(-363435148.0/4294967296.0,1,-nbitq), 
to_sfixed(316595776.0/4294967296.0,1,-nbitq), 
to_sfixed(834834841.0/4294967296.0,1,-nbitq), 
to_sfixed(-727582648.0/4294967296.0,1,-nbitq), 
to_sfixed(221760320.0/4294967296.0,1,-nbitq), 
to_sfixed(-691111468.0/4294967296.0,1,-nbitq), 
to_sfixed(293200613.0/4294967296.0,1,-nbitq), 
to_sfixed(266467237.0/4294967296.0,1,-nbitq), 
to_sfixed(-624656309.0/4294967296.0,1,-nbitq), 
to_sfixed(-713028368.0/4294967296.0,1,-nbitq), 
to_sfixed(-754545168.0/4294967296.0,1,-nbitq), 
to_sfixed(-253853176.0/4294967296.0,1,-nbitq), 
to_sfixed(-621597909.0/4294967296.0,1,-nbitq), 
to_sfixed(272241429.0/4294967296.0,1,-nbitq), 
to_sfixed(-511883687.0/4294967296.0,1,-nbitq), 
to_sfixed(-622723196.0/4294967296.0,1,-nbitq), 
to_sfixed(296554370.0/4294967296.0,1,-nbitq), 
to_sfixed(-709884601.0/4294967296.0,1,-nbitq), 
to_sfixed(-37547042.0/4294967296.0,1,-nbitq), 
to_sfixed(162117497.0/4294967296.0,1,-nbitq), 
to_sfixed(-6555172.0/4294967296.0,1,-nbitq), 
to_sfixed(274934906.0/4294967296.0,1,-nbitq), 
to_sfixed(-367211575.0/4294967296.0,1,-nbitq), 
to_sfixed(-37116255.0/4294967296.0,1,-nbitq), 
to_sfixed(527695624.0/4294967296.0,1,-nbitq), 
to_sfixed(56060543.0/4294967296.0,1,-nbitq), 
to_sfixed(291851414.0/4294967296.0,1,-nbitq), 
to_sfixed(180860427.0/4294967296.0,1,-nbitq), 
to_sfixed(3493325.0/4294967296.0,1,-nbitq), 
to_sfixed(21158927.0/4294967296.0,1,-nbitq), 
to_sfixed(345421031.0/4294967296.0,1,-nbitq), 
to_sfixed(-252038906.0/4294967296.0,1,-nbitq), 
to_sfixed(208835985.0/4294967296.0,1,-nbitq), 
to_sfixed(-304436941.0/4294967296.0,1,-nbitq), 
to_sfixed(297659029.0/4294967296.0,1,-nbitq), 
to_sfixed(-177829628.0/4294967296.0,1,-nbitq), 
to_sfixed(-41895726.0/4294967296.0,1,-nbitq), 
to_sfixed(-390721310.0/4294967296.0,1,-nbitq), 
to_sfixed(-112237242.0/4294967296.0,1,-nbitq), 
to_sfixed(-228474182.0/4294967296.0,1,-nbitq), 
to_sfixed(289865072.0/4294967296.0,1,-nbitq), 
to_sfixed(-80318722.0/4294967296.0,1,-nbitq), 
to_sfixed(258553087.0/4294967296.0,1,-nbitq), 
to_sfixed(-400139397.0/4294967296.0,1,-nbitq), 
to_sfixed(-346007992.0/4294967296.0,1,-nbitq), 
to_sfixed(-353465855.0/4294967296.0,1,-nbitq), 
to_sfixed(587630860.0/4294967296.0,1,-nbitq), 
to_sfixed(-432981441.0/4294967296.0,1,-nbitq), 
to_sfixed(-99182590.0/4294967296.0,1,-nbitq), 
to_sfixed(-431324962.0/4294967296.0,1,-nbitq), 
to_sfixed(-10037419.0/4294967296.0,1,-nbitq), 
to_sfixed(94905752.0/4294967296.0,1,-nbitq), 
to_sfixed(-271573358.0/4294967296.0,1,-nbitq), 
to_sfixed(137133586.0/4294967296.0,1,-nbitq), 
to_sfixed(-4714287.0/4294967296.0,1,-nbitq), 
to_sfixed(-321173728.0/4294967296.0,1,-nbitq), 
to_sfixed(453573376.0/4294967296.0,1,-nbitq), 
to_sfixed(-12852957.0/4294967296.0,1,-nbitq), 
to_sfixed(-9281339.0/4294967296.0,1,-nbitq), 
to_sfixed(-107889309.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-212950678.0/4294967296.0,1,-nbitq), 
to_sfixed(44694612.0/4294967296.0,1,-nbitq), 
to_sfixed(72741056.0/4294967296.0,1,-nbitq), 
to_sfixed(40257426.0/4294967296.0,1,-nbitq), 
to_sfixed(229884239.0/4294967296.0,1,-nbitq), 
to_sfixed(-117777314.0/4294967296.0,1,-nbitq), 
to_sfixed(-137206494.0/4294967296.0,1,-nbitq), 
to_sfixed(-530775909.0/4294967296.0,1,-nbitq), 
to_sfixed(-70123056.0/4294967296.0,1,-nbitq), 
to_sfixed(405365615.0/4294967296.0,1,-nbitq), 
to_sfixed(-120218707.0/4294967296.0,1,-nbitq), 
to_sfixed(458547333.0/4294967296.0,1,-nbitq), 
to_sfixed(-1218373565.0/4294967296.0,1,-nbitq), 
to_sfixed(-661822827.0/4294967296.0,1,-nbitq), 
to_sfixed(191696269.0/4294967296.0,1,-nbitq), 
to_sfixed(-146998500.0/4294967296.0,1,-nbitq), 
to_sfixed(-157639785.0/4294967296.0,1,-nbitq), 
to_sfixed(-346085911.0/4294967296.0,1,-nbitq), 
to_sfixed(624486372.0/4294967296.0,1,-nbitq), 
to_sfixed(337363788.0/4294967296.0,1,-nbitq), 
to_sfixed(-277648825.0/4294967296.0,1,-nbitq), 
to_sfixed(589285573.0/4294967296.0,1,-nbitq), 
to_sfixed(617287331.0/4294967296.0,1,-nbitq), 
to_sfixed(-789959414.0/4294967296.0,1,-nbitq), 
to_sfixed(422968002.0/4294967296.0,1,-nbitq), 
to_sfixed(-154985781.0/4294967296.0,1,-nbitq), 
to_sfixed(-180637410.0/4294967296.0,1,-nbitq), 
to_sfixed(44297660.0/4294967296.0,1,-nbitq), 
to_sfixed(104382099.0/4294967296.0,1,-nbitq), 
to_sfixed(-717059684.0/4294967296.0,1,-nbitq), 
to_sfixed(-251552106.0/4294967296.0,1,-nbitq), 
to_sfixed(203602255.0/4294967296.0,1,-nbitq), 
to_sfixed(112934703.0/4294967296.0,1,-nbitq), 
to_sfixed(446169081.0/4294967296.0,1,-nbitq), 
to_sfixed(-246318968.0/4294967296.0,1,-nbitq), 
to_sfixed(-678766651.0/4294967296.0,1,-nbitq), 
to_sfixed(363575890.0/4294967296.0,1,-nbitq), 
to_sfixed(-230648562.0/4294967296.0,1,-nbitq), 
to_sfixed(-321050668.0/4294967296.0,1,-nbitq), 
to_sfixed(69982722.0/4294967296.0,1,-nbitq), 
to_sfixed(-228908904.0/4294967296.0,1,-nbitq), 
to_sfixed(-164118138.0/4294967296.0,1,-nbitq), 
to_sfixed(187165719.0/4294967296.0,1,-nbitq), 
to_sfixed(-256005970.0/4294967296.0,1,-nbitq), 
to_sfixed(452723882.0/4294967296.0,1,-nbitq), 
to_sfixed(484332820.0/4294967296.0,1,-nbitq), 
to_sfixed(20507238.0/4294967296.0,1,-nbitq), 
to_sfixed(-203744547.0/4294967296.0,1,-nbitq), 
to_sfixed(269665369.0/4294967296.0,1,-nbitq), 
to_sfixed(677400997.0/4294967296.0,1,-nbitq), 
to_sfixed(71635943.0/4294967296.0,1,-nbitq), 
to_sfixed(-65956638.0/4294967296.0,1,-nbitq), 
to_sfixed(125787261.0/4294967296.0,1,-nbitq), 
to_sfixed(-488761342.0/4294967296.0,1,-nbitq), 
to_sfixed(-48587477.0/4294967296.0,1,-nbitq), 
to_sfixed(-176875570.0/4294967296.0,1,-nbitq), 
to_sfixed(-204001606.0/4294967296.0,1,-nbitq), 
to_sfixed(306499617.0/4294967296.0,1,-nbitq), 
to_sfixed(-319489251.0/4294967296.0,1,-nbitq), 
to_sfixed(-301801662.0/4294967296.0,1,-nbitq), 
to_sfixed(193788904.0/4294967296.0,1,-nbitq), 
to_sfixed(-307442871.0/4294967296.0,1,-nbitq), 
to_sfixed(440895983.0/4294967296.0,1,-nbitq), 
to_sfixed(-161599029.0/4294967296.0,1,-nbitq), 
to_sfixed(-231438907.0/4294967296.0,1,-nbitq), 
to_sfixed(228630471.0/4294967296.0,1,-nbitq), 
to_sfixed(221680905.0/4294967296.0,1,-nbitq), 
to_sfixed(-711896263.0/4294967296.0,1,-nbitq), 
to_sfixed(52142536.0/4294967296.0,1,-nbitq), 
to_sfixed(-116583104.0/4294967296.0,1,-nbitq), 
to_sfixed(-469762203.0/4294967296.0,1,-nbitq), 
to_sfixed(375403528.0/4294967296.0,1,-nbitq), 
to_sfixed(76831951.0/4294967296.0,1,-nbitq), 
to_sfixed(-132786296.0/4294967296.0,1,-nbitq), 
to_sfixed(256912277.0/4294967296.0,1,-nbitq), 
to_sfixed(-59992353.0/4294967296.0,1,-nbitq), 
to_sfixed(-66665855.0/4294967296.0,1,-nbitq), 
to_sfixed(-251488706.0/4294967296.0,1,-nbitq), 
to_sfixed(32435081.0/4294967296.0,1,-nbitq), 
to_sfixed(76725529.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-80266585.0/4294967296.0,1,-nbitq), 
to_sfixed(-191443300.0/4294967296.0,1,-nbitq), 
to_sfixed(379070236.0/4294967296.0,1,-nbitq), 
to_sfixed(-205110256.0/4294967296.0,1,-nbitq), 
to_sfixed(592607198.0/4294967296.0,1,-nbitq), 
to_sfixed(193893408.0/4294967296.0,1,-nbitq), 
to_sfixed(-183960317.0/4294967296.0,1,-nbitq), 
to_sfixed(-350158715.0/4294967296.0,1,-nbitq), 
to_sfixed(289957182.0/4294967296.0,1,-nbitq), 
to_sfixed(230286482.0/4294967296.0,1,-nbitq), 
to_sfixed(-273793879.0/4294967296.0,1,-nbitq), 
to_sfixed(12624568.0/4294967296.0,1,-nbitq), 
to_sfixed(-723727919.0/4294967296.0,1,-nbitq), 
to_sfixed(-130178566.0/4294967296.0,1,-nbitq), 
to_sfixed(-3895784.0/4294967296.0,1,-nbitq), 
to_sfixed(-71484162.0/4294967296.0,1,-nbitq), 
to_sfixed(131590303.0/4294967296.0,1,-nbitq), 
to_sfixed(-95501893.0/4294967296.0,1,-nbitq), 
to_sfixed(650746381.0/4294967296.0,1,-nbitq), 
to_sfixed(376175.0/4294967296.0,1,-nbitq), 
to_sfixed(-8133120.0/4294967296.0,1,-nbitq), 
to_sfixed(-36302869.0/4294967296.0,1,-nbitq), 
to_sfixed(119624486.0/4294967296.0,1,-nbitq), 
to_sfixed(-65737448.0/4294967296.0,1,-nbitq), 
to_sfixed(-319608375.0/4294967296.0,1,-nbitq), 
to_sfixed(-669268304.0/4294967296.0,1,-nbitq), 
to_sfixed(-309214072.0/4294967296.0,1,-nbitq), 
to_sfixed(-234691557.0/4294967296.0,1,-nbitq), 
to_sfixed(-293148485.0/4294967296.0,1,-nbitq), 
to_sfixed(-613667681.0/4294967296.0,1,-nbitq), 
to_sfixed(-13158418.0/4294967296.0,1,-nbitq), 
to_sfixed(-307214086.0/4294967296.0,1,-nbitq), 
to_sfixed(321193685.0/4294967296.0,1,-nbitq), 
to_sfixed(54233890.0/4294967296.0,1,-nbitq), 
to_sfixed(-314048278.0/4294967296.0,1,-nbitq), 
to_sfixed(-228406173.0/4294967296.0,1,-nbitq), 
to_sfixed(140937443.0/4294967296.0,1,-nbitq), 
to_sfixed(-739627877.0/4294967296.0,1,-nbitq), 
to_sfixed(-40940706.0/4294967296.0,1,-nbitq), 
to_sfixed(268613599.0/4294967296.0,1,-nbitq), 
to_sfixed(426358517.0/4294967296.0,1,-nbitq), 
to_sfixed(-175551113.0/4294967296.0,1,-nbitq), 
to_sfixed(-79225131.0/4294967296.0,1,-nbitq), 
to_sfixed(198430317.0/4294967296.0,1,-nbitq), 
to_sfixed(414514129.0/4294967296.0,1,-nbitq), 
to_sfixed(101985906.0/4294967296.0,1,-nbitq), 
to_sfixed(213652630.0/4294967296.0,1,-nbitq), 
to_sfixed(-66271337.0/4294967296.0,1,-nbitq), 
to_sfixed(405248277.0/4294967296.0,1,-nbitq), 
to_sfixed(566115977.0/4294967296.0,1,-nbitq), 
to_sfixed(104964823.0/4294967296.0,1,-nbitq), 
to_sfixed(-382814495.0/4294967296.0,1,-nbitq), 
to_sfixed(285645237.0/4294967296.0,1,-nbitq), 
to_sfixed(-361238776.0/4294967296.0,1,-nbitq), 
to_sfixed(139919887.0/4294967296.0,1,-nbitq), 
to_sfixed(-137888163.0/4294967296.0,1,-nbitq), 
to_sfixed(-141636773.0/4294967296.0,1,-nbitq), 
to_sfixed(-337835567.0/4294967296.0,1,-nbitq), 
to_sfixed(40344451.0/4294967296.0,1,-nbitq), 
to_sfixed(338150972.0/4294967296.0,1,-nbitq), 
to_sfixed(-181785360.0/4294967296.0,1,-nbitq), 
to_sfixed(-545341820.0/4294967296.0,1,-nbitq), 
to_sfixed(74150686.0/4294967296.0,1,-nbitq), 
to_sfixed(-149316599.0/4294967296.0,1,-nbitq), 
to_sfixed(61268079.0/4294967296.0,1,-nbitq), 
to_sfixed(-248533187.0/4294967296.0,1,-nbitq), 
to_sfixed(334184316.0/4294967296.0,1,-nbitq), 
to_sfixed(-176627501.0/4294967296.0,1,-nbitq), 
to_sfixed(236178630.0/4294967296.0,1,-nbitq), 
to_sfixed(197184777.0/4294967296.0,1,-nbitq), 
to_sfixed(-347083141.0/4294967296.0,1,-nbitq), 
to_sfixed(227640257.0/4294967296.0,1,-nbitq), 
to_sfixed(-115348411.0/4294967296.0,1,-nbitq), 
to_sfixed(129184796.0/4294967296.0,1,-nbitq), 
to_sfixed(-108986927.0/4294967296.0,1,-nbitq), 
to_sfixed(20135116.0/4294967296.0,1,-nbitq), 
to_sfixed(556551057.0/4294967296.0,1,-nbitq), 
to_sfixed(30210246.0/4294967296.0,1,-nbitq), 
to_sfixed(229821508.0/4294967296.0,1,-nbitq), 
to_sfixed(-191438867.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(49459511.0/4294967296.0,1,-nbitq), 
to_sfixed(-322199718.0/4294967296.0,1,-nbitq), 
to_sfixed(276374769.0/4294967296.0,1,-nbitq), 
to_sfixed(-815332352.0/4294967296.0,1,-nbitq), 
to_sfixed(329482846.0/4294967296.0,1,-nbitq), 
to_sfixed(56320266.0/4294967296.0,1,-nbitq), 
to_sfixed(316216158.0/4294967296.0,1,-nbitq), 
to_sfixed(-100840026.0/4294967296.0,1,-nbitq), 
to_sfixed(553168472.0/4294967296.0,1,-nbitq), 
to_sfixed(442173665.0/4294967296.0,1,-nbitq), 
to_sfixed(-62283472.0/4294967296.0,1,-nbitq), 
to_sfixed(356198612.0/4294967296.0,1,-nbitq), 
to_sfixed(-176419872.0/4294967296.0,1,-nbitq), 
to_sfixed(-284054942.0/4294967296.0,1,-nbitq), 
to_sfixed(-41851589.0/4294967296.0,1,-nbitq), 
to_sfixed(-277955117.0/4294967296.0,1,-nbitq), 
to_sfixed(362861471.0/4294967296.0,1,-nbitq), 
to_sfixed(-179637549.0/4294967296.0,1,-nbitq), 
to_sfixed(356859254.0/4294967296.0,1,-nbitq), 
to_sfixed(-479716109.0/4294967296.0,1,-nbitq), 
to_sfixed(-151823680.0/4294967296.0,1,-nbitq), 
to_sfixed(-12518758.0/4294967296.0,1,-nbitq), 
to_sfixed(125256518.0/4294967296.0,1,-nbitq), 
to_sfixed(-349618410.0/4294967296.0,1,-nbitq), 
to_sfixed(-1403333.0/4294967296.0,1,-nbitq), 
to_sfixed(-551732166.0/4294967296.0,1,-nbitq), 
to_sfixed(-139746931.0/4294967296.0,1,-nbitq), 
to_sfixed(-452333873.0/4294967296.0,1,-nbitq), 
to_sfixed(-488123633.0/4294967296.0,1,-nbitq), 
to_sfixed(-59605675.0/4294967296.0,1,-nbitq), 
to_sfixed(-204392988.0/4294967296.0,1,-nbitq), 
to_sfixed(173937811.0/4294967296.0,1,-nbitq), 
to_sfixed(385311754.0/4294967296.0,1,-nbitq), 
to_sfixed(-102561109.0/4294967296.0,1,-nbitq), 
to_sfixed(-91525787.0/4294967296.0,1,-nbitq), 
to_sfixed(-9020450.0/4294967296.0,1,-nbitq), 
to_sfixed(-97863213.0/4294967296.0,1,-nbitq), 
to_sfixed(-291185180.0/4294967296.0,1,-nbitq), 
to_sfixed(-3557066.0/4294967296.0,1,-nbitq), 
to_sfixed(397409499.0/4294967296.0,1,-nbitq), 
to_sfixed(-21109430.0/4294967296.0,1,-nbitq), 
to_sfixed(-45206901.0/4294967296.0,1,-nbitq), 
to_sfixed(-350374954.0/4294967296.0,1,-nbitq), 
to_sfixed(258735196.0/4294967296.0,1,-nbitq), 
to_sfixed(-178112739.0/4294967296.0,1,-nbitq), 
to_sfixed(65781480.0/4294967296.0,1,-nbitq), 
to_sfixed(-47854621.0/4294967296.0,1,-nbitq), 
to_sfixed(-420853253.0/4294967296.0,1,-nbitq), 
to_sfixed(-256789913.0/4294967296.0,1,-nbitq), 
to_sfixed(396683924.0/4294967296.0,1,-nbitq), 
to_sfixed(-41034295.0/4294967296.0,1,-nbitq), 
to_sfixed(-220485.0/4294967296.0,1,-nbitq), 
to_sfixed(-471700948.0/4294967296.0,1,-nbitq), 
to_sfixed(-680889924.0/4294967296.0,1,-nbitq), 
to_sfixed(-190170753.0/4294967296.0,1,-nbitq), 
to_sfixed(-334574341.0/4294967296.0,1,-nbitq), 
to_sfixed(-477849057.0/4294967296.0,1,-nbitq), 
to_sfixed(-268343044.0/4294967296.0,1,-nbitq), 
to_sfixed(-54280559.0/4294967296.0,1,-nbitq), 
to_sfixed(14703033.0/4294967296.0,1,-nbitq), 
to_sfixed(-255007619.0/4294967296.0,1,-nbitq), 
to_sfixed(138607310.0/4294967296.0,1,-nbitq), 
to_sfixed(241885609.0/4294967296.0,1,-nbitq), 
to_sfixed(-569695887.0/4294967296.0,1,-nbitq), 
to_sfixed(62654730.0/4294967296.0,1,-nbitq), 
to_sfixed(-256196727.0/4294967296.0,1,-nbitq), 
to_sfixed(273537120.0/4294967296.0,1,-nbitq), 
to_sfixed(-183212145.0/4294967296.0,1,-nbitq), 
to_sfixed(-13287595.0/4294967296.0,1,-nbitq), 
to_sfixed(117341448.0/4294967296.0,1,-nbitq), 
to_sfixed(244164066.0/4294967296.0,1,-nbitq), 
to_sfixed(16023253.0/4294967296.0,1,-nbitq), 
to_sfixed(-248505087.0/4294967296.0,1,-nbitq), 
to_sfixed(33174872.0/4294967296.0,1,-nbitq), 
to_sfixed(257971701.0/4294967296.0,1,-nbitq), 
to_sfixed(-419713127.0/4294967296.0,1,-nbitq), 
to_sfixed(307592034.0/4294967296.0,1,-nbitq), 
to_sfixed(136332165.0/4294967296.0,1,-nbitq), 
to_sfixed(503871485.0/4294967296.0,1,-nbitq), 
to_sfixed(-175974800.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-281125316.0/4294967296.0,1,-nbitq), 
to_sfixed(-129713489.0/4294967296.0,1,-nbitq), 
to_sfixed(635512399.0/4294967296.0,1,-nbitq), 
to_sfixed(-73425319.0/4294967296.0,1,-nbitq), 
to_sfixed(100927002.0/4294967296.0,1,-nbitq), 
to_sfixed(-910668786.0/4294967296.0,1,-nbitq), 
to_sfixed(302473257.0/4294967296.0,1,-nbitq), 
to_sfixed(139243788.0/4294967296.0,1,-nbitq), 
to_sfixed(650652490.0/4294967296.0,1,-nbitq), 
to_sfixed(-4096592.0/4294967296.0,1,-nbitq), 
to_sfixed(117543219.0/4294967296.0,1,-nbitq), 
to_sfixed(87595081.0/4294967296.0,1,-nbitq), 
to_sfixed(-456113614.0/4294967296.0,1,-nbitq), 
to_sfixed(222758662.0/4294967296.0,1,-nbitq), 
to_sfixed(75150942.0/4294967296.0,1,-nbitq), 
to_sfixed(-592876953.0/4294967296.0,1,-nbitq), 
to_sfixed(-139760223.0/4294967296.0,1,-nbitq), 
to_sfixed(229866963.0/4294967296.0,1,-nbitq), 
to_sfixed(594581611.0/4294967296.0,1,-nbitq), 
to_sfixed(-398613483.0/4294967296.0,1,-nbitq), 
to_sfixed(61013765.0/4294967296.0,1,-nbitq), 
to_sfixed(112372870.0/4294967296.0,1,-nbitq), 
to_sfixed(538094953.0/4294967296.0,1,-nbitq), 
to_sfixed(-435378501.0/4294967296.0,1,-nbitq), 
to_sfixed(-216542985.0/4294967296.0,1,-nbitq), 
to_sfixed(-759384487.0/4294967296.0,1,-nbitq), 
to_sfixed(-63098667.0/4294967296.0,1,-nbitq), 
to_sfixed(-250752008.0/4294967296.0,1,-nbitq), 
to_sfixed(-167476570.0/4294967296.0,1,-nbitq), 
to_sfixed(-86363697.0/4294967296.0,1,-nbitq), 
to_sfixed(-565584043.0/4294967296.0,1,-nbitq), 
to_sfixed(85946001.0/4294967296.0,1,-nbitq), 
to_sfixed(-98182183.0/4294967296.0,1,-nbitq), 
to_sfixed(-186217462.0/4294967296.0,1,-nbitq), 
to_sfixed(60549428.0/4294967296.0,1,-nbitq), 
to_sfixed(-7273906.0/4294967296.0,1,-nbitq), 
to_sfixed(404480923.0/4294967296.0,1,-nbitq), 
to_sfixed(-50388028.0/4294967296.0,1,-nbitq), 
to_sfixed(119391049.0/4294967296.0,1,-nbitq), 
to_sfixed(29884137.0/4294967296.0,1,-nbitq), 
to_sfixed(12573851.0/4294967296.0,1,-nbitq), 
to_sfixed(116672436.0/4294967296.0,1,-nbitq), 
to_sfixed(-284548799.0/4294967296.0,1,-nbitq), 
to_sfixed(-178577620.0/4294967296.0,1,-nbitq), 
to_sfixed(-318501963.0/4294967296.0,1,-nbitq), 
to_sfixed(608909917.0/4294967296.0,1,-nbitq), 
to_sfixed(73636261.0/4294967296.0,1,-nbitq), 
to_sfixed(-187324353.0/4294967296.0,1,-nbitq), 
to_sfixed(-262301771.0/4294967296.0,1,-nbitq), 
to_sfixed(296519031.0/4294967296.0,1,-nbitq), 
to_sfixed(365375638.0/4294967296.0,1,-nbitq), 
to_sfixed(92495873.0/4294967296.0,1,-nbitq), 
to_sfixed(-376079683.0/4294967296.0,1,-nbitq), 
to_sfixed(-616919659.0/4294967296.0,1,-nbitq), 
to_sfixed(-51183612.0/4294967296.0,1,-nbitq), 
to_sfixed(-185025112.0/4294967296.0,1,-nbitq), 
to_sfixed(-281249805.0/4294967296.0,1,-nbitq), 
to_sfixed(192569250.0/4294967296.0,1,-nbitq), 
to_sfixed(-187059611.0/4294967296.0,1,-nbitq), 
to_sfixed(-93931910.0/4294967296.0,1,-nbitq), 
to_sfixed(-309382467.0/4294967296.0,1,-nbitq), 
to_sfixed(436646613.0/4294967296.0,1,-nbitq), 
to_sfixed(-145277735.0/4294967296.0,1,-nbitq), 
to_sfixed(-767656656.0/4294967296.0,1,-nbitq), 
to_sfixed(-541601.0/4294967296.0,1,-nbitq), 
to_sfixed(130631641.0/4294967296.0,1,-nbitq), 
to_sfixed(160001815.0/4294967296.0,1,-nbitq), 
to_sfixed(-779735913.0/4294967296.0,1,-nbitq), 
to_sfixed(362527509.0/4294967296.0,1,-nbitq), 
to_sfixed(27510326.0/4294967296.0,1,-nbitq), 
to_sfixed(-261214846.0/4294967296.0,1,-nbitq), 
to_sfixed(-144353498.0/4294967296.0,1,-nbitq), 
to_sfixed(128525302.0/4294967296.0,1,-nbitq), 
to_sfixed(39586790.0/4294967296.0,1,-nbitq), 
to_sfixed(495265772.0/4294967296.0,1,-nbitq), 
to_sfixed(293895940.0/4294967296.0,1,-nbitq), 
to_sfixed(150360472.0/4294967296.0,1,-nbitq), 
to_sfixed(89886571.0/4294967296.0,1,-nbitq), 
to_sfixed(698707416.0/4294967296.0,1,-nbitq), 
to_sfixed(178638276.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-250338346.0/4294967296.0,1,-nbitq), 
to_sfixed(-72694305.0/4294967296.0,1,-nbitq), 
to_sfixed(502596977.0/4294967296.0,1,-nbitq), 
to_sfixed(-489266659.0/4294967296.0,1,-nbitq), 
to_sfixed(267983155.0/4294967296.0,1,-nbitq), 
to_sfixed(-803182771.0/4294967296.0,1,-nbitq), 
to_sfixed(-7587800.0/4294967296.0,1,-nbitq), 
to_sfixed(-412838176.0/4294967296.0,1,-nbitq), 
to_sfixed(404376746.0/4294967296.0,1,-nbitq), 
to_sfixed(148997103.0/4294967296.0,1,-nbitq), 
to_sfixed(-356279849.0/4294967296.0,1,-nbitq), 
to_sfixed(229380711.0/4294967296.0,1,-nbitq), 
to_sfixed(-852816660.0/4294967296.0,1,-nbitq), 
to_sfixed(-2560979.0/4294967296.0,1,-nbitq), 
to_sfixed(311677501.0/4294967296.0,1,-nbitq), 
to_sfixed(-307719449.0/4294967296.0,1,-nbitq), 
to_sfixed(68045737.0/4294967296.0,1,-nbitq), 
to_sfixed(-395589630.0/4294967296.0,1,-nbitq), 
to_sfixed(-68295460.0/4294967296.0,1,-nbitq), 
to_sfixed(-11044326.0/4294967296.0,1,-nbitq), 
to_sfixed(-148905321.0/4294967296.0,1,-nbitq), 
to_sfixed(330693407.0/4294967296.0,1,-nbitq), 
to_sfixed(10011015.0/4294967296.0,1,-nbitq), 
to_sfixed(37323426.0/4294967296.0,1,-nbitq), 
to_sfixed(-214306004.0/4294967296.0,1,-nbitq), 
to_sfixed(-415309582.0/4294967296.0,1,-nbitq), 
to_sfixed(346118494.0/4294967296.0,1,-nbitq), 
to_sfixed(-390901885.0/4294967296.0,1,-nbitq), 
to_sfixed(64627637.0/4294967296.0,1,-nbitq), 
to_sfixed(-451898957.0/4294967296.0,1,-nbitq), 
to_sfixed(-617740925.0/4294967296.0,1,-nbitq), 
to_sfixed(-16099040.0/4294967296.0,1,-nbitq), 
to_sfixed(254932835.0/4294967296.0,1,-nbitq), 
to_sfixed(-100816134.0/4294967296.0,1,-nbitq), 
to_sfixed(247712622.0/4294967296.0,1,-nbitq), 
to_sfixed(-286580442.0/4294967296.0,1,-nbitq), 
to_sfixed(38697798.0/4294967296.0,1,-nbitq), 
to_sfixed(62720958.0/4294967296.0,1,-nbitq), 
to_sfixed(51602351.0/4294967296.0,1,-nbitq), 
to_sfixed(-140001348.0/4294967296.0,1,-nbitq), 
to_sfixed(268457077.0/4294967296.0,1,-nbitq), 
to_sfixed(408900908.0/4294967296.0,1,-nbitq), 
to_sfixed(342458606.0/4294967296.0,1,-nbitq), 
to_sfixed(472245952.0/4294967296.0,1,-nbitq), 
to_sfixed(-161085351.0/4294967296.0,1,-nbitq), 
to_sfixed(263710412.0/4294967296.0,1,-nbitq), 
to_sfixed(141693069.0/4294967296.0,1,-nbitq), 
to_sfixed(-597107932.0/4294967296.0,1,-nbitq), 
to_sfixed(-263716331.0/4294967296.0,1,-nbitq), 
to_sfixed(152214035.0/4294967296.0,1,-nbitq), 
to_sfixed(-78868756.0/4294967296.0,1,-nbitq), 
to_sfixed(236690633.0/4294967296.0,1,-nbitq), 
to_sfixed(-307277720.0/4294967296.0,1,-nbitq), 
to_sfixed(-23081551.0/4294967296.0,1,-nbitq), 
to_sfixed(179058978.0/4294967296.0,1,-nbitq), 
to_sfixed(-96312212.0/4294967296.0,1,-nbitq), 
to_sfixed(-776332733.0/4294967296.0,1,-nbitq), 
to_sfixed(-162871839.0/4294967296.0,1,-nbitq), 
to_sfixed(-345772582.0/4294967296.0,1,-nbitq), 
to_sfixed(253780380.0/4294967296.0,1,-nbitq), 
to_sfixed(40909362.0/4294967296.0,1,-nbitq), 
to_sfixed(-88830518.0/4294967296.0,1,-nbitq), 
to_sfixed(2203197.0/4294967296.0,1,-nbitq), 
to_sfixed(-303310391.0/4294967296.0,1,-nbitq), 
to_sfixed(-23958819.0/4294967296.0,1,-nbitq), 
to_sfixed(-413651179.0/4294967296.0,1,-nbitq), 
to_sfixed(303536279.0/4294967296.0,1,-nbitq), 
to_sfixed(-642932128.0/4294967296.0,1,-nbitq), 
to_sfixed(418243819.0/4294967296.0,1,-nbitq), 
to_sfixed(353603272.0/4294967296.0,1,-nbitq), 
to_sfixed(-124810405.0/4294967296.0,1,-nbitq), 
to_sfixed(-141765084.0/4294967296.0,1,-nbitq), 
to_sfixed(222617338.0/4294967296.0,1,-nbitq), 
to_sfixed(75782840.0/4294967296.0,1,-nbitq), 
to_sfixed(68340257.0/4294967296.0,1,-nbitq), 
to_sfixed(223100868.0/4294967296.0,1,-nbitq), 
to_sfixed(-37344109.0/4294967296.0,1,-nbitq), 
to_sfixed(335427971.0/4294967296.0,1,-nbitq), 
to_sfixed(181154168.0/4294967296.0,1,-nbitq), 
to_sfixed(-112326240.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-190474654.0/4294967296.0,1,-nbitq), 
to_sfixed(-146994334.0/4294967296.0,1,-nbitq), 
to_sfixed(316426388.0/4294967296.0,1,-nbitq), 
to_sfixed(-275293783.0/4294967296.0,1,-nbitq), 
to_sfixed(-408546739.0/4294967296.0,1,-nbitq), 
to_sfixed(-52085164.0/4294967296.0,1,-nbitq), 
to_sfixed(275274473.0/4294967296.0,1,-nbitq), 
to_sfixed(-324784037.0/4294967296.0,1,-nbitq), 
to_sfixed(180438775.0/4294967296.0,1,-nbitq), 
to_sfixed(-174727464.0/4294967296.0,1,-nbitq), 
to_sfixed(-42635065.0/4294967296.0,1,-nbitq), 
to_sfixed(-278010921.0/4294967296.0,1,-nbitq), 
to_sfixed(-448259243.0/4294967296.0,1,-nbitq), 
to_sfixed(140614526.0/4294967296.0,1,-nbitq), 
to_sfixed(38815400.0/4294967296.0,1,-nbitq), 
to_sfixed(-397781542.0/4294967296.0,1,-nbitq), 
to_sfixed(-242607196.0/4294967296.0,1,-nbitq), 
to_sfixed(-233088225.0/4294967296.0,1,-nbitq), 
to_sfixed(172569833.0/4294967296.0,1,-nbitq), 
to_sfixed(149908521.0/4294967296.0,1,-nbitq), 
to_sfixed(19809987.0/4294967296.0,1,-nbitq), 
to_sfixed(53398072.0/4294967296.0,1,-nbitq), 
to_sfixed(266309944.0/4294967296.0,1,-nbitq), 
to_sfixed(-135681149.0/4294967296.0,1,-nbitq), 
to_sfixed(-84224465.0/4294967296.0,1,-nbitq), 
to_sfixed(-561187180.0/4294967296.0,1,-nbitq), 
to_sfixed(192347263.0/4294967296.0,1,-nbitq), 
to_sfixed(-57839815.0/4294967296.0,1,-nbitq), 
to_sfixed(-162019613.0/4294967296.0,1,-nbitq), 
to_sfixed(-40596092.0/4294967296.0,1,-nbitq), 
to_sfixed(-836173714.0/4294967296.0,1,-nbitq), 
to_sfixed(-188603845.0/4294967296.0,1,-nbitq), 
to_sfixed(-103927002.0/4294967296.0,1,-nbitq), 
to_sfixed(19382528.0/4294967296.0,1,-nbitq), 
to_sfixed(327274831.0/4294967296.0,1,-nbitq), 
to_sfixed(-34955678.0/4294967296.0,1,-nbitq), 
to_sfixed(-110194081.0/4294967296.0,1,-nbitq), 
to_sfixed(521308212.0/4294967296.0,1,-nbitq), 
to_sfixed(-279725186.0/4294967296.0,1,-nbitq), 
to_sfixed(405629313.0/4294967296.0,1,-nbitq), 
to_sfixed(48443368.0/4294967296.0,1,-nbitq), 
to_sfixed(88127901.0/4294967296.0,1,-nbitq), 
to_sfixed(-49033781.0/4294967296.0,1,-nbitq), 
to_sfixed(681306384.0/4294967296.0,1,-nbitq), 
to_sfixed(-521396059.0/4294967296.0,1,-nbitq), 
to_sfixed(653489517.0/4294967296.0,1,-nbitq), 
to_sfixed(160414297.0/4294967296.0,1,-nbitq), 
to_sfixed(-979683235.0/4294967296.0,1,-nbitq), 
to_sfixed(302603105.0/4294967296.0,1,-nbitq), 
to_sfixed(65405147.0/4294967296.0,1,-nbitq), 
to_sfixed(-110090856.0/4294967296.0,1,-nbitq), 
to_sfixed(-442633036.0/4294967296.0,1,-nbitq), 
to_sfixed(-220735565.0/4294967296.0,1,-nbitq), 
to_sfixed(47954959.0/4294967296.0,1,-nbitq), 
to_sfixed(-184819572.0/4294967296.0,1,-nbitq), 
to_sfixed(-443158662.0/4294967296.0,1,-nbitq), 
to_sfixed(-482158021.0/4294967296.0,1,-nbitq), 
to_sfixed(350410871.0/4294967296.0,1,-nbitq), 
to_sfixed(159593093.0/4294967296.0,1,-nbitq), 
to_sfixed(-158830617.0/4294967296.0,1,-nbitq), 
to_sfixed(273399992.0/4294967296.0,1,-nbitq), 
to_sfixed(-13637652.0/4294967296.0,1,-nbitq), 
to_sfixed(204361812.0/4294967296.0,1,-nbitq), 
to_sfixed(154665738.0/4294967296.0,1,-nbitq), 
to_sfixed(420284652.0/4294967296.0,1,-nbitq), 
to_sfixed(226118596.0/4294967296.0,1,-nbitq), 
to_sfixed(-209082179.0/4294967296.0,1,-nbitq), 
to_sfixed(-384539423.0/4294967296.0,1,-nbitq), 
to_sfixed(-8001884.0/4294967296.0,1,-nbitq), 
to_sfixed(-260366751.0/4294967296.0,1,-nbitq), 
to_sfixed(127685149.0/4294967296.0,1,-nbitq), 
to_sfixed(-101608467.0/4294967296.0,1,-nbitq), 
to_sfixed(-416051807.0/4294967296.0,1,-nbitq), 
to_sfixed(276796152.0/4294967296.0,1,-nbitq), 
to_sfixed(503333177.0/4294967296.0,1,-nbitq), 
to_sfixed(56759554.0/4294967296.0,1,-nbitq), 
to_sfixed(201354379.0/4294967296.0,1,-nbitq), 
to_sfixed(-91653629.0/4294967296.0,1,-nbitq), 
to_sfixed(540846965.0/4294967296.0,1,-nbitq), 
to_sfixed(-339525172.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-286487704.0/4294967296.0,1,-nbitq), 
to_sfixed(-545056764.0/4294967296.0,1,-nbitq), 
to_sfixed(276523612.0/4294967296.0,1,-nbitq), 
to_sfixed(-346245486.0/4294967296.0,1,-nbitq), 
to_sfixed(-405616779.0/4294967296.0,1,-nbitq), 
to_sfixed(371183386.0/4294967296.0,1,-nbitq), 
to_sfixed(-129138231.0/4294967296.0,1,-nbitq), 
to_sfixed(-214560905.0/4294967296.0,1,-nbitq), 
to_sfixed(126897845.0/4294967296.0,1,-nbitq), 
to_sfixed(-29530439.0/4294967296.0,1,-nbitq), 
to_sfixed(47783486.0/4294967296.0,1,-nbitq), 
to_sfixed(44585788.0/4294967296.0,1,-nbitq), 
to_sfixed(71179346.0/4294967296.0,1,-nbitq), 
to_sfixed(-28853036.0/4294967296.0,1,-nbitq), 
to_sfixed(-360657931.0/4294967296.0,1,-nbitq), 
to_sfixed(-424348568.0/4294967296.0,1,-nbitq), 
to_sfixed(37536298.0/4294967296.0,1,-nbitq), 
to_sfixed(237532594.0/4294967296.0,1,-nbitq), 
to_sfixed(424222037.0/4294967296.0,1,-nbitq), 
to_sfixed(236174357.0/4294967296.0,1,-nbitq), 
to_sfixed(-79394396.0/4294967296.0,1,-nbitq), 
to_sfixed(72084893.0/4294967296.0,1,-nbitq), 
to_sfixed(6895181.0/4294967296.0,1,-nbitq), 
to_sfixed(-77386343.0/4294967296.0,1,-nbitq), 
to_sfixed(393883819.0/4294967296.0,1,-nbitq), 
to_sfixed(-467912610.0/4294967296.0,1,-nbitq), 
to_sfixed(-195454717.0/4294967296.0,1,-nbitq), 
to_sfixed(-335461760.0/4294967296.0,1,-nbitq), 
to_sfixed(-213413950.0/4294967296.0,1,-nbitq), 
to_sfixed(-39110020.0/4294967296.0,1,-nbitq), 
to_sfixed(-520403234.0/4294967296.0,1,-nbitq), 
to_sfixed(61734609.0/4294967296.0,1,-nbitq), 
to_sfixed(371808938.0/4294967296.0,1,-nbitq), 
to_sfixed(22201710.0/4294967296.0,1,-nbitq), 
to_sfixed(380146099.0/4294967296.0,1,-nbitq), 
to_sfixed(176818621.0/4294967296.0,1,-nbitq), 
to_sfixed(-62437457.0/4294967296.0,1,-nbitq), 
to_sfixed(-113688329.0/4294967296.0,1,-nbitq), 
to_sfixed(-165770906.0/4294967296.0,1,-nbitq), 
to_sfixed(-33873735.0/4294967296.0,1,-nbitq), 
to_sfixed(-160750194.0/4294967296.0,1,-nbitq), 
to_sfixed(146213959.0/4294967296.0,1,-nbitq), 
to_sfixed(205772809.0/4294967296.0,1,-nbitq), 
to_sfixed(-92269183.0/4294967296.0,1,-nbitq), 
to_sfixed(-286918716.0/4294967296.0,1,-nbitq), 
to_sfixed(353004948.0/4294967296.0,1,-nbitq), 
to_sfixed(-336395487.0/4294967296.0,1,-nbitq), 
to_sfixed(-541206283.0/4294967296.0,1,-nbitq), 
to_sfixed(-61939095.0/4294967296.0,1,-nbitq), 
to_sfixed(359518049.0/4294967296.0,1,-nbitq), 
to_sfixed(-299840164.0/4294967296.0,1,-nbitq), 
to_sfixed(-629552030.0/4294967296.0,1,-nbitq), 
to_sfixed(324512240.0/4294967296.0,1,-nbitq), 
to_sfixed(-254256571.0/4294967296.0,1,-nbitq), 
to_sfixed(-149409455.0/4294967296.0,1,-nbitq), 
to_sfixed(-94368742.0/4294967296.0,1,-nbitq), 
to_sfixed(-501345366.0/4294967296.0,1,-nbitq), 
to_sfixed(361664120.0/4294967296.0,1,-nbitq), 
to_sfixed(-60084913.0/4294967296.0,1,-nbitq), 
to_sfixed(66925292.0/4294967296.0,1,-nbitq), 
to_sfixed(-248447508.0/4294967296.0,1,-nbitq), 
to_sfixed(-255373524.0/4294967296.0,1,-nbitq), 
to_sfixed(-224651357.0/4294967296.0,1,-nbitq), 
to_sfixed(-321338324.0/4294967296.0,1,-nbitq), 
to_sfixed(-95465067.0/4294967296.0,1,-nbitq), 
to_sfixed(-161914720.0/4294967296.0,1,-nbitq), 
to_sfixed(482628133.0/4294967296.0,1,-nbitq), 
to_sfixed(-74705436.0/4294967296.0,1,-nbitq), 
to_sfixed(-182029887.0/4294967296.0,1,-nbitq), 
to_sfixed(-443087856.0/4294967296.0,1,-nbitq), 
to_sfixed(-214535401.0/4294967296.0,1,-nbitq), 
to_sfixed(47970529.0/4294967296.0,1,-nbitq), 
to_sfixed(-92678900.0/4294967296.0,1,-nbitq), 
to_sfixed(413459364.0/4294967296.0,1,-nbitq), 
to_sfixed(104609358.0/4294967296.0,1,-nbitq), 
to_sfixed(-14390614.0/4294967296.0,1,-nbitq), 
to_sfixed(-375895987.0/4294967296.0,1,-nbitq), 
to_sfixed(-400222161.0/4294967296.0,1,-nbitq), 
to_sfixed(683277440.0/4294967296.0,1,-nbitq), 
to_sfixed(140684712.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(213753718.0/4294967296.0,1,-nbitq), 
to_sfixed(-185601077.0/4294967296.0,1,-nbitq), 
to_sfixed(99518368.0/4294967296.0,1,-nbitq), 
to_sfixed(-146306514.0/4294967296.0,1,-nbitq), 
to_sfixed(363309912.0/4294967296.0,1,-nbitq), 
to_sfixed(279676208.0/4294967296.0,1,-nbitq), 
to_sfixed(-163711745.0/4294967296.0,1,-nbitq), 
to_sfixed(-77693468.0/4294967296.0,1,-nbitq), 
to_sfixed(217166211.0/4294967296.0,1,-nbitq), 
to_sfixed(-255687266.0/4294967296.0,1,-nbitq), 
to_sfixed(-194677605.0/4294967296.0,1,-nbitq), 
to_sfixed(319326705.0/4294967296.0,1,-nbitq), 
to_sfixed(39180164.0/4294967296.0,1,-nbitq), 
to_sfixed(-58914466.0/4294967296.0,1,-nbitq), 
to_sfixed(384492756.0/4294967296.0,1,-nbitq), 
to_sfixed(-17626195.0/4294967296.0,1,-nbitq), 
to_sfixed(-60029023.0/4294967296.0,1,-nbitq), 
to_sfixed(-127061183.0/4294967296.0,1,-nbitq), 
to_sfixed(-81388883.0/4294967296.0,1,-nbitq), 
to_sfixed(98934679.0/4294967296.0,1,-nbitq), 
to_sfixed(-400240036.0/4294967296.0,1,-nbitq), 
to_sfixed(20365511.0/4294967296.0,1,-nbitq), 
to_sfixed(431696675.0/4294967296.0,1,-nbitq), 
to_sfixed(-162296692.0/4294967296.0,1,-nbitq), 
to_sfixed(272854972.0/4294967296.0,1,-nbitq), 
to_sfixed(-250005836.0/4294967296.0,1,-nbitq), 
to_sfixed(321669747.0/4294967296.0,1,-nbitq), 
to_sfixed(-311361855.0/4294967296.0,1,-nbitq), 
to_sfixed(-77958265.0/4294967296.0,1,-nbitq), 
to_sfixed(7551963.0/4294967296.0,1,-nbitq), 
to_sfixed(-398316564.0/4294967296.0,1,-nbitq), 
to_sfixed(-51457307.0/4294967296.0,1,-nbitq), 
to_sfixed(192663177.0/4294967296.0,1,-nbitq), 
to_sfixed(480554179.0/4294967296.0,1,-nbitq), 
to_sfixed(156998789.0/4294967296.0,1,-nbitq), 
to_sfixed(205288345.0/4294967296.0,1,-nbitq), 
to_sfixed(435842964.0/4294967296.0,1,-nbitq), 
to_sfixed(-441493869.0/4294967296.0,1,-nbitq), 
to_sfixed(-164500455.0/4294967296.0,1,-nbitq), 
to_sfixed(-99392389.0/4294967296.0,1,-nbitq), 
to_sfixed(-173136322.0/4294967296.0,1,-nbitq), 
to_sfixed(-191690196.0/4294967296.0,1,-nbitq), 
to_sfixed(340374818.0/4294967296.0,1,-nbitq), 
to_sfixed(-29688082.0/4294967296.0,1,-nbitq), 
to_sfixed(239801870.0/4294967296.0,1,-nbitq), 
to_sfixed(361166518.0/4294967296.0,1,-nbitq), 
to_sfixed(-249891617.0/4294967296.0,1,-nbitq), 
to_sfixed(-296679868.0/4294967296.0,1,-nbitq), 
to_sfixed(115316015.0/4294967296.0,1,-nbitq), 
to_sfixed(359805755.0/4294967296.0,1,-nbitq), 
to_sfixed(-29188044.0/4294967296.0,1,-nbitq), 
to_sfixed(4919934.0/4294967296.0,1,-nbitq), 
to_sfixed(-460464528.0/4294967296.0,1,-nbitq), 
to_sfixed(218125220.0/4294967296.0,1,-nbitq), 
to_sfixed(-405798668.0/4294967296.0,1,-nbitq), 
to_sfixed(-489501736.0/4294967296.0,1,-nbitq), 
to_sfixed(-282273362.0/4294967296.0,1,-nbitq), 
to_sfixed(-288440489.0/4294967296.0,1,-nbitq), 
to_sfixed(245988958.0/4294967296.0,1,-nbitq), 
to_sfixed(-281003285.0/4294967296.0,1,-nbitq), 
to_sfixed(-252983094.0/4294967296.0,1,-nbitq), 
to_sfixed(240437196.0/4294967296.0,1,-nbitq), 
to_sfixed(285585096.0/4294967296.0,1,-nbitq), 
to_sfixed(-380726586.0/4294967296.0,1,-nbitq), 
to_sfixed(-330027682.0/4294967296.0,1,-nbitq), 
to_sfixed(234791859.0/4294967296.0,1,-nbitq), 
to_sfixed(131443495.0/4294967296.0,1,-nbitq), 
to_sfixed(-290491400.0/4294967296.0,1,-nbitq), 
to_sfixed(-189283331.0/4294967296.0,1,-nbitq), 
to_sfixed(-144685337.0/4294967296.0,1,-nbitq), 
to_sfixed(-298511759.0/4294967296.0,1,-nbitq), 
to_sfixed(331513889.0/4294967296.0,1,-nbitq), 
to_sfixed(-97580897.0/4294967296.0,1,-nbitq), 
to_sfixed(160891902.0/4294967296.0,1,-nbitq), 
to_sfixed(-39729952.0/4294967296.0,1,-nbitq), 
to_sfixed(-234124915.0/4294967296.0,1,-nbitq), 
to_sfixed(-57284503.0/4294967296.0,1,-nbitq), 
to_sfixed(195275912.0/4294967296.0,1,-nbitq), 
to_sfixed(123357721.0/4294967296.0,1,-nbitq), 
to_sfixed(-160984236.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-55572482.0/4294967296.0,1,-nbitq), 
to_sfixed(-396695640.0/4294967296.0,1,-nbitq), 
to_sfixed(289426740.0/4294967296.0,1,-nbitq), 
to_sfixed(-8613763.0/4294967296.0,1,-nbitq), 
to_sfixed(-44436740.0/4294967296.0,1,-nbitq), 
to_sfixed(340314251.0/4294967296.0,1,-nbitq), 
to_sfixed(-99627257.0/4294967296.0,1,-nbitq), 
to_sfixed(-42907078.0/4294967296.0,1,-nbitq), 
to_sfixed(155827519.0/4294967296.0,1,-nbitq), 
to_sfixed(421995422.0/4294967296.0,1,-nbitq), 
to_sfixed(130103263.0/4294967296.0,1,-nbitq), 
to_sfixed(-183623259.0/4294967296.0,1,-nbitq), 
to_sfixed(249649382.0/4294967296.0,1,-nbitq), 
to_sfixed(-151888529.0/4294967296.0,1,-nbitq), 
to_sfixed(142145291.0/4294967296.0,1,-nbitq), 
to_sfixed(-370338878.0/4294967296.0,1,-nbitq), 
to_sfixed(-348913328.0/4294967296.0,1,-nbitq), 
to_sfixed(283582273.0/4294967296.0,1,-nbitq), 
to_sfixed(-114787959.0/4294967296.0,1,-nbitq), 
to_sfixed(-272867983.0/4294967296.0,1,-nbitq), 
to_sfixed(24854195.0/4294967296.0,1,-nbitq), 
to_sfixed(180213944.0/4294967296.0,1,-nbitq), 
to_sfixed(-14085207.0/4294967296.0,1,-nbitq), 
to_sfixed(335372531.0/4294967296.0,1,-nbitq), 
to_sfixed(-150274286.0/4294967296.0,1,-nbitq), 
to_sfixed(43445458.0/4294967296.0,1,-nbitq), 
to_sfixed(-9990762.0/4294967296.0,1,-nbitq), 
to_sfixed(35051082.0/4294967296.0,1,-nbitq), 
to_sfixed(-136699843.0/4294967296.0,1,-nbitq), 
to_sfixed(-27567725.0/4294967296.0,1,-nbitq), 
to_sfixed(-14155646.0/4294967296.0,1,-nbitq), 
to_sfixed(-519674215.0/4294967296.0,1,-nbitq), 
to_sfixed(-89966330.0/4294967296.0,1,-nbitq), 
to_sfixed(-44014205.0/4294967296.0,1,-nbitq), 
to_sfixed(173494612.0/4294967296.0,1,-nbitq), 
to_sfixed(260128135.0/4294967296.0,1,-nbitq), 
to_sfixed(165590068.0/4294967296.0,1,-nbitq), 
to_sfixed(133032868.0/4294967296.0,1,-nbitq), 
to_sfixed(224047549.0/4294967296.0,1,-nbitq), 
to_sfixed(303611593.0/4294967296.0,1,-nbitq), 
to_sfixed(-401078910.0/4294967296.0,1,-nbitq), 
to_sfixed(256278845.0/4294967296.0,1,-nbitq), 
to_sfixed(132889534.0/4294967296.0,1,-nbitq), 
to_sfixed(390007522.0/4294967296.0,1,-nbitq), 
to_sfixed(90319899.0/4294967296.0,1,-nbitq), 
to_sfixed(192530296.0/4294967296.0,1,-nbitq), 
to_sfixed(-390728653.0/4294967296.0,1,-nbitq), 
to_sfixed(-297077657.0/4294967296.0,1,-nbitq), 
to_sfixed(-47145270.0/4294967296.0,1,-nbitq), 
to_sfixed(-44195797.0/4294967296.0,1,-nbitq), 
to_sfixed(-80461859.0/4294967296.0,1,-nbitq), 
to_sfixed(403248003.0/4294967296.0,1,-nbitq), 
to_sfixed(-181221400.0/4294967296.0,1,-nbitq), 
to_sfixed(-28822034.0/4294967296.0,1,-nbitq), 
to_sfixed(422479751.0/4294967296.0,1,-nbitq), 
to_sfixed(123225844.0/4294967296.0,1,-nbitq), 
to_sfixed(-306098202.0/4294967296.0,1,-nbitq), 
to_sfixed(-401197210.0/4294967296.0,1,-nbitq), 
to_sfixed(-40903024.0/4294967296.0,1,-nbitq), 
to_sfixed(179356138.0/4294967296.0,1,-nbitq), 
to_sfixed(-326619187.0/4294967296.0,1,-nbitq), 
to_sfixed(-188078019.0/4294967296.0,1,-nbitq), 
to_sfixed(31873379.0/4294967296.0,1,-nbitq), 
to_sfixed(205010439.0/4294967296.0,1,-nbitq), 
to_sfixed(-390382.0/4294967296.0,1,-nbitq), 
to_sfixed(52012828.0/4294967296.0,1,-nbitq), 
to_sfixed(203351430.0/4294967296.0,1,-nbitq), 
to_sfixed(-126460309.0/4294967296.0,1,-nbitq), 
to_sfixed(399659842.0/4294967296.0,1,-nbitq), 
to_sfixed(425729910.0/4294967296.0,1,-nbitq), 
to_sfixed(-362279791.0/4294967296.0,1,-nbitq), 
to_sfixed(-192535502.0/4294967296.0,1,-nbitq), 
to_sfixed(92178698.0/4294967296.0,1,-nbitq), 
to_sfixed(-302690981.0/4294967296.0,1,-nbitq), 
to_sfixed(268884768.0/4294967296.0,1,-nbitq), 
to_sfixed(-589591783.0/4294967296.0,1,-nbitq), 
to_sfixed(-296327187.0/4294967296.0,1,-nbitq), 
to_sfixed(17144031.0/4294967296.0,1,-nbitq), 
to_sfixed(-256267749.0/4294967296.0,1,-nbitq), 
to_sfixed(146592147.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(88463952.0/4294967296.0,1,-nbitq), 
to_sfixed(-367235726.0/4294967296.0,1,-nbitq), 
to_sfixed(199457618.0/4294967296.0,1,-nbitq), 
to_sfixed(226944221.0/4294967296.0,1,-nbitq), 
to_sfixed(-139303867.0/4294967296.0,1,-nbitq), 
to_sfixed(95251704.0/4294967296.0,1,-nbitq), 
to_sfixed(281545423.0/4294967296.0,1,-nbitq), 
to_sfixed(-358138671.0/4294967296.0,1,-nbitq), 
to_sfixed(278074285.0/4294967296.0,1,-nbitq), 
to_sfixed(-296333603.0/4294967296.0,1,-nbitq), 
to_sfixed(100609459.0/4294967296.0,1,-nbitq), 
to_sfixed(563261285.0/4294967296.0,1,-nbitq), 
to_sfixed(-384959001.0/4294967296.0,1,-nbitq), 
to_sfixed(-184281222.0/4294967296.0,1,-nbitq), 
to_sfixed(-198558422.0/4294967296.0,1,-nbitq), 
to_sfixed(-227199229.0/4294967296.0,1,-nbitq), 
to_sfixed(81574285.0/4294967296.0,1,-nbitq), 
to_sfixed(-109709429.0/4294967296.0,1,-nbitq), 
to_sfixed(454937810.0/4294967296.0,1,-nbitq), 
to_sfixed(226201272.0/4294967296.0,1,-nbitq), 
to_sfixed(288171300.0/4294967296.0,1,-nbitq), 
to_sfixed(-38771355.0/4294967296.0,1,-nbitq), 
to_sfixed(22954517.0/4294967296.0,1,-nbitq), 
to_sfixed(310437626.0/4294967296.0,1,-nbitq), 
to_sfixed(70098802.0/4294967296.0,1,-nbitq), 
to_sfixed(-192775599.0/4294967296.0,1,-nbitq), 
to_sfixed(-188435277.0/4294967296.0,1,-nbitq), 
to_sfixed(-340550643.0/4294967296.0,1,-nbitq), 
to_sfixed(-78898514.0/4294967296.0,1,-nbitq), 
to_sfixed(68680505.0/4294967296.0,1,-nbitq), 
to_sfixed(-435075437.0/4294967296.0,1,-nbitq), 
to_sfixed(-498469346.0/4294967296.0,1,-nbitq), 
to_sfixed(3980088.0/4294967296.0,1,-nbitq), 
to_sfixed(-451197629.0/4294967296.0,1,-nbitq), 
to_sfixed(24753227.0/4294967296.0,1,-nbitq), 
to_sfixed(323313102.0/4294967296.0,1,-nbitq), 
to_sfixed(161129569.0/4294967296.0,1,-nbitq), 
to_sfixed(121311443.0/4294967296.0,1,-nbitq), 
to_sfixed(-44294205.0/4294967296.0,1,-nbitq), 
to_sfixed(-279070403.0/4294967296.0,1,-nbitq), 
to_sfixed(-421700971.0/4294967296.0,1,-nbitq), 
to_sfixed(158722364.0/4294967296.0,1,-nbitq), 
to_sfixed(-363012917.0/4294967296.0,1,-nbitq), 
to_sfixed(332473676.0/4294967296.0,1,-nbitq), 
to_sfixed(-66704338.0/4294967296.0,1,-nbitq), 
to_sfixed(48044646.0/4294967296.0,1,-nbitq), 
to_sfixed(138735948.0/4294967296.0,1,-nbitq), 
to_sfixed(-272886351.0/4294967296.0,1,-nbitq), 
to_sfixed(4034842.0/4294967296.0,1,-nbitq), 
to_sfixed(306060561.0/4294967296.0,1,-nbitq), 
to_sfixed(-327461657.0/4294967296.0,1,-nbitq), 
to_sfixed(112965078.0/4294967296.0,1,-nbitq), 
to_sfixed(-653246795.0/4294967296.0,1,-nbitq), 
to_sfixed(167147520.0/4294967296.0,1,-nbitq), 
to_sfixed(326450543.0/4294967296.0,1,-nbitq), 
to_sfixed(-6492779.0/4294967296.0,1,-nbitq), 
to_sfixed(421568879.0/4294967296.0,1,-nbitq), 
to_sfixed(-41374546.0/4294967296.0,1,-nbitq), 
to_sfixed(-41868206.0/4294967296.0,1,-nbitq), 
to_sfixed(-107133232.0/4294967296.0,1,-nbitq), 
to_sfixed(-67219189.0/4294967296.0,1,-nbitq), 
to_sfixed(246644400.0/4294967296.0,1,-nbitq), 
to_sfixed(-413197117.0/4294967296.0,1,-nbitq), 
to_sfixed(96849992.0/4294967296.0,1,-nbitq), 
to_sfixed(3532088.0/4294967296.0,1,-nbitq), 
to_sfixed(-421711929.0/4294967296.0,1,-nbitq), 
to_sfixed(399850797.0/4294967296.0,1,-nbitq), 
to_sfixed(300950902.0/4294967296.0,1,-nbitq), 
to_sfixed(-163683820.0/4294967296.0,1,-nbitq), 
to_sfixed(-153099806.0/4294967296.0,1,-nbitq), 
to_sfixed(-229211058.0/4294967296.0,1,-nbitq), 
to_sfixed(-110764936.0/4294967296.0,1,-nbitq), 
to_sfixed(128303414.0/4294967296.0,1,-nbitq), 
to_sfixed(124971364.0/4294967296.0,1,-nbitq), 
to_sfixed(124873335.0/4294967296.0,1,-nbitq), 
to_sfixed(-97618627.0/4294967296.0,1,-nbitq), 
to_sfixed(-218229229.0/4294967296.0,1,-nbitq), 
to_sfixed(-281422038.0/4294967296.0,1,-nbitq), 
to_sfixed(-390497817.0/4294967296.0,1,-nbitq), 
to_sfixed(389791254.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(194077921.0/4294967296.0,1,-nbitq), 
to_sfixed(76667970.0/4294967296.0,1,-nbitq), 
to_sfixed(379434830.0/4294967296.0,1,-nbitq), 
to_sfixed(81473246.0/4294967296.0,1,-nbitq), 
to_sfixed(400790333.0/4294967296.0,1,-nbitq), 
to_sfixed(-303898381.0/4294967296.0,1,-nbitq), 
to_sfixed(41351432.0/4294967296.0,1,-nbitq), 
to_sfixed(125701932.0/4294967296.0,1,-nbitq), 
to_sfixed(49053635.0/4294967296.0,1,-nbitq), 
to_sfixed(-298018831.0/4294967296.0,1,-nbitq), 
to_sfixed(6452710.0/4294967296.0,1,-nbitq), 
to_sfixed(-212622175.0/4294967296.0,1,-nbitq), 
to_sfixed(202199429.0/4294967296.0,1,-nbitq), 
to_sfixed(-192139467.0/4294967296.0,1,-nbitq), 
to_sfixed(-422022189.0/4294967296.0,1,-nbitq), 
to_sfixed(-410522384.0/4294967296.0,1,-nbitq), 
to_sfixed(363207746.0/4294967296.0,1,-nbitq), 
to_sfixed(-123631209.0/4294967296.0,1,-nbitq), 
to_sfixed(216359344.0/4294967296.0,1,-nbitq), 
to_sfixed(115693865.0/4294967296.0,1,-nbitq), 
to_sfixed(114668604.0/4294967296.0,1,-nbitq), 
to_sfixed(-72875624.0/4294967296.0,1,-nbitq), 
to_sfixed(-43725571.0/4294967296.0,1,-nbitq), 
to_sfixed(-76449569.0/4294967296.0,1,-nbitq), 
to_sfixed(163572245.0/4294967296.0,1,-nbitq), 
to_sfixed(-82176334.0/4294967296.0,1,-nbitq), 
to_sfixed(9263860.0/4294967296.0,1,-nbitq), 
to_sfixed(13251961.0/4294967296.0,1,-nbitq), 
to_sfixed(243484745.0/4294967296.0,1,-nbitq), 
to_sfixed(136426344.0/4294967296.0,1,-nbitq), 
to_sfixed(-345212367.0/4294967296.0,1,-nbitq), 
to_sfixed(-152767214.0/4294967296.0,1,-nbitq), 
to_sfixed(-195354713.0/4294967296.0,1,-nbitq), 
to_sfixed(-132259953.0/4294967296.0,1,-nbitq), 
to_sfixed(298485714.0/4294967296.0,1,-nbitq), 
to_sfixed(195860889.0/4294967296.0,1,-nbitq), 
to_sfixed(-304866352.0/4294967296.0,1,-nbitq), 
to_sfixed(-131012388.0/4294967296.0,1,-nbitq), 
to_sfixed(155556638.0/4294967296.0,1,-nbitq), 
to_sfixed(270362695.0/4294967296.0,1,-nbitq), 
to_sfixed(111406521.0/4294967296.0,1,-nbitq), 
to_sfixed(122794050.0/4294967296.0,1,-nbitq), 
to_sfixed(95971578.0/4294967296.0,1,-nbitq), 
to_sfixed(498479397.0/4294967296.0,1,-nbitq), 
to_sfixed(-213199509.0/4294967296.0,1,-nbitq), 
to_sfixed(390062599.0/4294967296.0,1,-nbitq), 
to_sfixed(184304893.0/4294967296.0,1,-nbitq), 
to_sfixed(-415334932.0/4294967296.0,1,-nbitq), 
to_sfixed(-190139436.0/4294967296.0,1,-nbitq), 
to_sfixed(364419180.0/4294967296.0,1,-nbitq), 
to_sfixed(12615446.0/4294967296.0,1,-nbitq), 
to_sfixed(289528587.0/4294967296.0,1,-nbitq), 
to_sfixed(-234969951.0/4294967296.0,1,-nbitq), 
to_sfixed(-1794464.0/4294967296.0,1,-nbitq), 
to_sfixed(251135175.0/4294967296.0,1,-nbitq), 
to_sfixed(-218914978.0/4294967296.0,1,-nbitq), 
to_sfixed(-82541149.0/4294967296.0,1,-nbitq), 
to_sfixed(-365469582.0/4294967296.0,1,-nbitq), 
to_sfixed(-368619166.0/4294967296.0,1,-nbitq), 
to_sfixed(104785724.0/4294967296.0,1,-nbitq), 
to_sfixed(-86591156.0/4294967296.0,1,-nbitq), 
to_sfixed(313521674.0/4294967296.0,1,-nbitq), 
to_sfixed(-430797248.0/4294967296.0,1,-nbitq), 
to_sfixed(482700993.0/4294967296.0,1,-nbitq), 
to_sfixed(393216199.0/4294967296.0,1,-nbitq), 
to_sfixed(76127839.0/4294967296.0,1,-nbitq), 
to_sfixed(714808125.0/4294967296.0,1,-nbitq), 
to_sfixed(-28176460.0/4294967296.0,1,-nbitq), 
to_sfixed(245079511.0/4294967296.0,1,-nbitq), 
to_sfixed(256029345.0/4294967296.0,1,-nbitq), 
to_sfixed(-435608909.0/4294967296.0,1,-nbitq), 
to_sfixed(99665440.0/4294967296.0,1,-nbitq), 
to_sfixed(95530911.0/4294967296.0,1,-nbitq), 
to_sfixed(-192994680.0/4294967296.0,1,-nbitq), 
to_sfixed(182157678.0/4294967296.0,1,-nbitq), 
to_sfixed(-462484070.0/4294967296.0,1,-nbitq), 
to_sfixed(310794964.0/4294967296.0,1,-nbitq), 
to_sfixed(-482546825.0/4294967296.0,1,-nbitq), 
to_sfixed(144229594.0/4294967296.0,1,-nbitq), 
to_sfixed(340917329.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(135872739.0/4294967296.0,1,-nbitq), 
to_sfixed(-138830896.0/4294967296.0,1,-nbitq), 
to_sfixed(315607083.0/4294967296.0,1,-nbitq), 
to_sfixed(-267544568.0/4294967296.0,1,-nbitq), 
to_sfixed(-226388787.0/4294967296.0,1,-nbitq), 
to_sfixed(227777395.0/4294967296.0,1,-nbitq), 
to_sfixed(12926232.0/4294967296.0,1,-nbitq), 
to_sfixed(14281564.0/4294967296.0,1,-nbitq), 
to_sfixed(108044760.0/4294967296.0,1,-nbitq), 
to_sfixed(347587209.0/4294967296.0,1,-nbitq), 
to_sfixed(69169350.0/4294967296.0,1,-nbitq), 
to_sfixed(247703995.0/4294967296.0,1,-nbitq), 
to_sfixed(-343062607.0/4294967296.0,1,-nbitq), 
to_sfixed(-40026450.0/4294967296.0,1,-nbitq), 
to_sfixed(163595247.0/4294967296.0,1,-nbitq), 
to_sfixed(215656912.0/4294967296.0,1,-nbitq), 
to_sfixed(266849565.0/4294967296.0,1,-nbitq), 
to_sfixed(-145315078.0/4294967296.0,1,-nbitq), 
to_sfixed(14852506.0/4294967296.0,1,-nbitq), 
to_sfixed(342114403.0/4294967296.0,1,-nbitq), 
to_sfixed(-344099038.0/4294967296.0,1,-nbitq), 
to_sfixed(285668539.0/4294967296.0,1,-nbitq), 
to_sfixed(164726353.0/4294967296.0,1,-nbitq), 
to_sfixed(-245124814.0/4294967296.0,1,-nbitq), 
to_sfixed(401087885.0/4294967296.0,1,-nbitq), 
to_sfixed(476065936.0/4294967296.0,1,-nbitq), 
to_sfixed(293091680.0/4294967296.0,1,-nbitq), 
to_sfixed(41650456.0/4294967296.0,1,-nbitq), 
to_sfixed(385397962.0/4294967296.0,1,-nbitq), 
to_sfixed(182325319.0/4294967296.0,1,-nbitq), 
to_sfixed(-44193572.0/4294967296.0,1,-nbitq), 
to_sfixed(256895455.0/4294967296.0,1,-nbitq), 
to_sfixed(280019641.0/4294967296.0,1,-nbitq), 
to_sfixed(-268357833.0/4294967296.0,1,-nbitq), 
to_sfixed(-33029288.0/4294967296.0,1,-nbitq), 
to_sfixed(32778752.0/4294967296.0,1,-nbitq), 
to_sfixed(-27729723.0/4294967296.0,1,-nbitq), 
to_sfixed(-301790279.0/4294967296.0,1,-nbitq), 
to_sfixed(-387618696.0/4294967296.0,1,-nbitq), 
to_sfixed(232106526.0/4294967296.0,1,-nbitq), 
to_sfixed(271896309.0/4294967296.0,1,-nbitq), 
to_sfixed(145951561.0/4294967296.0,1,-nbitq), 
to_sfixed(-198406063.0/4294967296.0,1,-nbitq), 
to_sfixed(-44294094.0/4294967296.0,1,-nbitq), 
to_sfixed(-117478942.0/4294967296.0,1,-nbitq), 
to_sfixed(286212072.0/4294967296.0,1,-nbitq), 
to_sfixed(189851560.0/4294967296.0,1,-nbitq), 
to_sfixed(-514875613.0/4294967296.0,1,-nbitq), 
to_sfixed(-125291645.0/4294967296.0,1,-nbitq), 
to_sfixed(74424937.0/4294967296.0,1,-nbitq), 
to_sfixed(-86102779.0/4294967296.0,1,-nbitq), 
to_sfixed(-61868245.0/4294967296.0,1,-nbitq), 
to_sfixed(-492341001.0/4294967296.0,1,-nbitq), 
to_sfixed(-18246760.0/4294967296.0,1,-nbitq), 
to_sfixed(173474521.0/4294967296.0,1,-nbitq), 
to_sfixed(-254461507.0/4294967296.0,1,-nbitq), 
to_sfixed(320305015.0/4294967296.0,1,-nbitq), 
to_sfixed(27526807.0/4294967296.0,1,-nbitq), 
to_sfixed(224543848.0/4294967296.0,1,-nbitq), 
to_sfixed(-49829005.0/4294967296.0,1,-nbitq), 
to_sfixed(252411308.0/4294967296.0,1,-nbitq), 
to_sfixed(304059896.0/4294967296.0,1,-nbitq), 
to_sfixed(-220127955.0/4294967296.0,1,-nbitq), 
to_sfixed(87629752.0/4294967296.0,1,-nbitq), 
to_sfixed(121478436.0/4294967296.0,1,-nbitq), 
to_sfixed(-461000108.0/4294967296.0,1,-nbitq), 
to_sfixed(93346439.0/4294967296.0,1,-nbitq), 
to_sfixed(288594414.0/4294967296.0,1,-nbitq), 
to_sfixed(24407205.0/4294967296.0,1,-nbitq), 
to_sfixed(477192772.0/4294967296.0,1,-nbitq), 
to_sfixed(-224038640.0/4294967296.0,1,-nbitq), 
to_sfixed(306631160.0/4294967296.0,1,-nbitq), 
to_sfixed(-308980191.0/4294967296.0,1,-nbitq), 
to_sfixed(448850832.0/4294967296.0,1,-nbitq), 
to_sfixed(222791016.0/4294967296.0,1,-nbitq), 
to_sfixed(-318895339.0/4294967296.0,1,-nbitq), 
to_sfixed(-7700885.0/4294967296.0,1,-nbitq), 
to_sfixed(114943967.0/4294967296.0,1,-nbitq), 
to_sfixed(21087588.0/4294967296.0,1,-nbitq), 
to_sfixed(-99511853.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-344387436.0/4294967296.0,1,-nbitq), 
to_sfixed(-578229542.0/4294967296.0,1,-nbitq), 
to_sfixed(-85276204.0/4294967296.0,1,-nbitq), 
to_sfixed(126760802.0/4294967296.0,1,-nbitq), 
to_sfixed(-8236298.0/4294967296.0,1,-nbitq), 
to_sfixed(25296451.0/4294967296.0,1,-nbitq), 
to_sfixed(-261544900.0/4294967296.0,1,-nbitq), 
to_sfixed(-463323816.0/4294967296.0,1,-nbitq), 
to_sfixed(-227407790.0/4294967296.0,1,-nbitq), 
to_sfixed(-366948436.0/4294967296.0,1,-nbitq), 
to_sfixed(142452716.0/4294967296.0,1,-nbitq), 
to_sfixed(-227712301.0/4294967296.0,1,-nbitq), 
to_sfixed(348153137.0/4294967296.0,1,-nbitq), 
to_sfixed(154215203.0/4294967296.0,1,-nbitq), 
to_sfixed(-247153444.0/4294967296.0,1,-nbitq), 
to_sfixed(199498488.0/4294967296.0,1,-nbitq), 
to_sfixed(-313256689.0/4294967296.0,1,-nbitq), 
to_sfixed(-102071703.0/4294967296.0,1,-nbitq), 
to_sfixed(162755741.0/4294967296.0,1,-nbitq), 
to_sfixed(-85694121.0/4294967296.0,1,-nbitq), 
to_sfixed(279600851.0/4294967296.0,1,-nbitq), 
to_sfixed(191219236.0/4294967296.0,1,-nbitq), 
to_sfixed(-163822217.0/4294967296.0,1,-nbitq), 
to_sfixed(86097548.0/4294967296.0,1,-nbitq), 
to_sfixed(215229668.0/4294967296.0,1,-nbitq), 
to_sfixed(-128393640.0/4294967296.0,1,-nbitq), 
to_sfixed(182646721.0/4294967296.0,1,-nbitq), 
to_sfixed(-582638612.0/4294967296.0,1,-nbitq), 
to_sfixed(456614175.0/4294967296.0,1,-nbitq), 
to_sfixed(176874500.0/4294967296.0,1,-nbitq), 
to_sfixed(-360303399.0/4294967296.0,1,-nbitq), 
to_sfixed(-30402788.0/4294967296.0,1,-nbitq), 
to_sfixed(-53249885.0/4294967296.0,1,-nbitq), 
to_sfixed(241024389.0/4294967296.0,1,-nbitq), 
to_sfixed(299590655.0/4294967296.0,1,-nbitq), 
to_sfixed(84660364.0/4294967296.0,1,-nbitq), 
to_sfixed(-167990853.0/4294967296.0,1,-nbitq), 
to_sfixed(155172725.0/4294967296.0,1,-nbitq), 
to_sfixed(61514573.0/4294967296.0,1,-nbitq), 
to_sfixed(-117667837.0/4294967296.0,1,-nbitq), 
to_sfixed(-143191701.0/4294967296.0,1,-nbitq), 
to_sfixed(375601261.0/4294967296.0,1,-nbitq), 
to_sfixed(-326740950.0/4294967296.0,1,-nbitq), 
to_sfixed(-179829574.0/4294967296.0,1,-nbitq), 
to_sfixed(191263689.0/4294967296.0,1,-nbitq), 
to_sfixed(101784876.0/4294967296.0,1,-nbitq), 
to_sfixed(333292471.0/4294967296.0,1,-nbitq), 
to_sfixed(-47439016.0/4294967296.0,1,-nbitq), 
to_sfixed(170275788.0/4294967296.0,1,-nbitq), 
to_sfixed(101421566.0/4294967296.0,1,-nbitq), 
to_sfixed(-53355039.0/4294967296.0,1,-nbitq), 
to_sfixed(-10251894.0/4294967296.0,1,-nbitq), 
to_sfixed(229508829.0/4294967296.0,1,-nbitq), 
to_sfixed(-16050594.0/4294967296.0,1,-nbitq), 
to_sfixed(380612999.0/4294967296.0,1,-nbitq), 
to_sfixed(90910342.0/4294967296.0,1,-nbitq), 
to_sfixed(13455426.0/4294967296.0,1,-nbitq), 
to_sfixed(83282643.0/4294967296.0,1,-nbitq), 
to_sfixed(-332072254.0/4294967296.0,1,-nbitq), 
to_sfixed(364457002.0/4294967296.0,1,-nbitq), 
to_sfixed(252079666.0/4294967296.0,1,-nbitq), 
to_sfixed(-182429358.0/4294967296.0,1,-nbitq), 
to_sfixed(171506934.0/4294967296.0,1,-nbitq), 
to_sfixed(51247460.0/4294967296.0,1,-nbitq), 
to_sfixed(421384463.0/4294967296.0,1,-nbitq), 
to_sfixed(203853347.0/4294967296.0,1,-nbitq), 
to_sfixed(172298957.0/4294967296.0,1,-nbitq), 
to_sfixed(-337313555.0/4294967296.0,1,-nbitq), 
to_sfixed(-199402408.0/4294967296.0,1,-nbitq), 
to_sfixed(97071518.0/4294967296.0,1,-nbitq), 
to_sfixed(-40868184.0/4294967296.0,1,-nbitq), 
to_sfixed(40442161.0/4294967296.0,1,-nbitq), 
to_sfixed(-482429891.0/4294967296.0,1,-nbitq), 
to_sfixed(-157945895.0/4294967296.0,1,-nbitq), 
to_sfixed(-124214867.0/4294967296.0,1,-nbitq), 
to_sfixed(81500493.0/4294967296.0,1,-nbitq), 
to_sfixed(-148706692.0/4294967296.0,1,-nbitq), 
to_sfixed(231965659.0/4294967296.0,1,-nbitq), 
to_sfixed(-477273675.0/4294967296.0,1,-nbitq), 
to_sfixed(-7880855.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(383198553.0/4294967296.0,1,-nbitq), 
to_sfixed(-115394666.0/4294967296.0,1,-nbitq), 
to_sfixed(-184692253.0/4294967296.0,1,-nbitq), 
to_sfixed(191942125.0/4294967296.0,1,-nbitq), 
to_sfixed(-23828262.0/4294967296.0,1,-nbitq), 
to_sfixed(206545444.0/4294967296.0,1,-nbitq), 
to_sfixed(-287019420.0/4294967296.0,1,-nbitq), 
to_sfixed(-69794875.0/4294967296.0,1,-nbitq), 
to_sfixed(-408289251.0/4294967296.0,1,-nbitq), 
to_sfixed(92125563.0/4294967296.0,1,-nbitq), 
to_sfixed(-183185570.0/4294967296.0,1,-nbitq), 
to_sfixed(255337832.0/4294967296.0,1,-nbitq), 
to_sfixed(-276357297.0/4294967296.0,1,-nbitq), 
to_sfixed(-57108254.0/4294967296.0,1,-nbitq), 
to_sfixed(-284634371.0/4294967296.0,1,-nbitq), 
to_sfixed(-70026628.0/4294967296.0,1,-nbitq), 
to_sfixed(310056202.0/4294967296.0,1,-nbitq), 
to_sfixed(158061242.0/4294967296.0,1,-nbitq), 
to_sfixed(187846866.0/4294967296.0,1,-nbitq), 
to_sfixed(-400567631.0/4294967296.0,1,-nbitq), 
to_sfixed(-80252000.0/4294967296.0,1,-nbitq), 
to_sfixed(-80554609.0/4294967296.0,1,-nbitq), 
to_sfixed(416722575.0/4294967296.0,1,-nbitq), 
to_sfixed(184159149.0/4294967296.0,1,-nbitq), 
to_sfixed(-162941989.0/4294967296.0,1,-nbitq), 
to_sfixed(-34650488.0/4294967296.0,1,-nbitq), 
to_sfixed(-146198942.0/4294967296.0,1,-nbitq), 
to_sfixed(-100941090.0/4294967296.0,1,-nbitq), 
to_sfixed(-225614793.0/4294967296.0,1,-nbitq), 
to_sfixed(257779189.0/4294967296.0,1,-nbitq), 
to_sfixed(-611049397.0/4294967296.0,1,-nbitq), 
to_sfixed(-330232669.0/4294967296.0,1,-nbitq), 
to_sfixed(-232270721.0/4294967296.0,1,-nbitq), 
to_sfixed(232716572.0/4294967296.0,1,-nbitq), 
to_sfixed(-125036684.0/4294967296.0,1,-nbitq), 
to_sfixed(348315120.0/4294967296.0,1,-nbitq), 
to_sfixed(-85184366.0/4294967296.0,1,-nbitq), 
to_sfixed(195078106.0/4294967296.0,1,-nbitq), 
to_sfixed(27383297.0/4294967296.0,1,-nbitq), 
to_sfixed(-269934583.0/4294967296.0,1,-nbitq), 
to_sfixed(-153380741.0/4294967296.0,1,-nbitq), 
to_sfixed(389463707.0/4294967296.0,1,-nbitq), 
to_sfixed(124967662.0/4294967296.0,1,-nbitq), 
to_sfixed(-74693094.0/4294967296.0,1,-nbitq), 
to_sfixed(107366799.0/4294967296.0,1,-nbitq), 
to_sfixed(-456661.0/4294967296.0,1,-nbitq), 
to_sfixed(-399503744.0/4294967296.0,1,-nbitq), 
to_sfixed(-187638489.0/4294967296.0,1,-nbitq), 
to_sfixed(90851776.0/4294967296.0,1,-nbitq), 
to_sfixed(-167711244.0/4294967296.0,1,-nbitq), 
to_sfixed(192326812.0/4294967296.0,1,-nbitq), 
to_sfixed(253256124.0/4294967296.0,1,-nbitq), 
to_sfixed(-413864843.0/4294967296.0,1,-nbitq), 
to_sfixed(33986146.0/4294967296.0,1,-nbitq), 
to_sfixed(-189326882.0/4294967296.0,1,-nbitq), 
to_sfixed(-312278128.0/4294967296.0,1,-nbitq), 
to_sfixed(458652029.0/4294967296.0,1,-nbitq), 
to_sfixed(-54755063.0/4294967296.0,1,-nbitq), 
to_sfixed(-252576828.0/4294967296.0,1,-nbitq), 
to_sfixed(-322136756.0/4294967296.0,1,-nbitq), 
to_sfixed(242980389.0/4294967296.0,1,-nbitq), 
to_sfixed(105765343.0/4294967296.0,1,-nbitq), 
to_sfixed(-391787303.0/4294967296.0,1,-nbitq), 
to_sfixed(347779614.0/4294967296.0,1,-nbitq), 
to_sfixed(-22811896.0/4294967296.0,1,-nbitq), 
to_sfixed(84746350.0/4294967296.0,1,-nbitq), 
to_sfixed(594687503.0/4294967296.0,1,-nbitq), 
to_sfixed(-100872882.0/4294967296.0,1,-nbitq), 
to_sfixed(230094324.0/4294967296.0,1,-nbitq), 
to_sfixed(198694694.0/4294967296.0,1,-nbitq), 
to_sfixed(-196665735.0/4294967296.0,1,-nbitq), 
to_sfixed(-344235389.0/4294967296.0,1,-nbitq), 
to_sfixed(-300677010.0/4294967296.0,1,-nbitq), 
to_sfixed(-317213948.0/4294967296.0,1,-nbitq), 
to_sfixed(214100711.0/4294967296.0,1,-nbitq), 
to_sfixed(-98675865.0/4294967296.0,1,-nbitq), 
to_sfixed(-291381008.0/4294967296.0,1,-nbitq), 
to_sfixed(40324447.0/4294967296.0,1,-nbitq), 
to_sfixed(-301972165.0/4294967296.0,1,-nbitq), 
to_sfixed(-43108359.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-103925446.0/4294967296.0,1,-nbitq), 
to_sfixed(-213406934.0/4294967296.0,1,-nbitq), 
to_sfixed(-109217977.0/4294967296.0,1,-nbitq), 
to_sfixed(-277303642.0/4294967296.0,1,-nbitq), 
to_sfixed(445718036.0/4294967296.0,1,-nbitq), 
to_sfixed(105781497.0/4294967296.0,1,-nbitq), 
to_sfixed(-399078633.0/4294967296.0,1,-nbitq), 
to_sfixed(-291627803.0/4294967296.0,1,-nbitq), 
to_sfixed(73805463.0/4294967296.0,1,-nbitq), 
to_sfixed(-324212655.0/4294967296.0,1,-nbitq), 
to_sfixed(-331430755.0/4294967296.0,1,-nbitq), 
to_sfixed(353510469.0/4294967296.0,1,-nbitq), 
to_sfixed(-80699723.0/4294967296.0,1,-nbitq), 
to_sfixed(153821086.0/4294967296.0,1,-nbitq), 
to_sfixed(3672076.0/4294967296.0,1,-nbitq), 
to_sfixed(316094605.0/4294967296.0,1,-nbitq), 
to_sfixed(113856920.0/4294967296.0,1,-nbitq), 
to_sfixed(-173892493.0/4294967296.0,1,-nbitq), 
to_sfixed(168742049.0/4294967296.0,1,-nbitq), 
to_sfixed(-64082238.0/4294967296.0,1,-nbitq), 
to_sfixed(-291933581.0/4294967296.0,1,-nbitq), 
to_sfixed(430687021.0/4294967296.0,1,-nbitq), 
to_sfixed(504258914.0/4294967296.0,1,-nbitq), 
to_sfixed(416550912.0/4294967296.0,1,-nbitq), 
to_sfixed(-253323910.0/4294967296.0,1,-nbitq), 
to_sfixed(466165237.0/4294967296.0,1,-nbitq), 
to_sfixed(-330713062.0/4294967296.0,1,-nbitq), 
to_sfixed(26272046.0/4294967296.0,1,-nbitq), 
to_sfixed(394744661.0/4294967296.0,1,-nbitq), 
to_sfixed(45777825.0/4294967296.0,1,-nbitq), 
to_sfixed(-361108706.0/4294967296.0,1,-nbitq), 
to_sfixed(-19777570.0/4294967296.0,1,-nbitq), 
to_sfixed(78530144.0/4294967296.0,1,-nbitq), 
to_sfixed(232779470.0/4294967296.0,1,-nbitq), 
to_sfixed(547706997.0/4294967296.0,1,-nbitq), 
to_sfixed(-68794544.0/4294967296.0,1,-nbitq), 
to_sfixed(424784591.0/4294967296.0,1,-nbitq), 
to_sfixed(304510150.0/4294967296.0,1,-nbitq), 
to_sfixed(211815574.0/4294967296.0,1,-nbitq), 
to_sfixed(420976607.0/4294967296.0,1,-nbitq), 
to_sfixed(-351239074.0/4294967296.0,1,-nbitq), 
to_sfixed(419231840.0/4294967296.0,1,-nbitq), 
to_sfixed(176226162.0/4294967296.0,1,-nbitq), 
to_sfixed(-327648981.0/4294967296.0,1,-nbitq), 
to_sfixed(-297141988.0/4294967296.0,1,-nbitq), 
to_sfixed(45762565.0/4294967296.0,1,-nbitq), 
to_sfixed(-285104944.0/4294967296.0,1,-nbitq), 
to_sfixed(208422931.0/4294967296.0,1,-nbitq), 
to_sfixed(320919003.0/4294967296.0,1,-nbitq), 
to_sfixed(185934411.0/4294967296.0,1,-nbitq), 
to_sfixed(142873913.0/4294967296.0,1,-nbitq), 
to_sfixed(468729065.0/4294967296.0,1,-nbitq), 
to_sfixed(198121665.0/4294967296.0,1,-nbitq), 
to_sfixed(-89356504.0/4294967296.0,1,-nbitq), 
to_sfixed(245662915.0/4294967296.0,1,-nbitq), 
to_sfixed(-157948639.0/4294967296.0,1,-nbitq), 
to_sfixed(318395626.0/4294967296.0,1,-nbitq), 
to_sfixed(-170714142.0/4294967296.0,1,-nbitq), 
to_sfixed(-307447717.0/4294967296.0,1,-nbitq), 
to_sfixed(237224609.0/4294967296.0,1,-nbitq), 
to_sfixed(-118932527.0/4294967296.0,1,-nbitq), 
to_sfixed(-169585437.0/4294967296.0,1,-nbitq), 
to_sfixed(-74552831.0/4294967296.0,1,-nbitq), 
to_sfixed(436026756.0/4294967296.0,1,-nbitq), 
to_sfixed(-73640655.0/4294967296.0,1,-nbitq), 
to_sfixed(-117638951.0/4294967296.0,1,-nbitq), 
to_sfixed(838372625.0/4294967296.0,1,-nbitq), 
to_sfixed(-214280416.0/4294967296.0,1,-nbitq), 
to_sfixed(-110282776.0/4294967296.0,1,-nbitq), 
to_sfixed(-39582439.0/4294967296.0,1,-nbitq), 
to_sfixed(259853603.0/4294967296.0,1,-nbitq), 
to_sfixed(132016931.0/4294967296.0,1,-nbitq), 
to_sfixed(-99238318.0/4294967296.0,1,-nbitq), 
to_sfixed(399074106.0/4294967296.0,1,-nbitq), 
to_sfixed(72865419.0/4294967296.0,1,-nbitq), 
to_sfixed(-18556245.0/4294967296.0,1,-nbitq), 
to_sfixed(-259325202.0/4294967296.0,1,-nbitq), 
to_sfixed(-473381384.0/4294967296.0,1,-nbitq), 
to_sfixed(-136030428.0/4294967296.0,1,-nbitq), 
to_sfixed(381030529.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-376711877.0/4294967296.0,1,-nbitq), 
to_sfixed(-11496080.0/4294967296.0,1,-nbitq), 
to_sfixed(445180284.0/4294967296.0,1,-nbitq), 
to_sfixed(194528045.0/4294967296.0,1,-nbitq), 
to_sfixed(346591735.0/4294967296.0,1,-nbitq), 
to_sfixed(193460922.0/4294967296.0,1,-nbitq), 
to_sfixed(-60095749.0/4294967296.0,1,-nbitq), 
to_sfixed(-103242841.0/4294967296.0,1,-nbitq), 
to_sfixed(6809176.0/4294967296.0,1,-nbitq), 
to_sfixed(154606436.0/4294967296.0,1,-nbitq), 
to_sfixed(-302758851.0/4294967296.0,1,-nbitq), 
to_sfixed(-32505678.0/4294967296.0,1,-nbitq), 
to_sfixed(237010252.0/4294967296.0,1,-nbitq), 
to_sfixed(454076748.0/4294967296.0,1,-nbitq), 
to_sfixed(-334175410.0/4294967296.0,1,-nbitq), 
to_sfixed(-354238199.0/4294967296.0,1,-nbitq), 
to_sfixed(231000559.0/4294967296.0,1,-nbitq), 
to_sfixed(-386086213.0/4294967296.0,1,-nbitq), 
to_sfixed(-89951950.0/4294967296.0,1,-nbitq), 
to_sfixed(226486484.0/4294967296.0,1,-nbitq), 
to_sfixed(207541854.0/4294967296.0,1,-nbitq), 
to_sfixed(431840112.0/4294967296.0,1,-nbitq), 
to_sfixed(337756724.0/4294967296.0,1,-nbitq), 
to_sfixed(202558935.0/4294967296.0,1,-nbitq), 
to_sfixed(282336454.0/4294967296.0,1,-nbitq), 
to_sfixed(-22091058.0/4294967296.0,1,-nbitq), 
to_sfixed(-29133054.0/4294967296.0,1,-nbitq), 
to_sfixed(22579120.0/4294967296.0,1,-nbitq), 
to_sfixed(186353501.0/4294967296.0,1,-nbitq), 
to_sfixed(389223512.0/4294967296.0,1,-nbitq), 
to_sfixed(-23754359.0/4294967296.0,1,-nbitq), 
to_sfixed(-376216995.0/4294967296.0,1,-nbitq), 
to_sfixed(180048241.0/4294967296.0,1,-nbitq), 
to_sfixed(254383813.0/4294967296.0,1,-nbitq), 
to_sfixed(-76390811.0/4294967296.0,1,-nbitq), 
to_sfixed(128870934.0/4294967296.0,1,-nbitq), 
to_sfixed(-196368129.0/4294967296.0,1,-nbitq), 
to_sfixed(-267985525.0/4294967296.0,1,-nbitq), 
to_sfixed(263008547.0/4294967296.0,1,-nbitq), 
to_sfixed(396002133.0/4294967296.0,1,-nbitq), 
to_sfixed(-346224815.0/4294967296.0,1,-nbitq), 
to_sfixed(-100860708.0/4294967296.0,1,-nbitq), 
to_sfixed(-254649825.0/4294967296.0,1,-nbitq), 
to_sfixed(335424290.0/4294967296.0,1,-nbitq), 
to_sfixed(185804689.0/4294967296.0,1,-nbitq), 
to_sfixed(434452191.0/4294967296.0,1,-nbitq), 
to_sfixed(269129355.0/4294967296.0,1,-nbitq), 
to_sfixed(170615189.0/4294967296.0,1,-nbitq), 
to_sfixed(-297673894.0/4294967296.0,1,-nbitq), 
to_sfixed(-138751362.0/4294967296.0,1,-nbitq), 
to_sfixed(-200791133.0/4294967296.0,1,-nbitq), 
to_sfixed(-212590554.0/4294967296.0,1,-nbitq), 
to_sfixed(-554958479.0/4294967296.0,1,-nbitq), 
to_sfixed(319002917.0/4294967296.0,1,-nbitq), 
to_sfixed(-175111033.0/4294967296.0,1,-nbitq), 
to_sfixed(-257497880.0/4294967296.0,1,-nbitq), 
to_sfixed(70747337.0/4294967296.0,1,-nbitq), 
to_sfixed(-276363226.0/4294967296.0,1,-nbitq), 
to_sfixed(118958559.0/4294967296.0,1,-nbitq), 
to_sfixed(11823179.0/4294967296.0,1,-nbitq), 
to_sfixed(299125864.0/4294967296.0,1,-nbitq), 
to_sfixed(371088167.0/4294967296.0,1,-nbitq), 
to_sfixed(298185415.0/4294967296.0,1,-nbitq), 
to_sfixed(190527066.0/4294967296.0,1,-nbitq), 
to_sfixed(-140821379.0/4294967296.0,1,-nbitq), 
to_sfixed(-248282839.0/4294967296.0,1,-nbitq), 
to_sfixed(361374737.0/4294967296.0,1,-nbitq), 
to_sfixed(-395289732.0/4294967296.0,1,-nbitq), 
to_sfixed(338173200.0/4294967296.0,1,-nbitq), 
to_sfixed(535874155.0/4294967296.0,1,-nbitq), 
to_sfixed(-163346424.0/4294967296.0,1,-nbitq), 
to_sfixed(-366492828.0/4294967296.0,1,-nbitq), 
to_sfixed(164333478.0/4294967296.0,1,-nbitq), 
to_sfixed(8293713.0/4294967296.0,1,-nbitq), 
to_sfixed(86796382.0/4294967296.0,1,-nbitq), 
to_sfixed(-202273386.0/4294967296.0,1,-nbitq), 
to_sfixed(-444358341.0/4294967296.0,1,-nbitq), 
to_sfixed(70461598.0/4294967296.0,1,-nbitq), 
to_sfixed(-463678948.0/4294967296.0,1,-nbitq), 
to_sfixed(-335617211.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-361222015.0/4294967296.0,1,-nbitq), 
to_sfixed(-39984956.0/4294967296.0,1,-nbitq), 
to_sfixed(-200776440.0/4294967296.0,1,-nbitq), 
to_sfixed(-138803195.0/4294967296.0,1,-nbitq), 
to_sfixed(373582914.0/4294967296.0,1,-nbitq), 
to_sfixed(295715956.0/4294967296.0,1,-nbitq), 
to_sfixed(179358853.0/4294967296.0,1,-nbitq), 
to_sfixed(317311888.0/4294967296.0,1,-nbitq), 
to_sfixed(-458901656.0/4294967296.0,1,-nbitq), 
to_sfixed(237838772.0/4294967296.0,1,-nbitq), 
to_sfixed(-164708070.0/4294967296.0,1,-nbitq), 
to_sfixed(-18808773.0/4294967296.0,1,-nbitq), 
to_sfixed(-234754418.0/4294967296.0,1,-nbitq), 
to_sfixed(-258688842.0/4294967296.0,1,-nbitq), 
to_sfixed(-189027809.0/4294967296.0,1,-nbitq), 
to_sfixed(-149989963.0/4294967296.0,1,-nbitq), 
to_sfixed(173824209.0/4294967296.0,1,-nbitq), 
to_sfixed(115136939.0/4294967296.0,1,-nbitq), 
to_sfixed(438788676.0/4294967296.0,1,-nbitq), 
to_sfixed(391758574.0/4294967296.0,1,-nbitq), 
to_sfixed(-91311908.0/4294967296.0,1,-nbitq), 
to_sfixed(145694570.0/4294967296.0,1,-nbitq), 
to_sfixed(512330499.0/4294967296.0,1,-nbitq), 
to_sfixed(288992062.0/4294967296.0,1,-nbitq), 
to_sfixed(160808837.0/4294967296.0,1,-nbitq), 
to_sfixed(232775755.0/4294967296.0,1,-nbitq), 
to_sfixed(52149233.0/4294967296.0,1,-nbitq), 
to_sfixed(-514326814.0/4294967296.0,1,-nbitq), 
to_sfixed(-88163803.0/4294967296.0,1,-nbitq), 
to_sfixed(-133389480.0/4294967296.0,1,-nbitq), 
to_sfixed(-535969281.0/4294967296.0,1,-nbitq), 
to_sfixed(-44977128.0/4294967296.0,1,-nbitq), 
to_sfixed(93006614.0/4294967296.0,1,-nbitq), 
to_sfixed(-294460419.0/4294967296.0,1,-nbitq), 
to_sfixed(124081477.0/4294967296.0,1,-nbitq), 
to_sfixed(-446795534.0/4294967296.0,1,-nbitq), 
to_sfixed(134811728.0/4294967296.0,1,-nbitq), 
to_sfixed(-11400523.0/4294967296.0,1,-nbitq), 
to_sfixed(-374682501.0/4294967296.0,1,-nbitq), 
to_sfixed(489083095.0/4294967296.0,1,-nbitq), 
to_sfixed(-158305174.0/4294967296.0,1,-nbitq), 
to_sfixed(-280783833.0/4294967296.0,1,-nbitq), 
to_sfixed(-48144626.0/4294967296.0,1,-nbitq), 
to_sfixed(307568174.0/4294967296.0,1,-nbitq), 
to_sfixed(-94780157.0/4294967296.0,1,-nbitq), 
to_sfixed(467473177.0/4294967296.0,1,-nbitq), 
to_sfixed(97978305.0/4294967296.0,1,-nbitq), 
to_sfixed(150123176.0/4294967296.0,1,-nbitq), 
to_sfixed(-364334652.0/4294967296.0,1,-nbitq), 
to_sfixed(156961894.0/4294967296.0,1,-nbitq), 
to_sfixed(-164944377.0/4294967296.0,1,-nbitq), 
to_sfixed(-337329411.0/4294967296.0,1,-nbitq), 
to_sfixed(158051293.0/4294967296.0,1,-nbitq), 
to_sfixed(444672761.0/4294967296.0,1,-nbitq), 
to_sfixed(-214402532.0/4294967296.0,1,-nbitq), 
to_sfixed(190099859.0/4294967296.0,1,-nbitq), 
to_sfixed(274305651.0/4294967296.0,1,-nbitq), 
to_sfixed(60888627.0/4294967296.0,1,-nbitq), 
to_sfixed(-220870037.0/4294967296.0,1,-nbitq), 
to_sfixed(-124653295.0/4294967296.0,1,-nbitq), 
to_sfixed(289573395.0/4294967296.0,1,-nbitq), 
to_sfixed(14647591.0/4294967296.0,1,-nbitq), 
to_sfixed(-11911109.0/4294967296.0,1,-nbitq), 
to_sfixed(171855969.0/4294967296.0,1,-nbitq), 
to_sfixed(-258948448.0/4294967296.0,1,-nbitq), 
to_sfixed(159514490.0/4294967296.0,1,-nbitq), 
to_sfixed(223788845.0/4294967296.0,1,-nbitq), 
to_sfixed(-348894756.0/4294967296.0,1,-nbitq), 
to_sfixed(103882558.0/4294967296.0,1,-nbitq), 
to_sfixed(-238441221.0/4294967296.0,1,-nbitq), 
to_sfixed(-379370549.0/4294967296.0,1,-nbitq), 
to_sfixed(-62356195.0/4294967296.0,1,-nbitq), 
to_sfixed(108255649.0/4294967296.0,1,-nbitq), 
to_sfixed(138975822.0/4294967296.0,1,-nbitq), 
to_sfixed(-252384219.0/4294967296.0,1,-nbitq), 
to_sfixed(-540041560.0/4294967296.0,1,-nbitq), 
to_sfixed(-251576059.0/4294967296.0,1,-nbitq), 
to_sfixed(16293334.0/4294967296.0,1,-nbitq), 
to_sfixed(80752281.0/4294967296.0,1,-nbitq), 
to_sfixed(-42242504.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(134084743.0/4294967296.0,1,-nbitq), 
to_sfixed(-350316253.0/4294967296.0,1,-nbitq), 
to_sfixed(-223552064.0/4294967296.0,1,-nbitq), 
to_sfixed(91987954.0/4294967296.0,1,-nbitq), 
to_sfixed(257225399.0/4294967296.0,1,-nbitq), 
to_sfixed(79250059.0/4294967296.0,1,-nbitq), 
to_sfixed(-123445618.0/4294967296.0,1,-nbitq), 
to_sfixed(205279191.0/4294967296.0,1,-nbitq), 
to_sfixed(-433348162.0/4294967296.0,1,-nbitq), 
to_sfixed(449896964.0/4294967296.0,1,-nbitq), 
to_sfixed(-218734607.0/4294967296.0,1,-nbitq), 
to_sfixed(318896517.0/4294967296.0,1,-nbitq), 
to_sfixed(192573013.0/4294967296.0,1,-nbitq), 
to_sfixed(-102387492.0/4294967296.0,1,-nbitq), 
to_sfixed(-260200980.0/4294967296.0,1,-nbitq), 
to_sfixed(-314379464.0/4294967296.0,1,-nbitq), 
to_sfixed(209036706.0/4294967296.0,1,-nbitq), 
to_sfixed(-341138029.0/4294967296.0,1,-nbitq), 
to_sfixed(8873080.0/4294967296.0,1,-nbitq), 
to_sfixed(-342082353.0/4294967296.0,1,-nbitq), 
to_sfixed(-344099608.0/4294967296.0,1,-nbitq), 
to_sfixed(379086998.0/4294967296.0,1,-nbitq), 
to_sfixed(19814568.0/4294967296.0,1,-nbitq), 
to_sfixed(85023922.0/4294967296.0,1,-nbitq), 
to_sfixed(-159472284.0/4294967296.0,1,-nbitq), 
to_sfixed(217082048.0/4294967296.0,1,-nbitq), 
to_sfixed(134628082.0/4294967296.0,1,-nbitq), 
to_sfixed(-176252203.0/4294967296.0,1,-nbitq), 
to_sfixed(-88188237.0/4294967296.0,1,-nbitq), 
to_sfixed(274625154.0/4294967296.0,1,-nbitq), 
to_sfixed(-95236599.0/4294967296.0,1,-nbitq), 
to_sfixed(133729551.0/4294967296.0,1,-nbitq), 
to_sfixed(277479155.0/4294967296.0,1,-nbitq), 
to_sfixed(-190262385.0/4294967296.0,1,-nbitq), 
to_sfixed(-193722374.0/4294967296.0,1,-nbitq), 
to_sfixed(-468933597.0/4294967296.0,1,-nbitq), 
to_sfixed(-210469398.0/4294967296.0,1,-nbitq), 
to_sfixed(44324529.0/4294967296.0,1,-nbitq), 
to_sfixed(-350626106.0/4294967296.0,1,-nbitq), 
to_sfixed(138195753.0/4294967296.0,1,-nbitq), 
to_sfixed(-183605414.0/4294967296.0,1,-nbitq), 
to_sfixed(-161816778.0/4294967296.0,1,-nbitq), 
to_sfixed(47780478.0/4294967296.0,1,-nbitq), 
to_sfixed(-395262473.0/4294967296.0,1,-nbitq), 
to_sfixed(197792294.0/4294967296.0,1,-nbitq), 
to_sfixed(386125957.0/4294967296.0,1,-nbitq), 
to_sfixed(-101939702.0/4294967296.0,1,-nbitq), 
to_sfixed(-209521277.0/4294967296.0,1,-nbitq), 
to_sfixed(287038358.0/4294967296.0,1,-nbitq), 
to_sfixed(102255003.0/4294967296.0,1,-nbitq), 
to_sfixed(322750817.0/4294967296.0,1,-nbitq), 
to_sfixed(-275636008.0/4294967296.0,1,-nbitq), 
to_sfixed(158914205.0/4294967296.0,1,-nbitq), 
to_sfixed(-247962705.0/4294967296.0,1,-nbitq), 
to_sfixed(457486303.0/4294967296.0,1,-nbitq), 
to_sfixed(-215754791.0/4294967296.0,1,-nbitq), 
to_sfixed(182917942.0/4294967296.0,1,-nbitq), 
to_sfixed(-291659008.0/4294967296.0,1,-nbitq), 
to_sfixed(-306865450.0/4294967296.0,1,-nbitq), 
to_sfixed(15416635.0/4294967296.0,1,-nbitq), 
to_sfixed(89306176.0/4294967296.0,1,-nbitq), 
to_sfixed(77770741.0/4294967296.0,1,-nbitq), 
to_sfixed(58964001.0/4294967296.0,1,-nbitq), 
to_sfixed(50482362.0/4294967296.0,1,-nbitq), 
to_sfixed(-231300667.0/4294967296.0,1,-nbitq), 
to_sfixed(-293179456.0/4294967296.0,1,-nbitq), 
to_sfixed(593363620.0/4294967296.0,1,-nbitq), 
to_sfixed(-278083453.0/4294967296.0,1,-nbitq), 
to_sfixed(-260654923.0/4294967296.0,1,-nbitq), 
to_sfixed(174805281.0/4294967296.0,1,-nbitq), 
to_sfixed(-406329797.0/4294967296.0,1,-nbitq), 
to_sfixed(-4457273.0/4294967296.0,1,-nbitq), 
to_sfixed(-12498893.0/4294967296.0,1,-nbitq), 
to_sfixed(-235754542.0/4294967296.0,1,-nbitq), 
to_sfixed(-87394393.0/4294967296.0,1,-nbitq), 
to_sfixed(-457149532.0/4294967296.0,1,-nbitq), 
to_sfixed(323433731.0/4294967296.0,1,-nbitq), 
to_sfixed(-305978139.0/4294967296.0,1,-nbitq), 
to_sfixed(99009416.0/4294967296.0,1,-nbitq), 
to_sfixed(249013519.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(245085150.0/4294967296.0,1,-nbitq), 
to_sfixed(117639385.0/4294967296.0,1,-nbitq), 
to_sfixed(308204012.0/4294967296.0,1,-nbitq), 
to_sfixed(-171436377.0/4294967296.0,1,-nbitq), 
to_sfixed(-136726400.0/4294967296.0,1,-nbitq), 
to_sfixed(176792990.0/4294967296.0,1,-nbitq), 
to_sfixed(26270903.0/4294967296.0,1,-nbitq), 
to_sfixed(259876695.0/4294967296.0,1,-nbitq), 
to_sfixed(-199601221.0/4294967296.0,1,-nbitq), 
to_sfixed(27882468.0/4294967296.0,1,-nbitq), 
to_sfixed(-788227.0/4294967296.0,1,-nbitq), 
to_sfixed(-350753850.0/4294967296.0,1,-nbitq), 
to_sfixed(-413803008.0/4294967296.0,1,-nbitq), 
to_sfixed(-8744427.0/4294967296.0,1,-nbitq), 
to_sfixed(-76133354.0/4294967296.0,1,-nbitq), 
to_sfixed(-267665474.0/4294967296.0,1,-nbitq), 
to_sfixed(355293053.0/4294967296.0,1,-nbitq), 
to_sfixed(-39300066.0/4294967296.0,1,-nbitq), 
to_sfixed(370690267.0/4294967296.0,1,-nbitq), 
to_sfixed(316709128.0/4294967296.0,1,-nbitq), 
to_sfixed(-329136900.0/4294967296.0,1,-nbitq), 
to_sfixed(496855744.0/4294967296.0,1,-nbitq), 
to_sfixed(82850192.0/4294967296.0,1,-nbitq), 
to_sfixed(42547037.0/4294967296.0,1,-nbitq), 
to_sfixed(198868661.0/4294967296.0,1,-nbitq), 
to_sfixed(477679882.0/4294967296.0,1,-nbitq), 
to_sfixed(192801239.0/4294967296.0,1,-nbitq), 
to_sfixed(-285201074.0/4294967296.0,1,-nbitq), 
to_sfixed(161457382.0/4294967296.0,1,-nbitq), 
to_sfixed(-67512617.0/4294967296.0,1,-nbitq), 
to_sfixed(-520924277.0/4294967296.0,1,-nbitq), 
to_sfixed(-101236682.0/4294967296.0,1,-nbitq), 
to_sfixed(158931546.0/4294967296.0,1,-nbitq), 
to_sfixed(-480753371.0/4294967296.0,1,-nbitq), 
to_sfixed(449320052.0/4294967296.0,1,-nbitq), 
to_sfixed(-13578706.0/4294967296.0,1,-nbitq), 
to_sfixed(-50021624.0/4294967296.0,1,-nbitq), 
to_sfixed(-345940693.0/4294967296.0,1,-nbitq), 
to_sfixed(-121398991.0/4294967296.0,1,-nbitq), 
to_sfixed(322126445.0/4294967296.0,1,-nbitq), 
to_sfixed(-156671019.0/4294967296.0,1,-nbitq), 
to_sfixed(312851546.0/4294967296.0,1,-nbitq), 
to_sfixed(-19486602.0/4294967296.0,1,-nbitq), 
to_sfixed(-64276724.0/4294967296.0,1,-nbitq), 
to_sfixed(597263856.0/4294967296.0,1,-nbitq), 
to_sfixed(354689283.0/4294967296.0,1,-nbitq), 
to_sfixed(-251419656.0/4294967296.0,1,-nbitq), 
to_sfixed(-387104125.0/4294967296.0,1,-nbitq), 
to_sfixed(-246114974.0/4294967296.0,1,-nbitq), 
to_sfixed(391199692.0/4294967296.0,1,-nbitq), 
to_sfixed(355115052.0/4294967296.0,1,-nbitq), 
to_sfixed(-366338986.0/4294967296.0,1,-nbitq), 
to_sfixed(-120815007.0/4294967296.0,1,-nbitq), 
to_sfixed(-298257659.0/4294967296.0,1,-nbitq), 
to_sfixed(214505249.0/4294967296.0,1,-nbitq), 
to_sfixed(-204391939.0/4294967296.0,1,-nbitq), 
to_sfixed(59264007.0/4294967296.0,1,-nbitq), 
to_sfixed(-550193796.0/4294967296.0,1,-nbitq), 
to_sfixed(-295388476.0/4294967296.0,1,-nbitq), 
to_sfixed(-166410687.0/4294967296.0,1,-nbitq), 
to_sfixed(-5066153.0/4294967296.0,1,-nbitq), 
to_sfixed(-417651254.0/4294967296.0,1,-nbitq), 
to_sfixed(-379305504.0/4294967296.0,1,-nbitq), 
to_sfixed(-342033508.0/4294967296.0,1,-nbitq), 
to_sfixed(7538925.0/4294967296.0,1,-nbitq), 
to_sfixed(-141551521.0/4294967296.0,1,-nbitq), 
to_sfixed(-11410331.0/4294967296.0,1,-nbitq), 
to_sfixed(285785491.0/4294967296.0,1,-nbitq), 
to_sfixed(-239796602.0/4294967296.0,1,-nbitq), 
to_sfixed(325102219.0/4294967296.0,1,-nbitq), 
to_sfixed(-345567174.0/4294967296.0,1,-nbitq), 
to_sfixed(223403573.0/4294967296.0,1,-nbitq), 
to_sfixed(-305737828.0/4294967296.0,1,-nbitq), 
to_sfixed(-139199511.0/4294967296.0,1,-nbitq), 
to_sfixed(-265068263.0/4294967296.0,1,-nbitq), 
to_sfixed(-470658291.0/4294967296.0,1,-nbitq), 
to_sfixed(-406164208.0/4294967296.0,1,-nbitq), 
to_sfixed(-468839194.0/4294967296.0,1,-nbitq), 
to_sfixed(-459059997.0/4294967296.0,1,-nbitq), 
to_sfixed(338929904.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-77197440.0/4294967296.0,1,-nbitq), 
to_sfixed(234582049.0/4294967296.0,1,-nbitq), 
to_sfixed(-128312964.0/4294967296.0,1,-nbitq), 
to_sfixed(-84214383.0/4294967296.0,1,-nbitq), 
to_sfixed(59775133.0/4294967296.0,1,-nbitq), 
to_sfixed(153298920.0/4294967296.0,1,-nbitq), 
to_sfixed(85727299.0/4294967296.0,1,-nbitq), 
to_sfixed(-274116919.0/4294967296.0,1,-nbitq), 
to_sfixed(-461930215.0/4294967296.0,1,-nbitq), 
to_sfixed(-115026042.0/4294967296.0,1,-nbitq), 
to_sfixed(164047062.0/4294967296.0,1,-nbitq), 
to_sfixed(153239540.0/4294967296.0,1,-nbitq), 
to_sfixed(-175229995.0/4294967296.0,1,-nbitq), 
to_sfixed(265482552.0/4294967296.0,1,-nbitq), 
to_sfixed(344223831.0/4294967296.0,1,-nbitq), 
to_sfixed(152521724.0/4294967296.0,1,-nbitq), 
to_sfixed(27627256.0/4294967296.0,1,-nbitq), 
to_sfixed(-283358327.0/4294967296.0,1,-nbitq), 
to_sfixed(212658133.0/4294967296.0,1,-nbitq), 
to_sfixed(-63462876.0/4294967296.0,1,-nbitq), 
to_sfixed(349379558.0/4294967296.0,1,-nbitq), 
to_sfixed(20210655.0/4294967296.0,1,-nbitq), 
to_sfixed(745104976.0/4294967296.0,1,-nbitq), 
to_sfixed(58806813.0/4294967296.0,1,-nbitq), 
to_sfixed(2582775.0/4294967296.0,1,-nbitq), 
to_sfixed(20351257.0/4294967296.0,1,-nbitq), 
to_sfixed(24445796.0/4294967296.0,1,-nbitq), 
to_sfixed(-291824626.0/4294967296.0,1,-nbitq), 
to_sfixed(228374876.0/4294967296.0,1,-nbitq), 
to_sfixed(-521266891.0/4294967296.0,1,-nbitq), 
to_sfixed(55097318.0/4294967296.0,1,-nbitq), 
to_sfixed(-29285304.0/4294967296.0,1,-nbitq), 
to_sfixed(-58430442.0/4294967296.0,1,-nbitq), 
to_sfixed(148692851.0/4294967296.0,1,-nbitq), 
to_sfixed(230828306.0/4294967296.0,1,-nbitq), 
to_sfixed(-673384757.0/4294967296.0,1,-nbitq), 
to_sfixed(-118694480.0/4294967296.0,1,-nbitq), 
to_sfixed(-198294641.0/4294967296.0,1,-nbitq), 
to_sfixed(245260001.0/4294967296.0,1,-nbitq), 
to_sfixed(50545813.0/4294967296.0,1,-nbitq), 
to_sfixed(-384136261.0/4294967296.0,1,-nbitq), 
to_sfixed(-125980447.0/4294967296.0,1,-nbitq), 
to_sfixed(-180432236.0/4294967296.0,1,-nbitq), 
to_sfixed(320129751.0/4294967296.0,1,-nbitq), 
to_sfixed(340650399.0/4294967296.0,1,-nbitq), 
to_sfixed(-245587650.0/4294967296.0,1,-nbitq), 
to_sfixed(231052109.0/4294967296.0,1,-nbitq), 
to_sfixed(315088216.0/4294967296.0,1,-nbitq), 
to_sfixed(-305504255.0/4294967296.0,1,-nbitq), 
to_sfixed(277531622.0/4294967296.0,1,-nbitq), 
to_sfixed(-227901668.0/4294967296.0,1,-nbitq), 
to_sfixed(189160171.0/4294967296.0,1,-nbitq), 
to_sfixed(-374540176.0/4294967296.0,1,-nbitq), 
to_sfixed(-127265285.0/4294967296.0,1,-nbitq), 
to_sfixed(-304734569.0/4294967296.0,1,-nbitq), 
to_sfixed(-2410891.0/4294967296.0,1,-nbitq), 
to_sfixed(71876221.0/4294967296.0,1,-nbitq), 
to_sfixed(-236234083.0/4294967296.0,1,-nbitq), 
to_sfixed(-153307035.0/4294967296.0,1,-nbitq), 
to_sfixed(201916441.0/4294967296.0,1,-nbitq), 
to_sfixed(116707802.0/4294967296.0,1,-nbitq), 
to_sfixed(49545987.0/4294967296.0,1,-nbitq), 
to_sfixed(191398812.0/4294967296.0,1,-nbitq), 
to_sfixed(70006698.0/4294967296.0,1,-nbitq), 
to_sfixed(124296851.0/4294967296.0,1,-nbitq), 
to_sfixed(-396729293.0/4294967296.0,1,-nbitq), 
to_sfixed(594051611.0/4294967296.0,1,-nbitq), 
to_sfixed(-105427080.0/4294967296.0,1,-nbitq), 
to_sfixed(312680404.0/4294967296.0,1,-nbitq), 
to_sfixed(19986086.0/4294967296.0,1,-nbitq), 
to_sfixed(-406225961.0/4294967296.0,1,-nbitq), 
to_sfixed(-98511398.0/4294967296.0,1,-nbitq), 
to_sfixed(-65858580.0/4294967296.0,1,-nbitq), 
to_sfixed(-99375829.0/4294967296.0,1,-nbitq), 
to_sfixed(107826062.0/4294967296.0,1,-nbitq), 
to_sfixed(-138958248.0/4294967296.0,1,-nbitq), 
to_sfixed(-157151127.0/4294967296.0,1,-nbitq), 
to_sfixed(-425457139.0/4294967296.0,1,-nbitq), 
to_sfixed(-81007617.0/4294967296.0,1,-nbitq), 
to_sfixed(-224838218.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-183585160.0/4294967296.0,1,-nbitq), 
to_sfixed(-183759712.0/4294967296.0,1,-nbitq), 
to_sfixed(158320811.0/4294967296.0,1,-nbitq), 
to_sfixed(430180517.0/4294967296.0,1,-nbitq), 
to_sfixed(312848181.0/4294967296.0,1,-nbitq), 
to_sfixed(18085342.0/4294967296.0,1,-nbitq), 
to_sfixed(378632303.0/4294967296.0,1,-nbitq), 
to_sfixed(-360931784.0/4294967296.0,1,-nbitq), 
to_sfixed(-298844115.0/4294967296.0,1,-nbitq), 
to_sfixed(-109564910.0/4294967296.0,1,-nbitq), 
to_sfixed(-169960040.0/4294967296.0,1,-nbitq), 
to_sfixed(-153238430.0/4294967296.0,1,-nbitq), 
to_sfixed(-493987657.0/4294967296.0,1,-nbitq), 
to_sfixed(-125655032.0/4294967296.0,1,-nbitq), 
to_sfixed(93621058.0/4294967296.0,1,-nbitq), 
to_sfixed(63827756.0/4294967296.0,1,-nbitq), 
to_sfixed(-384132046.0/4294967296.0,1,-nbitq), 
to_sfixed(-9627527.0/4294967296.0,1,-nbitq), 
to_sfixed(371007752.0/4294967296.0,1,-nbitq), 
to_sfixed(231649128.0/4294967296.0,1,-nbitq), 
to_sfixed(-212298512.0/4294967296.0,1,-nbitq), 
to_sfixed(267085979.0/4294967296.0,1,-nbitq), 
to_sfixed(188112941.0/4294967296.0,1,-nbitq), 
to_sfixed(313256964.0/4294967296.0,1,-nbitq), 
to_sfixed(172169143.0/4294967296.0,1,-nbitq), 
to_sfixed(328428495.0/4294967296.0,1,-nbitq), 
to_sfixed(105305674.0/4294967296.0,1,-nbitq), 
to_sfixed(-148199163.0/4294967296.0,1,-nbitq), 
to_sfixed(-12671387.0/4294967296.0,1,-nbitq), 
to_sfixed(-215637314.0/4294967296.0,1,-nbitq), 
to_sfixed(-421659905.0/4294967296.0,1,-nbitq), 
to_sfixed(-84380644.0/4294967296.0,1,-nbitq), 
to_sfixed(307127944.0/4294967296.0,1,-nbitq), 
to_sfixed(-349944414.0/4294967296.0,1,-nbitq), 
to_sfixed(512798392.0/4294967296.0,1,-nbitq), 
to_sfixed(-188097448.0/4294967296.0,1,-nbitq), 
to_sfixed(-243838158.0/4294967296.0,1,-nbitq), 
to_sfixed(-240190184.0/4294967296.0,1,-nbitq), 
to_sfixed(59564060.0/4294967296.0,1,-nbitq), 
to_sfixed(172886615.0/4294967296.0,1,-nbitq), 
to_sfixed(-255235079.0/4294967296.0,1,-nbitq), 
to_sfixed(-119128740.0/4294967296.0,1,-nbitq), 
to_sfixed(-304729927.0/4294967296.0,1,-nbitq), 
to_sfixed(139878665.0/4294967296.0,1,-nbitq), 
to_sfixed(721989477.0/4294967296.0,1,-nbitq), 
to_sfixed(92245741.0/4294967296.0,1,-nbitq), 
to_sfixed(-155546271.0/4294967296.0,1,-nbitq), 
to_sfixed(-378899798.0/4294967296.0,1,-nbitq), 
to_sfixed(-181369284.0/4294967296.0,1,-nbitq), 
to_sfixed(-280665907.0/4294967296.0,1,-nbitq), 
to_sfixed(152192333.0/4294967296.0,1,-nbitq), 
to_sfixed(502050443.0/4294967296.0,1,-nbitq), 
to_sfixed(-231407514.0/4294967296.0,1,-nbitq), 
to_sfixed(-751066.0/4294967296.0,1,-nbitq), 
to_sfixed(191534544.0/4294967296.0,1,-nbitq), 
to_sfixed(-67326895.0/4294967296.0,1,-nbitq), 
to_sfixed(-75110766.0/4294967296.0,1,-nbitq), 
to_sfixed(170647949.0/4294967296.0,1,-nbitq), 
to_sfixed(143918069.0/4294967296.0,1,-nbitq), 
to_sfixed(395130992.0/4294967296.0,1,-nbitq), 
to_sfixed(-301563849.0/4294967296.0,1,-nbitq), 
to_sfixed(-443862076.0/4294967296.0,1,-nbitq), 
to_sfixed(-80501711.0/4294967296.0,1,-nbitq), 
to_sfixed(-209592897.0/4294967296.0,1,-nbitq), 
to_sfixed(350498620.0/4294967296.0,1,-nbitq), 
to_sfixed(-5021187.0/4294967296.0,1,-nbitq), 
to_sfixed(122516610.0/4294967296.0,1,-nbitq), 
to_sfixed(211541498.0/4294967296.0,1,-nbitq), 
to_sfixed(-247410142.0/4294967296.0,1,-nbitq), 
to_sfixed(-187248831.0/4294967296.0,1,-nbitq), 
to_sfixed(244647290.0/4294967296.0,1,-nbitq), 
to_sfixed(312137898.0/4294967296.0,1,-nbitq), 
to_sfixed(-263576035.0/4294967296.0,1,-nbitq), 
to_sfixed(440936475.0/4294967296.0,1,-nbitq), 
to_sfixed(-49285880.0/4294967296.0,1,-nbitq), 
to_sfixed(-476389840.0/4294967296.0,1,-nbitq), 
to_sfixed(-307967478.0/4294967296.0,1,-nbitq), 
to_sfixed(-513552735.0/4294967296.0,1,-nbitq), 
to_sfixed(-294455900.0/4294967296.0,1,-nbitq), 
to_sfixed(108617225.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(130607458.0/4294967296.0,1,-nbitq), 
to_sfixed(-342521274.0/4294967296.0,1,-nbitq), 
to_sfixed(110059838.0/4294967296.0,1,-nbitq), 
to_sfixed(-292613756.0/4294967296.0,1,-nbitq), 
to_sfixed(-183237872.0/4294967296.0,1,-nbitq), 
to_sfixed(-483977247.0/4294967296.0,1,-nbitq), 
to_sfixed(-295899117.0/4294967296.0,1,-nbitq), 
to_sfixed(135184371.0/4294967296.0,1,-nbitq), 
to_sfixed(-262379227.0/4294967296.0,1,-nbitq), 
to_sfixed(-306897651.0/4294967296.0,1,-nbitq), 
to_sfixed(344250424.0/4294967296.0,1,-nbitq), 
to_sfixed(219574244.0/4294967296.0,1,-nbitq), 
to_sfixed(-301892595.0/4294967296.0,1,-nbitq), 
to_sfixed(104454138.0/4294967296.0,1,-nbitq), 
to_sfixed(373196812.0/4294967296.0,1,-nbitq), 
to_sfixed(-200294238.0/4294967296.0,1,-nbitq), 
to_sfixed(-133883720.0/4294967296.0,1,-nbitq), 
to_sfixed(296505842.0/4294967296.0,1,-nbitq), 
to_sfixed(358367024.0/4294967296.0,1,-nbitq), 
to_sfixed(336468636.0/4294967296.0,1,-nbitq), 
to_sfixed(87471885.0/4294967296.0,1,-nbitq), 
to_sfixed(431909920.0/4294967296.0,1,-nbitq), 
to_sfixed(479051331.0/4294967296.0,1,-nbitq), 
to_sfixed(204168335.0/4294967296.0,1,-nbitq), 
to_sfixed(426110400.0/4294967296.0,1,-nbitq), 
to_sfixed(446979523.0/4294967296.0,1,-nbitq), 
to_sfixed(388840863.0/4294967296.0,1,-nbitq), 
to_sfixed(-421435475.0/4294967296.0,1,-nbitq), 
to_sfixed(-282914153.0/4294967296.0,1,-nbitq), 
to_sfixed(210312865.0/4294967296.0,1,-nbitq), 
to_sfixed(181266051.0/4294967296.0,1,-nbitq), 
to_sfixed(-161594758.0/4294967296.0,1,-nbitq), 
to_sfixed(296369678.0/4294967296.0,1,-nbitq), 
to_sfixed(199043945.0/4294967296.0,1,-nbitq), 
to_sfixed(270050169.0/4294967296.0,1,-nbitq), 
to_sfixed(-535687333.0/4294967296.0,1,-nbitq), 
to_sfixed(362667217.0/4294967296.0,1,-nbitq), 
to_sfixed(-287335043.0/4294967296.0,1,-nbitq), 
to_sfixed(130022710.0/4294967296.0,1,-nbitq), 
to_sfixed(242801774.0/4294967296.0,1,-nbitq), 
to_sfixed(64697749.0/4294967296.0,1,-nbitq), 
to_sfixed(533558886.0/4294967296.0,1,-nbitq), 
to_sfixed(214433160.0/4294967296.0,1,-nbitq), 
to_sfixed(-292362225.0/4294967296.0,1,-nbitq), 
to_sfixed(224893966.0/4294967296.0,1,-nbitq), 
to_sfixed(506899781.0/4294967296.0,1,-nbitq), 
to_sfixed(310999255.0/4294967296.0,1,-nbitq), 
to_sfixed(-221132205.0/4294967296.0,1,-nbitq), 
to_sfixed(1005912.0/4294967296.0,1,-nbitq), 
to_sfixed(259688094.0/4294967296.0,1,-nbitq), 
to_sfixed(-266877292.0/4294967296.0,1,-nbitq), 
to_sfixed(-217519588.0/4294967296.0,1,-nbitq), 
to_sfixed(-276091692.0/4294967296.0,1,-nbitq), 
to_sfixed(-77468120.0/4294967296.0,1,-nbitq), 
to_sfixed(-95607264.0/4294967296.0,1,-nbitq), 
to_sfixed(79640540.0/4294967296.0,1,-nbitq), 
to_sfixed(-236392629.0/4294967296.0,1,-nbitq), 
to_sfixed(-138732099.0/4294967296.0,1,-nbitq), 
to_sfixed(-197673325.0/4294967296.0,1,-nbitq), 
to_sfixed(-48528571.0/4294967296.0,1,-nbitq), 
to_sfixed(93868917.0/4294967296.0,1,-nbitq), 
to_sfixed(-190677456.0/4294967296.0,1,-nbitq), 
to_sfixed(-331653227.0/4294967296.0,1,-nbitq), 
to_sfixed(-47268857.0/4294967296.0,1,-nbitq), 
to_sfixed(-106956823.0/4294967296.0,1,-nbitq), 
to_sfixed(-252690982.0/4294967296.0,1,-nbitq), 
to_sfixed(487323007.0/4294967296.0,1,-nbitq), 
to_sfixed(-254415410.0/4294967296.0,1,-nbitq), 
to_sfixed(-70195653.0/4294967296.0,1,-nbitq), 
to_sfixed(363004308.0/4294967296.0,1,-nbitq), 
to_sfixed(243692737.0/4294967296.0,1,-nbitq), 
to_sfixed(-223234065.0/4294967296.0,1,-nbitq), 
to_sfixed(-298078866.0/4294967296.0,1,-nbitq), 
to_sfixed(336593632.0/4294967296.0,1,-nbitq), 
to_sfixed(6883937.0/4294967296.0,1,-nbitq), 
to_sfixed(-516044320.0/4294967296.0,1,-nbitq), 
to_sfixed(333434419.0/4294967296.0,1,-nbitq), 
to_sfixed(-212913453.0/4294967296.0,1,-nbitq), 
to_sfixed(-386901674.0/4294967296.0,1,-nbitq), 
to_sfixed(-342094363.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-375734447.0/4294967296.0,1,-nbitq), 
to_sfixed(-454516792.0/4294967296.0,1,-nbitq), 
to_sfixed(128385047.0/4294967296.0,1,-nbitq), 
to_sfixed(10162550.0/4294967296.0,1,-nbitq), 
to_sfixed(-164645698.0/4294967296.0,1,-nbitq), 
to_sfixed(-115004681.0/4294967296.0,1,-nbitq), 
to_sfixed(148294196.0/4294967296.0,1,-nbitq), 
to_sfixed(107428954.0/4294967296.0,1,-nbitq), 
to_sfixed(346357805.0/4294967296.0,1,-nbitq), 
to_sfixed(140795994.0/4294967296.0,1,-nbitq), 
to_sfixed(242170229.0/4294967296.0,1,-nbitq), 
to_sfixed(444085370.0/4294967296.0,1,-nbitq), 
to_sfixed(-112118562.0/4294967296.0,1,-nbitq), 
to_sfixed(54902721.0/4294967296.0,1,-nbitq), 
to_sfixed(-169556115.0/4294967296.0,1,-nbitq), 
to_sfixed(-141243122.0/4294967296.0,1,-nbitq), 
to_sfixed(271093770.0/4294967296.0,1,-nbitq), 
to_sfixed(346703585.0/4294967296.0,1,-nbitq), 
to_sfixed(342140193.0/4294967296.0,1,-nbitq), 
to_sfixed(-333154469.0/4294967296.0,1,-nbitq), 
to_sfixed(-11182617.0/4294967296.0,1,-nbitq), 
to_sfixed(-217385533.0/4294967296.0,1,-nbitq), 
to_sfixed(797194824.0/4294967296.0,1,-nbitq), 
to_sfixed(-474735806.0/4294967296.0,1,-nbitq), 
to_sfixed(295646244.0/4294967296.0,1,-nbitq), 
to_sfixed(244478358.0/4294967296.0,1,-nbitq), 
to_sfixed(-85015928.0/4294967296.0,1,-nbitq), 
to_sfixed(-128130179.0/4294967296.0,1,-nbitq), 
to_sfixed(-163355661.0/4294967296.0,1,-nbitq), 
to_sfixed(-470305103.0/4294967296.0,1,-nbitq), 
to_sfixed(-593212118.0/4294967296.0,1,-nbitq), 
to_sfixed(-577122277.0/4294967296.0,1,-nbitq), 
to_sfixed(213081304.0/4294967296.0,1,-nbitq), 
to_sfixed(-80947817.0/4294967296.0,1,-nbitq), 
to_sfixed(322593535.0/4294967296.0,1,-nbitq), 
to_sfixed(-126661919.0/4294967296.0,1,-nbitq), 
to_sfixed(406745483.0/4294967296.0,1,-nbitq), 
to_sfixed(-343319360.0/4294967296.0,1,-nbitq), 
to_sfixed(-174636676.0/4294967296.0,1,-nbitq), 
to_sfixed(-36331069.0/4294967296.0,1,-nbitq), 
to_sfixed(69585523.0/4294967296.0,1,-nbitq), 
to_sfixed(83411430.0/4294967296.0,1,-nbitq), 
to_sfixed(322956808.0/4294967296.0,1,-nbitq), 
to_sfixed(182853785.0/4294967296.0,1,-nbitq), 
to_sfixed(-253095512.0/4294967296.0,1,-nbitq), 
to_sfixed(102117079.0/4294967296.0,1,-nbitq), 
to_sfixed(-364720445.0/4294967296.0,1,-nbitq), 
to_sfixed(-128497443.0/4294967296.0,1,-nbitq), 
to_sfixed(-281633595.0/4294967296.0,1,-nbitq), 
to_sfixed(453676908.0/4294967296.0,1,-nbitq), 
to_sfixed(-354402483.0/4294967296.0,1,-nbitq), 
to_sfixed(50971198.0/4294967296.0,1,-nbitq), 
to_sfixed(-373963198.0/4294967296.0,1,-nbitq), 
to_sfixed(168361220.0/4294967296.0,1,-nbitq), 
to_sfixed(32869172.0/4294967296.0,1,-nbitq), 
to_sfixed(-434050182.0/4294967296.0,1,-nbitq), 
to_sfixed(108274368.0/4294967296.0,1,-nbitq), 
to_sfixed(-353080509.0/4294967296.0,1,-nbitq), 
to_sfixed(101597601.0/4294967296.0,1,-nbitq), 
to_sfixed(-158059709.0/4294967296.0,1,-nbitq), 
to_sfixed(77638679.0/4294967296.0,1,-nbitq), 
to_sfixed(-92093149.0/4294967296.0,1,-nbitq), 
to_sfixed(-329288184.0/4294967296.0,1,-nbitq), 
to_sfixed(-377705517.0/4294967296.0,1,-nbitq), 
to_sfixed(293080054.0/4294967296.0,1,-nbitq), 
to_sfixed(158263811.0/4294967296.0,1,-nbitq), 
to_sfixed(651732587.0/4294967296.0,1,-nbitq), 
to_sfixed(-314356447.0/4294967296.0,1,-nbitq), 
to_sfixed(-273430453.0/4294967296.0,1,-nbitq), 
to_sfixed(59103254.0/4294967296.0,1,-nbitq), 
to_sfixed(-90955198.0/4294967296.0,1,-nbitq), 
to_sfixed(295632973.0/4294967296.0,1,-nbitq), 
to_sfixed(-368047907.0/4294967296.0,1,-nbitq), 
to_sfixed(47934528.0/4294967296.0,1,-nbitq), 
to_sfixed(215975598.0/4294967296.0,1,-nbitq), 
to_sfixed(-495210738.0/4294967296.0,1,-nbitq), 
to_sfixed(-336720810.0/4294967296.0,1,-nbitq), 
to_sfixed(-385833369.0/4294967296.0,1,-nbitq), 
to_sfixed(270915679.0/4294967296.0,1,-nbitq), 
to_sfixed(205581418.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-106734096.0/4294967296.0,1,-nbitq), 
to_sfixed(-30069772.0/4294967296.0,1,-nbitq), 
to_sfixed(-336313040.0/4294967296.0,1,-nbitq), 
to_sfixed(249721730.0/4294967296.0,1,-nbitq), 
to_sfixed(-35091023.0/4294967296.0,1,-nbitq), 
to_sfixed(309891784.0/4294967296.0,1,-nbitq), 
to_sfixed(-201391217.0/4294967296.0,1,-nbitq), 
to_sfixed(1004.0/4294967296.0,1,-nbitq), 
to_sfixed(-387550597.0/4294967296.0,1,-nbitq), 
to_sfixed(387856901.0/4294967296.0,1,-nbitq), 
to_sfixed(396455002.0/4294967296.0,1,-nbitq), 
to_sfixed(612394410.0/4294967296.0,1,-nbitq), 
to_sfixed(-505318182.0/4294967296.0,1,-nbitq), 
to_sfixed(140088314.0/4294967296.0,1,-nbitq), 
to_sfixed(413440917.0/4294967296.0,1,-nbitq), 
to_sfixed(-143742333.0/4294967296.0,1,-nbitq), 
to_sfixed(-97766296.0/4294967296.0,1,-nbitq), 
to_sfixed(-119066666.0/4294967296.0,1,-nbitq), 
to_sfixed(217354536.0/4294967296.0,1,-nbitq), 
to_sfixed(65627984.0/4294967296.0,1,-nbitq), 
to_sfixed(199952813.0/4294967296.0,1,-nbitq), 
to_sfixed(-10862538.0/4294967296.0,1,-nbitq), 
to_sfixed(130730990.0/4294967296.0,1,-nbitq), 
to_sfixed(-305635360.0/4294967296.0,1,-nbitq), 
to_sfixed(359960837.0/4294967296.0,1,-nbitq), 
to_sfixed(-89547480.0/4294967296.0,1,-nbitq), 
to_sfixed(63414335.0/4294967296.0,1,-nbitq), 
to_sfixed(-312694784.0/4294967296.0,1,-nbitq), 
to_sfixed(382782696.0/4294967296.0,1,-nbitq), 
to_sfixed(187516854.0/4294967296.0,1,-nbitq), 
to_sfixed(-491076012.0/4294967296.0,1,-nbitq), 
to_sfixed(-286245757.0/4294967296.0,1,-nbitq), 
to_sfixed(-29889243.0/4294967296.0,1,-nbitq), 
to_sfixed(-172981076.0/4294967296.0,1,-nbitq), 
to_sfixed(508686593.0/4294967296.0,1,-nbitq), 
to_sfixed(119057367.0/4294967296.0,1,-nbitq), 
to_sfixed(432674307.0/4294967296.0,1,-nbitq), 
to_sfixed(38507295.0/4294967296.0,1,-nbitq), 
to_sfixed(173731188.0/4294967296.0,1,-nbitq), 
to_sfixed(143808580.0/4294967296.0,1,-nbitq), 
to_sfixed(157128588.0/4294967296.0,1,-nbitq), 
to_sfixed(61093787.0/4294967296.0,1,-nbitq), 
to_sfixed(-46509276.0/4294967296.0,1,-nbitq), 
to_sfixed(-426748447.0/4294967296.0,1,-nbitq), 
to_sfixed(-502595701.0/4294967296.0,1,-nbitq), 
to_sfixed(-123173750.0/4294967296.0,1,-nbitq), 
to_sfixed(215752221.0/4294967296.0,1,-nbitq), 
to_sfixed(56454461.0/4294967296.0,1,-nbitq), 
to_sfixed(14132891.0/4294967296.0,1,-nbitq), 
to_sfixed(510878485.0/4294967296.0,1,-nbitq), 
to_sfixed(-108459280.0/4294967296.0,1,-nbitq), 
to_sfixed(111829028.0/4294967296.0,1,-nbitq), 
to_sfixed(-458131165.0/4294967296.0,1,-nbitq), 
to_sfixed(-40669391.0/4294967296.0,1,-nbitq), 
to_sfixed(365725219.0/4294967296.0,1,-nbitq), 
to_sfixed(-299414005.0/4294967296.0,1,-nbitq), 
to_sfixed(13564382.0/4294967296.0,1,-nbitq), 
to_sfixed(-32459080.0/4294967296.0,1,-nbitq), 
to_sfixed(140617711.0/4294967296.0,1,-nbitq), 
to_sfixed(315245332.0/4294967296.0,1,-nbitq), 
to_sfixed(-331942392.0/4294967296.0,1,-nbitq), 
to_sfixed(226969005.0/4294967296.0,1,-nbitq), 
to_sfixed(-268066163.0/4294967296.0,1,-nbitq), 
to_sfixed(79207929.0/4294967296.0,1,-nbitq), 
to_sfixed(412039789.0/4294967296.0,1,-nbitq), 
to_sfixed(-467637566.0/4294967296.0,1,-nbitq), 
to_sfixed(198627631.0/4294967296.0,1,-nbitq), 
to_sfixed(-195221504.0/4294967296.0,1,-nbitq), 
to_sfixed(256272367.0/4294967296.0,1,-nbitq), 
to_sfixed(-256146408.0/4294967296.0,1,-nbitq), 
to_sfixed(-427039625.0/4294967296.0,1,-nbitq), 
to_sfixed(250263103.0/4294967296.0,1,-nbitq), 
to_sfixed(-43423342.0/4294967296.0,1,-nbitq), 
to_sfixed(389366462.0/4294967296.0,1,-nbitq), 
to_sfixed(-154562899.0/4294967296.0,1,-nbitq), 
to_sfixed(-80812102.0/4294967296.0,1,-nbitq), 
to_sfixed(-131628610.0/4294967296.0,1,-nbitq), 
to_sfixed(212022108.0/4294967296.0,1,-nbitq), 
to_sfixed(297827781.0/4294967296.0,1,-nbitq), 
to_sfixed(-101287571.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-389130045.0/4294967296.0,1,-nbitq), 
to_sfixed(-129427411.0/4294967296.0,1,-nbitq), 
to_sfixed(294392763.0/4294967296.0,1,-nbitq), 
to_sfixed(180872447.0/4294967296.0,1,-nbitq), 
to_sfixed(325684881.0/4294967296.0,1,-nbitq), 
to_sfixed(-32773512.0/4294967296.0,1,-nbitq), 
to_sfixed(362253674.0/4294967296.0,1,-nbitq), 
to_sfixed(-425893116.0/4294967296.0,1,-nbitq), 
to_sfixed(-41146228.0/4294967296.0,1,-nbitq), 
to_sfixed(-145582102.0/4294967296.0,1,-nbitq), 
to_sfixed(-349288212.0/4294967296.0,1,-nbitq), 
to_sfixed(272030199.0/4294967296.0,1,-nbitq), 
to_sfixed(-38968963.0/4294967296.0,1,-nbitq), 
to_sfixed(-197795532.0/4294967296.0,1,-nbitq), 
to_sfixed(-251683871.0/4294967296.0,1,-nbitq), 
to_sfixed(250957813.0/4294967296.0,1,-nbitq), 
to_sfixed(-94590392.0/4294967296.0,1,-nbitq), 
to_sfixed(187926960.0/4294967296.0,1,-nbitq), 
to_sfixed(316557749.0/4294967296.0,1,-nbitq), 
to_sfixed(45728356.0/4294967296.0,1,-nbitq), 
to_sfixed(-208285577.0/4294967296.0,1,-nbitq), 
to_sfixed(-147761559.0/4294967296.0,1,-nbitq), 
to_sfixed(38149328.0/4294967296.0,1,-nbitq), 
to_sfixed(166712144.0/4294967296.0,1,-nbitq), 
to_sfixed(-306690748.0/4294967296.0,1,-nbitq), 
to_sfixed(-526700647.0/4294967296.0,1,-nbitq), 
to_sfixed(171009641.0/4294967296.0,1,-nbitq), 
to_sfixed(-324747281.0/4294967296.0,1,-nbitq), 
to_sfixed(152905195.0/4294967296.0,1,-nbitq), 
to_sfixed(-210548187.0/4294967296.0,1,-nbitq), 
to_sfixed(-193558802.0/4294967296.0,1,-nbitq), 
to_sfixed(-207319152.0/4294967296.0,1,-nbitq), 
to_sfixed(-205951399.0/4294967296.0,1,-nbitq), 
to_sfixed(273075141.0/4294967296.0,1,-nbitq), 
to_sfixed(5564210.0/4294967296.0,1,-nbitq), 
to_sfixed(342930665.0/4294967296.0,1,-nbitq), 
to_sfixed(149744232.0/4294967296.0,1,-nbitq), 
to_sfixed(379332974.0/4294967296.0,1,-nbitq), 
to_sfixed(404147756.0/4294967296.0,1,-nbitq), 
to_sfixed(-160131361.0/4294967296.0,1,-nbitq), 
to_sfixed(675615.0/4294967296.0,1,-nbitq), 
to_sfixed(556022945.0/4294967296.0,1,-nbitq), 
to_sfixed(-124386347.0/4294967296.0,1,-nbitq), 
to_sfixed(142787344.0/4294967296.0,1,-nbitq), 
to_sfixed(-17135219.0/4294967296.0,1,-nbitq), 
to_sfixed(195864090.0/4294967296.0,1,-nbitq), 
to_sfixed(-117933411.0/4294967296.0,1,-nbitq), 
to_sfixed(-427366702.0/4294967296.0,1,-nbitq), 
to_sfixed(99921961.0/4294967296.0,1,-nbitq), 
to_sfixed(499044684.0/4294967296.0,1,-nbitq), 
to_sfixed(301385287.0/4294967296.0,1,-nbitq), 
to_sfixed(-18763252.0/4294967296.0,1,-nbitq), 
to_sfixed(302440692.0/4294967296.0,1,-nbitq), 
to_sfixed(-322750220.0/4294967296.0,1,-nbitq), 
to_sfixed(24891609.0/4294967296.0,1,-nbitq), 
to_sfixed(158774467.0/4294967296.0,1,-nbitq), 
to_sfixed(402548972.0/4294967296.0,1,-nbitq), 
to_sfixed(20253457.0/4294967296.0,1,-nbitq), 
to_sfixed(434200938.0/4294967296.0,1,-nbitq), 
to_sfixed(-316102148.0/4294967296.0,1,-nbitq), 
to_sfixed(103492497.0/4294967296.0,1,-nbitq), 
to_sfixed(336284698.0/4294967296.0,1,-nbitq), 
to_sfixed(-21333345.0/4294967296.0,1,-nbitq), 
to_sfixed(-115381601.0/4294967296.0,1,-nbitq), 
to_sfixed(-303807731.0/4294967296.0,1,-nbitq), 
to_sfixed(227062914.0/4294967296.0,1,-nbitq), 
to_sfixed(616077748.0/4294967296.0,1,-nbitq), 
to_sfixed(-433303571.0/4294967296.0,1,-nbitq), 
to_sfixed(222485307.0/4294967296.0,1,-nbitq), 
to_sfixed(228234189.0/4294967296.0,1,-nbitq), 
to_sfixed(256482520.0/4294967296.0,1,-nbitq), 
to_sfixed(-200238882.0/4294967296.0,1,-nbitq), 
to_sfixed(70624289.0/4294967296.0,1,-nbitq), 
to_sfixed(379163908.0/4294967296.0,1,-nbitq), 
to_sfixed(12709905.0/4294967296.0,1,-nbitq), 
to_sfixed(-54135211.0/4294967296.0,1,-nbitq), 
to_sfixed(-214234478.0/4294967296.0,1,-nbitq), 
to_sfixed(-281327551.0/4294967296.0,1,-nbitq), 
to_sfixed(-29667190.0/4294967296.0,1,-nbitq), 
to_sfixed(-343192930.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(350600423.0/4294967296.0,1,-nbitq), 
to_sfixed(-89534334.0/4294967296.0,1,-nbitq), 
to_sfixed(-268086494.0/4294967296.0,1,-nbitq), 
to_sfixed(-233779932.0/4294967296.0,1,-nbitq), 
to_sfixed(198978658.0/4294967296.0,1,-nbitq), 
to_sfixed(-521531538.0/4294967296.0,1,-nbitq), 
to_sfixed(163323269.0/4294967296.0,1,-nbitq), 
to_sfixed(-227477291.0/4294967296.0,1,-nbitq), 
to_sfixed(-292730522.0/4294967296.0,1,-nbitq), 
to_sfixed(-103799882.0/4294967296.0,1,-nbitq), 
to_sfixed(-293712407.0/4294967296.0,1,-nbitq), 
to_sfixed(126254077.0/4294967296.0,1,-nbitq), 
to_sfixed(-130928650.0/4294967296.0,1,-nbitq), 
to_sfixed(139991027.0/4294967296.0,1,-nbitq), 
to_sfixed(46172136.0/4294967296.0,1,-nbitq), 
to_sfixed(-88843166.0/4294967296.0,1,-nbitq), 
to_sfixed(-419907880.0/4294967296.0,1,-nbitq), 
to_sfixed(327631213.0/4294967296.0,1,-nbitq), 
to_sfixed(15038543.0/4294967296.0,1,-nbitq), 
to_sfixed(-149984543.0/4294967296.0,1,-nbitq), 
to_sfixed(-386947727.0/4294967296.0,1,-nbitq), 
to_sfixed(427679286.0/4294967296.0,1,-nbitq), 
to_sfixed(426797866.0/4294967296.0,1,-nbitq), 
to_sfixed(231211571.0/4294967296.0,1,-nbitq), 
to_sfixed(281984846.0/4294967296.0,1,-nbitq), 
to_sfixed(-20889355.0/4294967296.0,1,-nbitq), 
to_sfixed(-86894883.0/4294967296.0,1,-nbitq), 
to_sfixed(-434879264.0/4294967296.0,1,-nbitq), 
to_sfixed(306595888.0/4294967296.0,1,-nbitq), 
to_sfixed(41685411.0/4294967296.0,1,-nbitq), 
to_sfixed(-497821958.0/4294967296.0,1,-nbitq), 
to_sfixed(-524333425.0/4294967296.0,1,-nbitq), 
to_sfixed(536566780.0/4294967296.0,1,-nbitq), 
to_sfixed(45703398.0/4294967296.0,1,-nbitq), 
to_sfixed(499953302.0/4294967296.0,1,-nbitq), 
to_sfixed(51041150.0/4294967296.0,1,-nbitq), 
to_sfixed(410568439.0/4294967296.0,1,-nbitq), 
to_sfixed(191779183.0/4294967296.0,1,-nbitq), 
to_sfixed(111495450.0/4294967296.0,1,-nbitq), 
to_sfixed(205293656.0/4294967296.0,1,-nbitq), 
to_sfixed(15435673.0/4294967296.0,1,-nbitq), 
to_sfixed(99902776.0/4294967296.0,1,-nbitq), 
to_sfixed(371834608.0/4294967296.0,1,-nbitq), 
to_sfixed(-322812721.0/4294967296.0,1,-nbitq), 
to_sfixed(-289559745.0/4294967296.0,1,-nbitq), 
to_sfixed(-84068017.0/4294967296.0,1,-nbitq), 
to_sfixed(-56481302.0/4294967296.0,1,-nbitq), 
to_sfixed(52607837.0/4294967296.0,1,-nbitq), 
to_sfixed(-187010814.0/4294967296.0,1,-nbitq), 
to_sfixed(-206739964.0/4294967296.0,1,-nbitq), 
to_sfixed(79551514.0/4294967296.0,1,-nbitq), 
to_sfixed(6028031.0/4294967296.0,1,-nbitq), 
to_sfixed(-309089882.0/4294967296.0,1,-nbitq), 
to_sfixed(-299067539.0/4294967296.0,1,-nbitq), 
to_sfixed(217363830.0/4294967296.0,1,-nbitq), 
to_sfixed(158081937.0/4294967296.0,1,-nbitq), 
to_sfixed(-244535391.0/4294967296.0,1,-nbitq), 
to_sfixed(139776578.0/4294967296.0,1,-nbitq), 
to_sfixed(-9830643.0/4294967296.0,1,-nbitq), 
to_sfixed(256503343.0/4294967296.0,1,-nbitq), 
to_sfixed(-163744742.0/4294967296.0,1,-nbitq), 
to_sfixed(227265653.0/4294967296.0,1,-nbitq), 
to_sfixed(402378471.0/4294967296.0,1,-nbitq), 
to_sfixed(-179488627.0/4294967296.0,1,-nbitq), 
to_sfixed(119755954.0/4294967296.0,1,-nbitq), 
to_sfixed(213832528.0/4294967296.0,1,-nbitq), 
to_sfixed(669762974.0/4294967296.0,1,-nbitq), 
to_sfixed(-389541964.0/4294967296.0,1,-nbitq), 
to_sfixed(92524406.0/4294967296.0,1,-nbitq), 
to_sfixed(173969922.0/4294967296.0,1,-nbitq), 
to_sfixed(-263330071.0/4294967296.0,1,-nbitq), 
to_sfixed(266364517.0/4294967296.0,1,-nbitq), 
to_sfixed(184246722.0/4294967296.0,1,-nbitq), 
to_sfixed(389430569.0/4294967296.0,1,-nbitq), 
to_sfixed(85240173.0/4294967296.0,1,-nbitq), 
to_sfixed(189424525.0/4294967296.0,1,-nbitq), 
to_sfixed(-426854465.0/4294967296.0,1,-nbitq), 
to_sfixed(263735679.0/4294967296.0,1,-nbitq), 
to_sfixed(359502191.0/4294967296.0,1,-nbitq), 
to_sfixed(147621202.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(191114402.0/4294967296.0,1,-nbitq), 
to_sfixed(-417546417.0/4294967296.0,1,-nbitq), 
to_sfixed(-44320642.0/4294967296.0,1,-nbitq), 
to_sfixed(-354721104.0/4294967296.0,1,-nbitq), 
to_sfixed(6375924.0/4294967296.0,1,-nbitq), 
to_sfixed(-60158679.0/4294967296.0,1,-nbitq), 
to_sfixed(-338936639.0/4294967296.0,1,-nbitq), 
to_sfixed(121900003.0/4294967296.0,1,-nbitq), 
to_sfixed(348764579.0/4294967296.0,1,-nbitq), 
to_sfixed(-195954780.0/4294967296.0,1,-nbitq), 
to_sfixed(-45220749.0/4294967296.0,1,-nbitq), 
to_sfixed(394257860.0/4294967296.0,1,-nbitq), 
to_sfixed(-180999549.0/4294967296.0,1,-nbitq), 
to_sfixed(224413062.0/4294967296.0,1,-nbitq), 
to_sfixed(139326162.0/4294967296.0,1,-nbitq), 
to_sfixed(172587143.0/4294967296.0,1,-nbitq), 
to_sfixed(-63167541.0/4294967296.0,1,-nbitq), 
to_sfixed(-253583461.0/4294967296.0,1,-nbitq), 
to_sfixed(632193680.0/4294967296.0,1,-nbitq), 
to_sfixed(-293257669.0/4294967296.0,1,-nbitq), 
to_sfixed(251718995.0/4294967296.0,1,-nbitq), 
to_sfixed(99419632.0/4294967296.0,1,-nbitq), 
to_sfixed(-105027125.0/4294967296.0,1,-nbitq), 
to_sfixed(225632068.0/4294967296.0,1,-nbitq), 
to_sfixed(-253158578.0/4294967296.0,1,-nbitq), 
to_sfixed(-451424869.0/4294967296.0,1,-nbitq), 
to_sfixed(334201757.0/4294967296.0,1,-nbitq), 
to_sfixed(-233478171.0/4294967296.0,1,-nbitq), 
to_sfixed(339151003.0/4294967296.0,1,-nbitq), 
to_sfixed(46201816.0/4294967296.0,1,-nbitq), 
to_sfixed(-117080396.0/4294967296.0,1,-nbitq), 
to_sfixed(-438141069.0/4294967296.0,1,-nbitq), 
to_sfixed(595260247.0/4294967296.0,1,-nbitq), 
to_sfixed(-83334037.0/4294967296.0,1,-nbitq), 
to_sfixed(547428576.0/4294967296.0,1,-nbitq), 
to_sfixed(-253993840.0/4294967296.0,1,-nbitq), 
to_sfixed(-193003569.0/4294967296.0,1,-nbitq), 
to_sfixed(66964267.0/4294967296.0,1,-nbitq), 
to_sfixed(-214011894.0/4294967296.0,1,-nbitq), 
to_sfixed(3231880.0/4294967296.0,1,-nbitq), 
to_sfixed(146333490.0/4294967296.0,1,-nbitq), 
to_sfixed(-152282969.0/4294967296.0,1,-nbitq), 
to_sfixed(59094630.0/4294967296.0,1,-nbitq), 
to_sfixed(-307439544.0/4294967296.0,1,-nbitq), 
to_sfixed(11570074.0/4294967296.0,1,-nbitq), 
to_sfixed(-49351761.0/4294967296.0,1,-nbitq), 
to_sfixed(-157473235.0/4294967296.0,1,-nbitq), 
to_sfixed(-636733963.0/4294967296.0,1,-nbitq), 
to_sfixed(-292889150.0/4294967296.0,1,-nbitq), 
to_sfixed(-70401241.0/4294967296.0,1,-nbitq), 
to_sfixed(208529049.0/4294967296.0,1,-nbitq), 
to_sfixed(216423634.0/4294967296.0,1,-nbitq), 
to_sfixed(90814401.0/4294967296.0,1,-nbitq), 
to_sfixed(-382958933.0/4294967296.0,1,-nbitq), 
to_sfixed(-325055477.0/4294967296.0,1,-nbitq), 
to_sfixed(93242133.0/4294967296.0,1,-nbitq), 
to_sfixed(-148456017.0/4294967296.0,1,-nbitq), 
to_sfixed(51065360.0/4294967296.0,1,-nbitq), 
to_sfixed(233594754.0/4294967296.0,1,-nbitq), 
to_sfixed(256967065.0/4294967296.0,1,-nbitq), 
to_sfixed(-211371438.0/4294967296.0,1,-nbitq), 
to_sfixed(361293155.0/4294967296.0,1,-nbitq), 
to_sfixed(378330738.0/4294967296.0,1,-nbitq), 
to_sfixed(27404951.0/4294967296.0,1,-nbitq), 
to_sfixed(37529277.0/4294967296.0,1,-nbitq), 
to_sfixed(1858834.0/4294967296.0,1,-nbitq), 
to_sfixed(188684723.0/4294967296.0,1,-nbitq), 
to_sfixed(-506272385.0/4294967296.0,1,-nbitq), 
to_sfixed(278507752.0/4294967296.0,1,-nbitq), 
to_sfixed(-50650522.0/4294967296.0,1,-nbitq), 
to_sfixed(-336886489.0/4294967296.0,1,-nbitq), 
to_sfixed(381236073.0/4294967296.0,1,-nbitq), 
to_sfixed(7722946.0/4294967296.0,1,-nbitq), 
to_sfixed(-305081485.0/4294967296.0,1,-nbitq), 
to_sfixed(609204018.0/4294967296.0,1,-nbitq), 
to_sfixed(-192563306.0/4294967296.0,1,-nbitq), 
to_sfixed(201108316.0/4294967296.0,1,-nbitq), 
to_sfixed(74023459.0/4294967296.0,1,-nbitq), 
to_sfixed(1734697.0/4294967296.0,1,-nbitq), 
to_sfixed(34540228.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(416626125.0/4294967296.0,1,-nbitq), 
to_sfixed(-464923091.0/4294967296.0,1,-nbitq), 
to_sfixed(24962992.0/4294967296.0,1,-nbitq), 
to_sfixed(-98635580.0/4294967296.0,1,-nbitq), 
to_sfixed(-293111488.0/4294967296.0,1,-nbitq), 
to_sfixed(-156685737.0/4294967296.0,1,-nbitq), 
to_sfixed(173323821.0/4294967296.0,1,-nbitq), 
to_sfixed(114966399.0/4294967296.0,1,-nbitq), 
to_sfixed(-120351764.0/4294967296.0,1,-nbitq), 
to_sfixed(251188795.0/4294967296.0,1,-nbitq), 
to_sfixed(12621322.0/4294967296.0,1,-nbitq), 
to_sfixed(297994071.0/4294967296.0,1,-nbitq), 
to_sfixed(-582385845.0/4294967296.0,1,-nbitq), 
to_sfixed(-162615878.0/4294967296.0,1,-nbitq), 
to_sfixed(386603225.0/4294967296.0,1,-nbitq), 
to_sfixed(-381660261.0/4294967296.0,1,-nbitq), 
to_sfixed(-405610971.0/4294967296.0,1,-nbitq), 
to_sfixed(-392340272.0/4294967296.0,1,-nbitq), 
to_sfixed(503932111.0/4294967296.0,1,-nbitq), 
to_sfixed(28123205.0/4294967296.0,1,-nbitq), 
to_sfixed(371371677.0/4294967296.0,1,-nbitq), 
to_sfixed(296349811.0/4294967296.0,1,-nbitq), 
to_sfixed(515430964.0/4294967296.0,1,-nbitq), 
to_sfixed(-197454537.0/4294967296.0,1,-nbitq), 
to_sfixed(118405935.0/4294967296.0,1,-nbitq), 
to_sfixed(-45589939.0/4294967296.0,1,-nbitq), 
to_sfixed(-12653831.0/4294967296.0,1,-nbitq), 
to_sfixed(-531874878.0/4294967296.0,1,-nbitq), 
to_sfixed(256247939.0/4294967296.0,1,-nbitq), 
to_sfixed(517242378.0/4294967296.0,1,-nbitq), 
to_sfixed(-319737617.0/4294967296.0,1,-nbitq), 
to_sfixed(-376461266.0/4294967296.0,1,-nbitq), 
to_sfixed(146230831.0/4294967296.0,1,-nbitq), 
to_sfixed(553721846.0/4294967296.0,1,-nbitq), 
to_sfixed(517843730.0/4294967296.0,1,-nbitq), 
to_sfixed(367436025.0/4294967296.0,1,-nbitq), 
to_sfixed(421308622.0/4294967296.0,1,-nbitq), 
to_sfixed(-64130592.0/4294967296.0,1,-nbitq), 
to_sfixed(263706881.0/4294967296.0,1,-nbitq), 
to_sfixed(306288236.0/4294967296.0,1,-nbitq), 
to_sfixed(-193175728.0/4294967296.0,1,-nbitq), 
to_sfixed(271685638.0/4294967296.0,1,-nbitq), 
to_sfixed(-250854400.0/4294967296.0,1,-nbitq), 
to_sfixed(-308423521.0/4294967296.0,1,-nbitq), 
to_sfixed(-42718135.0/4294967296.0,1,-nbitq), 
to_sfixed(66292378.0/4294967296.0,1,-nbitq), 
to_sfixed(-20879546.0/4294967296.0,1,-nbitq), 
to_sfixed(-130781994.0/4294967296.0,1,-nbitq), 
to_sfixed(166689011.0/4294967296.0,1,-nbitq), 
to_sfixed(-294825446.0/4294967296.0,1,-nbitq), 
to_sfixed(162806944.0/4294967296.0,1,-nbitq), 
to_sfixed(47565090.0/4294967296.0,1,-nbitq), 
to_sfixed(61098831.0/4294967296.0,1,-nbitq), 
to_sfixed(-7780300.0/4294967296.0,1,-nbitq), 
to_sfixed(-286574590.0/4294967296.0,1,-nbitq), 
to_sfixed(40720553.0/4294967296.0,1,-nbitq), 
to_sfixed(113963272.0/4294967296.0,1,-nbitq), 
to_sfixed(-140561160.0/4294967296.0,1,-nbitq), 
to_sfixed(-219945299.0/4294967296.0,1,-nbitq), 
to_sfixed(-18020700.0/4294967296.0,1,-nbitq), 
to_sfixed(-394425961.0/4294967296.0,1,-nbitq), 
to_sfixed(475089325.0/4294967296.0,1,-nbitq), 
to_sfixed(-176528548.0/4294967296.0,1,-nbitq), 
to_sfixed(248017821.0/4294967296.0,1,-nbitq), 
to_sfixed(-146830721.0/4294967296.0,1,-nbitq), 
to_sfixed(-132850366.0/4294967296.0,1,-nbitq), 
to_sfixed(26898986.0/4294967296.0,1,-nbitq), 
to_sfixed(-432811250.0/4294967296.0,1,-nbitq), 
to_sfixed(92563781.0/4294967296.0,1,-nbitq), 
to_sfixed(-397672249.0/4294967296.0,1,-nbitq), 
to_sfixed(-484733411.0/4294967296.0,1,-nbitq), 
to_sfixed(-246616585.0/4294967296.0,1,-nbitq), 
to_sfixed(-137137062.0/4294967296.0,1,-nbitq), 
to_sfixed(-313356424.0/4294967296.0,1,-nbitq), 
to_sfixed(381360411.0/4294967296.0,1,-nbitq), 
to_sfixed(-467533513.0/4294967296.0,1,-nbitq), 
to_sfixed(-23019670.0/4294967296.0,1,-nbitq), 
to_sfixed(-163979621.0/4294967296.0,1,-nbitq), 
to_sfixed(383522163.0/4294967296.0,1,-nbitq), 
to_sfixed(109469420.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(14392640.0/4294967296.0,1,-nbitq), 
to_sfixed(-191569190.0/4294967296.0,1,-nbitq), 
to_sfixed(-242815936.0/4294967296.0,1,-nbitq), 
to_sfixed(-405802623.0/4294967296.0,1,-nbitq), 
to_sfixed(-145127580.0/4294967296.0,1,-nbitq), 
to_sfixed(89178857.0/4294967296.0,1,-nbitq), 
to_sfixed(-97419187.0/4294967296.0,1,-nbitq), 
to_sfixed(214202523.0/4294967296.0,1,-nbitq), 
to_sfixed(-78668603.0/4294967296.0,1,-nbitq), 
to_sfixed(140343167.0/4294967296.0,1,-nbitq), 
to_sfixed(-393701391.0/4294967296.0,1,-nbitq), 
to_sfixed(279434410.0/4294967296.0,1,-nbitq), 
to_sfixed(298967227.0/4294967296.0,1,-nbitq), 
to_sfixed(376766460.0/4294967296.0,1,-nbitq), 
to_sfixed(-35197878.0/4294967296.0,1,-nbitq), 
to_sfixed(-120497391.0/4294967296.0,1,-nbitq), 
to_sfixed(294861548.0/4294967296.0,1,-nbitq), 
to_sfixed(-180271795.0/4294967296.0,1,-nbitq), 
to_sfixed(512501697.0/4294967296.0,1,-nbitq), 
to_sfixed(-65923869.0/4294967296.0,1,-nbitq), 
to_sfixed(230227041.0/4294967296.0,1,-nbitq), 
to_sfixed(20835014.0/4294967296.0,1,-nbitq), 
to_sfixed(-179599515.0/4294967296.0,1,-nbitq), 
to_sfixed(-253900235.0/4294967296.0,1,-nbitq), 
to_sfixed(-289902160.0/4294967296.0,1,-nbitq), 
to_sfixed(37472683.0/4294967296.0,1,-nbitq), 
to_sfixed(-249185034.0/4294967296.0,1,-nbitq), 
to_sfixed(-5758463.0/4294967296.0,1,-nbitq), 
to_sfixed(-252180825.0/4294967296.0,1,-nbitq), 
to_sfixed(267090433.0/4294967296.0,1,-nbitq), 
to_sfixed(118354163.0/4294967296.0,1,-nbitq), 
to_sfixed(-222339719.0/4294967296.0,1,-nbitq), 
to_sfixed(-225644249.0/4294967296.0,1,-nbitq), 
to_sfixed(222403832.0/4294967296.0,1,-nbitq), 
to_sfixed(342027107.0/4294967296.0,1,-nbitq), 
to_sfixed(-54846051.0/4294967296.0,1,-nbitq), 
to_sfixed(-295908786.0/4294967296.0,1,-nbitq), 
to_sfixed(4201665.0/4294967296.0,1,-nbitq), 
to_sfixed(133429087.0/4294967296.0,1,-nbitq), 
to_sfixed(393065013.0/4294967296.0,1,-nbitq), 
to_sfixed(-165307146.0/4294967296.0,1,-nbitq), 
to_sfixed(350391348.0/4294967296.0,1,-nbitq), 
to_sfixed(201424980.0/4294967296.0,1,-nbitq), 
to_sfixed(34418778.0/4294967296.0,1,-nbitq), 
to_sfixed(-199960292.0/4294967296.0,1,-nbitq), 
to_sfixed(234718907.0/4294967296.0,1,-nbitq), 
to_sfixed(-65356188.0/4294967296.0,1,-nbitq), 
to_sfixed(-68594907.0/4294967296.0,1,-nbitq), 
to_sfixed(334170237.0/4294967296.0,1,-nbitq), 
to_sfixed(-108745234.0/4294967296.0,1,-nbitq), 
to_sfixed(200802731.0/4294967296.0,1,-nbitq), 
to_sfixed(459602607.0/4294967296.0,1,-nbitq), 
to_sfixed(-161461730.0/4294967296.0,1,-nbitq), 
to_sfixed(-161908463.0/4294967296.0,1,-nbitq), 
to_sfixed(-219922735.0/4294967296.0,1,-nbitq), 
to_sfixed(49041397.0/4294967296.0,1,-nbitq), 
to_sfixed(-331449758.0/4294967296.0,1,-nbitq), 
to_sfixed(-360344412.0/4294967296.0,1,-nbitq), 
to_sfixed(-179940308.0/4294967296.0,1,-nbitq), 
to_sfixed(132628321.0/4294967296.0,1,-nbitq), 
to_sfixed(-303848957.0/4294967296.0,1,-nbitq), 
to_sfixed(253100837.0/4294967296.0,1,-nbitq), 
to_sfixed(-362899203.0/4294967296.0,1,-nbitq), 
to_sfixed(213931219.0/4294967296.0,1,-nbitq), 
to_sfixed(447800236.0/4294967296.0,1,-nbitq), 
to_sfixed(-182502815.0/4294967296.0,1,-nbitq), 
to_sfixed(552015099.0/4294967296.0,1,-nbitq), 
to_sfixed(161929374.0/4294967296.0,1,-nbitq), 
to_sfixed(283465639.0/4294967296.0,1,-nbitq), 
to_sfixed(41850375.0/4294967296.0,1,-nbitq), 
to_sfixed(-381411782.0/4294967296.0,1,-nbitq), 
to_sfixed(-223677346.0/4294967296.0,1,-nbitq), 
to_sfixed(-496929678.0/4294967296.0,1,-nbitq), 
to_sfixed(434823592.0/4294967296.0,1,-nbitq), 
to_sfixed(388077596.0/4294967296.0,1,-nbitq), 
to_sfixed(83225245.0/4294967296.0,1,-nbitq), 
to_sfixed(-352632328.0/4294967296.0,1,-nbitq), 
to_sfixed(-366986498.0/4294967296.0,1,-nbitq), 
to_sfixed(185002821.0/4294967296.0,1,-nbitq), 
to_sfixed(-216493303.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-241424556.0/4294967296.0,1,-nbitq), 
to_sfixed(209838489.0/4294967296.0,1,-nbitq), 
to_sfixed(-279962966.0/4294967296.0,1,-nbitq), 
to_sfixed(-378810767.0/4294967296.0,1,-nbitq), 
to_sfixed(138905367.0/4294967296.0,1,-nbitq), 
to_sfixed(-239915215.0/4294967296.0,1,-nbitq), 
to_sfixed(262805807.0/4294967296.0,1,-nbitq), 
to_sfixed(-92875510.0/4294967296.0,1,-nbitq), 
to_sfixed(157209673.0/4294967296.0,1,-nbitq), 
to_sfixed(-20441001.0/4294967296.0,1,-nbitq), 
to_sfixed(-2513802.0/4294967296.0,1,-nbitq), 
to_sfixed(-38793967.0/4294967296.0,1,-nbitq), 
to_sfixed(254690139.0/4294967296.0,1,-nbitq), 
to_sfixed(-271685579.0/4294967296.0,1,-nbitq), 
to_sfixed(-154552662.0/4294967296.0,1,-nbitq), 
to_sfixed(-475666575.0/4294967296.0,1,-nbitq), 
to_sfixed(-7515062.0/4294967296.0,1,-nbitq), 
to_sfixed(-299683311.0/4294967296.0,1,-nbitq), 
to_sfixed(621267473.0/4294967296.0,1,-nbitq), 
to_sfixed(-422315850.0/4294967296.0,1,-nbitq), 
to_sfixed(-156202704.0/4294967296.0,1,-nbitq), 
to_sfixed(232024742.0/4294967296.0,1,-nbitq), 
to_sfixed(319208382.0/4294967296.0,1,-nbitq), 
to_sfixed(-367693393.0/4294967296.0,1,-nbitq), 
to_sfixed(212941816.0/4294967296.0,1,-nbitq), 
to_sfixed(-63275017.0/4294967296.0,1,-nbitq), 
to_sfixed(-261715881.0/4294967296.0,1,-nbitq), 
to_sfixed(-145009777.0/4294967296.0,1,-nbitq), 
to_sfixed(-26447797.0/4294967296.0,1,-nbitq), 
to_sfixed(68560895.0/4294967296.0,1,-nbitq), 
to_sfixed(-246639596.0/4294967296.0,1,-nbitq), 
to_sfixed(-231219938.0/4294967296.0,1,-nbitq), 
to_sfixed(-194718970.0/4294967296.0,1,-nbitq), 
to_sfixed(-312451281.0/4294967296.0,1,-nbitq), 
to_sfixed(380955063.0/4294967296.0,1,-nbitq), 
to_sfixed(-38866743.0/4294967296.0,1,-nbitq), 
to_sfixed(-265974227.0/4294967296.0,1,-nbitq), 
to_sfixed(-418226351.0/4294967296.0,1,-nbitq), 
to_sfixed(194650725.0/4294967296.0,1,-nbitq), 
to_sfixed(-108286252.0/4294967296.0,1,-nbitq), 
to_sfixed(172264097.0/4294967296.0,1,-nbitq), 
to_sfixed(269930098.0/4294967296.0,1,-nbitq), 
to_sfixed(-50491708.0/4294967296.0,1,-nbitq), 
to_sfixed(438237950.0/4294967296.0,1,-nbitq), 
to_sfixed(321493090.0/4294967296.0,1,-nbitq), 
to_sfixed(248275725.0/4294967296.0,1,-nbitq), 
to_sfixed(-211097918.0/4294967296.0,1,-nbitq), 
to_sfixed(-121725067.0/4294967296.0,1,-nbitq), 
to_sfixed(-175425958.0/4294967296.0,1,-nbitq), 
to_sfixed(119392698.0/4294967296.0,1,-nbitq), 
to_sfixed(72052147.0/4294967296.0,1,-nbitq), 
to_sfixed(413271858.0/4294967296.0,1,-nbitq), 
to_sfixed(-95903628.0/4294967296.0,1,-nbitq), 
to_sfixed(286575345.0/4294967296.0,1,-nbitq), 
to_sfixed(13203779.0/4294967296.0,1,-nbitq), 
to_sfixed(-413009117.0/4294967296.0,1,-nbitq), 
to_sfixed(-307686989.0/4294967296.0,1,-nbitq), 
to_sfixed(55205430.0/4294967296.0,1,-nbitq), 
to_sfixed(-16578007.0/4294967296.0,1,-nbitq), 
to_sfixed(-326741380.0/4294967296.0,1,-nbitq), 
to_sfixed(279285561.0/4294967296.0,1,-nbitq), 
to_sfixed(-217610274.0/4294967296.0,1,-nbitq), 
to_sfixed(-413942728.0/4294967296.0,1,-nbitq), 
to_sfixed(-103984975.0/4294967296.0,1,-nbitq), 
to_sfixed(-266543321.0/4294967296.0,1,-nbitq), 
to_sfixed(-99502453.0/4294967296.0,1,-nbitq), 
to_sfixed(437121361.0/4294967296.0,1,-nbitq), 
to_sfixed(32150137.0/4294967296.0,1,-nbitq), 
to_sfixed(299017320.0/4294967296.0,1,-nbitq), 
to_sfixed(-54557010.0/4294967296.0,1,-nbitq), 
to_sfixed(-539855927.0/4294967296.0,1,-nbitq), 
to_sfixed(-105633523.0/4294967296.0,1,-nbitq), 
to_sfixed(-487581988.0/4294967296.0,1,-nbitq), 
to_sfixed(98052030.0/4294967296.0,1,-nbitq), 
to_sfixed(179758050.0/4294967296.0,1,-nbitq), 
to_sfixed(-156229377.0/4294967296.0,1,-nbitq), 
to_sfixed(232139153.0/4294967296.0,1,-nbitq), 
to_sfixed(-416238286.0/4294967296.0,1,-nbitq), 
to_sfixed(123289079.0/4294967296.0,1,-nbitq), 
to_sfixed(84807580.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-97501897.0/4294967296.0,1,-nbitq), 
to_sfixed(21561192.0/4294967296.0,1,-nbitq), 
to_sfixed(87194467.0/4294967296.0,1,-nbitq), 
to_sfixed(129569250.0/4294967296.0,1,-nbitq), 
to_sfixed(34785318.0/4294967296.0,1,-nbitq), 
to_sfixed(-155128097.0/4294967296.0,1,-nbitq), 
to_sfixed(233772076.0/4294967296.0,1,-nbitq), 
to_sfixed(-175203371.0/4294967296.0,1,-nbitq), 
to_sfixed(191646769.0/4294967296.0,1,-nbitq), 
to_sfixed(442839798.0/4294967296.0,1,-nbitq), 
to_sfixed(-335352170.0/4294967296.0,1,-nbitq), 
to_sfixed(192308248.0/4294967296.0,1,-nbitq), 
to_sfixed(251021495.0/4294967296.0,1,-nbitq), 
to_sfixed(245860357.0/4294967296.0,1,-nbitq), 
to_sfixed(314499818.0/4294967296.0,1,-nbitq), 
to_sfixed(-217203059.0/4294967296.0,1,-nbitq), 
to_sfixed(312034242.0/4294967296.0,1,-nbitq), 
to_sfixed(412437937.0/4294967296.0,1,-nbitq), 
to_sfixed(97062666.0/4294967296.0,1,-nbitq), 
to_sfixed(-181240819.0/4294967296.0,1,-nbitq), 
to_sfixed(351313553.0/4294967296.0,1,-nbitq), 
to_sfixed(70306525.0/4294967296.0,1,-nbitq), 
to_sfixed(262655751.0/4294967296.0,1,-nbitq), 
to_sfixed(6244173.0/4294967296.0,1,-nbitq), 
to_sfixed(256218969.0/4294967296.0,1,-nbitq), 
to_sfixed(16901037.0/4294967296.0,1,-nbitq), 
to_sfixed(-366280805.0/4294967296.0,1,-nbitq), 
to_sfixed(5208055.0/4294967296.0,1,-nbitq), 
to_sfixed(211338495.0/4294967296.0,1,-nbitq), 
to_sfixed(176162116.0/4294967296.0,1,-nbitq), 
to_sfixed(-499731844.0/4294967296.0,1,-nbitq), 
to_sfixed(-491721788.0/4294967296.0,1,-nbitq), 
to_sfixed(325991966.0/4294967296.0,1,-nbitq), 
to_sfixed(-373400324.0/4294967296.0,1,-nbitq), 
to_sfixed(464679846.0/4294967296.0,1,-nbitq), 
to_sfixed(-162887249.0/4294967296.0,1,-nbitq), 
to_sfixed(309563374.0/4294967296.0,1,-nbitq), 
to_sfixed(-289091354.0/4294967296.0,1,-nbitq), 
to_sfixed(350615726.0/4294967296.0,1,-nbitq), 
to_sfixed(435892593.0/4294967296.0,1,-nbitq), 
to_sfixed(-151453664.0/4294967296.0,1,-nbitq), 
to_sfixed(-77236711.0/4294967296.0,1,-nbitq), 
to_sfixed(-47661112.0/4294967296.0,1,-nbitq), 
to_sfixed(283890169.0/4294967296.0,1,-nbitq), 
to_sfixed(199126243.0/4294967296.0,1,-nbitq), 
to_sfixed(-176182829.0/4294967296.0,1,-nbitq), 
to_sfixed(327569180.0/4294967296.0,1,-nbitq), 
to_sfixed(-444903739.0/4294967296.0,1,-nbitq), 
to_sfixed(-49396045.0/4294967296.0,1,-nbitq), 
to_sfixed(420617395.0/4294967296.0,1,-nbitq), 
to_sfixed(-232786511.0/4294967296.0,1,-nbitq), 
to_sfixed(178745461.0/4294967296.0,1,-nbitq), 
to_sfixed(-623252177.0/4294967296.0,1,-nbitq), 
to_sfixed(-224056422.0/4294967296.0,1,-nbitq), 
to_sfixed(-102840309.0/4294967296.0,1,-nbitq), 
to_sfixed(-141303550.0/4294967296.0,1,-nbitq), 
to_sfixed(164852688.0/4294967296.0,1,-nbitq), 
to_sfixed(-294897617.0/4294967296.0,1,-nbitq), 
to_sfixed(-127777625.0/4294967296.0,1,-nbitq), 
to_sfixed(325404050.0/4294967296.0,1,-nbitq), 
to_sfixed(-263530984.0/4294967296.0,1,-nbitq), 
to_sfixed(52976660.0/4294967296.0,1,-nbitq), 
to_sfixed(-377607384.0/4294967296.0,1,-nbitq), 
to_sfixed(-287605306.0/4294967296.0,1,-nbitq), 
to_sfixed(267812526.0/4294967296.0,1,-nbitq), 
to_sfixed(255162175.0/4294967296.0,1,-nbitq), 
to_sfixed(285015748.0/4294967296.0,1,-nbitq), 
to_sfixed(-247041366.0/4294967296.0,1,-nbitq), 
to_sfixed(114615626.0/4294967296.0,1,-nbitq), 
to_sfixed(400807439.0/4294967296.0,1,-nbitq), 
to_sfixed(-191843199.0/4294967296.0,1,-nbitq), 
to_sfixed(198441703.0/4294967296.0,1,-nbitq), 
to_sfixed(119225234.0/4294967296.0,1,-nbitq), 
to_sfixed(-333395925.0/4294967296.0,1,-nbitq), 
to_sfixed(497665942.0/4294967296.0,1,-nbitq), 
to_sfixed(-554687334.0/4294967296.0,1,-nbitq), 
to_sfixed(-428104561.0/4294967296.0,1,-nbitq), 
to_sfixed(173457484.0/4294967296.0,1,-nbitq), 
to_sfixed(197164919.0/4294967296.0,1,-nbitq), 
to_sfixed(250155307.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-51201556.0/4294967296.0,1,-nbitq), 
to_sfixed(47917472.0/4294967296.0,1,-nbitq), 
to_sfixed(-355578891.0/4294967296.0,1,-nbitq), 
to_sfixed(-440784905.0/4294967296.0,1,-nbitq), 
to_sfixed(-29248081.0/4294967296.0,1,-nbitq), 
to_sfixed(-467317948.0/4294967296.0,1,-nbitq), 
to_sfixed(66664902.0/4294967296.0,1,-nbitq), 
to_sfixed(305481115.0/4294967296.0,1,-nbitq), 
to_sfixed(-14940664.0/4294967296.0,1,-nbitq), 
to_sfixed(-263203755.0/4294967296.0,1,-nbitq), 
to_sfixed(-244578126.0/4294967296.0,1,-nbitq), 
to_sfixed(3356560.0/4294967296.0,1,-nbitq), 
to_sfixed(-234695902.0/4294967296.0,1,-nbitq), 
to_sfixed(-328836542.0/4294967296.0,1,-nbitq), 
to_sfixed(291141095.0/4294967296.0,1,-nbitq), 
to_sfixed(130619099.0/4294967296.0,1,-nbitq), 
to_sfixed(175806557.0/4294967296.0,1,-nbitq), 
to_sfixed(288108207.0/4294967296.0,1,-nbitq), 
to_sfixed(617484080.0/4294967296.0,1,-nbitq), 
to_sfixed(232118072.0/4294967296.0,1,-nbitq), 
to_sfixed(-365222385.0/4294967296.0,1,-nbitq), 
to_sfixed(182052075.0/4294967296.0,1,-nbitq), 
to_sfixed(410182635.0/4294967296.0,1,-nbitq), 
to_sfixed(385814685.0/4294967296.0,1,-nbitq), 
to_sfixed(-156191952.0/4294967296.0,1,-nbitq), 
to_sfixed(-12444668.0/4294967296.0,1,-nbitq), 
to_sfixed(198566031.0/4294967296.0,1,-nbitq), 
to_sfixed(-226275966.0/4294967296.0,1,-nbitq), 
to_sfixed(264280755.0/4294967296.0,1,-nbitq), 
to_sfixed(353737943.0/4294967296.0,1,-nbitq), 
to_sfixed(-586009492.0/4294967296.0,1,-nbitq), 
to_sfixed(-360902807.0/4294967296.0,1,-nbitq), 
to_sfixed(31372054.0/4294967296.0,1,-nbitq), 
to_sfixed(-88829713.0/4294967296.0,1,-nbitq), 
to_sfixed(10041562.0/4294967296.0,1,-nbitq), 
to_sfixed(-180729708.0/4294967296.0,1,-nbitq), 
to_sfixed(194831230.0/4294967296.0,1,-nbitq), 
to_sfixed(-217490895.0/4294967296.0,1,-nbitq), 
to_sfixed(128153828.0/4294967296.0,1,-nbitq), 
to_sfixed(373280637.0/4294967296.0,1,-nbitq), 
to_sfixed(-5781846.0/4294967296.0,1,-nbitq), 
to_sfixed(70110684.0/4294967296.0,1,-nbitq), 
to_sfixed(194246028.0/4294967296.0,1,-nbitq), 
to_sfixed(347480160.0/4294967296.0,1,-nbitq), 
to_sfixed(185811802.0/4294967296.0,1,-nbitq), 
to_sfixed(336533109.0/4294967296.0,1,-nbitq), 
to_sfixed(56636770.0/4294967296.0,1,-nbitq), 
to_sfixed(-323865782.0/4294967296.0,1,-nbitq), 
to_sfixed(362978510.0/4294967296.0,1,-nbitq), 
to_sfixed(305112277.0/4294967296.0,1,-nbitq), 
to_sfixed(-191146533.0/4294967296.0,1,-nbitq), 
to_sfixed(-279881977.0/4294967296.0,1,-nbitq), 
to_sfixed(-199149060.0/4294967296.0,1,-nbitq), 
to_sfixed(326307285.0/4294967296.0,1,-nbitq), 
to_sfixed(297560925.0/4294967296.0,1,-nbitq), 
to_sfixed(332126364.0/4294967296.0,1,-nbitq), 
to_sfixed(300195774.0/4294967296.0,1,-nbitq), 
to_sfixed(19811729.0/4294967296.0,1,-nbitq), 
to_sfixed(222163803.0/4294967296.0,1,-nbitq), 
to_sfixed(-17684423.0/4294967296.0,1,-nbitq), 
to_sfixed(-277738931.0/4294967296.0,1,-nbitq), 
to_sfixed(475989307.0/4294967296.0,1,-nbitq), 
to_sfixed(-152919799.0/4294967296.0,1,-nbitq), 
to_sfixed(224125363.0/4294967296.0,1,-nbitq), 
to_sfixed(-220105453.0/4294967296.0,1,-nbitq), 
to_sfixed(290659062.0/4294967296.0,1,-nbitq), 
to_sfixed(506400802.0/4294967296.0,1,-nbitq), 
to_sfixed(-347848955.0/4294967296.0,1,-nbitq), 
to_sfixed(-252416832.0/4294967296.0,1,-nbitq), 
to_sfixed(551098957.0/4294967296.0,1,-nbitq), 
to_sfixed(-160992812.0/4294967296.0,1,-nbitq), 
to_sfixed(311852489.0/4294967296.0,1,-nbitq), 
to_sfixed(155186887.0/4294967296.0,1,-nbitq), 
to_sfixed(355015659.0/4294967296.0,1,-nbitq), 
to_sfixed(-214782714.0/4294967296.0,1,-nbitq), 
to_sfixed(-216148914.0/4294967296.0,1,-nbitq), 
to_sfixed(32017814.0/4294967296.0,1,-nbitq), 
to_sfixed(-366750264.0/4294967296.0,1,-nbitq), 
to_sfixed(-140413735.0/4294967296.0,1,-nbitq), 
to_sfixed(-240000862.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(278185752.0/4294967296.0,1,-nbitq), 
to_sfixed(-280031427.0/4294967296.0,1,-nbitq), 
to_sfixed(-29677964.0/4294967296.0,1,-nbitq), 
to_sfixed(67769487.0/4294967296.0,1,-nbitq), 
to_sfixed(26304605.0/4294967296.0,1,-nbitq), 
to_sfixed(-122902921.0/4294967296.0,1,-nbitq), 
to_sfixed(308533430.0/4294967296.0,1,-nbitq), 
to_sfixed(362926015.0/4294967296.0,1,-nbitq), 
to_sfixed(-157092729.0/4294967296.0,1,-nbitq), 
to_sfixed(-97373522.0/4294967296.0,1,-nbitq), 
to_sfixed(-82242448.0/4294967296.0,1,-nbitq), 
to_sfixed(258007208.0/4294967296.0,1,-nbitq), 
to_sfixed(-151181371.0/4294967296.0,1,-nbitq), 
to_sfixed(430293667.0/4294967296.0,1,-nbitq), 
to_sfixed(-158647835.0/4294967296.0,1,-nbitq), 
to_sfixed(-311313184.0/4294967296.0,1,-nbitq), 
to_sfixed(80095856.0/4294967296.0,1,-nbitq), 
to_sfixed(83629571.0/4294967296.0,1,-nbitq), 
to_sfixed(447521747.0/4294967296.0,1,-nbitq), 
to_sfixed(-216173475.0/4294967296.0,1,-nbitq), 
to_sfixed(318388816.0/4294967296.0,1,-nbitq), 
to_sfixed(225335143.0/4294967296.0,1,-nbitq), 
to_sfixed(406265590.0/4294967296.0,1,-nbitq), 
to_sfixed(54921699.0/4294967296.0,1,-nbitq), 
to_sfixed(20555999.0/4294967296.0,1,-nbitq), 
to_sfixed(303003983.0/4294967296.0,1,-nbitq), 
to_sfixed(-186029749.0/4294967296.0,1,-nbitq), 
to_sfixed(-333400962.0/4294967296.0,1,-nbitq), 
to_sfixed(320122232.0/4294967296.0,1,-nbitq), 
to_sfixed(-283360302.0/4294967296.0,1,-nbitq), 
to_sfixed(-248828185.0/4294967296.0,1,-nbitq), 
to_sfixed(196798556.0/4294967296.0,1,-nbitq), 
to_sfixed(331668024.0/4294967296.0,1,-nbitq), 
to_sfixed(-65054455.0/4294967296.0,1,-nbitq), 
to_sfixed(-139072262.0/4294967296.0,1,-nbitq), 
to_sfixed(-5344646.0/4294967296.0,1,-nbitq), 
to_sfixed(156789175.0/4294967296.0,1,-nbitq), 
to_sfixed(-125793157.0/4294967296.0,1,-nbitq), 
to_sfixed(-39281005.0/4294967296.0,1,-nbitq), 
to_sfixed(-265605076.0/4294967296.0,1,-nbitq), 
to_sfixed(-30863238.0/4294967296.0,1,-nbitq), 
to_sfixed(-35235825.0/4294967296.0,1,-nbitq), 
to_sfixed(-258971030.0/4294967296.0,1,-nbitq), 
to_sfixed(-72449449.0/4294967296.0,1,-nbitq), 
to_sfixed(81265506.0/4294967296.0,1,-nbitq), 
to_sfixed(401096694.0/4294967296.0,1,-nbitq), 
to_sfixed(96621930.0/4294967296.0,1,-nbitq), 
to_sfixed(-15247198.0/4294967296.0,1,-nbitq), 
to_sfixed(-101059316.0/4294967296.0,1,-nbitq), 
to_sfixed(-115599115.0/4294967296.0,1,-nbitq), 
to_sfixed(-356088851.0/4294967296.0,1,-nbitq), 
to_sfixed(35504966.0/4294967296.0,1,-nbitq), 
to_sfixed(76457830.0/4294967296.0,1,-nbitq), 
to_sfixed(-207387097.0/4294967296.0,1,-nbitq), 
to_sfixed(-200793665.0/4294967296.0,1,-nbitq), 
to_sfixed(385312843.0/4294967296.0,1,-nbitq), 
to_sfixed(382935913.0/4294967296.0,1,-nbitq), 
to_sfixed(8220840.0/4294967296.0,1,-nbitq), 
to_sfixed(169907324.0/4294967296.0,1,-nbitq), 
to_sfixed(146362181.0/4294967296.0,1,-nbitq), 
to_sfixed(-325777256.0/4294967296.0,1,-nbitq), 
to_sfixed(303806363.0/4294967296.0,1,-nbitq), 
to_sfixed(55639635.0/4294967296.0,1,-nbitq), 
to_sfixed(-235673430.0/4294967296.0,1,-nbitq), 
to_sfixed(-102762357.0/4294967296.0,1,-nbitq), 
to_sfixed(229294398.0/4294967296.0,1,-nbitq), 
to_sfixed(575938198.0/4294967296.0,1,-nbitq), 
to_sfixed(314531643.0/4294967296.0,1,-nbitq), 
to_sfixed(-314156687.0/4294967296.0,1,-nbitq), 
to_sfixed(374946749.0/4294967296.0,1,-nbitq), 
to_sfixed(88454394.0/4294967296.0,1,-nbitq), 
to_sfixed(-356860308.0/4294967296.0,1,-nbitq), 
to_sfixed(-551604228.0/4294967296.0,1,-nbitq), 
to_sfixed(104862762.0/4294967296.0,1,-nbitq), 
to_sfixed(278714605.0/4294967296.0,1,-nbitq), 
to_sfixed(-362113428.0/4294967296.0,1,-nbitq), 
to_sfixed(-167075423.0/4294967296.0,1,-nbitq), 
to_sfixed(-399190979.0/4294967296.0,1,-nbitq), 
to_sfixed(5478252.0/4294967296.0,1,-nbitq), 
to_sfixed(331114314.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-185480330.0/4294967296.0,1,-nbitq), 
to_sfixed(76422508.0/4294967296.0,1,-nbitq), 
to_sfixed(86167229.0/4294967296.0,1,-nbitq), 
to_sfixed(-297473306.0/4294967296.0,1,-nbitq), 
to_sfixed(92922989.0/4294967296.0,1,-nbitq), 
to_sfixed(181586338.0/4294967296.0,1,-nbitq), 
to_sfixed(-234489653.0/4294967296.0,1,-nbitq), 
to_sfixed(-224279635.0/4294967296.0,1,-nbitq), 
to_sfixed(102591164.0/4294967296.0,1,-nbitq), 
to_sfixed(326215596.0/4294967296.0,1,-nbitq), 
to_sfixed(-112554119.0/4294967296.0,1,-nbitq), 
to_sfixed(118453862.0/4294967296.0,1,-nbitq), 
to_sfixed(-258147361.0/4294967296.0,1,-nbitq), 
to_sfixed(161013417.0/4294967296.0,1,-nbitq), 
to_sfixed(-178952867.0/4294967296.0,1,-nbitq), 
to_sfixed(-179010867.0/4294967296.0,1,-nbitq), 
to_sfixed(-118704235.0/4294967296.0,1,-nbitq), 
to_sfixed(-339672984.0/4294967296.0,1,-nbitq), 
to_sfixed(77773191.0/4294967296.0,1,-nbitq), 
to_sfixed(-445271160.0/4294967296.0,1,-nbitq), 
to_sfixed(296737549.0/4294967296.0,1,-nbitq), 
to_sfixed(284381333.0/4294967296.0,1,-nbitq), 
to_sfixed(-120637185.0/4294967296.0,1,-nbitq), 
to_sfixed(115404311.0/4294967296.0,1,-nbitq), 
to_sfixed(337562378.0/4294967296.0,1,-nbitq), 
to_sfixed(-159163001.0/4294967296.0,1,-nbitq), 
to_sfixed(327465008.0/4294967296.0,1,-nbitq), 
to_sfixed(-379285395.0/4294967296.0,1,-nbitq), 
to_sfixed(331.0/4294967296.0,1,-nbitq), 
to_sfixed(181616993.0/4294967296.0,1,-nbitq), 
to_sfixed(-283228182.0/4294967296.0,1,-nbitq), 
to_sfixed(-386245692.0/4294967296.0,1,-nbitq), 
to_sfixed(362379618.0/4294967296.0,1,-nbitq), 
to_sfixed(-410346895.0/4294967296.0,1,-nbitq), 
to_sfixed(365626991.0/4294967296.0,1,-nbitq), 
to_sfixed(159240642.0/4294967296.0,1,-nbitq), 
to_sfixed(331320327.0/4294967296.0,1,-nbitq), 
to_sfixed(-311230152.0/4294967296.0,1,-nbitq), 
to_sfixed(45742755.0/4294967296.0,1,-nbitq), 
to_sfixed(127091536.0/4294967296.0,1,-nbitq), 
to_sfixed(-394146086.0/4294967296.0,1,-nbitq), 
to_sfixed(121569823.0/4294967296.0,1,-nbitq), 
to_sfixed(-15981871.0/4294967296.0,1,-nbitq), 
to_sfixed(-16165666.0/4294967296.0,1,-nbitq), 
to_sfixed(-328186639.0/4294967296.0,1,-nbitq), 
to_sfixed(-37660649.0/4294967296.0,1,-nbitq), 
to_sfixed(-359366137.0/4294967296.0,1,-nbitq), 
to_sfixed(34860834.0/4294967296.0,1,-nbitq), 
to_sfixed(-367140533.0/4294967296.0,1,-nbitq), 
to_sfixed(504173896.0/4294967296.0,1,-nbitq), 
to_sfixed(114770992.0/4294967296.0,1,-nbitq), 
to_sfixed(459204885.0/4294967296.0,1,-nbitq), 
to_sfixed(-50616148.0/4294967296.0,1,-nbitq), 
to_sfixed(336739314.0/4294967296.0,1,-nbitq), 
to_sfixed(222201562.0/4294967296.0,1,-nbitq), 
to_sfixed(-363906392.0/4294967296.0,1,-nbitq), 
to_sfixed(-4020584.0/4294967296.0,1,-nbitq), 
to_sfixed(-58084805.0/4294967296.0,1,-nbitq), 
to_sfixed(-270162058.0/4294967296.0,1,-nbitq), 
to_sfixed(-316553210.0/4294967296.0,1,-nbitq), 
to_sfixed(292318517.0/4294967296.0,1,-nbitq), 
to_sfixed(110683311.0/4294967296.0,1,-nbitq), 
to_sfixed(-36238036.0/4294967296.0,1,-nbitq), 
to_sfixed(317109704.0/4294967296.0,1,-nbitq), 
to_sfixed(8010498.0/4294967296.0,1,-nbitq), 
to_sfixed(-69909050.0/4294967296.0,1,-nbitq), 
to_sfixed(211904616.0/4294967296.0,1,-nbitq), 
to_sfixed(-251199831.0/4294967296.0,1,-nbitq), 
to_sfixed(-136724397.0/4294967296.0,1,-nbitq), 
to_sfixed(-125587496.0/4294967296.0,1,-nbitq), 
to_sfixed(-153830764.0/4294967296.0,1,-nbitq), 
to_sfixed(267408336.0/4294967296.0,1,-nbitq), 
to_sfixed(103219601.0/4294967296.0,1,-nbitq), 
to_sfixed(-114411358.0/4294967296.0,1,-nbitq), 
to_sfixed(454665916.0/4294967296.0,1,-nbitq), 
to_sfixed(-257539095.0/4294967296.0,1,-nbitq), 
to_sfixed(289490465.0/4294967296.0,1,-nbitq), 
to_sfixed(-66918201.0/4294967296.0,1,-nbitq), 
to_sfixed(-46521208.0/4294967296.0,1,-nbitq), 
to_sfixed(169113458.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(107915451.0/4294967296.0,1,-nbitq), 
to_sfixed(42508125.0/4294967296.0,1,-nbitq), 
to_sfixed(207039498.0/4294967296.0,1,-nbitq), 
to_sfixed(166279140.0/4294967296.0,1,-nbitq), 
to_sfixed(-146755760.0/4294967296.0,1,-nbitq), 
to_sfixed(-3853977.0/4294967296.0,1,-nbitq), 
to_sfixed(11780283.0/4294967296.0,1,-nbitq), 
to_sfixed(-143161132.0/4294967296.0,1,-nbitq), 
to_sfixed(149244756.0/4294967296.0,1,-nbitq), 
to_sfixed(-279401295.0/4294967296.0,1,-nbitq), 
to_sfixed(-346322785.0/4294967296.0,1,-nbitq), 
to_sfixed(364250639.0/4294967296.0,1,-nbitq), 
to_sfixed(417436947.0/4294967296.0,1,-nbitq), 
to_sfixed(-177929721.0/4294967296.0,1,-nbitq), 
to_sfixed(-246219376.0/4294967296.0,1,-nbitq), 
to_sfixed(161970101.0/4294967296.0,1,-nbitq), 
to_sfixed(356479074.0/4294967296.0,1,-nbitq), 
to_sfixed(251892482.0/4294967296.0,1,-nbitq), 
to_sfixed(523055080.0/4294967296.0,1,-nbitq), 
to_sfixed(29516768.0/4294967296.0,1,-nbitq), 
to_sfixed(-362635614.0/4294967296.0,1,-nbitq), 
to_sfixed(-113889701.0/4294967296.0,1,-nbitq), 
to_sfixed(506843254.0/4294967296.0,1,-nbitq), 
to_sfixed(286800820.0/4294967296.0,1,-nbitq), 
to_sfixed(27305523.0/4294967296.0,1,-nbitq), 
to_sfixed(419095485.0/4294967296.0,1,-nbitq), 
to_sfixed(166264537.0/4294967296.0,1,-nbitq), 
to_sfixed(-578461169.0/4294967296.0,1,-nbitq), 
to_sfixed(-86294784.0/4294967296.0,1,-nbitq), 
to_sfixed(377900938.0/4294967296.0,1,-nbitq), 
to_sfixed(174867063.0/4294967296.0,1,-nbitq), 
to_sfixed(133949274.0/4294967296.0,1,-nbitq), 
to_sfixed(-223320217.0/4294967296.0,1,-nbitq), 
to_sfixed(215385809.0/4294967296.0,1,-nbitq), 
to_sfixed(-92321564.0/4294967296.0,1,-nbitq), 
to_sfixed(-180782168.0/4294967296.0,1,-nbitq), 
to_sfixed(-193737773.0/4294967296.0,1,-nbitq), 
to_sfixed(-103025035.0/4294967296.0,1,-nbitq), 
to_sfixed(-107685558.0/4294967296.0,1,-nbitq), 
to_sfixed(-160600721.0/4294967296.0,1,-nbitq), 
to_sfixed(-294855616.0/4294967296.0,1,-nbitq), 
to_sfixed(309590104.0/4294967296.0,1,-nbitq), 
to_sfixed(216112199.0/4294967296.0,1,-nbitq), 
to_sfixed(26774603.0/4294967296.0,1,-nbitq), 
to_sfixed(233136680.0/4294967296.0,1,-nbitq), 
to_sfixed(-151240828.0/4294967296.0,1,-nbitq), 
to_sfixed(-14701920.0/4294967296.0,1,-nbitq), 
to_sfixed(-536529258.0/4294967296.0,1,-nbitq), 
to_sfixed(137726193.0/4294967296.0,1,-nbitq), 
to_sfixed(137488302.0/4294967296.0,1,-nbitq), 
to_sfixed(-75767484.0/4294967296.0,1,-nbitq), 
to_sfixed(252714029.0/4294967296.0,1,-nbitq), 
to_sfixed(-51125335.0/4294967296.0,1,-nbitq), 
to_sfixed(142591269.0/4294967296.0,1,-nbitq), 
to_sfixed(64746167.0/4294967296.0,1,-nbitq), 
to_sfixed(-366926388.0/4294967296.0,1,-nbitq), 
to_sfixed(165208442.0/4294967296.0,1,-nbitq), 
to_sfixed(-55051988.0/4294967296.0,1,-nbitq), 
to_sfixed(269862277.0/4294967296.0,1,-nbitq), 
to_sfixed(13696514.0/4294967296.0,1,-nbitq), 
to_sfixed(-385625466.0/4294967296.0,1,-nbitq), 
to_sfixed(-246283826.0/4294967296.0,1,-nbitq), 
to_sfixed(137629617.0/4294967296.0,1,-nbitq), 
to_sfixed(-4279940.0/4294967296.0,1,-nbitq), 
to_sfixed(202324009.0/4294967296.0,1,-nbitq), 
to_sfixed(-63554091.0/4294967296.0,1,-nbitq), 
to_sfixed(824139672.0/4294967296.0,1,-nbitq), 
to_sfixed(-398387097.0/4294967296.0,1,-nbitq), 
to_sfixed(173010583.0/4294967296.0,1,-nbitq), 
to_sfixed(-117244121.0/4294967296.0,1,-nbitq), 
to_sfixed(-416635581.0/4294967296.0,1,-nbitq), 
to_sfixed(58263802.0/4294967296.0,1,-nbitq), 
to_sfixed(-22542826.0/4294967296.0,1,-nbitq), 
to_sfixed(392004790.0/4294967296.0,1,-nbitq), 
to_sfixed(-225469865.0/4294967296.0,1,-nbitq), 
to_sfixed(-607477110.0/4294967296.0,1,-nbitq), 
to_sfixed(-34100256.0/4294967296.0,1,-nbitq), 
to_sfixed(290621362.0/4294967296.0,1,-nbitq), 
to_sfixed(179768507.0/4294967296.0,1,-nbitq), 
to_sfixed(-218086407.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(304047478.0/4294967296.0,1,-nbitq), 
to_sfixed(-213930931.0/4294967296.0,1,-nbitq), 
to_sfixed(-169172116.0/4294967296.0,1,-nbitq), 
to_sfixed(314956089.0/4294967296.0,1,-nbitq), 
to_sfixed(397518515.0/4294967296.0,1,-nbitq), 
to_sfixed(275126879.0/4294967296.0,1,-nbitq), 
to_sfixed(102614155.0/4294967296.0,1,-nbitq), 
to_sfixed(356310287.0/4294967296.0,1,-nbitq), 
to_sfixed(184852898.0/4294967296.0,1,-nbitq), 
to_sfixed(-368142343.0/4294967296.0,1,-nbitq), 
to_sfixed(119072218.0/4294967296.0,1,-nbitq), 
to_sfixed(-235179152.0/4294967296.0,1,-nbitq), 
to_sfixed(-137498651.0/4294967296.0,1,-nbitq), 
to_sfixed(-290556819.0/4294967296.0,1,-nbitq), 
to_sfixed(-307205971.0/4294967296.0,1,-nbitq), 
to_sfixed(-189147834.0/4294967296.0,1,-nbitq), 
to_sfixed(-424838911.0/4294967296.0,1,-nbitq), 
to_sfixed(-121774875.0/4294967296.0,1,-nbitq), 
to_sfixed(586520387.0/4294967296.0,1,-nbitq), 
to_sfixed(165363553.0/4294967296.0,1,-nbitq), 
to_sfixed(-397191177.0/4294967296.0,1,-nbitq), 
to_sfixed(-87801351.0/4294967296.0,1,-nbitq), 
to_sfixed(365299100.0/4294967296.0,1,-nbitq), 
to_sfixed(-341828027.0/4294967296.0,1,-nbitq), 
to_sfixed(262848229.0/4294967296.0,1,-nbitq), 
to_sfixed(497984768.0/4294967296.0,1,-nbitq), 
to_sfixed(344066264.0/4294967296.0,1,-nbitq), 
to_sfixed(-341910375.0/4294967296.0,1,-nbitq), 
to_sfixed(204137692.0/4294967296.0,1,-nbitq), 
to_sfixed(-383520420.0/4294967296.0,1,-nbitq), 
to_sfixed(8983721.0/4294967296.0,1,-nbitq), 
to_sfixed(11530670.0/4294967296.0,1,-nbitq), 
to_sfixed(204725629.0/4294967296.0,1,-nbitq), 
to_sfixed(-453497249.0/4294967296.0,1,-nbitq), 
to_sfixed(270090817.0/4294967296.0,1,-nbitq), 
to_sfixed(-292802556.0/4294967296.0,1,-nbitq), 
to_sfixed(-263407227.0/4294967296.0,1,-nbitq), 
to_sfixed(190678702.0/4294967296.0,1,-nbitq), 
to_sfixed(-1551070.0/4294967296.0,1,-nbitq), 
to_sfixed(361334701.0/4294967296.0,1,-nbitq), 
to_sfixed(-57447621.0/4294967296.0,1,-nbitq), 
to_sfixed(22556039.0/4294967296.0,1,-nbitq), 
to_sfixed(-191836284.0/4294967296.0,1,-nbitq), 
to_sfixed(-308434187.0/4294967296.0,1,-nbitq), 
to_sfixed(546079372.0/4294967296.0,1,-nbitq), 
to_sfixed(-221165353.0/4294967296.0,1,-nbitq), 
to_sfixed(180422600.0/4294967296.0,1,-nbitq), 
to_sfixed(19963385.0/4294967296.0,1,-nbitq), 
to_sfixed(-180182343.0/4294967296.0,1,-nbitq), 
to_sfixed(-247088684.0/4294967296.0,1,-nbitq), 
to_sfixed(-108346077.0/4294967296.0,1,-nbitq), 
to_sfixed(148709621.0/4294967296.0,1,-nbitq), 
to_sfixed(80759230.0/4294967296.0,1,-nbitq), 
to_sfixed(-92165416.0/4294967296.0,1,-nbitq), 
to_sfixed(166315772.0/4294967296.0,1,-nbitq), 
to_sfixed(-368211848.0/4294967296.0,1,-nbitq), 
to_sfixed(202222459.0/4294967296.0,1,-nbitq), 
to_sfixed(56759767.0/4294967296.0,1,-nbitq), 
to_sfixed(149647595.0/4294967296.0,1,-nbitq), 
to_sfixed(150624600.0/4294967296.0,1,-nbitq), 
to_sfixed(-286407064.0/4294967296.0,1,-nbitq), 
to_sfixed(14551939.0/4294967296.0,1,-nbitq), 
to_sfixed(-238753743.0/4294967296.0,1,-nbitq), 
to_sfixed(-224869696.0/4294967296.0,1,-nbitq), 
to_sfixed(30385077.0/4294967296.0,1,-nbitq), 
to_sfixed(-203326799.0/4294967296.0,1,-nbitq), 
to_sfixed(259815772.0/4294967296.0,1,-nbitq), 
to_sfixed(-384495363.0/4294967296.0,1,-nbitq), 
to_sfixed(41443052.0/4294967296.0,1,-nbitq), 
to_sfixed(-207425477.0/4294967296.0,1,-nbitq), 
to_sfixed(-244945801.0/4294967296.0,1,-nbitq), 
to_sfixed(-272625401.0/4294967296.0,1,-nbitq), 
to_sfixed(-328977034.0/4294967296.0,1,-nbitq), 
to_sfixed(-245659719.0/4294967296.0,1,-nbitq), 
to_sfixed(174755132.0/4294967296.0,1,-nbitq), 
to_sfixed(-19001617.0/4294967296.0,1,-nbitq), 
to_sfixed(99055138.0/4294967296.0,1,-nbitq), 
to_sfixed(-392334173.0/4294967296.0,1,-nbitq), 
to_sfixed(-260776558.0/4294967296.0,1,-nbitq), 
to_sfixed(354664804.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(132945796.0/4294967296.0,1,-nbitq), 
to_sfixed(-330285543.0/4294967296.0,1,-nbitq), 
to_sfixed(-276940294.0/4294967296.0,1,-nbitq), 
to_sfixed(-187522545.0/4294967296.0,1,-nbitq), 
to_sfixed(30157389.0/4294967296.0,1,-nbitq), 
to_sfixed(86393272.0/4294967296.0,1,-nbitq), 
to_sfixed(-344310076.0/4294967296.0,1,-nbitq), 
to_sfixed(370473464.0/4294967296.0,1,-nbitq), 
to_sfixed(210942061.0/4294967296.0,1,-nbitq), 
to_sfixed(-125549821.0/4294967296.0,1,-nbitq), 
to_sfixed(-31033593.0/4294967296.0,1,-nbitq), 
to_sfixed(-101307116.0/4294967296.0,1,-nbitq), 
to_sfixed(-222745275.0/4294967296.0,1,-nbitq), 
to_sfixed(28172529.0/4294967296.0,1,-nbitq), 
to_sfixed(-305941835.0/4294967296.0,1,-nbitq), 
to_sfixed(217289060.0/4294967296.0,1,-nbitq), 
to_sfixed(375606952.0/4294967296.0,1,-nbitq), 
to_sfixed(82605260.0/4294967296.0,1,-nbitq), 
to_sfixed(134014.0/4294967296.0,1,-nbitq), 
to_sfixed(76322184.0/4294967296.0,1,-nbitq), 
to_sfixed(120380821.0/4294967296.0,1,-nbitq), 
to_sfixed(409176664.0/4294967296.0,1,-nbitq), 
to_sfixed(629349615.0/4294967296.0,1,-nbitq), 
to_sfixed(32673266.0/4294967296.0,1,-nbitq), 
to_sfixed(75119491.0/4294967296.0,1,-nbitq), 
to_sfixed(116174630.0/4294967296.0,1,-nbitq), 
to_sfixed(173747285.0/4294967296.0,1,-nbitq), 
to_sfixed(191029143.0/4294967296.0,1,-nbitq), 
to_sfixed(274099274.0/4294967296.0,1,-nbitq), 
to_sfixed(-443045454.0/4294967296.0,1,-nbitq), 
to_sfixed(62335511.0/4294967296.0,1,-nbitq), 
to_sfixed(220468682.0/4294967296.0,1,-nbitq), 
to_sfixed(-18175614.0/4294967296.0,1,-nbitq), 
to_sfixed(173000757.0/4294967296.0,1,-nbitq), 
to_sfixed(337660946.0/4294967296.0,1,-nbitq), 
to_sfixed(-440604133.0/4294967296.0,1,-nbitq), 
to_sfixed(267466861.0/4294967296.0,1,-nbitq), 
to_sfixed(199787407.0/4294967296.0,1,-nbitq), 
to_sfixed(-19977419.0/4294967296.0,1,-nbitq), 
to_sfixed(-90654.0/4294967296.0,1,-nbitq), 
to_sfixed(-319571668.0/4294967296.0,1,-nbitq), 
to_sfixed(273470689.0/4294967296.0,1,-nbitq), 
to_sfixed(207020382.0/4294967296.0,1,-nbitq), 
to_sfixed(78807909.0/4294967296.0,1,-nbitq), 
to_sfixed(24437402.0/4294967296.0,1,-nbitq), 
to_sfixed(326416752.0/4294967296.0,1,-nbitq), 
to_sfixed(-424247677.0/4294967296.0,1,-nbitq), 
to_sfixed(-204949874.0/4294967296.0,1,-nbitq), 
to_sfixed(309694541.0/4294967296.0,1,-nbitq), 
to_sfixed(344326285.0/4294967296.0,1,-nbitq), 
to_sfixed(259377416.0/4294967296.0,1,-nbitq), 
to_sfixed(410749634.0/4294967296.0,1,-nbitq), 
to_sfixed(-390937440.0/4294967296.0,1,-nbitq), 
to_sfixed(478096485.0/4294967296.0,1,-nbitq), 
to_sfixed(46838020.0/4294967296.0,1,-nbitq), 
to_sfixed(-289481759.0/4294967296.0,1,-nbitq), 
to_sfixed(-157376850.0/4294967296.0,1,-nbitq), 
to_sfixed(-491402723.0/4294967296.0,1,-nbitq), 
to_sfixed(-303293908.0/4294967296.0,1,-nbitq), 
to_sfixed(-252949244.0/4294967296.0,1,-nbitq), 
to_sfixed(-89621763.0/4294967296.0,1,-nbitq), 
to_sfixed(346394878.0/4294967296.0,1,-nbitq), 
to_sfixed(-294082219.0/4294967296.0,1,-nbitq), 
to_sfixed(-412981123.0/4294967296.0,1,-nbitq), 
to_sfixed(404056866.0/4294967296.0,1,-nbitq), 
to_sfixed(128913538.0/4294967296.0,1,-nbitq), 
to_sfixed(376692302.0/4294967296.0,1,-nbitq), 
to_sfixed(309770198.0/4294967296.0,1,-nbitq), 
to_sfixed(-235771625.0/4294967296.0,1,-nbitq), 
to_sfixed(196203807.0/4294967296.0,1,-nbitq), 
to_sfixed(-320951699.0/4294967296.0,1,-nbitq), 
to_sfixed(-272807274.0/4294967296.0,1,-nbitq), 
to_sfixed(-115022185.0/4294967296.0,1,-nbitq), 
to_sfixed(618482.0/4294967296.0,1,-nbitq), 
to_sfixed(523376478.0/4294967296.0,1,-nbitq), 
to_sfixed(-444385806.0/4294967296.0,1,-nbitq), 
to_sfixed(-366816679.0/4294967296.0,1,-nbitq), 
to_sfixed(-169371608.0/4294967296.0,1,-nbitq), 
to_sfixed(-504348838.0/4294967296.0,1,-nbitq), 
to_sfixed(-195165068.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-187649142.0/4294967296.0,1,-nbitq), 
to_sfixed(-239260615.0/4294967296.0,1,-nbitq), 
to_sfixed(-231094311.0/4294967296.0,1,-nbitq), 
to_sfixed(-251596024.0/4294967296.0,1,-nbitq), 
to_sfixed(-46871086.0/4294967296.0,1,-nbitq), 
to_sfixed(-322475989.0/4294967296.0,1,-nbitq), 
to_sfixed(-331640114.0/4294967296.0,1,-nbitq), 
to_sfixed(-90991717.0/4294967296.0,1,-nbitq), 
to_sfixed(-315725900.0/4294967296.0,1,-nbitq), 
to_sfixed(139551560.0/4294967296.0,1,-nbitq), 
to_sfixed(-352697131.0/4294967296.0,1,-nbitq), 
to_sfixed(-49831715.0/4294967296.0,1,-nbitq), 
to_sfixed(128843444.0/4294967296.0,1,-nbitq), 
to_sfixed(365498906.0/4294967296.0,1,-nbitq), 
to_sfixed(-14131437.0/4294967296.0,1,-nbitq), 
to_sfixed(175501182.0/4294967296.0,1,-nbitq), 
to_sfixed(-419809429.0/4294967296.0,1,-nbitq), 
to_sfixed(-334196806.0/4294967296.0,1,-nbitq), 
to_sfixed(614776639.0/4294967296.0,1,-nbitq), 
to_sfixed(-449683626.0/4294967296.0,1,-nbitq), 
to_sfixed(-196545340.0/4294967296.0,1,-nbitq), 
to_sfixed(158771854.0/4294967296.0,1,-nbitq), 
to_sfixed(502653996.0/4294967296.0,1,-nbitq), 
to_sfixed(33900564.0/4294967296.0,1,-nbitq), 
to_sfixed(260728892.0/4294967296.0,1,-nbitq), 
to_sfixed(372578901.0/4294967296.0,1,-nbitq), 
to_sfixed(184289802.0/4294967296.0,1,-nbitq), 
to_sfixed(-202211059.0/4294967296.0,1,-nbitq), 
to_sfixed(-221960602.0/4294967296.0,1,-nbitq), 
to_sfixed(211584146.0/4294967296.0,1,-nbitq), 
to_sfixed(45142209.0/4294967296.0,1,-nbitq), 
to_sfixed(-311777379.0/4294967296.0,1,-nbitq), 
to_sfixed(-134856387.0/4294967296.0,1,-nbitq), 
to_sfixed(213268229.0/4294967296.0,1,-nbitq), 
to_sfixed(408412523.0/4294967296.0,1,-nbitq), 
to_sfixed(54033968.0/4294967296.0,1,-nbitq), 
to_sfixed(235166953.0/4294967296.0,1,-nbitq), 
to_sfixed(61979040.0/4294967296.0,1,-nbitq), 
to_sfixed(-173822960.0/4294967296.0,1,-nbitq), 
to_sfixed(433121192.0/4294967296.0,1,-nbitq), 
to_sfixed(141931719.0/4294967296.0,1,-nbitq), 
to_sfixed(117236002.0/4294967296.0,1,-nbitq), 
to_sfixed(383478744.0/4294967296.0,1,-nbitq), 
to_sfixed(-2549668.0/4294967296.0,1,-nbitq), 
to_sfixed(-27194144.0/4294967296.0,1,-nbitq), 
to_sfixed(-45584553.0/4294967296.0,1,-nbitq), 
to_sfixed(-319014343.0/4294967296.0,1,-nbitq), 
to_sfixed(-206634780.0/4294967296.0,1,-nbitq), 
to_sfixed(150419009.0/4294967296.0,1,-nbitq), 
to_sfixed(-195437016.0/4294967296.0,1,-nbitq), 
to_sfixed(-12566981.0/4294967296.0,1,-nbitq), 
to_sfixed(-49073109.0/4294967296.0,1,-nbitq), 
to_sfixed(-602693948.0/4294967296.0,1,-nbitq), 
to_sfixed(222079421.0/4294967296.0,1,-nbitq), 
to_sfixed(-149816047.0/4294967296.0,1,-nbitq), 
to_sfixed(-128126801.0/4294967296.0,1,-nbitq), 
to_sfixed(369632123.0/4294967296.0,1,-nbitq), 
to_sfixed(-466986683.0/4294967296.0,1,-nbitq), 
to_sfixed(-359825169.0/4294967296.0,1,-nbitq), 
to_sfixed(-355542635.0/4294967296.0,1,-nbitq), 
to_sfixed(119174277.0/4294967296.0,1,-nbitq), 
to_sfixed(313043347.0/4294967296.0,1,-nbitq), 
to_sfixed(-45314312.0/4294967296.0,1,-nbitq), 
to_sfixed(-380902098.0/4294967296.0,1,-nbitq), 
to_sfixed(-261361504.0/4294967296.0,1,-nbitq), 
to_sfixed(-54048074.0/4294967296.0,1,-nbitq), 
to_sfixed(111977962.0/4294967296.0,1,-nbitq), 
to_sfixed(73663872.0/4294967296.0,1,-nbitq), 
to_sfixed(-319406830.0/4294967296.0,1,-nbitq), 
to_sfixed(138630713.0/4294967296.0,1,-nbitq), 
to_sfixed(-15367535.0/4294967296.0,1,-nbitq), 
to_sfixed(199711616.0/4294967296.0,1,-nbitq), 
to_sfixed(58553651.0/4294967296.0,1,-nbitq), 
to_sfixed(177940244.0/4294967296.0,1,-nbitq), 
to_sfixed(-27674459.0/4294967296.0,1,-nbitq), 
to_sfixed(-261718460.0/4294967296.0,1,-nbitq), 
to_sfixed(-126263684.0/4294967296.0,1,-nbitq), 
to_sfixed(255794147.0/4294967296.0,1,-nbitq), 
to_sfixed(-74934118.0/4294967296.0,1,-nbitq), 
to_sfixed(526186.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(214368097.0/4294967296.0,1,-nbitq), 
to_sfixed(151737188.0/4294967296.0,1,-nbitq), 
to_sfixed(-74746821.0/4294967296.0,1,-nbitq), 
to_sfixed(-84729745.0/4294967296.0,1,-nbitq), 
to_sfixed(-86435596.0/4294967296.0,1,-nbitq), 
to_sfixed(-395361416.0/4294967296.0,1,-nbitq), 
to_sfixed(-296998039.0/4294967296.0,1,-nbitq), 
to_sfixed(-271286599.0/4294967296.0,1,-nbitq), 
to_sfixed(272771105.0/4294967296.0,1,-nbitq), 
to_sfixed(233989607.0/4294967296.0,1,-nbitq), 
to_sfixed(-107880895.0/4294967296.0,1,-nbitq), 
to_sfixed(307966062.0/4294967296.0,1,-nbitq), 
to_sfixed(-124558413.0/4294967296.0,1,-nbitq), 
to_sfixed(-12263023.0/4294967296.0,1,-nbitq), 
to_sfixed(303600269.0/4294967296.0,1,-nbitq), 
to_sfixed(-202132133.0/4294967296.0,1,-nbitq), 
to_sfixed(-314238869.0/4294967296.0,1,-nbitq), 
to_sfixed(198734371.0/4294967296.0,1,-nbitq), 
to_sfixed(-53500401.0/4294967296.0,1,-nbitq), 
to_sfixed(62772855.0/4294967296.0,1,-nbitq), 
to_sfixed(354757285.0/4294967296.0,1,-nbitq), 
to_sfixed(503145589.0/4294967296.0,1,-nbitq), 
to_sfixed(500363399.0/4294967296.0,1,-nbitq), 
to_sfixed(236554434.0/4294967296.0,1,-nbitq), 
to_sfixed(-86427287.0/4294967296.0,1,-nbitq), 
to_sfixed(183425673.0/4294967296.0,1,-nbitq), 
to_sfixed(-279558246.0/4294967296.0,1,-nbitq), 
to_sfixed(-339728093.0/4294967296.0,1,-nbitq), 
to_sfixed(-162595944.0/4294967296.0,1,-nbitq), 
to_sfixed(327606994.0/4294967296.0,1,-nbitq), 
to_sfixed(-508181996.0/4294967296.0,1,-nbitq), 
to_sfixed(-468815343.0/4294967296.0,1,-nbitq), 
to_sfixed(289371350.0/4294967296.0,1,-nbitq), 
to_sfixed(-398611863.0/4294967296.0,1,-nbitq), 
to_sfixed(-102154236.0/4294967296.0,1,-nbitq), 
to_sfixed(-276639691.0/4294967296.0,1,-nbitq), 
to_sfixed(-243657264.0/4294967296.0,1,-nbitq), 
to_sfixed(-235529118.0/4294967296.0,1,-nbitq), 
to_sfixed(305695813.0/4294967296.0,1,-nbitq), 
to_sfixed(152640138.0/4294967296.0,1,-nbitq), 
to_sfixed(-207001483.0/4294967296.0,1,-nbitq), 
to_sfixed(-48129891.0/4294967296.0,1,-nbitq), 
to_sfixed(-393221775.0/4294967296.0,1,-nbitq), 
to_sfixed(16906052.0/4294967296.0,1,-nbitq), 
to_sfixed(185567601.0/4294967296.0,1,-nbitq), 
to_sfixed(-30189060.0/4294967296.0,1,-nbitq), 
to_sfixed(289199951.0/4294967296.0,1,-nbitq), 
to_sfixed(-283024223.0/4294967296.0,1,-nbitq), 
to_sfixed(-103506301.0/4294967296.0,1,-nbitq), 
to_sfixed(-200760028.0/4294967296.0,1,-nbitq), 
to_sfixed(-17426110.0/4294967296.0,1,-nbitq), 
to_sfixed(400645027.0/4294967296.0,1,-nbitq), 
to_sfixed(-556098126.0/4294967296.0,1,-nbitq), 
to_sfixed(-38082863.0/4294967296.0,1,-nbitq), 
to_sfixed(199210538.0/4294967296.0,1,-nbitq), 
to_sfixed(146936963.0/4294967296.0,1,-nbitq), 
to_sfixed(342175700.0/4294967296.0,1,-nbitq), 
to_sfixed(-165803866.0/4294967296.0,1,-nbitq), 
to_sfixed(41856519.0/4294967296.0,1,-nbitq), 
to_sfixed(401535505.0/4294967296.0,1,-nbitq), 
to_sfixed(-296662204.0/4294967296.0,1,-nbitq), 
to_sfixed(271014202.0/4294967296.0,1,-nbitq), 
to_sfixed(-265222953.0/4294967296.0,1,-nbitq), 
to_sfixed(23228863.0/4294967296.0,1,-nbitq), 
to_sfixed(-140317279.0/4294967296.0,1,-nbitq), 
to_sfixed(-87095295.0/4294967296.0,1,-nbitq), 
to_sfixed(747377727.0/4294967296.0,1,-nbitq), 
to_sfixed(-57084978.0/4294967296.0,1,-nbitq), 
to_sfixed(-140050293.0/4294967296.0,1,-nbitq), 
to_sfixed(33027264.0/4294967296.0,1,-nbitq), 
to_sfixed(51127820.0/4294967296.0,1,-nbitq), 
to_sfixed(-30946104.0/4294967296.0,1,-nbitq), 
to_sfixed(-342087530.0/4294967296.0,1,-nbitq), 
to_sfixed(341131908.0/4294967296.0,1,-nbitq), 
to_sfixed(52559535.0/4294967296.0,1,-nbitq), 
to_sfixed(-398742062.0/4294967296.0,1,-nbitq), 
to_sfixed(61648559.0/4294967296.0,1,-nbitq), 
to_sfixed(235980813.0/4294967296.0,1,-nbitq), 
to_sfixed(-469879008.0/4294967296.0,1,-nbitq), 
to_sfixed(215637185.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-189669970.0/4294967296.0,1,-nbitq), 
to_sfixed(153540073.0/4294967296.0,1,-nbitq), 
to_sfixed(35044692.0/4294967296.0,1,-nbitq), 
to_sfixed(81985947.0/4294967296.0,1,-nbitq), 
to_sfixed(244544871.0/4294967296.0,1,-nbitq), 
to_sfixed(240949071.0/4294967296.0,1,-nbitq), 
to_sfixed(255593926.0/4294967296.0,1,-nbitq), 
to_sfixed(135225292.0/4294967296.0,1,-nbitq), 
to_sfixed(-430860039.0/4294967296.0,1,-nbitq), 
to_sfixed(48711820.0/4294967296.0,1,-nbitq), 
to_sfixed(-348665018.0/4294967296.0,1,-nbitq), 
to_sfixed(122227332.0/4294967296.0,1,-nbitq), 
to_sfixed(-132582843.0/4294967296.0,1,-nbitq), 
to_sfixed(383028179.0/4294967296.0,1,-nbitq), 
to_sfixed(147356916.0/4294967296.0,1,-nbitq), 
to_sfixed(322036325.0/4294967296.0,1,-nbitq), 
to_sfixed(-74833689.0/4294967296.0,1,-nbitq), 
to_sfixed(-165651628.0/4294967296.0,1,-nbitq), 
to_sfixed(367376540.0/4294967296.0,1,-nbitq), 
to_sfixed(-243483587.0/4294967296.0,1,-nbitq), 
to_sfixed(-336372729.0/4294967296.0,1,-nbitq), 
to_sfixed(307710848.0/4294967296.0,1,-nbitq), 
to_sfixed(59496584.0/4294967296.0,1,-nbitq), 
to_sfixed(271537915.0/4294967296.0,1,-nbitq), 
to_sfixed(197535328.0/4294967296.0,1,-nbitq), 
to_sfixed(51462019.0/4294967296.0,1,-nbitq), 
to_sfixed(-24298162.0/4294967296.0,1,-nbitq), 
to_sfixed(-184507966.0/4294967296.0,1,-nbitq), 
to_sfixed(-190451086.0/4294967296.0,1,-nbitq), 
to_sfixed(-124423318.0/4294967296.0,1,-nbitq), 
to_sfixed(-471649580.0/4294967296.0,1,-nbitq), 
to_sfixed(-377661182.0/4294967296.0,1,-nbitq), 
to_sfixed(135650296.0/4294967296.0,1,-nbitq), 
to_sfixed(-512339772.0/4294967296.0,1,-nbitq), 
to_sfixed(445771170.0/4294967296.0,1,-nbitq), 
to_sfixed(273144190.0/4294967296.0,1,-nbitq), 
to_sfixed(140277685.0/4294967296.0,1,-nbitq), 
to_sfixed(20985935.0/4294967296.0,1,-nbitq), 
to_sfixed(252410742.0/4294967296.0,1,-nbitq), 
to_sfixed(218818597.0/4294967296.0,1,-nbitq), 
to_sfixed(-149981059.0/4294967296.0,1,-nbitq), 
to_sfixed(16114701.0/4294967296.0,1,-nbitq), 
to_sfixed(378910287.0/4294967296.0,1,-nbitq), 
to_sfixed(-368949984.0/4294967296.0,1,-nbitq), 
to_sfixed(-71492988.0/4294967296.0,1,-nbitq), 
to_sfixed(188159880.0/4294967296.0,1,-nbitq), 
to_sfixed(141779332.0/4294967296.0,1,-nbitq), 
to_sfixed(-265592110.0/4294967296.0,1,-nbitq), 
to_sfixed(-102541193.0/4294967296.0,1,-nbitq), 
to_sfixed(358887041.0/4294967296.0,1,-nbitq), 
to_sfixed(-323486571.0/4294967296.0,1,-nbitq), 
to_sfixed(-48515843.0/4294967296.0,1,-nbitq), 
to_sfixed(-586841493.0/4294967296.0,1,-nbitq), 
to_sfixed(-92240337.0/4294967296.0,1,-nbitq), 
to_sfixed(373003449.0/4294967296.0,1,-nbitq), 
to_sfixed(153745382.0/4294967296.0,1,-nbitq), 
to_sfixed(-74144827.0/4294967296.0,1,-nbitq), 
to_sfixed(-369962004.0/4294967296.0,1,-nbitq), 
to_sfixed(-224902267.0/4294967296.0,1,-nbitq), 
to_sfixed(-360605874.0/4294967296.0,1,-nbitq), 
to_sfixed(154778855.0/4294967296.0,1,-nbitq), 
to_sfixed(224040540.0/4294967296.0,1,-nbitq), 
to_sfixed(-51581806.0/4294967296.0,1,-nbitq), 
to_sfixed(410078961.0/4294967296.0,1,-nbitq), 
to_sfixed(34541703.0/4294967296.0,1,-nbitq), 
to_sfixed(-370836138.0/4294967296.0,1,-nbitq), 
to_sfixed(633133215.0/4294967296.0,1,-nbitq), 
to_sfixed(253206007.0/4294967296.0,1,-nbitq), 
to_sfixed(182668540.0/4294967296.0,1,-nbitq), 
to_sfixed(542300026.0/4294967296.0,1,-nbitq), 
to_sfixed(-313069430.0/4294967296.0,1,-nbitq), 
to_sfixed(155679970.0/4294967296.0,1,-nbitq), 
to_sfixed(251647835.0/4294967296.0,1,-nbitq), 
to_sfixed(146141816.0/4294967296.0,1,-nbitq), 
to_sfixed(180779349.0/4294967296.0,1,-nbitq), 
to_sfixed(-213829182.0/4294967296.0,1,-nbitq), 
to_sfixed(3797351.0/4294967296.0,1,-nbitq), 
to_sfixed(110280473.0/4294967296.0,1,-nbitq), 
to_sfixed(-120983615.0/4294967296.0,1,-nbitq), 
to_sfixed(-221529664.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(312561542.0/4294967296.0,1,-nbitq), 
to_sfixed(58338396.0/4294967296.0,1,-nbitq), 
to_sfixed(-35773734.0/4294967296.0,1,-nbitq), 
to_sfixed(-151575483.0/4294967296.0,1,-nbitq), 
to_sfixed(288682430.0/4294967296.0,1,-nbitq), 
to_sfixed(-186883851.0/4294967296.0,1,-nbitq), 
to_sfixed(242684092.0/4294967296.0,1,-nbitq), 
to_sfixed(283574216.0/4294967296.0,1,-nbitq), 
to_sfixed(-415472888.0/4294967296.0,1,-nbitq), 
to_sfixed(-325205854.0/4294967296.0,1,-nbitq), 
to_sfixed(130693725.0/4294967296.0,1,-nbitq), 
to_sfixed(94868577.0/4294967296.0,1,-nbitq), 
to_sfixed(-168964923.0/4294967296.0,1,-nbitq), 
to_sfixed(401214162.0/4294967296.0,1,-nbitq), 
to_sfixed(64007632.0/4294967296.0,1,-nbitq), 
to_sfixed(-401863461.0/4294967296.0,1,-nbitq), 
to_sfixed(80119376.0/4294967296.0,1,-nbitq), 
to_sfixed(-339961186.0/4294967296.0,1,-nbitq), 
to_sfixed(489228669.0/4294967296.0,1,-nbitq), 
to_sfixed(260334341.0/4294967296.0,1,-nbitq), 
to_sfixed(-37521905.0/4294967296.0,1,-nbitq), 
to_sfixed(417570814.0/4294967296.0,1,-nbitq), 
to_sfixed(242273244.0/4294967296.0,1,-nbitq), 
to_sfixed(-200072783.0/4294967296.0,1,-nbitq), 
to_sfixed(17040778.0/4294967296.0,1,-nbitq), 
to_sfixed(8162347.0/4294967296.0,1,-nbitq), 
to_sfixed(181862593.0/4294967296.0,1,-nbitq), 
to_sfixed(-120928499.0/4294967296.0,1,-nbitq), 
to_sfixed(7993340.0/4294967296.0,1,-nbitq), 
to_sfixed(-33893171.0/4294967296.0,1,-nbitq), 
to_sfixed(-223848043.0/4294967296.0,1,-nbitq), 
to_sfixed(-356944249.0/4294967296.0,1,-nbitq), 
to_sfixed(-230513126.0/4294967296.0,1,-nbitq), 
to_sfixed(-367404933.0/4294967296.0,1,-nbitq), 
to_sfixed(290117702.0/4294967296.0,1,-nbitq), 
to_sfixed(-392516318.0/4294967296.0,1,-nbitq), 
to_sfixed(-254391318.0/4294967296.0,1,-nbitq), 
to_sfixed(25770083.0/4294967296.0,1,-nbitq), 
to_sfixed(-33030284.0/4294967296.0,1,-nbitq), 
to_sfixed(186655155.0/4294967296.0,1,-nbitq), 
to_sfixed(-157182739.0/4294967296.0,1,-nbitq), 
to_sfixed(-11365726.0/4294967296.0,1,-nbitq), 
to_sfixed(172826314.0/4294967296.0,1,-nbitq), 
to_sfixed(181963054.0/4294967296.0,1,-nbitq), 
to_sfixed(423033281.0/4294967296.0,1,-nbitq), 
to_sfixed(398571790.0/4294967296.0,1,-nbitq), 
to_sfixed(-162830622.0/4294967296.0,1,-nbitq), 
to_sfixed(-233009523.0/4294967296.0,1,-nbitq), 
to_sfixed(-420347924.0/4294967296.0,1,-nbitq), 
to_sfixed(377887633.0/4294967296.0,1,-nbitq), 
to_sfixed(-84911514.0/4294967296.0,1,-nbitq), 
to_sfixed(-77169640.0/4294967296.0,1,-nbitq), 
to_sfixed(70244413.0/4294967296.0,1,-nbitq), 
to_sfixed(64412557.0/4294967296.0,1,-nbitq), 
to_sfixed(7308608.0/4294967296.0,1,-nbitq), 
to_sfixed(148753660.0/4294967296.0,1,-nbitq), 
to_sfixed(269695749.0/4294967296.0,1,-nbitq), 
to_sfixed(-557334065.0/4294967296.0,1,-nbitq), 
to_sfixed(-313182700.0/4294967296.0,1,-nbitq), 
to_sfixed(166999491.0/4294967296.0,1,-nbitq), 
to_sfixed(191084863.0/4294967296.0,1,-nbitq), 
to_sfixed(30785315.0/4294967296.0,1,-nbitq), 
to_sfixed(-291008118.0/4294967296.0,1,-nbitq), 
to_sfixed(216631949.0/4294967296.0,1,-nbitq), 
to_sfixed(-226666259.0/4294967296.0,1,-nbitq), 
to_sfixed(224749863.0/4294967296.0,1,-nbitq), 
to_sfixed(199584705.0/4294967296.0,1,-nbitq), 
to_sfixed(-185183976.0/4294967296.0,1,-nbitq), 
to_sfixed(127526451.0/4294967296.0,1,-nbitq), 
to_sfixed(238919926.0/4294967296.0,1,-nbitq), 
to_sfixed(153069302.0/4294967296.0,1,-nbitq), 
to_sfixed(-150644884.0/4294967296.0,1,-nbitq), 
to_sfixed(-414296885.0/4294967296.0,1,-nbitq), 
to_sfixed(-201043948.0/4294967296.0,1,-nbitq), 
to_sfixed(99291928.0/4294967296.0,1,-nbitq), 
to_sfixed(-528662267.0/4294967296.0,1,-nbitq), 
to_sfixed(210091807.0/4294967296.0,1,-nbitq), 
to_sfixed(-353175585.0/4294967296.0,1,-nbitq), 
to_sfixed(-326752011.0/4294967296.0,1,-nbitq), 
to_sfixed(318869184.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(293389809.0/4294967296.0,1,-nbitq), 
to_sfixed(-379347799.0/4294967296.0,1,-nbitq), 
to_sfixed(355583633.0/4294967296.0,1,-nbitq), 
to_sfixed(272280020.0/4294967296.0,1,-nbitq), 
to_sfixed(-29061340.0/4294967296.0,1,-nbitq), 
to_sfixed(-348485651.0/4294967296.0,1,-nbitq), 
to_sfixed(140704931.0/4294967296.0,1,-nbitq), 
to_sfixed(-111963170.0/4294967296.0,1,-nbitq), 
to_sfixed(222689751.0/4294967296.0,1,-nbitq), 
to_sfixed(-342538651.0/4294967296.0,1,-nbitq), 
to_sfixed(357358252.0/4294967296.0,1,-nbitq), 
to_sfixed(138915536.0/4294967296.0,1,-nbitq), 
to_sfixed(-65233538.0/4294967296.0,1,-nbitq), 
to_sfixed(-93092260.0/4294967296.0,1,-nbitq), 
to_sfixed(-398406955.0/4294967296.0,1,-nbitq), 
to_sfixed(42354185.0/4294967296.0,1,-nbitq), 
to_sfixed(35848354.0/4294967296.0,1,-nbitq), 
to_sfixed(-254565872.0/4294967296.0,1,-nbitq), 
to_sfixed(303169911.0/4294967296.0,1,-nbitq), 
to_sfixed(348592008.0/4294967296.0,1,-nbitq), 
to_sfixed(152257410.0/4294967296.0,1,-nbitq), 
to_sfixed(217133463.0/4294967296.0,1,-nbitq), 
to_sfixed(562465634.0/4294967296.0,1,-nbitq), 
to_sfixed(-109032048.0/4294967296.0,1,-nbitq), 
to_sfixed(-45252786.0/4294967296.0,1,-nbitq), 
to_sfixed(504831935.0/4294967296.0,1,-nbitq), 
to_sfixed(327319244.0/4294967296.0,1,-nbitq), 
to_sfixed(-619220284.0/4294967296.0,1,-nbitq), 
to_sfixed(156421429.0/4294967296.0,1,-nbitq), 
to_sfixed(-135583988.0/4294967296.0,1,-nbitq), 
to_sfixed(-83913747.0/4294967296.0,1,-nbitq), 
to_sfixed(-16330871.0/4294967296.0,1,-nbitq), 
to_sfixed(17216436.0/4294967296.0,1,-nbitq), 
to_sfixed(191443839.0/4294967296.0,1,-nbitq), 
to_sfixed(80793269.0/4294967296.0,1,-nbitq), 
to_sfixed(202389044.0/4294967296.0,1,-nbitq), 
to_sfixed(30451054.0/4294967296.0,1,-nbitq), 
to_sfixed(-59102364.0/4294967296.0,1,-nbitq), 
to_sfixed(137264570.0/4294967296.0,1,-nbitq), 
to_sfixed(396011595.0/4294967296.0,1,-nbitq), 
to_sfixed(-210185267.0/4294967296.0,1,-nbitq), 
to_sfixed(309178971.0/4294967296.0,1,-nbitq), 
to_sfixed(11312643.0/4294967296.0,1,-nbitq), 
to_sfixed(-73930602.0/4294967296.0,1,-nbitq), 
to_sfixed(44086623.0/4294967296.0,1,-nbitq), 
to_sfixed(259894352.0/4294967296.0,1,-nbitq), 
to_sfixed(-403127296.0/4294967296.0,1,-nbitq), 
to_sfixed(-192723606.0/4294967296.0,1,-nbitq), 
to_sfixed(-73180797.0/4294967296.0,1,-nbitq), 
to_sfixed(150633776.0/4294967296.0,1,-nbitq), 
to_sfixed(-79337362.0/4294967296.0,1,-nbitq), 
to_sfixed(-227188588.0/4294967296.0,1,-nbitq), 
to_sfixed(-622677692.0/4294967296.0,1,-nbitq), 
to_sfixed(-215947962.0/4294967296.0,1,-nbitq), 
to_sfixed(338088813.0/4294967296.0,1,-nbitq), 
to_sfixed(350780086.0/4294967296.0,1,-nbitq), 
to_sfixed(-109623040.0/4294967296.0,1,-nbitq), 
to_sfixed(-57223434.0/4294967296.0,1,-nbitq), 
to_sfixed(113444654.0/4294967296.0,1,-nbitq), 
to_sfixed(-215733702.0/4294967296.0,1,-nbitq), 
to_sfixed(90418117.0/4294967296.0,1,-nbitq), 
to_sfixed(219248833.0/4294967296.0,1,-nbitq), 
to_sfixed(-409395365.0/4294967296.0,1,-nbitq), 
to_sfixed(-143419871.0/4294967296.0,1,-nbitq), 
to_sfixed(-69403472.0/4294967296.0,1,-nbitq), 
to_sfixed(-113396867.0/4294967296.0,1,-nbitq), 
to_sfixed(723006128.0/4294967296.0,1,-nbitq), 
to_sfixed(168533523.0/4294967296.0,1,-nbitq), 
to_sfixed(143937895.0/4294967296.0,1,-nbitq), 
to_sfixed(-17917884.0/4294967296.0,1,-nbitq), 
to_sfixed(158290906.0/4294967296.0,1,-nbitq), 
to_sfixed(-346090463.0/4294967296.0,1,-nbitq), 
to_sfixed(-150989174.0/4294967296.0,1,-nbitq), 
to_sfixed(-259966592.0/4294967296.0,1,-nbitq), 
to_sfixed(-264634281.0/4294967296.0,1,-nbitq), 
to_sfixed(-244632796.0/4294967296.0,1,-nbitq), 
to_sfixed(-184608280.0/4294967296.0,1,-nbitq), 
to_sfixed(-211034780.0/4294967296.0,1,-nbitq), 
to_sfixed(-399338286.0/4294967296.0,1,-nbitq), 
to_sfixed(-181155640.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(8878476.0/4294967296.0,1,-nbitq), 
to_sfixed(-355866221.0/4294967296.0,1,-nbitq), 
to_sfixed(-133160799.0/4294967296.0,1,-nbitq), 
to_sfixed(211183099.0/4294967296.0,1,-nbitq), 
to_sfixed(-160067646.0/4294967296.0,1,-nbitq), 
to_sfixed(-112417181.0/4294967296.0,1,-nbitq), 
to_sfixed(109271295.0/4294967296.0,1,-nbitq), 
to_sfixed(378304022.0/4294967296.0,1,-nbitq), 
to_sfixed(-435551468.0/4294967296.0,1,-nbitq), 
to_sfixed(215133099.0/4294967296.0,1,-nbitq), 
to_sfixed(-363370079.0/4294967296.0,1,-nbitq), 
to_sfixed(239482908.0/4294967296.0,1,-nbitq), 
to_sfixed(-35659811.0/4294967296.0,1,-nbitq), 
to_sfixed(324825145.0/4294967296.0,1,-nbitq), 
to_sfixed(-274567723.0/4294967296.0,1,-nbitq), 
to_sfixed(-267650114.0/4294967296.0,1,-nbitq), 
to_sfixed(-99803897.0/4294967296.0,1,-nbitq), 
to_sfixed(85267348.0/4294967296.0,1,-nbitq), 
to_sfixed(153967297.0/4294967296.0,1,-nbitq), 
to_sfixed(311776105.0/4294967296.0,1,-nbitq), 
to_sfixed(363012101.0/4294967296.0,1,-nbitq), 
to_sfixed(85433559.0/4294967296.0,1,-nbitq), 
to_sfixed(-137031779.0/4294967296.0,1,-nbitq), 
to_sfixed(276601849.0/4294967296.0,1,-nbitq), 
to_sfixed(229052863.0/4294967296.0,1,-nbitq), 
to_sfixed(132434628.0/4294967296.0,1,-nbitq), 
to_sfixed(312584278.0/4294967296.0,1,-nbitq), 
to_sfixed(-519756893.0/4294967296.0,1,-nbitq), 
to_sfixed(471440045.0/4294967296.0,1,-nbitq), 
to_sfixed(4390492.0/4294967296.0,1,-nbitq), 
to_sfixed(-38804482.0/4294967296.0,1,-nbitq), 
to_sfixed(-157700857.0/4294967296.0,1,-nbitq), 
to_sfixed(364694463.0/4294967296.0,1,-nbitq), 
to_sfixed(-283345602.0/4294967296.0,1,-nbitq), 
to_sfixed(89318410.0/4294967296.0,1,-nbitq), 
to_sfixed(-236776211.0/4294967296.0,1,-nbitq), 
to_sfixed(-290147976.0/4294967296.0,1,-nbitq), 
to_sfixed(442418462.0/4294967296.0,1,-nbitq), 
to_sfixed(79379386.0/4294967296.0,1,-nbitq), 
to_sfixed(483990958.0/4294967296.0,1,-nbitq), 
to_sfixed(-191722818.0/4294967296.0,1,-nbitq), 
to_sfixed(-290787127.0/4294967296.0,1,-nbitq), 
to_sfixed(-48802412.0/4294967296.0,1,-nbitq), 
to_sfixed(96752615.0/4294967296.0,1,-nbitq), 
to_sfixed(-99541371.0/4294967296.0,1,-nbitq), 
to_sfixed(213582437.0/4294967296.0,1,-nbitq), 
to_sfixed(-417885951.0/4294967296.0,1,-nbitq), 
to_sfixed(-336064857.0/4294967296.0,1,-nbitq), 
to_sfixed(-52102632.0/4294967296.0,1,-nbitq), 
to_sfixed(113519847.0/4294967296.0,1,-nbitq), 
to_sfixed(-188004193.0/4294967296.0,1,-nbitq), 
to_sfixed(-94262841.0/4294967296.0,1,-nbitq), 
to_sfixed(-229490341.0/4294967296.0,1,-nbitq), 
to_sfixed(-218869880.0/4294967296.0,1,-nbitq), 
to_sfixed(40451526.0/4294967296.0,1,-nbitq), 
to_sfixed(-428661844.0/4294967296.0,1,-nbitq), 
to_sfixed(-258306037.0/4294967296.0,1,-nbitq), 
to_sfixed(-92884618.0/4294967296.0,1,-nbitq), 
to_sfixed(-146461088.0/4294967296.0,1,-nbitq), 
to_sfixed(43764532.0/4294967296.0,1,-nbitq), 
to_sfixed(-331149159.0/4294967296.0,1,-nbitq), 
to_sfixed(-91576873.0/4294967296.0,1,-nbitq), 
to_sfixed(-309873419.0/4294967296.0,1,-nbitq), 
to_sfixed(213267716.0/4294967296.0,1,-nbitq), 
to_sfixed(389619617.0/4294967296.0,1,-nbitq), 
to_sfixed(242647983.0/4294967296.0,1,-nbitq), 
to_sfixed(72678710.0/4294967296.0,1,-nbitq), 
to_sfixed(-83921613.0/4294967296.0,1,-nbitq), 
to_sfixed(-47518069.0/4294967296.0,1,-nbitq), 
to_sfixed(129022026.0/4294967296.0,1,-nbitq), 
to_sfixed(-234397144.0/4294967296.0,1,-nbitq), 
to_sfixed(-230453202.0/4294967296.0,1,-nbitq), 
to_sfixed(-209824890.0/4294967296.0,1,-nbitq), 
to_sfixed(458360489.0/4294967296.0,1,-nbitq), 
to_sfixed(305204288.0/4294967296.0,1,-nbitq), 
to_sfixed(-212782667.0/4294967296.0,1,-nbitq), 
to_sfixed(-85795145.0/4294967296.0,1,-nbitq), 
to_sfixed(-135053291.0/4294967296.0,1,-nbitq), 
to_sfixed(-389755227.0/4294967296.0,1,-nbitq), 
to_sfixed(102226576.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(64894728.0/4294967296.0,1,-nbitq), 
to_sfixed(162328864.0/4294967296.0,1,-nbitq), 
to_sfixed(83534269.0/4294967296.0,1,-nbitq), 
to_sfixed(11842868.0/4294967296.0,1,-nbitq), 
to_sfixed(174686402.0/4294967296.0,1,-nbitq), 
to_sfixed(231351183.0/4294967296.0,1,-nbitq), 
to_sfixed(255766893.0/4294967296.0,1,-nbitq), 
to_sfixed(22809073.0/4294967296.0,1,-nbitq), 
to_sfixed(-402668485.0/4294967296.0,1,-nbitq), 
to_sfixed(-141830832.0/4294967296.0,1,-nbitq), 
to_sfixed(136836881.0/4294967296.0,1,-nbitq), 
to_sfixed(156442258.0/4294967296.0,1,-nbitq), 
to_sfixed(21300365.0/4294967296.0,1,-nbitq), 
to_sfixed(428599900.0/4294967296.0,1,-nbitq), 
to_sfixed(-10244878.0/4294967296.0,1,-nbitq), 
to_sfixed(198555932.0/4294967296.0,1,-nbitq), 
to_sfixed(-333756131.0/4294967296.0,1,-nbitq), 
to_sfixed(-326163865.0/4294967296.0,1,-nbitq), 
to_sfixed(355366269.0/4294967296.0,1,-nbitq), 
to_sfixed(207215086.0/4294967296.0,1,-nbitq), 
to_sfixed(8876246.0/4294967296.0,1,-nbitq), 
to_sfixed(364733001.0/4294967296.0,1,-nbitq), 
to_sfixed(-11587703.0/4294967296.0,1,-nbitq), 
to_sfixed(1823031.0/4294967296.0,1,-nbitq), 
to_sfixed(332129212.0/4294967296.0,1,-nbitq), 
to_sfixed(184267361.0/4294967296.0,1,-nbitq), 
to_sfixed(404934434.0/4294967296.0,1,-nbitq), 
to_sfixed(97521592.0/4294967296.0,1,-nbitq), 
to_sfixed(-206273856.0/4294967296.0,1,-nbitq), 
to_sfixed(94667703.0/4294967296.0,1,-nbitq), 
to_sfixed(-494913823.0/4294967296.0,1,-nbitq), 
to_sfixed(232180866.0/4294967296.0,1,-nbitq), 
to_sfixed(91458497.0/4294967296.0,1,-nbitq), 
to_sfixed(-399318805.0/4294967296.0,1,-nbitq), 
to_sfixed(-98895372.0/4294967296.0,1,-nbitq), 
to_sfixed(-87226334.0/4294967296.0,1,-nbitq), 
to_sfixed(250798359.0/4294967296.0,1,-nbitq), 
to_sfixed(237211919.0/4294967296.0,1,-nbitq), 
to_sfixed(91093960.0/4294967296.0,1,-nbitq), 
to_sfixed(-158745893.0/4294967296.0,1,-nbitq), 
to_sfixed(103085378.0/4294967296.0,1,-nbitq), 
to_sfixed(-107858856.0/4294967296.0,1,-nbitq), 
to_sfixed(105165890.0/4294967296.0,1,-nbitq), 
to_sfixed(-35249525.0/4294967296.0,1,-nbitq), 
to_sfixed(-181467044.0/4294967296.0,1,-nbitq), 
to_sfixed(177285730.0/4294967296.0,1,-nbitq), 
to_sfixed(219175540.0/4294967296.0,1,-nbitq), 
to_sfixed(-123737913.0/4294967296.0,1,-nbitq), 
to_sfixed(386562683.0/4294967296.0,1,-nbitq), 
to_sfixed(487419618.0/4294967296.0,1,-nbitq), 
to_sfixed(24756603.0/4294967296.0,1,-nbitq), 
to_sfixed(-185702152.0/4294967296.0,1,-nbitq), 
to_sfixed(-303991529.0/4294967296.0,1,-nbitq), 
to_sfixed(-243670115.0/4294967296.0,1,-nbitq), 
to_sfixed(374484069.0/4294967296.0,1,-nbitq), 
to_sfixed(-183054733.0/4294967296.0,1,-nbitq), 
to_sfixed(-69181699.0/4294967296.0,1,-nbitq), 
to_sfixed(-261443235.0/4294967296.0,1,-nbitq), 
to_sfixed(-4986114.0/4294967296.0,1,-nbitq), 
to_sfixed(51980716.0/4294967296.0,1,-nbitq), 
to_sfixed(365246259.0/4294967296.0,1,-nbitq), 
to_sfixed(387285624.0/4294967296.0,1,-nbitq), 
to_sfixed(-328797491.0/4294967296.0,1,-nbitq), 
to_sfixed(434218064.0/4294967296.0,1,-nbitq), 
to_sfixed(86659130.0/4294967296.0,1,-nbitq), 
to_sfixed(304467414.0/4294967296.0,1,-nbitq), 
to_sfixed(136243054.0/4294967296.0,1,-nbitq), 
to_sfixed(-126286796.0/4294967296.0,1,-nbitq), 
to_sfixed(429392587.0/4294967296.0,1,-nbitq), 
to_sfixed(543911520.0/4294967296.0,1,-nbitq), 
to_sfixed(-303589523.0/4294967296.0,1,-nbitq), 
to_sfixed(309340611.0/4294967296.0,1,-nbitq), 
to_sfixed(154282806.0/4294967296.0,1,-nbitq), 
to_sfixed(159506564.0/4294967296.0,1,-nbitq), 
to_sfixed(-10937756.0/4294967296.0,1,-nbitq), 
to_sfixed(-339018170.0/4294967296.0,1,-nbitq), 
to_sfixed(-43699119.0/4294967296.0,1,-nbitq), 
to_sfixed(-449582864.0/4294967296.0,1,-nbitq), 
to_sfixed(57219517.0/4294967296.0,1,-nbitq), 
to_sfixed(278640923.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-339005085.0/4294967296.0,1,-nbitq), 
to_sfixed(-233638118.0/4294967296.0,1,-nbitq), 
to_sfixed(325782567.0/4294967296.0,1,-nbitq), 
to_sfixed(-55013235.0/4294967296.0,1,-nbitq), 
to_sfixed(-229041580.0/4294967296.0,1,-nbitq), 
to_sfixed(-369204401.0/4294967296.0,1,-nbitq), 
to_sfixed(359291566.0/4294967296.0,1,-nbitq), 
to_sfixed(-99990200.0/4294967296.0,1,-nbitq), 
to_sfixed(-130083993.0/4294967296.0,1,-nbitq), 
to_sfixed(-38341055.0/4294967296.0,1,-nbitq), 
to_sfixed(203825326.0/4294967296.0,1,-nbitq), 
to_sfixed(278498727.0/4294967296.0,1,-nbitq), 
to_sfixed(-349835550.0/4294967296.0,1,-nbitq), 
to_sfixed(221307199.0/4294967296.0,1,-nbitq), 
to_sfixed(-37786599.0/4294967296.0,1,-nbitq), 
to_sfixed(279253816.0/4294967296.0,1,-nbitq), 
to_sfixed(-77614511.0/4294967296.0,1,-nbitq), 
to_sfixed(374691293.0/4294967296.0,1,-nbitq), 
to_sfixed(-215435566.0/4294967296.0,1,-nbitq), 
to_sfixed(-113683131.0/4294967296.0,1,-nbitq), 
to_sfixed(-57605199.0/4294967296.0,1,-nbitq), 
to_sfixed(132120038.0/4294967296.0,1,-nbitq), 
to_sfixed(294055155.0/4294967296.0,1,-nbitq), 
to_sfixed(431520414.0/4294967296.0,1,-nbitq), 
to_sfixed(-307773520.0/4294967296.0,1,-nbitq), 
to_sfixed(-98407284.0/4294967296.0,1,-nbitq), 
to_sfixed(-66395715.0/4294967296.0,1,-nbitq), 
to_sfixed(-13579956.0/4294967296.0,1,-nbitq), 
to_sfixed(461289205.0/4294967296.0,1,-nbitq), 
to_sfixed(303183185.0/4294967296.0,1,-nbitq), 
to_sfixed(140506355.0/4294967296.0,1,-nbitq), 
to_sfixed(-370796451.0/4294967296.0,1,-nbitq), 
to_sfixed(-105926251.0/4294967296.0,1,-nbitq), 
to_sfixed(-255406814.0/4294967296.0,1,-nbitq), 
to_sfixed(-177338775.0/4294967296.0,1,-nbitq), 
to_sfixed(-330928435.0/4294967296.0,1,-nbitq), 
to_sfixed(32635838.0/4294967296.0,1,-nbitq), 
to_sfixed(-169862555.0/4294967296.0,1,-nbitq), 
to_sfixed(-381625713.0/4294967296.0,1,-nbitq), 
to_sfixed(-143358190.0/4294967296.0,1,-nbitq), 
to_sfixed(161982299.0/4294967296.0,1,-nbitq), 
to_sfixed(-107858297.0/4294967296.0,1,-nbitq), 
to_sfixed(51618242.0/4294967296.0,1,-nbitq), 
to_sfixed(-1493524.0/4294967296.0,1,-nbitq), 
to_sfixed(194819707.0/4294967296.0,1,-nbitq), 
to_sfixed(176357490.0/4294967296.0,1,-nbitq), 
to_sfixed(-312476791.0/4294967296.0,1,-nbitq), 
to_sfixed(-40729710.0/4294967296.0,1,-nbitq), 
to_sfixed(-46666714.0/4294967296.0,1,-nbitq), 
to_sfixed(308713202.0/4294967296.0,1,-nbitq), 
to_sfixed(377684951.0/4294967296.0,1,-nbitq), 
to_sfixed(-268252665.0/4294967296.0,1,-nbitq), 
to_sfixed(-181782568.0/4294967296.0,1,-nbitq), 
to_sfixed(-101704502.0/4294967296.0,1,-nbitq), 
to_sfixed(-93142518.0/4294967296.0,1,-nbitq), 
to_sfixed(232753729.0/4294967296.0,1,-nbitq), 
to_sfixed(-38498468.0/4294967296.0,1,-nbitq), 
to_sfixed(-60625651.0/4294967296.0,1,-nbitq), 
to_sfixed(-121303214.0/4294967296.0,1,-nbitq), 
to_sfixed(403812742.0/4294967296.0,1,-nbitq), 
to_sfixed(374085785.0/4294967296.0,1,-nbitq), 
to_sfixed(20367497.0/4294967296.0,1,-nbitq), 
to_sfixed(-327377168.0/4294967296.0,1,-nbitq), 
to_sfixed(187228354.0/4294967296.0,1,-nbitq), 
to_sfixed(-100911610.0/4294967296.0,1,-nbitq), 
to_sfixed(-360691684.0/4294967296.0,1,-nbitq), 
to_sfixed(674283694.0/4294967296.0,1,-nbitq), 
to_sfixed(-29878674.0/4294967296.0,1,-nbitq), 
to_sfixed(439425287.0/4294967296.0,1,-nbitq), 
to_sfixed(-335898.0/4294967296.0,1,-nbitq), 
to_sfixed(121452840.0/4294967296.0,1,-nbitq), 
to_sfixed(-374287223.0/4294967296.0,1,-nbitq), 
to_sfixed(-224560507.0/4294967296.0,1,-nbitq), 
to_sfixed(107414710.0/4294967296.0,1,-nbitq), 
to_sfixed(320536131.0/4294967296.0,1,-nbitq), 
to_sfixed(-456848741.0/4294967296.0,1,-nbitq), 
to_sfixed(-157440140.0/4294967296.0,1,-nbitq), 
to_sfixed(-500731811.0/4294967296.0,1,-nbitq), 
to_sfixed(-245379889.0/4294967296.0,1,-nbitq), 
to_sfixed(338568716.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-61275038.0/4294967296.0,1,-nbitq), 
to_sfixed(-68932351.0/4294967296.0,1,-nbitq), 
to_sfixed(81863246.0/4294967296.0,1,-nbitq), 
to_sfixed(241911926.0/4294967296.0,1,-nbitq), 
to_sfixed(-110248644.0/4294967296.0,1,-nbitq), 
to_sfixed(-395446067.0/4294967296.0,1,-nbitq), 
to_sfixed(84635240.0/4294967296.0,1,-nbitq), 
to_sfixed(226343381.0/4294967296.0,1,-nbitq), 
to_sfixed(-85209232.0/4294967296.0,1,-nbitq), 
to_sfixed(21094831.0/4294967296.0,1,-nbitq), 
to_sfixed(-278651103.0/4294967296.0,1,-nbitq), 
to_sfixed(-129648505.0/4294967296.0,1,-nbitq), 
to_sfixed(-307546398.0/4294967296.0,1,-nbitq), 
to_sfixed(-241669650.0/4294967296.0,1,-nbitq), 
to_sfixed(-375730612.0/4294967296.0,1,-nbitq), 
to_sfixed(229221395.0/4294967296.0,1,-nbitq), 
to_sfixed(297368577.0/4294967296.0,1,-nbitq), 
to_sfixed(-80308653.0/4294967296.0,1,-nbitq), 
to_sfixed(291938067.0/4294967296.0,1,-nbitq), 
to_sfixed(-273597469.0/4294967296.0,1,-nbitq), 
to_sfixed(-353643938.0/4294967296.0,1,-nbitq), 
to_sfixed(27054406.0/4294967296.0,1,-nbitq), 
to_sfixed(439156754.0/4294967296.0,1,-nbitq), 
to_sfixed(180726786.0/4294967296.0,1,-nbitq), 
to_sfixed(243203268.0/4294967296.0,1,-nbitq), 
to_sfixed(361316220.0/4294967296.0,1,-nbitq), 
to_sfixed(-129982583.0/4294967296.0,1,-nbitq), 
to_sfixed(48457682.0/4294967296.0,1,-nbitq), 
to_sfixed(439551986.0/4294967296.0,1,-nbitq), 
to_sfixed(250776080.0/4294967296.0,1,-nbitq), 
to_sfixed(-464089854.0/4294967296.0,1,-nbitq), 
to_sfixed(227998423.0/4294967296.0,1,-nbitq), 
to_sfixed(-222857432.0/4294967296.0,1,-nbitq), 
to_sfixed(-187121325.0/4294967296.0,1,-nbitq), 
to_sfixed(119267697.0/4294967296.0,1,-nbitq), 
to_sfixed(156653802.0/4294967296.0,1,-nbitq), 
to_sfixed(-318287110.0/4294967296.0,1,-nbitq), 
to_sfixed(63742352.0/4294967296.0,1,-nbitq), 
to_sfixed(-381475323.0/4294967296.0,1,-nbitq), 
to_sfixed(-88446586.0/4294967296.0,1,-nbitq), 
to_sfixed(-200593428.0/4294967296.0,1,-nbitq), 
to_sfixed(377856523.0/4294967296.0,1,-nbitq), 
to_sfixed(-243738379.0/4294967296.0,1,-nbitq), 
to_sfixed(-195544534.0/4294967296.0,1,-nbitq), 
to_sfixed(-285027419.0/4294967296.0,1,-nbitq), 
to_sfixed(193371598.0/4294967296.0,1,-nbitq), 
to_sfixed(-436900435.0/4294967296.0,1,-nbitq), 
to_sfixed(-152728355.0/4294967296.0,1,-nbitq), 
to_sfixed(-255852009.0/4294967296.0,1,-nbitq), 
to_sfixed(536286837.0/4294967296.0,1,-nbitq), 
to_sfixed(-155457321.0/4294967296.0,1,-nbitq), 
to_sfixed(292248174.0/4294967296.0,1,-nbitq), 
to_sfixed(-151144633.0/4294967296.0,1,-nbitq), 
to_sfixed(116076981.0/4294967296.0,1,-nbitq), 
to_sfixed(-371959856.0/4294967296.0,1,-nbitq), 
to_sfixed(258792452.0/4294967296.0,1,-nbitq), 
to_sfixed(335346757.0/4294967296.0,1,-nbitq), 
to_sfixed(150717168.0/4294967296.0,1,-nbitq), 
to_sfixed(324628442.0/4294967296.0,1,-nbitq), 
to_sfixed(124504081.0/4294967296.0,1,-nbitq), 
to_sfixed(-359208267.0/4294967296.0,1,-nbitq), 
to_sfixed(-36849611.0/4294967296.0,1,-nbitq), 
to_sfixed(-31450758.0/4294967296.0,1,-nbitq), 
to_sfixed(98711369.0/4294967296.0,1,-nbitq), 
to_sfixed(-292806761.0/4294967296.0,1,-nbitq), 
to_sfixed(187872722.0/4294967296.0,1,-nbitq), 
to_sfixed(674634268.0/4294967296.0,1,-nbitq), 
to_sfixed(-280740323.0/4294967296.0,1,-nbitq), 
to_sfixed(370675330.0/4294967296.0,1,-nbitq), 
to_sfixed(417271377.0/4294967296.0,1,-nbitq), 
to_sfixed(-43702724.0/4294967296.0,1,-nbitq), 
to_sfixed(-364073929.0/4294967296.0,1,-nbitq), 
to_sfixed(-307315328.0/4294967296.0,1,-nbitq), 
to_sfixed(365703843.0/4294967296.0,1,-nbitq), 
to_sfixed(161828262.0/4294967296.0,1,-nbitq), 
to_sfixed(-133336414.0/4294967296.0,1,-nbitq), 
to_sfixed(136324453.0/4294967296.0,1,-nbitq), 
to_sfixed(-394722283.0/4294967296.0,1,-nbitq), 
to_sfixed(-55390941.0/4294967296.0,1,-nbitq), 
to_sfixed(215403792.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(160465278.0/4294967296.0,1,-nbitq), 
to_sfixed(-385888946.0/4294967296.0,1,-nbitq), 
to_sfixed(-58226640.0/4294967296.0,1,-nbitq), 
to_sfixed(193145022.0/4294967296.0,1,-nbitq), 
to_sfixed(295962741.0/4294967296.0,1,-nbitq), 
to_sfixed(170502274.0/4294967296.0,1,-nbitq), 
to_sfixed(-109579177.0/4294967296.0,1,-nbitq), 
to_sfixed(-333525430.0/4294967296.0,1,-nbitq), 
to_sfixed(-162767498.0/4294967296.0,1,-nbitq), 
to_sfixed(-189028335.0/4294967296.0,1,-nbitq), 
to_sfixed(102877915.0/4294967296.0,1,-nbitq), 
to_sfixed(294275127.0/4294967296.0,1,-nbitq), 
to_sfixed(167599204.0/4294967296.0,1,-nbitq), 
to_sfixed(435547711.0/4294967296.0,1,-nbitq), 
to_sfixed(-249220173.0/4294967296.0,1,-nbitq), 
to_sfixed(-240361636.0/4294967296.0,1,-nbitq), 
to_sfixed(137246051.0/4294967296.0,1,-nbitq), 
to_sfixed(233455103.0/4294967296.0,1,-nbitq), 
to_sfixed(-141588063.0/4294967296.0,1,-nbitq), 
to_sfixed(112252276.0/4294967296.0,1,-nbitq), 
to_sfixed(195118758.0/4294967296.0,1,-nbitq), 
to_sfixed(-145107491.0/4294967296.0,1,-nbitq), 
to_sfixed(51527384.0/4294967296.0,1,-nbitq), 
to_sfixed(-61974838.0/4294967296.0,1,-nbitq), 
to_sfixed(265204889.0/4294967296.0,1,-nbitq), 
to_sfixed(481848341.0/4294967296.0,1,-nbitq), 
to_sfixed(-139996242.0/4294967296.0,1,-nbitq), 
to_sfixed(57896022.0/4294967296.0,1,-nbitq), 
to_sfixed(51769470.0/4294967296.0,1,-nbitq), 
to_sfixed(-136853284.0/4294967296.0,1,-nbitq), 
to_sfixed(-559903553.0/4294967296.0,1,-nbitq), 
to_sfixed(-44311290.0/4294967296.0,1,-nbitq), 
to_sfixed(116620887.0/4294967296.0,1,-nbitq), 
to_sfixed(186670224.0/4294967296.0,1,-nbitq), 
to_sfixed(231446176.0/4294967296.0,1,-nbitq), 
to_sfixed(-30254877.0/4294967296.0,1,-nbitq), 
to_sfixed(-217622090.0/4294967296.0,1,-nbitq), 
to_sfixed(-418982235.0/4294967296.0,1,-nbitq), 
to_sfixed(-28848400.0/4294967296.0,1,-nbitq), 
to_sfixed(-29660054.0/4294967296.0,1,-nbitq), 
to_sfixed(-101921570.0/4294967296.0,1,-nbitq), 
to_sfixed(477610614.0/4294967296.0,1,-nbitq), 
to_sfixed(24615003.0/4294967296.0,1,-nbitq), 
to_sfixed(305593017.0/4294967296.0,1,-nbitq), 
to_sfixed(-235197883.0/4294967296.0,1,-nbitq), 
to_sfixed(-8025629.0/4294967296.0,1,-nbitq), 
to_sfixed(196580244.0/4294967296.0,1,-nbitq), 
to_sfixed(57534870.0/4294967296.0,1,-nbitq), 
to_sfixed(-32069490.0/4294967296.0,1,-nbitq), 
to_sfixed(207581739.0/4294967296.0,1,-nbitq), 
to_sfixed(379481728.0/4294967296.0,1,-nbitq), 
to_sfixed(98842210.0/4294967296.0,1,-nbitq), 
to_sfixed(-511778573.0/4294967296.0,1,-nbitq), 
to_sfixed(182661537.0/4294967296.0,1,-nbitq), 
to_sfixed(89823256.0/4294967296.0,1,-nbitq), 
to_sfixed(-340309143.0/4294967296.0,1,-nbitq), 
to_sfixed(186672344.0/4294967296.0,1,-nbitq), 
to_sfixed(-29094974.0/4294967296.0,1,-nbitq), 
to_sfixed(-185439754.0/4294967296.0,1,-nbitq), 
to_sfixed(-11239139.0/4294967296.0,1,-nbitq), 
to_sfixed(157507473.0/4294967296.0,1,-nbitq), 
to_sfixed(108827918.0/4294967296.0,1,-nbitq), 
to_sfixed(-488516909.0/4294967296.0,1,-nbitq), 
to_sfixed(-9001454.0/4294967296.0,1,-nbitq), 
to_sfixed(208525614.0/4294967296.0,1,-nbitq), 
to_sfixed(-110201898.0/4294967296.0,1,-nbitq), 
to_sfixed(690942356.0/4294967296.0,1,-nbitq), 
to_sfixed(122244831.0/4294967296.0,1,-nbitq), 
to_sfixed(7425950.0/4294967296.0,1,-nbitq), 
to_sfixed(467417497.0/4294967296.0,1,-nbitq), 
to_sfixed(-240741918.0/4294967296.0,1,-nbitq), 
to_sfixed(-222416981.0/4294967296.0,1,-nbitq), 
to_sfixed(129954920.0/4294967296.0,1,-nbitq), 
to_sfixed(405439093.0/4294967296.0,1,-nbitq), 
to_sfixed(172840910.0/4294967296.0,1,-nbitq), 
to_sfixed(-377095880.0/4294967296.0,1,-nbitq), 
to_sfixed(-196383858.0/4294967296.0,1,-nbitq), 
to_sfixed(134896236.0/4294967296.0,1,-nbitq), 
to_sfixed(458142652.0/4294967296.0,1,-nbitq), 
to_sfixed(-156874490.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-103267865.0/4294967296.0,1,-nbitq), 
to_sfixed(-270674682.0/4294967296.0,1,-nbitq), 
to_sfixed(310793538.0/4294967296.0,1,-nbitq), 
to_sfixed(-435045307.0/4294967296.0,1,-nbitq), 
to_sfixed(273647237.0/4294967296.0,1,-nbitq), 
to_sfixed(-430833051.0/4294967296.0,1,-nbitq), 
to_sfixed(28666516.0/4294967296.0,1,-nbitq), 
to_sfixed(-106379913.0/4294967296.0,1,-nbitq), 
to_sfixed(-289986430.0/4294967296.0,1,-nbitq), 
to_sfixed(141401010.0/4294967296.0,1,-nbitq), 
to_sfixed(258333101.0/4294967296.0,1,-nbitq), 
to_sfixed(-112841743.0/4294967296.0,1,-nbitq), 
to_sfixed(-85460928.0/4294967296.0,1,-nbitq), 
to_sfixed(-248428979.0/4294967296.0,1,-nbitq), 
to_sfixed(-169063997.0/4294967296.0,1,-nbitq), 
to_sfixed(114770809.0/4294967296.0,1,-nbitq), 
to_sfixed(-306196083.0/4294967296.0,1,-nbitq), 
to_sfixed(-249521831.0/4294967296.0,1,-nbitq), 
to_sfixed(335759497.0/4294967296.0,1,-nbitq), 
to_sfixed(335353914.0/4294967296.0,1,-nbitq), 
to_sfixed(102537557.0/4294967296.0,1,-nbitq), 
to_sfixed(59414357.0/4294967296.0,1,-nbitq), 
to_sfixed(-127056200.0/4294967296.0,1,-nbitq), 
to_sfixed(147921519.0/4294967296.0,1,-nbitq), 
to_sfixed(177996982.0/4294967296.0,1,-nbitq), 
to_sfixed(240977366.0/4294967296.0,1,-nbitq), 
to_sfixed(8378238.0/4294967296.0,1,-nbitq), 
to_sfixed(-128990211.0/4294967296.0,1,-nbitq), 
to_sfixed(338118690.0/4294967296.0,1,-nbitq), 
to_sfixed(-220825720.0/4294967296.0,1,-nbitq), 
to_sfixed(-154106695.0/4294967296.0,1,-nbitq), 
to_sfixed(9746955.0/4294967296.0,1,-nbitq), 
to_sfixed(160483333.0/4294967296.0,1,-nbitq), 
to_sfixed(54773060.0/4294967296.0,1,-nbitq), 
to_sfixed(90926267.0/4294967296.0,1,-nbitq), 
to_sfixed(442389639.0/4294967296.0,1,-nbitq), 
to_sfixed(-36607981.0/4294967296.0,1,-nbitq), 
to_sfixed(141200399.0/4294967296.0,1,-nbitq), 
to_sfixed(-176086601.0/4294967296.0,1,-nbitq), 
to_sfixed(-116078805.0/4294967296.0,1,-nbitq), 
to_sfixed(232543119.0/4294967296.0,1,-nbitq), 
to_sfixed(-78814907.0/4294967296.0,1,-nbitq), 
to_sfixed(-305299847.0/4294967296.0,1,-nbitq), 
to_sfixed(14247004.0/4294967296.0,1,-nbitq), 
to_sfixed(-55803564.0/4294967296.0,1,-nbitq), 
to_sfixed(-162247009.0/4294967296.0,1,-nbitq), 
to_sfixed(24149767.0/4294967296.0,1,-nbitq), 
to_sfixed(-297066985.0/4294967296.0,1,-nbitq), 
to_sfixed(-196806783.0/4294967296.0,1,-nbitq), 
to_sfixed(-29300089.0/4294967296.0,1,-nbitq), 
to_sfixed(-233125272.0/4294967296.0,1,-nbitq), 
to_sfixed(10271462.0/4294967296.0,1,-nbitq), 
to_sfixed(154259926.0/4294967296.0,1,-nbitq), 
to_sfixed(-34495935.0/4294967296.0,1,-nbitq), 
to_sfixed(203272314.0/4294967296.0,1,-nbitq), 
to_sfixed(54932727.0/4294967296.0,1,-nbitq), 
to_sfixed(132766340.0/4294967296.0,1,-nbitq), 
to_sfixed(-430097985.0/4294967296.0,1,-nbitq), 
to_sfixed(-316877088.0/4294967296.0,1,-nbitq), 
to_sfixed(31716955.0/4294967296.0,1,-nbitq), 
to_sfixed(394693551.0/4294967296.0,1,-nbitq), 
to_sfixed(42427661.0/4294967296.0,1,-nbitq), 
to_sfixed(-301018002.0/4294967296.0,1,-nbitq), 
to_sfixed(221695373.0/4294967296.0,1,-nbitq), 
to_sfixed(94543778.0/4294967296.0,1,-nbitq), 
to_sfixed(225771921.0/4294967296.0,1,-nbitq), 
to_sfixed(553655806.0/4294967296.0,1,-nbitq), 
to_sfixed(-425729667.0/4294967296.0,1,-nbitq), 
to_sfixed(-92071093.0/4294967296.0,1,-nbitq), 
to_sfixed(258693225.0/4294967296.0,1,-nbitq), 
to_sfixed(62109370.0/4294967296.0,1,-nbitq), 
to_sfixed(38440218.0/4294967296.0,1,-nbitq), 
to_sfixed(-258264374.0/4294967296.0,1,-nbitq), 
to_sfixed(-224828534.0/4294967296.0,1,-nbitq), 
to_sfixed(108131146.0/4294967296.0,1,-nbitq), 
to_sfixed(-506662962.0/4294967296.0,1,-nbitq), 
to_sfixed(367818508.0/4294967296.0,1,-nbitq), 
to_sfixed(22584009.0/4294967296.0,1,-nbitq), 
to_sfixed(285180184.0/4294967296.0,1,-nbitq), 
to_sfixed(215154042.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq), 
to_sfixed(0.0/4294967296.0,1,-nbitq)  ) 
 ) ;

constant coef2 : typtabcnf2 := ( ( to_sfixed(510345655.0/4294967296.0,1,-nbitq), 
to_sfixed(481262387.0/4294967296.0,1,-nbitq), 
to_sfixed(-880876840.0/4294967296.0,1,-nbitq), 
to_sfixed(-740381076.0/4294967296.0,1,-nbitq), 
to_sfixed(552223413.0/4294967296.0,1,-nbitq), 
to_sfixed(-644759981.0/4294967296.0,1,-nbitq), 
to_sfixed(508581876.0/4294967296.0,1,-nbitq), 
to_sfixed(-88322714.0/4294967296.0,1,-nbitq), 
to_sfixed(-855382299.0/4294967296.0,1,-nbitq), 
to_sfixed(779846809.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-1967822058.0/4294967296.0,1,-nbitq), 
to_sfixed(-997420102.0/4294967296.0,1,-nbitq), 
to_sfixed(165086289.0/4294967296.0,1,-nbitq), 
to_sfixed(-573830493.0/4294967296.0,1,-nbitq), 
to_sfixed(1094162481.0/4294967296.0,1,-nbitq), 
to_sfixed(1831049747.0/4294967296.0,1,-nbitq), 
to_sfixed(-1352688536.0/4294967296.0,1,-nbitq), 
to_sfixed(-343966684.0/4294967296.0,1,-nbitq), 
to_sfixed(-633580759.0/4294967296.0,1,-nbitq), 
to_sfixed(81024205.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-140576633.0/4294967296.0,1,-nbitq), 
to_sfixed(1380158524.0/4294967296.0,1,-nbitq), 
to_sfixed(-1503003841.0/4294967296.0,1,-nbitq), 
to_sfixed(-1160624254.0/4294967296.0,1,-nbitq), 
to_sfixed(-1607915204.0/4294967296.0,1,-nbitq), 
to_sfixed(281992920.0/4294967296.0,1,-nbitq), 
to_sfixed(1927941293.0/4294967296.0,1,-nbitq), 
to_sfixed(-1597250443.0/4294967296.0,1,-nbitq), 
to_sfixed(-441050336.0/4294967296.0,1,-nbitq), 
to_sfixed(321951657.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(550412425.0/4294967296.0,1,-nbitq), 
to_sfixed(-450696930.0/4294967296.0,1,-nbitq), 
to_sfixed(1461308244.0/4294967296.0,1,-nbitq), 
to_sfixed(-716506242.0/4294967296.0,1,-nbitq), 
to_sfixed(-1074654480.0/4294967296.0,1,-nbitq), 
to_sfixed(-1224804137.0/4294967296.0,1,-nbitq), 
to_sfixed(598810368.0/4294967296.0,1,-nbitq), 
to_sfixed(1943096370.0/4294967296.0,1,-nbitq), 
to_sfixed(-1150347122.0/4294967296.0,1,-nbitq), 
to_sfixed(-814690308.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(417481410.0/4294967296.0,1,-nbitq), 
to_sfixed(-1321835937.0/4294967296.0,1,-nbitq), 
to_sfixed(1043381801.0/4294967296.0,1,-nbitq), 
to_sfixed(-319590477.0/4294967296.0,1,-nbitq), 
to_sfixed(853359395.0/4294967296.0,1,-nbitq), 
to_sfixed(113411374.0/4294967296.0,1,-nbitq), 
to_sfixed(479298347.0/4294967296.0,1,-nbitq), 
to_sfixed(913692422.0/4294967296.0,1,-nbitq), 
to_sfixed(-508885478.0/4294967296.0,1,-nbitq), 
to_sfixed(-2285965770.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-2219318509.0/4294967296.0,1,-nbitq), 
to_sfixed(452343780.0/4294967296.0,1,-nbitq), 
to_sfixed(525066905.0/4294967296.0,1,-nbitq), 
to_sfixed(1701634583.0/4294967296.0,1,-nbitq), 
to_sfixed(464160935.0/4294967296.0,1,-nbitq), 
to_sfixed(-1261014034.0/4294967296.0,1,-nbitq), 
to_sfixed(110613081.0/4294967296.0,1,-nbitq), 
to_sfixed(97797902.0/4294967296.0,1,-nbitq), 
to_sfixed(-290200576.0/4294967296.0,1,-nbitq), 
to_sfixed(-1648231894.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-181169297.0/4294967296.0,1,-nbitq), 
to_sfixed(-262548870.0/4294967296.0,1,-nbitq), 
to_sfixed(114610915.0/4294967296.0,1,-nbitq), 
to_sfixed(17518742.0/4294967296.0,1,-nbitq), 
to_sfixed(-542233175.0/4294967296.0,1,-nbitq), 
to_sfixed(-272032907.0/4294967296.0,1,-nbitq), 
to_sfixed(813042547.0/4294967296.0,1,-nbitq), 
to_sfixed(616580243.0/4294967296.0,1,-nbitq), 
to_sfixed(955876700.0/4294967296.0,1,-nbitq), 
to_sfixed(934342429.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(1126871603.0/4294967296.0,1,-nbitq), 
to_sfixed(-1590248796.0/4294967296.0,1,-nbitq), 
to_sfixed(-819361470.0/4294967296.0,1,-nbitq), 
to_sfixed(-905662292.0/4294967296.0,1,-nbitq), 
to_sfixed(432669163.0/4294967296.0,1,-nbitq), 
to_sfixed(1164871769.0/4294967296.0,1,-nbitq), 
to_sfixed(1049193721.0/4294967296.0,1,-nbitq), 
to_sfixed(930177897.0/4294967296.0,1,-nbitq), 
to_sfixed(948610472.0/4294967296.0,1,-nbitq), 
to_sfixed(1119505172.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(1154303187.0/4294967296.0,1,-nbitq), 
to_sfixed(-549874814.0/4294967296.0,1,-nbitq), 
to_sfixed(893927118.0/4294967296.0,1,-nbitq), 
to_sfixed(-1300839732.0/4294967296.0,1,-nbitq), 
to_sfixed(-1118502113.0/4294967296.0,1,-nbitq), 
to_sfixed(12145018.0/4294967296.0,1,-nbitq), 
to_sfixed(993366253.0/4294967296.0,1,-nbitq), 
to_sfixed(-1519609776.0/4294967296.0,1,-nbitq), 
to_sfixed(-877416461.0/4294967296.0,1,-nbitq), 
to_sfixed(-706102881.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-349597992.0/4294967296.0,1,-nbitq), 
to_sfixed(-106643830.0/4294967296.0,1,-nbitq), 
to_sfixed(1045590781.0/4294967296.0,1,-nbitq), 
to_sfixed(-787648168.0/4294967296.0,1,-nbitq), 
to_sfixed(124673066.0/4294967296.0,1,-nbitq), 
to_sfixed(795537482.0/4294967296.0,1,-nbitq), 
to_sfixed(186365523.0/4294967296.0,1,-nbitq), 
to_sfixed(-910724981.0/4294967296.0,1,-nbitq), 
to_sfixed(1090403512.0/4294967296.0,1,-nbitq), 
to_sfixed(201736924.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-1363495938.0/4294967296.0,1,-nbitq), 
to_sfixed(-901014330.0/4294967296.0,1,-nbitq), 
to_sfixed(1384784214.0/4294967296.0,1,-nbitq), 
to_sfixed(-1437828225.0/4294967296.0,1,-nbitq), 
to_sfixed(1135734128.0/4294967296.0,1,-nbitq), 
to_sfixed(-25199412.0/4294967296.0,1,-nbitq), 
to_sfixed(411185946.0/4294967296.0,1,-nbitq), 
to_sfixed(50495471.0/4294967296.0,1,-nbitq), 
to_sfixed(-82334242.0/4294967296.0,1,-nbitq), 
to_sfixed(240618276.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-346706062.0/4294967296.0,1,-nbitq), 
to_sfixed(-590610058.0/4294967296.0,1,-nbitq), 
to_sfixed(839185563.0/4294967296.0,1,-nbitq), 
to_sfixed(-973894712.0/4294967296.0,1,-nbitq), 
to_sfixed(1494537704.0/4294967296.0,1,-nbitq), 
to_sfixed(-367514324.0/4294967296.0,1,-nbitq), 
to_sfixed(1230697141.0/4294967296.0,1,-nbitq), 
to_sfixed(1448024834.0/4294967296.0,1,-nbitq), 
to_sfixed(571540122.0/4294967296.0,1,-nbitq), 
to_sfixed(-1428708244.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-237292238.0/4294967296.0,1,-nbitq), 
to_sfixed(-416883199.0/4294967296.0,1,-nbitq), 
to_sfixed(640413270.0/4294967296.0,1,-nbitq), 
to_sfixed(1534802697.0/4294967296.0,1,-nbitq), 
to_sfixed(-1040848608.0/4294967296.0,1,-nbitq), 
to_sfixed(1479261716.0/4294967296.0,1,-nbitq), 
to_sfixed(-992399801.0/4294967296.0,1,-nbitq), 
to_sfixed(1922238714.0/4294967296.0,1,-nbitq), 
to_sfixed(97398611.0/4294967296.0,1,-nbitq), 
to_sfixed(848659943.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(502142981.0/4294967296.0,1,-nbitq), 
to_sfixed(426127910.0/4294967296.0,1,-nbitq), 
to_sfixed(-1153509452.0/4294967296.0,1,-nbitq), 
to_sfixed(1178701637.0/4294967296.0,1,-nbitq), 
to_sfixed(300608058.0/4294967296.0,1,-nbitq), 
to_sfixed(-1614100596.0/4294967296.0,1,-nbitq), 
to_sfixed(-324096380.0/4294967296.0,1,-nbitq), 
to_sfixed(-504620296.0/4294967296.0,1,-nbitq), 
to_sfixed(-1910374340.0/4294967296.0,1,-nbitq), 
to_sfixed(1946147950.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(405031251.0/4294967296.0,1,-nbitq), 
to_sfixed(770993081.0/4294967296.0,1,-nbitq), 
to_sfixed(-917222276.0/4294967296.0,1,-nbitq), 
to_sfixed(-412014296.0/4294967296.0,1,-nbitq), 
to_sfixed(740270187.0/4294967296.0,1,-nbitq), 
to_sfixed(-935991413.0/4294967296.0,1,-nbitq), 
to_sfixed(-682402518.0/4294967296.0,1,-nbitq), 
to_sfixed(-328138406.0/4294967296.0,1,-nbitq), 
to_sfixed(50532511.0/4294967296.0,1,-nbitq), 
to_sfixed(-807809428.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(409693202.0/4294967296.0,1,-nbitq), 
to_sfixed(-1565837861.0/4294967296.0,1,-nbitq), 
to_sfixed(-986560092.0/4294967296.0,1,-nbitq), 
to_sfixed(-1211914110.0/4294967296.0,1,-nbitq), 
to_sfixed(165154054.0/4294967296.0,1,-nbitq), 
to_sfixed(573899832.0/4294967296.0,1,-nbitq), 
to_sfixed(1417207861.0/4294967296.0,1,-nbitq), 
to_sfixed(-107273849.0/4294967296.0,1,-nbitq), 
to_sfixed(136360951.0/4294967296.0,1,-nbitq), 
to_sfixed(202116963.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(547658394.0/4294967296.0,1,-nbitq), 
to_sfixed(204680429.0/4294967296.0,1,-nbitq), 
to_sfixed(589413687.0/4294967296.0,1,-nbitq), 
to_sfixed(516117654.0/4294967296.0,1,-nbitq), 
to_sfixed(-616723173.0/4294967296.0,1,-nbitq), 
to_sfixed(-860456249.0/4294967296.0,1,-nbitq), 
to_sfixed(-843947373.0/4294967296.0,1,-nbitq), 
to_sfixed(-135263306.0/4294967296.0,1,-nbitq), 
to_sfixed(-922240340.0/4294967296.0,1,-nbitq), 
to_sfixed(33606690.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-453192026.0/4294967296.0,1,-nbitq), 
to_sfixed(914085052.0/4294967296.0,1,-nbitq), 
to_sfixed(-444782136.0/4294967296.0,1,-nbitq), 
to_sfixed(414055735.0/4294967296.0,1,-nbitq), 
to_sfixed(643683031.0/4294967296.0,1,-nbitq), 
to_sfixed(-631530365.0/4294967296.0,1,-nbitq), 
to_sfixed(1026907510.0/4294967296.0,1,-nbitq), 
to_sfixed(864759925.0/4294967296.0,1,-nbitq), 
to_sfixed(116327093.0/4294967296.0,1,-nbitq), 
to_sfixed(-1045364137.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(1405857336.0/4294967296.0,1,-nbitq), 
to_sfixed(85985123.0/4294967296.0,1,-nbitq), 
to_sfixed(65514460.0/4294967296.0,1,-nbitq), 
to_sfixed(-475167255.0/4294967296.0,1,-nbitq), 
to_sfixed(1375016558.0/4294967296.0,1,-nbitq), 
to_sfixed(355853933.0/4294967296.0,1,-nbitq), 
to_sfixed(-1032238370.0/4294967296.0,1,-nbitq), 
to_sfixed(-2085559120.0/4294967296.0,1,-nbitq), 
to_sfixed(-868901136.0/4294967296.0,1,-nbitq), 
to_sfixed(786164945.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-254840463.0/4294967296.0,1,-nbitq), 
to_sfixed(-445715300.0/4294967296.0,1,-nbitq), 
to_sfixed(-380628569.0/4294967296.0,1,-nbitq), 
to_sfixed(-378983399.0/4294967296.0,1,-nbitq), 
to_sfixed(1257236629.0/4294967296.0,1,-nbitq), 
to_sfixed(1193315567.0/4294967296.0,1,-nbitq), 
to_sfixed(653353561.0/4294967296.0,1,-nbitq), 
to_sfixed(1246732047.0/4294967296.0,1,-nbitq), 
to_sfixed(418478878.0/4294967296.0,1,-nbitq), 
to_sfixed(801230355.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(604620098.0/4294967296.0,1,-nbitq), 
to_sfixed(-471686867.0/4294967296.0,1,-nbitq), 
to_sfixed(283428465.0/4294967296.0,1,-nbitq), 
to_sfixed(-827505616.0/4294967296.0,1,-nbitq), 
to_sfixed(227344324.0/4294967296.0,1,-nbitq), 
to_sfixed(-1046017163.0/4294967296.0,1,-nbitq), 
to_sfixed(595678232.0/4294967296.0,1,-nbitq), 
to_sfixed(100969738.0/4294967296.0,1,-nbitq), 
to_sfixed(-701015515.0/4294967296.0,1,-nbitq), 
to_sfixed(-528611691.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-671188680.0/4294967296.0,1,-nbitq), 
to_sfixed(820592681.0/4294967296.0,1,-nbitq), 
to_sfixed(-246734667.0/4294967296.0,1,-nbitq), 
to_sfixed(-263277230.0/4294967296.0,1,-nbitq), 
to_sfixed(-830053484.0/4294967296.0,1,-nbitq), 
to_sfixed(503183343.0/4294967296.0,1,-nbitq), 
to_sfixed(1200707227.0/4294967296.0,1,-nbitq), 
to_sfixed(-357874407.0/4294967296.0,1,-nbitq), 
to_sfixed(-1117794433.0/4294967296.0,1,-nbitq), 
to_sfixed(-944928874.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(474739331.0/4294967296.0,1,-nbitq), 
to_sfixed(-713734653.0/4294967296.0,1,-nbitq), 
to_sfixed(906056429.0/4294967296.0,1,-nbitq), 
to_sfixed(871170699.0/4294967296.0,1,-nbitq), 
to_sfixed(1085161145.0/4294967296.0,1,-nbitq), 
to_sfixed(-1800473968.0/4294967296.0,1,-nbitq), 
to_sfixed(215846386.0/4294967296.0,1,-nbitq), 
to_sfixed(107296721.0/4294967296.0,1,-nbitq), 
to_sfixed(-1089189053.0/4294967296.0,1,-nbitq), 
to_sfixed(-583677033.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(658826386.0/4294967296.0,1,-nbitq), 
to_sfixed(1240139672.0/4294967296.0,1,-nbitq), 
to_sfixed(-943371268.0/4294967296.0,1,-nbitq), 
to_sfixed(-778846817.0/4294967296.0,1,-nbitq), 
to_sfixed(-503065691.0/4294967296.0,1,-nbitq), 
to_sfixed(1174913466.0/4294967296.0,1,-nbitq), 
to_sfixed(-230232688.0/4294967296.0,1,-nbitq), 
to_sfixed(919168492.0/4294967296.0,1,-nbitq), 
to_sfixed(-1432287909.0/4294967296.0,1,-nbitq), 
to_sfixed(1603587536.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(618350970.0/4294967296.0,1,-nbitq), 
to_sfixed(-267483038.0/4294967296.0,1,-nbitq), 
to_sfixed(-781000757.0/4294967296.0,1,-nbitq), 
to_sfixed(-180560057.0/4294967296.0,1,-nbitq), 
to_sfixed(97510279.0/4294967296.0,1,-nbitq), 
to_sfixed(577720669.0/4294967296.0,1,-nbitq), 
to_sfixed(-626526718.0/4294967296.0,1,-nbitq), 
to_sfixed(-698169919.0/4294967296.0,1,-nbitq), 
to_sfixed(-372146700.0/4294967296.0,1,-nbitq), 
to_sfixed(971630836.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-370885190.0/4294967296.0,1,-nbitq), 
to_sfixed(433915147.0/4294967296.0,1,-nbitq), 
to_sfixed(87772591.0/4294967296.0,1,-nbitq), 
to_sfixed(1045795407.0/4294967296.0,1,-nbitq), 
to_sfixed(1215851247.0/4294967296.0,1,-nbitq), 
to_sfixed(-524663155.0/4294967296.0,1,-nbitq), 
to_sfixed(-1012480196.0/4294967296.0,1,-nbitq), 
to_sfixed(825429868.0/4294967296.0,1,-nbitq), 
to_sfixed(-1532654054.0/4294967296.0,1,-nbitq), 
to_sfixed(-38796898.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-325025134.0/4294967296.0,1,-nbitq), 
to_sfixed(-15407496.0/4294967296.0,1,-nbitq), 
to_sfixed(-763618729.0/4294967296.0,1,-nbitq), 
to_sfixed(-645291540.0/4294967296.0,1,-nbitq), 
to_sfixed(-588655134.0/4294967296.0,1,-nbitq), 
to_sfixed(912580807.0/4294967296.0,1,-nbitq), 
to_sfixed(-605691996.0/4294967296.0,1,-nbitq), 
to_sfixed(-965046557.0/4294967296.0,1,-nbitq), 
to_sfixed(451897671.0/4294967296.0,1,-nbitq), 
to_sfixed(58562157.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-2095735682.0/4294967296.0,1,-nbitq), 
to_sfixed(307596888.0/4294967296.0,1,-nbitq), 
to_sfixed(-1032930084.0/4294967296.0,1,-nbitq), 
to_sfixed(-343126443.0/4294967296.0,1,-nbitq), 
to_sfixed(1272250385.0/4294967296.0,1,-nbitq), 
to_sfixed(346674424.0/4294967296.0,1,-nbitq), 
to_sfixed(942945781.0/4294967296.0,1,-nbitq), 
to_sfixed(493369020.0/4294967296.0,1,-nbitq), 
to_sfixed(566056334.0/4294967296.0,1,-nbitq), 
to_sfixed(-1114598957.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(1410911983.0/4294967296.0,1,-nbitq), 
to_sfixed(-699658224.0/4294967296.0,1,-nbitq), 
to_sfixed(-960266231.0/4294967296.0,1,-nbitq), 
to_sfixed(-882161475.0/4294967296.0,1,-nbitq), 
to_sfixed(-841441916.0/4294967296.0,1,-nbitq), 
to_sfixed(761791239.0/4294967296.0,1,-nbitq), 
to_sfixed(-982555444.0/4294967296.0,1,-nbitq), 
to_sfixed(559297291.0/4294967296.0,1,-nbitq), 
to_sfixed(-1762880303.0/4294967296.0,1,-nbitq), 
to_sfixed(1405402072.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-1169354486.0/4294967296.0,1,-nbitq), 
to_sfixed(-496032716.0/4294967296.0,1,-nbitq), 
to_sfixed(-911798258.0/4294967296.0,1,-nbitq), 
to_sfixed(886004742.0/4294967296.0,1,-nbitq), 
to_sfixed(-1711367841.0/4294967296.0,1,-nbitq), 
to_sfixed(447747492.0/4294967296.0,1,-nbitq), 
to_sfixed(164371606.0/4294967296.0,1,-nbitq), 
to_sfixed(1232799168.0/4294967296.0,1,-nbitq), 
to_sfixed(1245059603.0/4294967296.0,1,-nbitq), 
to_sfixed(471958268.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-1417253970.0/4294967296.0,1,-nbitq), 
to_sfixed(1192336948.0/4294967296.0,1,-nbitq), 
to_sfixed(-958982477.0/4294967296.0,1,-nbitq), 
to_sfixed(-1061091188.0/4294967296.0,1,-nbitq), 
to_sfixed(1572037183.0/4294967296.0,1,-nbitq), 
to_sfixed(1550357536.0/4294967296.0,1,-nbitq), 
to_sfixed(467942608.0/4294967296.0,1,-nbitq), 
to_sfixed(1567763464.0/4294967296.0,1,-nbitq), 
to_sfixed(513897296.0/4294967296.0,1,-nbitq), 
to_sfixed(-729016063.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(68219442.0/4294967296.0,1,-nbitq), 
to_sfixed(-1108985754.0/4294967296.0,1,-nbitq), 
to_sfixed(234200400.0/4294967296.0,1,-nbitq), 
to_sfixed(454696051.0/4294967296.0,1,-nbitq), 
to_sfixed(1529512585.0/4294967296.0,1,-nbitq), 
to_sfixed(757386066.0/4294967296.0,1,-nbitq), 
to_sfixed(-1272410900.0/4294967296.0,1,-nbitq), 
to_sfixed(905339295.0/4294967296.0,1,-nbitq), 
to_sfixed(-1887856630.0/4294967296.0,1,-nbitq), 
to_sfixed(1441971657.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-244878179.0/4294967296.0,1,-nbitq), 
to_sfixed(-518884873.0/4294967296.0,1,-nbitq), 
to_sfixed(-604214274.0/4294967296.0,1,-nbitq), 
to_sfixed(-590445902.0/4294967296.0,1,-nbitq), 
to_sfixed(518118482.0/4294967296.0,1,-nbitq), 
to_sfixed(1358320537.0/4294967296.0,1,-nbitq), 
to_sfixed(253299071.0/4294967296.0,1,-nbitq), 
to_sfixed(-235351585.0/4294967296.0,1,-nbitq), 
to_sfixed(-775553509.0/4294967296.0,1,-nbitq), 
to_sfixed(-445640893.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-307358763.0/4294967296.0,1,-nbitq), 
to_sfixed(453201554.0/4294967296.0,1,-nbitq), 
to_sfixed(-974377505.0/4294967296.0,1,-nbitq), 
to_sfixed(-651531775.0/4294967296.0,1,-nbitq), 
to_sfixed(-240948423.0/4294967296.0,1,-nbitq), 
to_sfixed(369677880.0/4294967296.0,1,-nbitq), 
to_sfixed(-1110268130.0/4294967296.0,1,-nbitq), 
to_sfixed(1143321556.0/4294967296.0,1,-nbitq), 
to_sfixed(1235305381.0/4294967296.0,1,-nbitq), 
to_sfixed(-884665984.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(1391491287.0/4294967296.0,1,-nbitq), 
to_sfixed(-179780311.0/4294967296.0,1,-nbitq), 
to_sfixed(-1082749470.0/4294967296.0,1,-nbitq), 
to_sfixed(204988447.0/4294967296.0,1,-nbitq), 
to_sfixed(591404682.0/4294967296.0,1,-nbitq), 
to_sfixed(-769898983.0/4294967296.0,1,-nbitq), 
to_sfixed(-547030439.0/4294967296.0,1,-nbitq), 
to_sfixed(59112352.0/4294967296.0,1,-nbitq), 
to_sfixed(-980736425.0/4294967296.0,1,-nbitq), 
to_sfixed(-819701707.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-2188852662.0/4294967296.0,1,-nbitq), 
to_sfixed(332264810.0/4294967296.0,1,-nbitq), 
to_sfixed(498527989.0/4294967296.0,1,-nbitq), 
to_sfixed(319060200.0/4294967296.0,1,-nbitq), 
to_sfixed(-1552961514.0/4294967296.0,1,-nbitq), 
to_sfixed(136423230.0/4294967296.0,1,-nbitq), 
to_sfixed(995377419.0/4294967296.0,1,-nbitq), 
to_sfixed(573375988.0/4294967296.0,1,-nbitq), 
to_sfixed(-1234116701.0/4294967296.0,1,-nbitq), 
to_sfixed(-1195709081.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-998444241.0/4294967296.0,1,-nbitq), 
to_sfixed(-25968131.0/4294967296.0,1,-nbitq), 
to_sfixed(727337886.0/4294967296.0,1,-nbitq), 
to_sfixed(-824142983.0/4294967296.0,1,-nbitq), 
to_sfixed(-623398085.0/4294967296.0,1,-nbitq), 
to_sfixed(913271759.0/4294967296.0,1,-nbitq), 
to_sfixed(1439503778.0/4294967296.0,1,-nbitq), 
to_sfixed(-536194890.0/4294967296.0,1,-nbitq), 
to_sfixed(-7713172.0/4294967296.0,1,-nbitq), 
to_sfixed(-924148955.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(965766931.0/4294967296.0,1,-nbitq), 
to_sfixed(-1509829932.0/4294967296.0,1,-nbitq), 
to_sfixed(-790268073.0/4294967296.0,1,-nbitq), 
to_sfixed(155465663.0/4294967296.0,1,-nbitq), 
to_sfixed(-638590199.0/4294967296.0,1,-nbitq), 
to_sfixed(-533845429.0/4294967296.0,1,-nbitq), 
to_sfixed(364681333.0/4294967296.0,1,-nbitq), 
to_sfixed(797159541.0/4294967296.0,1,-nbitq), 
to_sfixed(955912538.0/4294967296.0,1,-nbitq), 
to_sfixed(-1016575807.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(1339874741.0/4294967296.0,1,-nbitq), 
to_sfixed(1001440369.0/4294967296.0,1,-nbitq), 
to_sfixed(-1052865777.0/4294967296.0,1,-nbitq), 
to_sfixed(418099158.0/4294967296.0,1,-nbitq), 
to_sfixed(1003372266.0/4294967296.0,1,-nbitq), 
to_sfixed(-1011232890.0/4294967296.0,1,-nbitq), 
to_sfixed(-805172130.0/4294967296.0,1,-nbitq), 
to_sfixed(-41918936.0/4294967296.0,1,-nbitq), 
to_sfixed(816665072.0/4294967296.0,1,-nbitq), 
to_sfixed(130470109.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-642637569.0/4294967296.0,1,-nbitq), 
to_sfixed(73077305.0/4294967296.0,1,-nbitq), 
to_sfixed(-306430737.0/4294967296.0,1,-nbitq), 
to_sfixed(-863443365.0/4294967296.0,1,-nbitq), 
to_sfixed(-875701935.0/4294967296.0,1,-nbitq), 
to_sfixed(-749155805.0/4294967296.0,1,-nbitq), 
to_sfixed(98860791.0/4294967296.0,1,-nbitq), 
to_sfixed(782429383.0/4294967296.0,1,-nbitq), 
to_sfixed(-239972140.0/4294967296.0,1,-nbitq), 
to_sfixed(-482680283.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-459412992.0/4294967296.0,1,-nbitq), 
to_sfixed(-204716491.0/4294967296.0,1,-nbitq), 
to_sfixed(791653885.0/4294967296.0,1,-nbitq), 
to_sfixed(-538884521.0/4294967296.0,1,-nbitq), 
to_sfixed(-179093601.0/4294967296.0,1,-nbitq), 
to_sfixed(-770672645.0/4294967296.0,1,-nbitq), 
to_sfixed(-1806336998.0/4294967296.0,1,-nbitq), 
to_sfixed(430631758.0/4294967296.0,1,-nbitq), 
to_sfixed(-504616525.0/4294967296.0,1,-nbitq), 
to_sfixed(-507252424.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(443848988.0/4294967296.0,1,-nbitq), 
to_sfixed(-418472903.0/4294967296.0,1,-nbitq), 
to_sfixed(-81546796.0/4294967296.0,1,-nbitq), 
to_sfixed(-479216620.0/4294967296.0,1,-nbitq), 
to_sfixed(-1123799370.0/4294967296.0,1,-nbitq), 
to_sfixed(-979854049.0/4294967296.0,1,-nbitq), 
to_sfixed(372944842.0/4294967296.0,1,-nbitq), 
to_sfixed(195002057.0/4294967296.0,1,-nbitq), 
to_sfixed(-1426717454.0/4294967296.0,1,-nbitq), 
to_sfixed(-1736956060.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(797882238.0/4294967296.0,1,-nbitq), 
to_sfixed(1260176401.0/4294967296.0,1,-nbitq), 
to_sfixed(-321782427.0/4294967296.0,1,-nbitq), 
to_sfixed(1266282021.0/4294967296.0,1,-nbitq), 
to_sfixed(1228315852.0/4294967296.0,1,-nbitq), 
to_sfixed(140907911.0/4294967296.0,1,-nbitq), 
to_sfixed(270381890.0/4294967296.0,1,-nbitq), 
to_sfixed(-898680557.0/4294967296.0,1,-nbitq), 
to_sfixed(-642369528.0/4294967296.0,1,-nbitq), 
to_sfixed(-1384885843.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(721237192.0/4294967296.0,1,-nbitq), 
to_sfixed(389335052.0/4294967296.0,1,-nbitq), 
to_sfixed(-963073893.0/4294967296.0,1,-nbitq), 
to_sfixed(1293463030.0/4294967296.0,1,-nbitq), 
to_sfixed(732209390.0/4294967296.0,1,-nbitq), 
to_sfixed(886722805.0/4294967296.0,1,-nbitq), 
to_sfixed(283192735.0/4294967296.0,1,-nbitq), 
to_sfixed(-954817343.0/4294967296.0,1,-nbitq), 
to_sfixed(-1895885541.0/4294967296.0,1,-nbitq), 
to_sfixed(-450313392.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(79167939.0/4294967296.0,1,-nbitq), 
to_sfixed(717130179.0/4294967296.0,1,-nbitq), 
to_sfixed(488067592.0/4294967296.0,1,-nbitq), 
to_sfixed(-410627719.0/4294967296.0,1,-nbitq), 
to_sfixed(787967063.0/4294967296.0,1,-nbitq), 
to_sfixed(-1096380682.0/4294967296.0,1,-nbitq), 
to_sfixed(288999286.0/4294967296.0,1,-nbitq), 
to_sfixed(-45606777.0/4294967296.0,1,-nbitq), 
to_sfixed(-1631416459.0/4294967296.0,1,-nbitq), 
to_sfixed(992612841.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(395003319.0/4294967296.0,1,-nbitq), 
to_sfixed(846977384.0/4294967296.0,1,-nbitq), 
to_sfixed(1156215808.0/4294967296.0,1,-nbitq), 
to_sfixed(-1118651797.0/4294967296.0,1,-nbitq), 
to_sfixed(101068275.0/4294967296.0,1,-nbitq), 
to_sfixed(886545464.0/4294967296.0,1,-nbitq), 
to_sfixed(325237571.0/4294967296.0,1,-nbitq), 
to_sfixed(-1119462246.0/4294967296.0,1,-nbitq), 
to_sfixed(-1002458802.0/4294967296.0,1,-nbitq), 
to_sfixed(-1114267629.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-39595001.0/4294967296.0,1,-nbitq), 
to_sfixed(-608444704.0/4294967296.0,1,-nbitq), 
to_sfixed(-228134830.0/4294967296.0,1,-nbitq), 
to_sfixed(517568123.0/4294967296.0,1,-nbitq), 
to_sfixed(-37232471.0/4294967296.0,1,-nbitq), 
to_sfixed(-179968320.0/4294967296.0,1,-nbitq), 
to_sfixed(272417410.0/4294967296.0,1,-nbitq), 
to_sfixed(109372558.0/4294967296.0,1,-nbitq), 
to_sfixed(-850415195.0/4294967296.0,1,-nbitq), 
to_sfixed(360317394.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-583439429.0/4294967296.0,1,-nbitq), 
to_sfixed(-1049822742.0/4294967296.0,1,-nbitq), 
to_sfixed(1315940606.0/4294967296.0,1,-nbitq), 
to_sfixed(-1014085080.0/4294967296.0,1,-nbitq), 
to_sfixed(1556935.0/4294967296.0,1,-nbitq), 
to_sfixed(-818469110.0/4294967296.0,1,-nbitq), 
to_sfixed(1159378501.0/4294967296.0,1,-nbitq), 
to_sfixed(777019553.0/4294967296.0,1,-nbitq), 
to_sfixed(482529581.0/4294967296.0,1,-nbitq), 
to_sfixed(-671354441.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(106575840.0/4294967296.0,1,-nbitq), 
to_sfixed(464179102.0/4294967296.0,1,-nbitq), 
to_sfixed(-491485483.0/4294967296.0,1,-nbitq), 
to_sfixed(1044489648.0/4294967296.0,1,-nbitq), 
to_sfixed(1088549206.0/4294967296.0,1,-nbitq), 
to_sfixed(480672769.0/4294967296.0,1,-nbitq), 
to_sfixed(-7931600.0/4294967296.0,1,-nbitq), 
to_sfixed(-1168470915.0/4294967296.0,1,-nbitq), 
to_sfixed(347909923.0/4294967296.0,1,-nbitq), 
to_sfixed(323137680.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(213946185.0/4294967296.0,1,-nbitq), 
to_sfixed(220748210.0/4294967296.0,1,-nbitq), 
to_sfixed(1986200501.0/4294967296.0,1,-nbitq), 
to_sfixed(973533229.0/4294967296.0,1,-nbitq), 
to_sfixed(-315531571.0/4294967296.0,1,-nbitq), 
to_sfixed(-1008974837.0/4294967296.0,1,-nbitq), 
to_sfixed(-1080879823.0/4294967296.0,1,-nbitq), 
to_sfixed(-1249281001.0/4294967296.0,1,-nbitq), 
to_sfixed(402896469.0/4294967296.0,1,-nbitq), 
to_sfixed(-816189574.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-400209534.0/4294967296.0,1,-nbitq), 
to_sfixed(507757491.0/4294967296.0,1,-nbitq), 
to_sfixed(-312234281.0/4294967296.0,1,-nbitq), 
to_sfixed(-40792828.0/4294967296.0,1,-nbitq), 
to_sfixed(-1175723607.0/4294967296.0,1,-nbitq), 
to_sfixed(-1107287709.0/4294967296.0,1,-nbitq), 
to_sfixed(121125267.0/4294967296.0,1,-nbitq), 
to_sfixed(-681601319.0/4294967296.0,1,-nbitq), 
to_sfixed(692126442.0/4294967296.0,1,-nbitq), 
to_sfixed(964502448.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(1149114805.0/4294967296.0,1,-nbitq), 
to_sfixed(747060164.0/4294967296.0,1,-nbitq), 
to_sfixed(264186055.0/4294967296.0,1,-nbitq), 
to_sfixed(-355406485.0/4294967296.0,1,-nbitq), 
to_sfixed(839125242.0/4294967296.0,1,-nbitq), 
to_sfixed(-1194640461.0/4294967296.0,1,-nbitq), 
to_sfixed(818695115.0/4294967296.0,1,-nbitq), 
to_sfixed(792920992.0/4294967296.0,1,-nbitq), 
to_sfixed(511121817.0/4294967296.0,1,-nbitq), 
to_sfixed(-95506318.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-1195629042.0/4294967296.0,1,-nbitq), 
to_sfixed(180313211.0/4294967296.0,1,-nbitq), 
to_sfixed(1302980012.0/4294967296.0,1,-nbitq), 
to_sfixed(315922560.0/4294967296.0,1,-nbitq), 
to_sfixed(-1162298173.0/4294967296.0,1,-nbitq), 
to_sfixed(1174682893.0/4294967296.0,1,-nbitq), 
to_sfixed(-1304977383.0/4294967296.0,1,-nbitq), 
to_sfixed(-1245306624.0/4294967296.0,1,-nbitq), 
to_sfixed(823886303.0/4294967296.0,1,-nbitq), 
to_sfixed(584673484.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(838353311.0/4294967296.0,1,-nbitq), 
to_sfixed(-878007390.0/4294967296.0,1,-nbitq), 
to_sfixed(32971386.0/4294967296.0,1,-nbitq), 
to_sfixed(1320263746.0/4294967296.0,1,-nbitq), 
to_sfixed(727417398.0/4294967296.0,1,-nbitq), 
to_sfixed(580411934.0/4294967296.0,1,-nbitq), 
to_sfixed(1276621630.0/4294967296.0,1,-nbitq), 
to_sfixed(-247286161.0/4294967296.0,1,-nbitq), 
to_sfixed(-1305350259.0/4294967296.0,1,-nbitq), 
to_sfixed(12215060.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(262829814.0/4294967296.0,1,-nbitq), 
to_sfixed(-555519607.0/4294967296.0,1,-nbitq), 
to_sfixed(1075143846.0/4294967296.0,1,-nbitq), 
to_sfixed(1147783279.0/4294967296.0,1,-nbitq), 
to_sfixed(186502505.0/4294967296.0,1,-nbitq), 
to_sfixed(1568811037.0/4294967296.0,1,-nbitq), 
to_sfixed(-259770412.0/4294967296.0,1,-nbitq), 
to_sfixed(999631690.0/4294967296.0,1,-nbitq), 
to_sfixed(-990695264.0/4294967296.0,1,-nbitq), 
to_sfixed(-1909030230.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-203700821.0/4294967296.0,1,-nbitq), 
to_sfixed(-154898498.0/4294967296.0,1,-nbitq), 
to_sfixed(1236074099.0/4294967296.0,1,-nbitq), 
to_sfixed(-273763503.0/4294967296.0,1,-nbitq), 
to_sfixed(531454040.0/4294967296.0,1,-nbitq), 
to_sfixed(-1271173183.0/4294967296.0,1,-nbitq), 
to_sfixed(840894505.0/4294967296.0,1,-nbitq), 
to_sfixed(-269484454.0/4294967296.0,1,-nbitq), 
to_sfixed(-439469206.0/4294967296.0,1,-nbitq), 
to_sfixed(738125453.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-191397610.0/4294967296.0,1,-nbitq), 
to_sfixed(85797766.0/4294967296.0,1,-nbitq), 
to_sfixed(1434262122.0/4294967296.0,1,-nbitq), 
to_sfixed(952161321.0/4294967296.0,1,-nbitq), 
to_sfixed(66199310.0/4294967296.0,1,-nbitq), 
to_sfixed(-930525167.0/4294967296.0,1,-nbitq), 
to_sfixed(96847946.0/4294967296.0,1,-nbitq), 
to_sfixed(-1004847862.0/4294967296.0,1,-nbitq), 
to_sfixed(1067766509.0/4294967296.0,1,-nbitq), 
to_sfixed(736141005.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(657247924.0/4294967296.0,1,-nbitq), 
to_sfixed(456483261.0/4294967296.0,1,-nbitq), 
to_sfixed(-12733777.0/4294967296.0,1,-nbitq), 
to_sfixed(-1431953666.0/4294967296.0,1,-nbitq), 
to_sfixed(-567345251.0/4294967296.0,1,-nbitq), 
to_sfixed(-233215701.0/4294967296.0,1,-nbitq), 
to_sfixed(-667004941.0/4294967296.0,1,-nbitq), 
to_sfixed(886761049.0/4294967296.0,1,-nbitq), 
to_sfixed(935715390.0/4294967296.0,1,-nbitq), 
to_sfixed(-175436240.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(134279748.0/4294967296.0,1,-nbitq), 
to_sfixed(391611466.0/4294967296.0,1,-nbitq), 
to_sfixed(-451427631.0/4294967296.0,1,-nbitq), 
to_sfixed(796570189.0/4294967296.0,1,-nbitq), 
to_sfixed(194108147.0/4294967296.0,1,-nbitq), 
to_sfixed(-120024414.0/4294967296.0,1,-nbitq), 
to_sfixed(-83822262.0/4294967296.0,1,-nbitq), 
to_sfixed(-201766250.0/4294967296.0,1,-nbitq), 
to_sfixed(-87909127.0/4294967296.0,1,-nbitq), 
to_sfixed(-428449010.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-663863538.0/4294967296.0,1,-nbitq), 
to_sfixed(-233311948.0/4294967296.0,1,-nbitq), 
to_sfixed(-702440199.0/4294967296.0,1,-nbitq), 
to_sfixed(377495986.0/4294967296.0,1,-nbitq), 
to_sfixed(-874402840.0/4294967296.0,1,-nbitq), 
to_sfixed(394475522.0/4294967296.0,1,-nbitq), 
to_sfixed(-741501067.0/4294967296.0,1,-nbitq), 
to_sfixed(1142612157.0/4294967296.0,1,-nbitq), 
to_sfixed(-838964181.0/4294967296.0,1,-nbitq), 
to_sfixed(-289980471.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-317852182.0/4294967296.0,1,-nbitq), 
to_sfixed(321139865.0/4294967296.0,1,-nbitq), 
to_sfixed(-794436437.0/4294967296.0,1,-nbitq), 
to_sfixed(444412197.0/4294967296.0,1,-nbitq), 
to_sfixed(-565630953.0/4294967296.0,1,-nbitq), 
to_sfixed(-1018971891.0/4294967296.0,1,-nbitq), 
to_sfixed(-533557379.0/4294967296.0,1,-nbitq), 
to_sfixed(169626857.0/4294967296.0,1,-nbitq), 
to_sfixed(40268230.0/4294967296.0,1,-nbitq), 
to_sfixed(371503686.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(1120523551.0/4294967296.0,1,-nbitq), 
to_sfixed(-731203944.0/4294967296.0,1,-nbitq), 
to_sfixed(-1581775411.0/4294967296.0,1,-nbitq), 
to_sfixed(44847142.0/4294967296.0,1,-nbitq), 
to_sfixed(-895846647.0/4294967296.0,1,-nbitq), 
to_sfixed(-714489636.0/4294967296.0,1,-nbitq), 
to_sfixed(-428640722.0/4294967296.0,1,-nbitq), 
to_sfixed(-883480610.0/4294967296.0,1,-nbitq), 
to_sfixed(-137323975.0/4294967296.0,1,-nbitq), 
to_sfixed(-829781859.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(998240906.0/4294967296.0,1,-nbitq), 
to_sfixed(-1445069213.0/4294967296.0,1,-nbitq), 
to_sfixed(-1100602241.0/4294967296.0,1,-nbitq), 
to_sfixed(-114218302.0/4294967296.0,1,-nbitq), 
to_sfixed(772299114.0/4294967296.0,1,-nbitq), 
to_sfixed(1415216769.0/4294967296.0,1,-nbitq), 
to_sfixed(-919164792.0/4294967296.0,1,-nbitq), 
to_sfixed(461480726.0/4294967296.0,1,-nbitq), 
to_sfixed(523489703.0/4294967296.0,1,-nbitq), 
to_sfixed(399720370.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-391823085.0/4294967296.0,1,-nbitq), 
to_sfixed(1158849258.0/4294967296.0,1,-nbitq), 
to_sfixed(-907186495.0/4294967296.0,1,-nbitq), 
to_sfixed(695450536.0/4294967296.0,1,-nbitq), 
to_sfixed(-1040016417.0/4294967296.0,1,-nbitq), 
to_sfixed(-445414905.0/4294967296.0,1,-nbitq), 
to_sfixed(-509725126.0/4294967296.0,1,-nbitq), 
to_sfixed(1581540461.0/4294967296.0,1,-nbitq), 
to_sfixed(-89761985.0/4294967296.0,1,-nbitq), 
to_sfixed(-16803626.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(1129112607.0/4294967296.0,1,-nbitq), 
to_sfixed(-120243808.0/4294967296.0,1,-nbitq), 
to_sfixed(234236890.0/4294967296.0,1,-nbitq), 
to_sfixed(-555100450.0/4294967296.0,1,-nbitq), 
to_sfixed(290383699.0/4294967296.0,1,-nbitq), 
to_sfixed(306138328.0/4294967296.0,1,-nbitq), 
to_sfixed(1049506435.0/4294967296.0,1,-nbitq), 
to_sfixed(-1055217111.0/4294967296.0,1,-nbitq), 
to_sfixed(-489372058.0/4294967296.0,1,-nbitq), 
to_sfixed(-685421738.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(203688173.0/4294967296.0,1,-nbitq), 
to_sfixed(-894955781.0/4294967296.0,1,-nbitq), 
to_sfixed(544492935.0/4294967296.0,1,-nbitq), 
to_sfixed(-705116346.0/4294967296.0,1,-nbitq), 
to_sfixed(-44755640.0/4294967296.0,1,-nbitq), 
to_sfixed(-276291500.0/4294967296.0,1,-nbitq), 
to_sfixed(-883208301.0/4294967296.0,1,-nbitq), 
to_sfixed(873099501.0/4294967296.0,1,-nbitq), 
to_sfixed(284965735.0/4294967296.0,1,-nbitq), 
to_sfixed(750120168.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(2219625653.0/4294967296.0,1,-nbitq), 
to_sfixed(-1915848674.0/4294967296.0,1,-nbitq), 
to_sfixed(1252779977.0/4294967296.0,1,-nbitq), 
to_sfixed(1338054385.0/4294967296.0,1,-nbitq), 
to_sfixed(-1888651873.0/4294967296.0,1,-nbitq), 
to_sfixed(-1152389035.0/4294967296.0,1,-nbitq), 
to_sfixed(-1014560311.0/4294967296.0,1,-nbitq), 
to_sfixed(-1285086929.0/4294967296.0,1,-nbitq), 
to_sfixed(4080540.0/4294967296.0,1,-nbitq), 
to_sfixed(1769782401.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-91405190.0/4294967296.0,1,-nbitq), 
to_sfixed(312825944.0/4294967296.0,1,-nbitq), 
to_sfixed(-18740514.0/4294967296.0,1,-nbitq), 
to_sfixed(243158280.0/4294967296.0,1,-nbitq), 
to_sfixed(-623517538.0/4294967296.0,1,-nbitq), 
to_sfixed(1899366586.0/4294967296.0,1,-nbitq), 
to_sfixed(-1624652682.0/4294967296.0,1,-nbitq), 
to_sfixed(426887179.0/4294967296.0,1,-nbitq), 
to_sfixed(-675876963.0/4294967296.0,1,-nbitq), 
to_sfixed(-873876018.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(737296861.0/4294967296.0,1,-nbitq), 
to_sfixed(945623640.0/4294967296.0,1,-nbitq), 
to_sfixed(-777639363.0/4294967296.0,1,-nbitq), 
to_sfixed(824281123.0/4294967296.0,1,-nbitq), 
to_sfixed(195822905.0/4294967296.0,1,-nbitq), 
to_sfixed(178109259.0/4294967296.0,1,-nbitq), 
to_sfixed(-740295505.0/4294967296.0,1,-nbitq), 
to_sfixed(-558441444.0/4294967296.0,1,-nbitq), 
to_sfixed(247492564.0/4294967296.0,1,-nbitq), 
to_sfixed(1000025759.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-786598726.0/4294967296.0,1,-nbitq), 
to_sfixed(-1662094370.0/4294967296.0,1,-nbitq), 
to_sfixed(311591769.0/4294967296.0,1,-nbitq), 
to_sfixed(776928438.0/4294967296.0,1,-nbitq), 
to_sfixed(-973241814.0/4294967296.0,1,-nbitq), 
to_sfixed(1069111593.0/4294967296.0,1,-nbitq), 
to_sfixed(734339777.0/4294967296.0,1,-nbitq), 
to_sfixed(268687110.0/4294967296.0,1,-nbitq), 
to_sfixed(1627808017.0/4294967296.0,1,-nbitq), 
to_sfixed(764211718.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-562836800.0/4294967296.0,1,-nbitq), 
to_sfixed(-931611205.0/4294967296.0,1,-nbitq), 
to_sfixed(-961195560.0/4294967296.0,1,-nbitq), 
to_sfixed(443652156.0/4294967296.0,1,-nbitq), 
to_sfixed(-1199488588.0/4294967296.0,1,-nbitq), 
to_sfixed(904528448.0/4294967296.0,1,-nbitq), 
to_sfixed(-172960197.0/4294967296.0,1,-nbitq), 
to_sfixed(2100028974.0/4294967296.0,1,-nbitq), 
to_sfixed(-178516578.0/4294967296.0,1,-nbitq), 
to_sfixed(115621978.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(950827032.0/4294967296.0,1,-nbitq), 
to_sfixed(308192011.0/4294967296.0,1,-nbitq), 
to_sfixed(-545119355.0/4294967296.0,1,-nbitq), 
to_sfixed(413624063.0/4294967296.0,1,-nbitq), 
to_sfixed(488531317.0/4294967296.0,1,-nbitq), 
to_sfixed(773776687.0/4294967296.0,1,-nbitq), 
to_sfixed(716441261.0/4294967296.0,1,-nbitq), 
to_sfixed(417538015.0/4294967296.0,1,-nbitq), 
to_sfixed(-1018503848.0/4294967296.0,1,-nbitq), 
to_sfixed(-239449559.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-1603022977.0/4294967296.0,1,-nbitq), 
to_sfixed(686775165.0/4294967296.0,1,-nbitq), 
to_sfixed(-190229460.0/4294967296.0,1,-nbitq), 
to_sfixed(-1300803965.0/4294967296.0,1,-nbitq), 
to_sfixed(-358902312.0/4294967296.0,1,-nbitq), 
to_sfixed(335550156.0/4294967296.0,1,-nbitq), 
to_sfixed(-965076761.0/4294967296.0,1,-nbitq), 
to_sfixed(-421463082.0/4294967296.0,1,-nbitq), 
to_sfixed(1244351412.0/4294967296.0,1,-nbitq), 
to_sfixed(1157220713.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(369658475.0/4294967296.0,1,-nbitq), 
to_sfixed(711422544.0/4294967296.0,1,-nbitq), 
to_sfixed(-50748442.0/4294967296.0,1,-nbitq), 
to_sfixed(603509935.0/4294967296.0,1,-nbitq), 
to_sfixed(820736842.0/4294967296.0,1,-nbitq), 
to_sfixed(-829421680.0/4294967296.0,1,-nbitq), 
to_sfixed(-225596213.0/4294967296.0,1,-nbitq), 
to_sfixed(530586534.0/4294967296.0,1,-nbitq), 
to_sfixed(-813880989.0/4294967296.0,1,-nbitq), 
to_sfixed(629228631.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(679668017.0/4294967296.0,1,-nbitq), 
to_sfixed(-905831244.0/4294967296.0,1,-nbitq), 
to_sfixed(-587089814.0/4294967296.0,1,-nbitq), 
to_sfixed(-1046894416.0/4294967296.0,1,-nbitq), 
to_sfixed(-59681453.0/4294967296.0,1,-nbitq), 
to_sfixed(-87766028.0/4294967296.0,1,-nbitq), 
to_sfixed(713027262.0/4294967296.0,1,-nbitq), 
to_sfixed(-786646086.0/4294967296.0,1,-nbitq), 
to_sfixed(947898006.0/4294967296.0,1,-nbitq), 
to_sfixed(-320234202.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(710421428.0/4294967296.0,1,-nbitq), 
to_sfixed(-1256756064.0/4294967296.0,1,-nbitq), 
to_sfixed(-1450119962.0/4294967296.0,1,-nbitq), 
to_sfixed(-550904379.0/4294967296.0,1,-nbitq), 
to_sfixed(-236128983.0/4294967296.0,1,-nbitq), 
to_sfixed(1305113264.0/4294967296.0,1,-nbitq), 
to_sfixed(956212842.0/4294967296.0,1,-nbitq), 
to_sfixed(-581370387.0/4294967296.0,1,-nbitq), 
to_sfixed(572824807.0/4294967296.0,1,-nbitq), 
to_sfixed(744128258.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(-468392431.0/4294967296.0,1,-nbitq), 
to_sfixed(574076521.0/4294967296.0,1,-nbitq), 
to_sfixed(1184926321.0/4294967296.0,1,-nbitq), 
to_sfixed(-637384917.0/4294967296.0,1,-nbitq), 
to_sfixed(-888275719.0/4294967296.0,1,-nbitq), 
to_sfixed(-1920574403.0/4294967296.0,1,-nbitq), 
to_sfixed(924627810.0/4294967296.0,1,-nbitq), 
to_sfixed(-971506202.0/4294967296.0,1,-nbitq), 
to_sfixed(-1431529258.0/4294967296.0,1,-nbitq), 
to_sfixed(-619712604.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(505454804.0/4294967296.0,1,-nbitq), 
to_sfixed(627475243.0/4294967296.0,1,-nbitq), 
to_sfixed(220449406.0/4294967296.0,1,-nbitq), 
to_sfixed(100548409.0/4294967296.0,1,-nbitq), 
to_sfixed(-936769918.0/4294967296.0,1,-nbitq), 
to_sfixed(841801676.0/4294967296.0,1,-nbitq), 
to_sfixed(887363081.0/4294967296.0,1,-nbitq), 
to_sfixed(469039882.0/4294967296.0,1,-nbitq), 
to_sfixed(648720101.0/4294967296.0,1,-nbitq), 
to_sfixed(-151125614.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(1077519827.0/4294967296.0,1,-nbitq), 
to_sfixed(639105248.0/4294967296.0,1,-nbitq), 
to_sfixed(-871060534.0/4294967296.0,1,-nbitq), 
to_sfixed(407027695.0/4294967296.0,1,-nbitq), 
to_sfixed(-1338026190.0/4294967296.0,1,-nbitq), 
to_sfixed(1092873630.0/4294967296.0,1,-nbitq), 
to_sfixed(593598906.0/4294967296.0,1,-nbitq), 
to_sfixed(-673593459.0/4294967296.0,1,-nbitq), 
to_sfixed(-804215026.0/4294967296.0,1,-nbitq), 
to_sfixed(1302968502.0/4294967296.0,1,-nbitq)  ), 
( to_sfixed(464710766.0/4294967296.0,1,-nbitq), 
to_sfixed(-130348645.0/4294967296.0,1,-nbitq), 
to_sfixed(-521694683.0/4294967296.0,1,-nbitq), 
to_sfixed(-694275462.0/4294967296.0,1,-nbitq), 
to_sfixed(-10316148.0/4294967296.0,1,-nbitq), 
to_sfixed(-413227483.0/4294967296.0,1,-nbitq), 
to_sfixed(560102646.0/4294967296.0,1,-nbitq), 
to_sfixed(1070252290.0/4294967296.0,1,-nbitq), 
to_sfixed(-88633277.0/4294967296.0,1,-nbitq), 
to_sfixed(253096180.0/4294967296.0,1,-nbitq)  ) 
 ) ;

end package coeff;